

module iir_core_obf(inData, clk, reset, outData);
  input [31:0] inData;
  input clk, reset;
  output [31:0] outData;
  wire [31:0] inData;
  wire clk, reset;
  wire [31:0] outData;
  wire __0, __9_, __9_00, __9_00__29804, __9_00__29896, __9_00__29993,
       __9_00__30083, __9_00__30177;
  wire __9_00__30272, __9_00__30366, __9_0_, __9_0___29724,
       __9_0___29725, __9_0___29726, __9_0___29727, __9_0___29728;
  wire __9_0___29729, __9_0___29805, __9_0___29806, __9_0___29807,
       __9_0___29808, __9_0___29809, __9_0___29810, __9_0___29811;
  wire __9_0___29812, __9_0___29897, __9_0___29898, __9_0___29899,
       __9_0___29900, __9_0___29901, __9_0___29902, __9_0___29903;
  wire __9_0___29904, __9_0___29994, __9_0___29995, __9_0___29996,
       __9_0___29997, __9_0___29998, __9_0___29999, __9_0___30000;
  wire __9_0___30001, __9_0___30084, __9_0___30085, __9_0___30086,
       __9_0___30087, __9_0___30088, __9_0___30089, __9_0___30090;
  wire __9_0___30091, __9_0___30178, __9_0___30179, __9_0___30180,
       __9_0___30181, __9_0___30182, __9_0___30183, __9_0___30184;
  wire __9_0___30273, __9_0___30274, __9_0___30275, __9_0___30276,
       __9_0___30277, __9_0___30278, __9_0___30279, __9_0___30280;
  wire __9_0___30367, __9_0___30368, __9_0___30369, __9_0___30370,
       __9_0___30371, __9_0___30372, __9_0___30373, __9_09;
  wire __9_09__29813, __9_09__29905, __9_09__30002, __9_09__30092,
       __9_09__30185, __9_09__30281, __9_09__30374, __9_9_;
  wire __9_9___29797, __9_9___29798, __9_9___29799, __9_9___29800,
       __9_9___29801, __9_9___29802, __9_9___29803, __9_9___29888;
  wire __9_9___29889, __9_9___29890, __9_9___29891, __9_9___29892,
       __9_9___29893, __9_9___29894, __9_9___29986, __9_9___29987;
  wire __9_9___29988, __9_9___29989, __9_9___29990, __9_9___29991,
       __9_9___30075, __9_9___30076, __9_9___30077, __9_9___30078;
  wire __9_9___30079, __9_9___30080, __9_9___30081, __9_9___30170,
       __9_9___30171, __9_9___30172, __9_9___30173, __9_9___30174;
  wire __9_9___30175, __9_9___30264, __9_9___30265, __9_9___30266,
       __9_9___30267, __9_9___30268, __9_9___30269, __9_9___30270;
  wire __9_9___30358, __9_9___30359, __9_9___30360, __9_9___30361,
       __9_9___30362, __9_9___30363, __9_9___30364, __9_9___30365;
  wire __9_9___30446, __9_9___30447, __9_9___30448, __9_9___30449,
       __9_9___30450, __9_9___30451, __9_9___30452, __9_9___30453;
  wire __9_90, __9_90__29887, __9_90__29985, __9_90__30074,
       __9_90__30169, __9_90__30263, __9_90__30357, __9_90__30445;
  wire __9_99, __9_99__29895, __9_99__29992, __9_99__30082,
       __9_99__30176, __9_99__30271, __9_99__30454, __9__;
  wire __9__0, __9__0__29744, __9__0__29752, __9__0__29760,
       __9__0__29770, __9__0__29780, __9__0__29789, __9__0__29814;
  wire __9__0__29824, __9__0__29832, __9__0__29841, __9__0__29850,
       __9__0__29868, __9__0__29878, __9__0__29906, __9__0__29916;
  wire __9__0__29926, __9__0__29936, __9__0__29946, __9__0__29956,
       __9__0__29966, __9__0__29975, __9__0__30003, __9__0__30011;
  wire __9__0__30038, __9__0__30048, __9__0__30064, __9__0__30093,
       __9__0__30102, __9__0__30111, __9__0__30120, __9__0__30130;
  wire __9__0__30140, __9__0__30150, __9__0__30159, __9__0__30186,
       __9__0__30196, __9__0__30206, __9__0__30216, __9__0__30226;
  wire __9__0__30234, __9__0__30244, __9__0__30254, __9__0__30282,
       __9__0__30291, __9__0__30310, __9__0__30320, __9__0__30330;
  wire __9__0__30338, __9__0__30347, __9__0__30375, __9__0__30394,
       __9__0__30403, __9__0__30411, __9__0__30420, __9__0__30429;
  wire __9__0__30438, __9__9, __9__9__29743, __9__9__29751,
       __9__9__29759, __9__9__29769, __9__9__29779, __9__9__29788;
  wire __9__9__29796, __9__9__29823, __9__9__29831, __9__9__29840,
       __9__9__29849, __9__9__29859, __9__9__29867, __9__9__29877;
  wire __9__9__29886, __9__9__29915, __9__9__29925, __9__9__29935,
       __9__9__29945, __9__9__29955, __9__9__29965, __9__9__29974;
  wire __9__9__29984, __9__9__30010, __9__9__30020, __9__9__30029,
       __9__9__30047, __9__9__30056, __9__9__30063, __9__9__30073;
  wire __9__9__30101, __9__9__30110, __9__9__30119, __9__9__30129,
       __9__9__30139, __9__9__30149, __9__9__30158, __9__9__30168;
  wire __9__9__30195, __9__9__30205, __9__9__30215, __9__9__30225,
       __9__9__30233, __9__9__30243, __9__9__30253, __9__9__30262;
  wire __9__9__30290, __9__9__30300, __9__9__30309, __9__9__30319,
       __9__9__30329, __9__9__30337, __9__9__30356, __9__9__30384;
  wire __9__9__30393, __9__9__30402, __9__9__30410, __9__9__30419,
       __9__9__30437, __9__9__30444, __9___, __9___22166;
  wire __9___22167, __9___22168, __9___22169, __9____22287,
       __9_____29730, __9_____29731, __9_____29732, __9_____29733;
  wire __9_____29734, __9_____29735, __9_____29736, __9_____29737,
       __9_____29738, __9_____29739, __9_____29740, __9_____29741;
  wire __9_____29742, __9_____29745, __9_____29746, __9_____29747,
       __9_____29748, __9_____29749, __9_____29750, __9_____29753;
  wire __9_____29754, __9_____29755, __9_____29756, __9_____29757,
       __9_____29758, __9_____29761, __9_____29762, __9_____29763;
  wire __9_____29764, __9_____29765, __9_____29766, __9_____29767,
       __9_____29768, __9_____29771, __9_____29772, __9_____29773;
  wire __9_____29774, __9_____29775, __9_____29776, __9_____29777,
       __9_____29778, __9_____29781, __9_____29782, __9_____29783;
  wire __9_____29784, __9_____29785, __9_____29786, __9_____29787,
       __9_____29790, __9_____29791, __9_____29792, __9_____29793;
  wire __9_____29794, __9_____29795, __9_____29815, __9_____29816,
       __9_____29817, __9_____29818, __9_____29819, __9_____29820;
  wire __9_____29821, __9_____29822, __9_____29825, __9_____29826,
       __9_____29827, __9_____29828, __9_____29829, __9_____29830;
  wire __9_____29833, __9_____29834, __9_____29835, __9_____29836,
       __9_____29837, __9_____29838, __9_____29839, __9_____29842;
  wire __9_____29843, __9_____29844, __9_____29845, __9_____29846,
       __9_____29847, __9_____29848, __9_____29851, __9_____29852;
  wire __9_____29853, __9_____29854, __9_____29855, __9_____29856,
       __9_____29857, __9_____29858, __9_____29860, __9_____29861;
  wire __9_____29862, __9_____29863, __9_____29864, __9_____29865,
       __9_____29866, __9_____29869, __9_____29870, __9_____29871;
  wire __9_____29872, __9_____29873, __9_____29874, __9_____29875,
       __9_____29876, __9_____29879, __9_____29880, __9_____29881;
  wire __9_____29882, __9_____29883, __9_____29884, __9_____29885,
       __9_____29907, __9_____29908, __9_____29909, __9_____29910;
  wire __9_____29911, __9_____29912, __9_____29913, __9_____29914,
       __9_____29917, __9_____29918, __9_____29919, __9_____29920;
  wire __9_____29921, __9_____29922, __9_____29923, __9_____29924,
       __9_____29927, __9_____29928, __9_____29929, __9_____29930;
  wire __9_____29931, __9_____29932, __9_____29933, __9_____29934,
       __9_____29937, __9_____29938, __9_____29939, __9_____29940;
  wire __9_____29941, __9_____29942, __9_____29943, __9_____29944,
       __9_____29947, __9_____29948, __9_____29949, __9_____29950;
  wire __9_____29951, __9_____29952, __9_____29953, __9_____29954,
       __9_____29957, __9_____29958, __9_____29959, __9_____29960;
  wire __9_____29961, __9_____29962, __9_____29963, __9_____29964,
       __9_____29967, __9_____29968, __9_____29969, __9_____29970;
  wire __9_____29971, __9_____29972, __9_____29973, __9_____29976,
       __9_____29977, __9_____29978, __9_____29979, __9_____29980;
  wire __9_____29981, __9_____29982, __9_____29983, __9_____30004,
       __9_____30005, __9_____30006, __9_____30007, __9_____30008;
  wire __9_____30009, __9_____30012, __9_____30013, __9_____30014,
       __9_____30015, __9_____30016, __9_____30017, __9_____30018;
  wire __9_____30019, __9_____30021, __9_____30022, __9_____30023,
       __9_____30024, __9_____30025, __9_____30026, __9_____30027;
  wire __9_____30028, __9_____30030, __9_____30031, __9_____30032,
       __9_____30033, __9_____30034, __9_____30035, __9_____30036;
  wire __9_____30037, __9_____30039, __9_____30040, __9_____30041,
       __9_____30042, __9_____30043, __9_____30044, __9_____30045;
  wire __9_____30046, __9_____30049, __9_____30050, __9_____30051,
       __9_____30052, __9_____30053, __9_____30054, __9_____30055;
  wire __9_____30057, __9_____30058, __9_____30059, __9_____30060,
       __9_____30061, __9_____30062, __9_____30065, __9_____30066;
  wire __9_____30067, __9_____30068, __9_____30069, __9_____30070,
       __9_____30071, __9_____30072, __9_____30094, __9_____30095;
  wire __9_____30096, __9_____30097, __9_____30098, __9_____30099,
       __9_____30100, __9_____30103, __9_____30104, __9_____30105;
  wire __9_____30106, __9_____30107, __9_____30108, __9_____30109,
       __9_____30112, __9_____30113, __9_____30114, __9_____30115;
  wire __9_____30116, __9_____30117, __9_____30118, __9_____30121,
       __9_____30122, __9_____30123, __9_____30124, __9_____30125;
  wire __9_____30126, __9_____30127, __9_____30128, __9_____30131,
       __9_____30132, __9_____30133, __9_____30134, __9_____30135;
  wire __9_____30136, __9_____30137, __9_____30138, __9_____30141,
       __9_____30142, __9_____30143, __9_____30144, __9_____30145;
  wire __9_____30146, __9_____30147, __9_____30148, __9_____30151,
       __9_____30152, __9_____30153, __9_____30154, __9_____30155;
  wire __9_____30156, __9_____30157, __9_____30160, __9_____30161,
       __9_____30162, __9_____30163, __9_____30164, __9_____30165;
  wire __9_____30166, __9_____30167, __9_____30187, __9_____30188,
       __9_____30189, __9_____30190, __9_____30191, __9_____30192;
  wire __9_____30193, __9_____30194, __9_____30197, __9_____30198,
       __9_____30199, __9_____30200, __9_____30201, __9_____30202;
  wire __9_____30203, __9_____30204, __9_____30207, __9_____30208,
       __9_____30209, __9_____30210, __9_____30211, __9_____30212;
  wire __9_____30213, __9_____30214, __9_____30217, __9_____30218,
       __9_____30219, __9_____30220, __9_____30221, __9_____30222;
  wire __9_____30223, __9_____30224, __9_____30227, __9_____30228,
       __9_____30229, __9_____30230, __9_____30231, __9_____30232;
  wire __9_____30235, __9_____30236, __9_____30237, __9_____30238,
       __9_____30239, __9_____30240, __9_____30241, __9_____30242;
  wire __9_____30245, __9_____30246, __9_____30247, __9_____30248,
       __9_____30249, __9_____30250, __9_____30251, __9_____30252;
  wire __9_____30255, __9_____30256, __9_____30257, __9_____30258,
       __9_____30259, __9_____30260, __9_____30261, __9_____30283;
  wire __9_____30284, __9_____30285, __9_____30286, __9_____30287,
       __9_____30288, __9_____30289, __9_____30292, __9_____30293;
  wire __9_____30294, __9_____30295, __9_____30296, __9_____30297,
       __9_____30298, __9_____30299, __9_____30301, __9_____30302;
  wire __9_____30303, __9_____30304, __9_____30305, __9_____30306,
       __9_____30307, __9_____30308, __9_____30311, __9_____30312;
  wire __9_____30313, __9_____30314, __9_____30315, __9_____30316,
       __9_____30317, __9_____30318, __9_____30321, __9_____30322;
  wire __9_____30323, __9_____30324, __9_____30325, __9_____30326,
       __9_____30327, __9_____30328, __9_____30331, __9_____30332;
  wire __9_____30333, __9_____30334, __9_____30335, __9_____30336,
       __9_____30339, __9_____30340, __9_____30341, __9_____30342;
  wire __9_____30343, __9_____30344, __9_____30345, __9_____30346,
       __9_____30348, __9_____30349, __9_____30350, __9_____30351;
  wire __9_____30352, __9_____30353, __9_____30354, __9_____30355,
       __9_____30376, __9_____30377, __9_____30378, __9_____30379;
  wire __9_____30380, __9_____30381, __9_____30382, __9_____30383,
       __9_____30385, __9_____30386, __9_____30387, __9_____30388;
  wire __9_____30389, __9_____30390, __9_____30391, __9_____30392,
       __9_____30395, __9_____30396, __9_____30397, __9_____30398;
  wire __9_____30399, __9_____30400, __9_____30401, __9_____30404,
       __9_____30405, __9_____30406, __9_____30407, __9_____30408;
  wire __9_____30409, __9_____30412, __9_____30413, __9_____30414,
       __9_____30415, __9_____30416, __9_____30417, __9_____30418;
  wire __9_____30421, __9_____30422, __9_____30423, __9_____30424,
       __9_____30425, __9_____30426, __9_____30427, __9_____30428;
  wire __9_____30430, __9_____30431, __9_____30432, __9_____30433,
       __9_____30434, __9_____30435, __9_____30436, __9_____30439;
  wire __9_____30440, __9_____30441, __9_____30442, __9_____30443,
       __90, __90_0, __90_0__29650, __90_0__29660;
  wire __90_0__29670, __90_0__29680, __90_0__29689, __90_0__29699,
       __90_0__29709, __90_9, __90_9__29659, __90_9__29669;
  wire __90_9__29679, __90_9__29688, __90_9__29698, __90_9__29708,
       __90_9__29717, __90__, __90____29645, __90____29646;
  wire __90____29647, __90____29648, __90____29649, __90____29651,
       __90____29652, __90____29653, __90____29654, __90____29655;
  wire __90____29656, __90____29657, __90____29658, __90____29661,
       __90____29662, __90____29663, __90____29664, __90____29665;
  wire __90____29666, __90____29667, __90____29668, __90____29671,
       __90____29672, __90____29673, __90____29674, __90____29675;
  wire __90____29676, __90____29677, __90____29678, __90____29681,
       __90____29682, __90____29683, __90____29684, __90____29685;
  wire __90____29686, __90____29687, __90____29690, __90____29691,
       __90____29692, __90____29693, __90____29694, __90____29695;
  wire __90____29696, __90____29697, __90____29700, __90____29701,
       __90____29702, __90____29703, __90____29704, __90____29705;
  wire __90____29706, __90____29707, __90____29710, __90____29711,
       __90____29712, __90____29713, __90____29714, __90____29715;
  wire __90____29716, __99_0, __99_0__30469, __99_0__30479,
       __99_0__30489, __99_0__30499, __99_0__30509, __99_0__30518;
  wire __99_0__30528, __99_9, __99_9__30478, __99_9__30488,
       __99_9__30498, __99_9__30508, __99_9__30517, __99_9__30527;
  wire __99_9__30537, __99__, __99____30462, __99____30463,
       __99____30464, __99____30465, __99____30466, __99____30467;
  wire __99____30468, __99____30470, __99____30471, __99____30472,
       __99____30473, __99____30474, __99____30475, __99____30476;
  wire __99____30477, __99____30480, __99____30481, __99____30482,
       __99____30483, __99____30484, __99____30485, __99____30486;
  wire __99____30487, __99____30490, __99____30491, __99____30492,
       __99____30493, __99____30494, __99____30495, __99____30496;
  wire __99____30497, __99____30500, __99____30501, __99____30502,
       __99____30503, __99____30504, __99____30505, __99____30506;
  wire __99____30507, __99____30510, __99____30511, __99____30512,
       __99____30513, __99____30514, __99____30515, __99____30516;
  wire __99____30519, __99____30520, __99____30521, __99____30522,
       __99____30523, __99____30524, __99____30525, __99____30526;
  wire __99____30529, __99____30530, __99____30531, __99____30532,
       __99____30533, __99____30534, __99____30535, __99____30536;
  wire __900_, __900___29638, __900___29639, __900___29640,
       __900___29641, __900___29642, __900___29643, __900___29644;
  wire __909_, __909___29718, __909___29719, __909___29720,
       __909___29721, __909___29722, __909___29723, __990_;
  wire __990___30455, __990___30456, __990___30457, __990___30458,
       __990___30459, __990___30460, __990___30461, __999_;
  wire __999___30538, __999___30539, __999___30540, __999___30541,
       __999___30542, __999___30543, __999___30544, __9090;
  wire __9099, __9900, __9909, __9990, __9999, ___, ___0, ___00;
  wire ___000, ___0000__30545, ___0000__39892, ___000__24168,
       ___000__25125, ___000__26051, ___000__28736, ___000___30546;
  wire ___000___30547, ___000___30548, ___000___30549, ___000___30550,
       ___000___30551, ___000___30552, ___000___30553, ___000___39893;
  wire ___000___39894, ___000___39895, ___000___39896, ___000___39897,
       ___000___39898, ___000___39899, ___000___39900, ___00_;
  wire ___00_0__30555, ___00_0__30565, ___00_0__30574, ___00_0__30584,
       ___00_0__30593, ___00_0__30603, ___00_0__30612, ___00_0__30622;
  wire ___00_0__39902, ___00_0__39912, ___00_0__39922, ___00_0__39930,
       ___00_0__39939, ___00_0__39949, ___00_0__39956, ___00_0__39964;
  wire ___00_9__30564, ___00_9__30573, ___00_9__30583, ___00_9__30592,
       ___00_9__30602, ___00_9__30611, ___00_9__30621, ___00_9__30631;
  wire ___00_9__39911, ___00_9__39921, ___00_9__39948, ___00_9__39955,
       ___00_9__39963, ___00_9__39972, ___00__22196, ___00__22272;
  wire ___00___22288, ___00___22289, ___00___23216, ___00___23217,
       ___00___23218, ___00___23219, ___00___23220, ___00___23221;
  wire ___00___23222, ___00___23223, ___00___24169, ___00___24170,
       ___00___24171, ___00___24172, ___00___24173, ___00___24174;
  wire ___00___24175, ___00___24176, ___00___25126, ___00___25127,
       ___00___25128, ___00___25129, ___00___25130, ___00___25131;
  wire ___00___25132, ___00___25133, ___00___26052, ___00___26053,
       ___00___26054, ___00___26055, ___00___26056, ___00___26057;
  wire ___00___26058, ___00___26954, ___00___26955, ___00___26956,
       ___00___26957, ___00___26958, ___00___27827, ___00___27828;
  wire ___00___27829, ___00___27830, ___00___27831, ___00___27832,
       ___00___27833, ___00___27834, ___00___28737, ___00___28738;
  wire ___00___28739, ___00___28740, ___00___28741, ___00___28742,
       ___00___28743, ___00___28744, ___00____30556, ___00____30557;
  wire ___00____30558, ___00____30559, ___00____30560, ___00____30561,
       ___00____30562, ___00____30563, ___00____30566, ___00____30567;
  wire ___00____30568, ___00____30569, ___00____30570, ___00____30571,
       ___00____30572, ___00____30575, ___00____30576, ___00____30577;
  wire ___00____30578, ___00____30579, ___00____30580, ___00____30581,
       ___00____30582, ___00____30585, ___00____30586, ___00____30587;
  wire ___00____30588, ___00____30589, ___00____30590, ___00____30591,
       ___00____30594, ___00____30595, ___00____30596, ___00____30597;
  wire ___00____30598, ___00____30599, ___00____30600, ___00____30601,
       ___00____30604, ___00____30605, ___00____30606, ___00____30607;
  wire ___00____30608, ___00____30609, ___00____30610, ___00____30613,
       ___00____30614, ___00____30615, ___00____30616, ___00____30617;
  wire ___00____30618, ___00____30619, ___00____30620, ___00____30623,
       ___00____30624, ___00____30625, ___00____30626, ___00____30627;
  wire ___00____30628, ___00____30629, ___00____30630, ___00____39903,
       ___00____39904, ___00____39905, ___00____39906, ___00____39907;
  wire ___00____39908, ___00____39909, ___00____39910, ___00____39913,
       ___00____39914, ___00____39915, ___00____39916, ___00____39917;
  wire ___00____39918, ___00____39919, ___00____39920, ___00____39923,
       ___00____39924, ___00____39925, ___00____39926, ___00____39927;
  wire ___00____39928, ___00____39929, ___00____39931, ___00____39932,
       ___00____39933, ___00____39934, ___00____39935, ___00____39936;
  wire ___00____39937, ___00____39938, ___00____39940, ___00____39941,
       ___00____39942, ___00____39943, ___00____39944, ___00____39945;
  wire ___00____39946, ___00____39947, ___00____39950, ___00____39951,
       ___00____39952, ___00____39953, ___00____39954, ___00____39957;
  wire ___00____39958, ___00____39959, ___00____39960, ___00____39961,
       ___00____39962, ___00____39965, ___00____39966, ___00____39967;
  wire ___00____39968, ___00____39969, ___00____39970, ___00____39971,
       ___00____41368, ___0_, ___0_0, ___0_00__30642;
  wire ___0_00__30740, ___0_00__30833, ___0_00__30927, ___0_00__31023,
       ___0_00__31118, ___0_00__31216, ___0_00__31310, ___0_00__39983;
  wire ___0_00__40079, ___0_00__40177, ___0_00__40273, ___0_00__40363,
       ___0_00__40461, ___0_00__40561, ___0_0__22297, ___0_0__22307;
  wire ___0_0__22324, ___0_0__22334, ___0_0__22344, ___0_0__23225,
       ___0_0__23235, ___0_0__23244, ___0_0__23253, ___0_0__23263;
  wire ___0_0__23273, ___0_0__23281, ___0_0__23291, ___0_0__24178,
       ___0_0__24188, ___0_0__24198, ___0_0__24208, ___0_0__24218;
  wire ___0_0__24228, ___0_0__24238, ___0_0__24248, ___0_0__25135,
       ___0_0__25145, ___0_0__25155, ___0_0__25165, ___0_0__25175;
  wire ___0_0__25185, ___0_0__25194, ___0_0__25203, ___0_0__26060,
       ___0_0__26069, ___0_0__26082, ___0_0__26092, ___0_0__26102;
  wire ___0_0__26112, ___0_0__26122, ___0_0__26960, ___0_0__26967,
       ___0_0__26999, ___0_0__27009, ___0_0__27018, ___0_0__27836;
  wire ___0_0__27845, ___0_0__27855, ___0_0__27865, ___0_0__27875,
       ___0_0__27884, ___0_0__27894, ___0_0__28746, ___0_0__28756;
  wire ___0_0__28766, ___0_0__28776, ___0_0__28786, ___0_0__28796,
       ___0_0__28805, ___0_0__28815, ___0_0___30643, ___0_0___30644;
  wire ___0_0___30645, ___0_0___30646, ___0_0___30647, ___0_0___30648,
       ___0_0___30649, ___0_0___30650, ___0_0___30741, ___0_0___30742;
  wire ___0_0___30743, ___0_0___30744, ___0_0___30745, ___0_0___30746,
       ___0_0___30747, ___0_0___30748, ___0_0___30834, ___0_0___30835;
  wire ___0_0___30836, ___0_0___30837, ___0_0___30838, ___0_0___30839,
       ___0_0___30840, ___0_0___30928, ___0_0___30929, ___0_0___30930;
  wire ___0_0___30931, ___0_0___30932, ___0_0___30933, ___0_0___31024,
       ___0_0___31025, ___0_0___31026, ___0_0___31027, ___0_0___31028;
  wire ___0_0___31029, ___0_0___31030, ___0_0___31031, ___0_0___31119,
       ___0_0___31120, ___0_0___31121, ___0_0___31122, ___0_0___31123;
  wire ___0_0___31124, ___0_0___31125, ___0_0___31126, ___0_0___31217,
       ___0_0___31218, ___0_0___31219, ___0_0___31220, ___0_0___31311;
  wire ___0_0___31312, ___0_0___31313, ___0_0___31314, ___0_0___31315,
       ___0_0___31316, ___0_0___31317, ___0_0___31318, ___0_0___39984;
  wire ___0_0___39985, ___0_0___39986, ___0_0___39987, ___0_0___39988,
       ___0_0___39989, ___0_0___39990, ___0_0___39991, ___0_0___40080;
  wire ___0_0___40081, ___0_0___40082, ___0_0___40083, ___0_0___40084,
       ___0_0___40085, ___0_0___40086, ___0_0___40087, ___0_0___40178;
  wire ___0_0___40179, ___0_0___40180, ___0_0___40181, ___0_0___40182,
       ___0_0___40183, ___0_0___40184, ___0_0___40185, ___0_0___40274;
  wire ___0_0___40275, ___0_0___40276, ___0_0___40277, ___0_0___40278,
       ___0_0___40279, ___0_0___40280, ___0_0___40281, ___0_0___40364;
  wire ___0_0___40365, ___0_0___40366, ___0_0___40367, ___0_0___40368,
       ___0_0___40369, ___0_0___40370, ___0_0___40371, ___0_0___40462;
  wire ___0_0___40463, ___0_0___40464, ___0_0___40465, ___0_0___40466,
       ___0_0___40467, ___0_0___40468, ___0_0___40469, ___0_0___40562;
  wire ___0_0___40563, ___0_0___40564, ___0_0___40565, ___0_0___40566,
       ___0_0___40567, ___0_0___40568, ___0_0___40569, ___0_09__30651;
  wire ___0_09__30749, ___0_09__30841, ___0_09__30934, ___0_09__31032,
       ___0_09__31127, ___0_09__31221, ___0_09__31319, ___0_09__39992;
  wire ___0_09__40088, ___0_09__40186, ___0_09__40282, ___0_09__40372,
       ___0_09__40470, ___0_09__40570, ___0_9, ___0_9__22306;
  wire ___0_9__22316, ___0_9__22323, ___0_9__22333, ___0_9__22343,
       ___0_9__22353, ___0_9__23234, ___0_9__23243, ___0_9__23262;
  wire ___0_9__23272, ___0_9__23290, ___0_9__23300, ___0_9__24187,
       ___0_9__24197, ___0_9__24207, ___0_9__24217, ___0_9__24227;
  wire ___0_9__24237, ___0_9__24247, ___0_9__24256, ___0_9__25144,
       ___0_9__25154, ___0_9__25164, ___0_9__25174, ___0_9__25184;
  wire ___0_9__25193, ___0_9__25202, ___0_9__25212, ___0_9__26081,
       ___0_9__26091, ___0_9__26101, ___0_9__26111, ___0_9__26121;
  wire ___0_9__26131, ___0_9__26966, ___0_9__26976, ___0_9__26991,
       ___0_9__26998, ___0_9__27008, ___0_9__27017, ___0_9__27844;
  wire ___0_9__27854, ___0_9__27864, ___0_9__27874, ___0_9__27883,
       ___0_9__27893, ___0_9__27902, ___0_9__27911, ___0_9__28755;
  wire ___0_9__28765, ___0_9__28775, ___0_9__28785, ___0_9__28795,
       ___0_9__28804, ___0_9__28814, ___0_9__28824, ___0_9___30731;
  wire ___0_9___30732, ___0_9___30733, ___0_9___30734, ___0_9___30735,
       ___0_9___30736, ___0_9___30737, ___0_9___30738, ___0_9___30824;
  wire ___0_9___30825, ___0_9___30826, ___0_9___30827, ___0_9___30828,
       ___0_9___30829, ___0_9___30830, ___0_9___30831, ___0_9___30920;
  wire ___0_9___30921, ___0_9___30922, ___0_9___30923, ___0_9___30924,
       ___0_9___30925, ___0_9___31014, ___0_9___31015, ___0_9___31016;
  wire ___0_9___31017, ___0_9___31018, ___0_9___31019, ___0_9___31020,
       ___0_9___31021, ___0_9___31109, ___0_9___31110, ___0_9___31111;
  wire ___0_9___31112, ___0_9___31113, ___0_9___31114, ___0_9___31115,
       ___0_9___31116, ___0_9___31207, ___0_9___31208, ___0_9___31209;
  wire ___0_9___31210, ___0_9___31211, ___0_9___31212, ___0_9___31213,
       ___0_9___31214, ___0_9___31301, ___0_9___31302, ___0_9___31303;
  wire ___0_9___31304, ___0_9___31305, ___0_9___31306, ___0_9___31307,
       ___0_9___31308, ___0_9___31399, ___0_9___31400, ___0_9___31401;
  wire ___0_9___31402, ___0_9___31403, ___0_9___31404, ___0_9___31405,
       ___0_9___31406, ___0_9___40070, ___0_9___40071, ___0_9___40072;
  wire ___0_9___40073, ___0_9___40074, ___0_9___40075, ___0_9___40076,
       ___0_9___40077, ___0_9___40169, ___0_9___40170, ___0_9___40171;
  wire ___0_9___40172, ___0_9___40173, ___0_9___40174, ___0_9___40175,
       ___0_9___40264, ___0_9___40265, ___0_9___40266, ___0_9___40267;
  wire ___0_9___40268, ___0_9___40269, ___0_9___40270, ___0_9___40271,
       ___0_9___40354, ___0_9___40355, ___0_9___40356, ___0_9___40357;
  wire ___0_9___40358, ___0_9___40359, ___0_9___40360, ___0_9___40361,
       ___0_9___40452, ___0_9___40453, ___0_9___40454, ___0_9___40455;
  wire ___0_9___40456, ___0_9___40457, ___0_9___40458, ___0_9___40459,
       ___0_9___40552, ___0_9___40553, ___0_9___40554, ___0_9___40555;
  wire ___0_9___40556, ___0_9___40557, ___0_9___40558, ___0_9___40559,
       ___0_9___40645, ___0_9___40653, ___0_9___40654, ___0_90__30730;
  wire ___0_90__30823, ___0_90__30919, ___0_90__31013, ___0_90__31108,
       ___0_90__31206, ___0_90__31300, ___0_90__31398, ___0_90__40069;
  wire ___0_90__40168, ___0_90__40263, ___0_90__40353, ___0_90__40451,
       ___0_90__40551, ___0_99__30739, ___0_99__30832, ___0_99__30926;
  wire ___0_99__31022, ___0_99__31117, ___0_99__31215, ___0_99__31309,
       ___0_99__31407, ___0_99__40078, ___0_99__40176, ___0_99__40272;
  wire ___0_99__40362, ___0_99__40460, ___0_99__40560, ___0__,
       ___0__0__30652, ___0__0__30662, ___0__0__30672, ___0__0__30682;
  wire ___0__0__30692, ___0__0__30701, ___0__0__30711, ___0__0__30721,
       ___0__0__30750, ___0__0__30759, ___0__0__30769, ___0__0__30778;
  wire ___0__0__30787, ___0__0__30796, ___0__0__30804, ___0__0__30814,
       ___0__0__30842, ___0__0__30852, ___0__0__30862, ___0__0__30872;
  wire ___0__0__30881, ___0__0__30891, ___0__0__30899, ___0__0__30909,
       ___0__0__30935, ___0__0__30945, ___0__0__30955, ___0__0__30965;
  wire ___0__0__30975, ___0__0__30985, ___0__0__30994, ___0__0__31003,
       ___0__0__31033, ___0__0__31042, ___0__0__31051, ___0__0__31061;
  wire ___0__0__31071, ___0__0__31080, ___0__0__31090, ___0__0__31099,
       ___0__0__31128, ___0__0__31138, ___0__0__31148, ___0__0__31158;
  wire ___0__0__31168, ___0__0__31178, ___0__0__31188, ___0__0__31197,
       ___0__0__31222, ___0__0__31232, ___0__0__31241, ___0__0__31251;
  wire ___0__0__31261, ___0__0__31271, ___0__0__31281, ___0__0__31290,
       ___0__0__31320, ___0__0__31330, ___0__0__31339, ___0__0__31348;
  wire ___0__0__31358, ___0__0__31368, ___0__0__31378, ___0__0__31388,
       ___0__0__39993, ___0__0__40002, ___0__0__40012, ___0__0__40021;
  wire ___0__0__40039, ___0__0__40049, ___0__0__40059, ___0__0__40089,
       ___0__0__40099, ___0__0__40109, ___0__0__40119, ___0__0__40129;
  wire ___0__0__40139, ___0__0__40149, ___0__0__40159, ___0__0__40187,
       ___0__0__40197, ___0__0__40206, ___0__0__40215, ___0__0__40233;
  wire ___0__0__40243, ___0__0__40253, ___0__0__40283, ___0__0__40291,
       ___0__0__40301, ___0__0__40309, ___0__0__40318, ___0__0__40325;
  wire ___0__0__40333, ___0__0__40343, ___0__0__40373, ___0__0__40383,
       ___0__0__40393, ___0__0__40403, ___0__0__40413, ___0__0__40421;
  wire ___0__0__40431, ___0__0__40441, ___0__0__40471, ___0__0__40481,
       ___0__0__40491, ___0__0__40501, ___0__0__40511, ___0__0__40521;
  wire ___0__0__40531, ___0__0__40541, ___0__0__40571, ___0__0__40581,
       ___0__0__40591, ___0__0__40599, ___0__0__40609, ___0__0__40619;
  wire ___0__0__40629, ___0__0__40639, ___0__0__40648, ___0__9__30661,
       ___0__9__30671, ___0__9__30681, ___0__9__30691, ___0__9__30710;
  wire ___0__9__30720, ___0__9__30729, ___0__9__30758, ___0__9__30768,
       ___0__9__30777, ___0__9__30786, ___0__9__30795, ___0__9__30813;
  wire ___0__9__30822, ___0__9__30851, ___0__9__30861, ___0__9__30871,
       ___0__9__30880, ___0__9__30890, ___0__9__30898, ___0__9__30908;
  wire ___0__9__30918, ___0__9__30944, ___0__9__30954, ___0__9__30964,
       ___0__9__30974, ___0__9__30984, ___0__9__30993, ___0__9__31012;
  wire ___0__9__31041, ___0__9__31050, ___0__9__31060, ___0__9__31070,
       ___0__9__31089, ___0__9__31098, ___0__9__31107, ___0__9__31137;
  wire ___0__9__31147, ___0__9__31157, ___0__9__31167, ___0__9__31177,
       ___0__9__31187, ___0__9__31196, ___0__9__31205, ___0__9__31231;
  wire ___0__9__31240, ___0__9__31250, ___0__9__31260, ___0__9__31270,
       ___0__9__31280, ___0__9__31289, ___0__9__31299, ___0__9__31329;
  wire ___0__9__31347, ___0__9__31357, ___0__9__31367, ___0__9__31377,
       ___0__9__31387, ___0__9__31397, ___0__9__40001, ___0__9__40011;
  wire ___0__9__40020, ___0__9__40029, ___0__9__40038, ___0__9__40048,
       ___0__9__40058, ___0__9__40068, ___0__9__40098, ___0__9__40108;
  wire ___0__9__40118, ___0__9__40128, ___0__9__40138, ___0__9__40148,
       ___0__9__40158, ___0__9__40167, ___0__9__40196, ___0__9__40214;
  wire ___0__9__40223, ___0__9__40232, ___0__9__40242, ___0__9__40252,
       ___0__9__40262, ___0__9__40290, ___0__9__40300, ___0__9__40317;
  wire ___0__9__40332, ___0__9__40342, ___0__9__40352, ___0__9__40382,
       ___0__9__40392, ___0__9__40402, ___0__9__40412, ___0__9__40420;
  wire ___0__9__40430, ___0__9__40440, ___0__9__40450, ___0__9__40480,
       ___0__9__40490, ___0__9__40500, ___0__9__40510, ___0__9__40520;
  wire ___0__9__40530, ___0__9__40540, ___0__9__40550, ___0__9__40580,
       ___0__9__40590, ___0__9__40608, ___0__9__40618, ___0__9__40628;
  wire ___0__9__40638, ___0__22134, ___0__22149, ___0__22157,
       ___0___22170, ___0___22171, ___0___22197, ___0___22198;
  wire ___0___22199, ___0___22200, ___0___22201, ___0___22202,
       ___0___22203, ___0___22204, ___0___22273, ___0___22274;
  wire ___0___22275, ___0___22276, ___0____22290, ___0____22291,
       ___0____22292, ___0____22293, ___0____22294, ___0____22295;
  wire ___0____22296, ___0____22298, ___0____22299, ___0____22300,
       ___0____22301, ___0____22302, ___0____22303, ___0____22304;
  wire ___0____22305, ___0____22308, ___0____22309, ___0____22310,
       ___0____22311, ___0____22312, ___0____22313, ___0____22314;
  wire ___0____22315, ___0____22317, ___0____22318, ___0____22319,
       ___0____22320, ___0____22321, ___0____22322, ___0____22325;
  wire ___0____22326, ___0____22327, ___0____22328, ___0____22329,
       ___0____22330, ___0____22331, ___0____22332, ___0____22335;
  wire ___0____22336, ___0____22337, ___0____22338, ___0____22339,
       ___0____22340, ___0____22341, ___0____22342, ___0____22345;
  wire ___0____22346, ___0____22347, ___0____22348, ___0____22349,
       ___0____22350, ___0____22351, ___0____22352, ___0____23226;
  wire ___0____23227, ___0____23228, ___0____23229, ___0____23230,
       ___0____23231, ___0____23232, ___0____23233, ___0____23236;
  wire ___0____23237, ___0____23238, ___0____23239, ___0____23240,
       ___0____23241, ___0____23242, ___0____23245, ___0____23246;
  wire ___0____23247, ___0____23248, ___0____23249, ___0____23250,
       ___0____23251, ___0____23252, ___0____23254, ___0____23255;
  wire ___0____23256, ___0____23257, ___0____23258, ___0____23259,
       ___0____23260, ___0____23261, ___0____23264, ___0____23265;
  wire ___0____23266, ___0____23267, ___0____23268, ___0____23269,
       ___0____23270, ___0____23271, ___0____23274, ___0____23275;
  wire ___0____23276, ___0____23277, ___0____23278, ___0____23279,
       ___0____23280, ___0____23282, ___0____23283, ___0____23284;
  wire ___0____23285, ___0____23286, ___0____23287, ___0____23288,
       ___0____23289, ___0____23292, ___0____23293, ___0____23294;
  wire ___0____23295, ___0____23296, ___0____23297, ___0____23298,
       ___0____23299, ___0____24179, ___0____24180, ___0____24181;
  wire ___0____24182, ___0____24183, ___0____24184, ___0____24185,
       ___0____24186, ___0____24189, ___0____24190, ___0____24191;
  wire ___0____24192, ___0____24193, ___0____24194, ___0____24195,
       ___0____24196, ___0____24199, ___0____24200, ___0____24201;
  wire ___0____24202, ___0____24203, ___0____24204, ___0____24205,
       ___0____24206, ___0____24209, ___0____24210, ___0____24211;
  wire ___0____24212, ___0____24213, ___0____24214, ___0____24215,
       ___0____24216, ___0____24219, ___0____24220, ___0____24221;
  wire ___0____24222, ___0____24223, ___0____24224, ___0____24225,
       ___0____24226, ___0____24229, ___0____24230, ___0____24231;
  wire ___0____24232, ___0____24233, ___0____24234, ___0____24235,
       ___0____24236, ___0____24239, ___0____24240, ___0____24241;
  wire ___0____24242, ___0____24243, ___0____24244, ___0____24245,
       ___0____24246, ___0____24249, ___0____24250, ___0____24251;
  wire ___0____24252, ___0____24253, ___0____24254, ___0____24255,
       ___0____25136, ___0____25137, ___0____25138, ___0____25139;
  wire ___0____25140, ___0____25141, ___0____25142, ___0____25143,
       ___0____25146, ___0____25147, ___0____25148, ___0____25149;
  wire ___0____25150, ___0____25151, ___0____25152, ___0____25153,
       ___0____25156, ___0____25157, ___0____25158, ___0____25159;
  wire ___0____25160, ___0____25161, ___0____25162, ___0____25163,
       ___0____25166, ___0____25167, ___0____25168, ___0____25169;
  wire ___0____25170, ___0____25171, ___0____25172, ___0____25173,
       ___0____25176, ___0____25177, ___0____25178, ___0____25179;
  wire ___0____25180, ___0____25181, ___0____25182, ___0____25183,
       ___0____25186, ___0____25187, ___0____25188, ___0____25189;
  wire ___0____25190, ___0____25191, ___0____25192, ___0____25195,
       ___0____25196, ___0____25197, ___0____25198, ___0____25199;
  wire ___0____25200, ___0____25201, ___0____25204, ___0____25205,
       ___0____25206, ___0____25207, ___0____25208, ___0____25209;
  wire ___0____25210, ___0____25211, ___0____26061, ___0____26062,
       ___0____26063, ___0____26064, ___0____26065, ___0____26066;
  wire ___0____26067, ___0____26068, ___0____26070, ___0____26071,
       ___0____26072, ___0____26073, ___0____26074, ___0____26075;
  wire ___0____26076, ___0____26077, ___0____26078, ___0____26079,
       ___0____26080, ___0____26083, ___0____26084, ___0____26085;
  wire ___0____26086, ___0____26087, ___0____26088, ___0____26089,
       ___0____26090, ___0____26093, ___0____26094, ___0____26095;
  wire ___0____26096, ___0____26097, ___0____26098, ___0____26099,
       ___0____26100, ___0____26103, ___0____26104, ___0____26105;
  wire ___0____26106, ___0____26107, ___0____26108, ___0____26109,
       ___0____26110, ___0____26113, ___0____26114, ___0____26115;
  wire ___0____26116, ___0____26117, ___0____26118, ___0____26119,
       ___0____26120, ___0____26123, ___0____26124, ___0____26125;
  wire ___0____26126, ___0____26127, ___0____26128, ___0____26129,
       ___0____26130, ___0____26961, ___0____26962, ___0____26963;
  wire ___0____26964, ___0____26965, ___0____26968, ___0____26969,
       ___0____26970, ___0____26971, ___0____26972, ___0____26973;
  wire ___0____26974, ___0____26975, ___0____26977, ___0____26978,
       ___0____26979, ___0____26980, ___0____26981, ___0____26982;
  wire ___0____26983, ___0____26984, ___0____26985, ___0____26986,
       ___0____26987, ___0____26988, ___0____26989, ___0____26990;
  wire ___0____26992, ___0____26993, ___0____26994, ___0____26995,
       ___0____26996, ___0____26997, ___0____27000, ___0____27001;
  wire ___0____27002, ___0____27003, ___0____27004, ___0____27005,
       ___0____27006, ___0____27007, ___0____27010, ___0____27011;
  wire ___0____27012, ___0____27013, ___0____27014, ___0____27015,
       ___0____27016, ___0____27019, ___0____27020, ___0____27021;
  wire ___0____27022, ___0____27023, ___0____27024, ___0____27025,
       ___0____27837, ___0____27838, ___0____27839, ___0____27840;
  wire ___0____27841, ___0____27842, ___0____27843, ___0____27846,
       ___0____27847, ___0____27848, ___0____27849, ___0____27850;
  wire ___0____27851, ___0____27852, ___0____27853, ___0____27856,
       ___0____27857, ___0____27858, ___0____27859, ___0____27860;
  wire ___0____27861, ___0____27862, ___0____27863, ___0____27866,
       ___0____27867, ___0____27868, ___0____27869, ___0____27870;
  wire ___0____27871, ___0____27872, ___0____27873, ___0____27876,
       ___0____27877, ___0____27878, ___0____27879, ___0____27880;
  wire ___0____27881, ___0____27882, ___0____27885, ___0____27886,
       ___0____27887, ___0____27888, ___0____27889, ___0____27890;
  wire ___0____27891, ___0____27892, ___0____27895, ___0____27896,
       ___0____27897, ___0____27898, ___0____27899, ___0____27900;
  wire ___0____27901, ___0____27903, ___0____27904, ___0____27905,
       ___0____27906, ___0____27907, ___0____27908, ___0____27909;
  wire ___0____27910, ___0____28747, ___0____28748, ___0____28749,
       ___0____28750, ___0____28751, ___0____28752, ___0____28753;
  wire ___0____28754, ___0____28757, ___0____28758, ___0____28759,
       ___0____28760, ___0____28761, ___0____28762, ___0____28763;
  wire ___0____28764, ___0____28767, ___0____28768, ___0____28769,
       ___0____28770, ___0____28771, ___0____28772, ___0____28773;
  wire ___0____28774, ___0____28777, ___0____28778, ___0____28779,
       ___0____28780, ___0____28781, ___0____28782, ___0____28783;
  wire ___0____28784, ___0____28787, ___0____28788, ___0____28789,
       ___0____28790, ___0____28791, ___0____28792, ___0____28793;
  wire ___0____28794, ___0____28797, ___0____28798, ___0____28799,
       ___0____28800, ___0____28801, ___0____28802, ___0____28803;
  wire ___0____28806, ___0____28807, ___0____28808, ___0____28809,
       ___0____28810, ___0____28811, ___0____28812, ___0____28813;
  wire ___0____28816, ___0____28817, ___0____28818, ___0____28819,
       ___0____28820, ___0____28821, ___0____28822, ___0____28823;
  wire ___0_____30653, ___0_____30654, ___0_____30655, ___0_____30656,
       ___0_____30657, ___0_____30658, ___0_____30659, ___0_____30660;
  wire ___0_____30663, ___0_____30664, ___0_____30665, ___0_____30666,
       ___0_____30667, ___0_____30668, ___0_____30669, ___0_____30670;
  wire ___0_____30673, ___0_____30674, ___0_____30675, ___0_____30676,
       ___0_____30677, ___0_____30678, ___0_____30679, ___0_____30680;
  wire ___0_____30683, ___0_____30684, ___0_____30685, ___0_____30686,
       ___0_____30687, ___0_____30688, ___0_____30689, ___0_____30690;
  wire ___0_____30693, ___0_____30694, ___0_____30695, ___0_____30696,
       ___0_____30697, ___0_____30698, ___0_____30699, ___0_____30700;
  wire ___0_____30702, ___0_____30703, ___0_____30704, ___0_____30705,
       ___0_____30706, ___0_____30707, ___0_____30708, ___0_____30709;
  wire ___0_____30712, ___0_____30713, ___0_____30714, ___0_____30715,
       ___0_____30716, ___0_____30717, ___0_____30718, ___0_____30719;
  wire ___0_____30722, ___0_____30723, ___0_____30724, ___0_____30725,
       ___0_____30726, ___0_____30727, ___0_____30728, ___0_____30751;
  wire ___0_____30752, ___0_____30753, ___0_____30754, ___0_____30755,
       ___0_____30756, ___0_____30757, ___0_____30760, ___0_____30761;
  wire ___0_____30762, ___0_____30763, ___0_____30764, ___0_____30765,
       ___0_____30766, ___0_____30767, ___0_____30770, ___0_____30771;
  wire ___0_____30772, ___0_____30773, ___0_____30774, ___0_____30775,
       ___0_____30776, ___0_____30779, ___0_____30780, ___0_____30781;
  wire ___0_____30782, ___0_____30783, ___0_____30784, ___0_____30785,
       ___0_____30788, ___0_____30789, ___0_____30790, ___0_____30791;
  wire ___0_____30792, ___0_____30793, ___0_____30794, ___0_____30797,
       ___0_____30798, ___0_____30799, ___0_____30800, ___0_____30801;
  wire ___0_____30802, ___0_____30803, ___0_____30805, ___0_____30806,
       ___0_____30807, ___0_____30808, ___0_____30809, ___0_____30810;
  wire ___0_____30811, ___0_____30812, ___0_____30815, ___0_____30816,
       ___0_____30817, ___0_____30818, ___0_____30819, ___0_____30820;
  wire ___0_____30821, ___0_____30843, ___0_____30844, ___0_____30845,
       ___0_____30846, ___0_____30847, ___0_____30848, ___0_____30849;
  wire ___0_____30850, ___0_____30853, ___0_____30854, ___0_____30855,
       ___0_____30856, ___0_____30857, ___0_____30858, ___0_____30859;
  wire ___0_____30860, ___0_____30863, ___0_____30864, ___0_____30865,
       ___0_____30866, ___0_____30867, ___0_____30868, ___0_____30869;
  wire ___0_____30870, ___0_____30873, ___0_____30874, ___0_____30875,
       ___0_____30876, ___0_____30877, ___0_____30878, ___0_____30879;
  wire ___0_____30882, ___0_____30883, ___0_____30884, ___0_____30885,
       ___0_____30886, ___0_____30887, ___0_____30888, ___0_____30889;
  wire ___0_____30892, ___0_____30893, ___0_____30894, ___0_____30895,
       ___0_____30896, ___0_____30897, ___0_____30900, ___0_____30901;
  wire ___0_____30902, ___0_____30903, ___0_____30904, ___0_____30905,
       ___0_____30906, ___0_____30907, ___0_____30910, ___0_____30911;
  wire ___0_____30912, ___0_____30913, ___0_____30914, ___0_____30915,
       ___0_____30916, ___0_____30917, ___0_____30936, ___0_____30937;
  wire ___0_____30938, ___0_____30939, ___0_____30940, ___0_____30941,
       ___0_____30942, ___0_____30943, ___0_____30946, ___0_____30947;
  wire ___0_____30948, ___0_____30949, ___0_____30950, ___0_____30951,
       ___0_____30952, ___0_____30953, ___0_____30956, ___0_____30957;
  wire ___0_____30958, ___0_____30959, ___0_____30960, ___0_____30961,
       ___0_____30962, ___0_____30963, ___0_____30966, ___0_____30967;
  wire ___0_____30968, ___0_____30969, ___0_____30970, ___0_____30971,
       ___0_____30972, ___0_____30973, ___0_____30976, ___0_____30977;
  wire ___0_____30978, ___0_____30979, ___0_____30980, ___0_____30981,
       ___0_____30982, ___0_____30983, ___0_____30986, ___0_____30987;
  wire ___0_____30988, ___0_____30989, ___0_____30990, ___0_____30991,
       ___0_____30992, ___0_____30995, ___0_____30996, ___0_____30997;
  wire ___0_____30998, ___0_____30999, ___0_____31000, ___0_____31001,
       ___0_____31002, ___0_____31004, ___0_____31005, ___0_____31006;
  wire ___0_____31007, ___0_____31008, ___0_____31009, ___0_____31010,
       ___0_____31011, ___0_____31034, ___0_____31035, ___0_____31036;
  wire ___0_____31037, ___0_____31038, ___0_____31039, ___0_____31040,
       ___0_____31043, ___0_____31044, ___0_____31045, ___0_____31046;
  wire ___0_____31047, ___0_____31048, ___0_____31049, ___0_____31052,
       ___0_____31053, ___0_____31054, ___0_____31055, ___0_____31056;
  wire ___0_____31057, ___0_____31058, ___0_____31059, ___0_____31062,
       ___0_____31063, ___0_____31064, ___0_____31065, ___0_____31066;
  wire ___0_____31067, ___0_____31068, ___0_____31069, ___0_____31072,
       ___0_____31073, ___0_____31074, ___0_____31075, ___0_____31076;
  wire ___0_____31077, ___0_____31078, ___0_____31079, ___0_____31081,
       ___0_____31082, ___0_____31083, ___0_____31084, ___0_____31085;
  wire ___0_____31086, ___0_____31087, ___0_____31088, ___0_____31091,
       ___0_____31092, ___0_____31093, ___0_____31094, ___0_____31095;
  wire ___0_____31096, ___0_____31097, ___0_____31100, ___0_____31101,
       ___0_____31102, ___0_____31103, ___0_____31104, ___0_____31105;
  wire ___0_____31106, ___0_____31129, ___0_____31130, ___0_____31131,
       ___0_____31132, ___0_____31133, ___0_____31134, ___0_____31135;
  wire ___0_____31136, ___0_____31139, ___0_____31140, ___0_____31141,
       ___0_____31142, ___0_____31143, ___0_____31144, ___0_____31145;
  wire ___0_____31146, ___0_____31149, ___0_____31150, ___0_____31151,
       ___0_____31152, ___0_____31153, ___0_____31154, ___0_____31155;
  wire ___0_____31156, ___0_____31159, ___0_____31160, ___0_____31161,
       ___0_____31162, ___0_____31163, ___0_____31164, ___0_____31165;
  wire ___0_____31166, ___0_____31169, ___0_____31170, ___0_____31171,
       ___0_____31172, ___0_____31173, ___0_____31174, ___0_____31175;
  wire ___0_____31176, ___0_____31179, ___0_____31180, ___0_____31181,
       ___0_____31182, ___0_____31183, ___0_____31184, ___0_____31185;
  wire ___0_____31186, ___0_____31189, ___0_____31190, ___0_____31191,
       ___0_____31192, ___0_____31193, ___0_____31194, ___0_____31195;
  wire ___0_____31198, ___0_____31199, ___0_____31200, ___0_____31201,
       ___0_____31202, ___0_____31203, ___0_____31204, ___0_____31223;
  wire ___0_____31224, ___0_____31225, ___0_____31226, ___0_____31227,
       ___0_____31228, ___0_____31229, ___0_____31230, ___0_____31233;
  wire ___0_____31234, ___0_____31235, ___0_____31236, ___0_____31237,
       ___0_____31238, ___0_____31239, ___0_____31242, ___0_____31243;
  wire ___0_____31244, ___0_____31245, ___0_____31246, ___0_____31247,
       ___0_____31248, ___0_____31249, ___0_____31252, ___0_____31253;
  wire ___0_____31254, ___0_____31255, ___0_____31256, ___0_____31257,
       ___0_____31258, ___0_____31259, ___0_____31262, ___0_____31263;
  wire ___0_____31264, ___0_____31265, ___0_____31266, ___0_____31267,
       ___0_____31268, ___0_____31269, ___0_____31272, ___0_____31273;
  wire ___0_____31274, ___0_____31275, ___0_____31276, ___0_____31277,
       ___0_____31278, ___0_____31279, ___0_____31282, ___0_____31283;
  wire ___0_____31284, ___0_____31285, ___0_____31286, ___0_____31287,
       ___0_____31288, ___0_____31291, ___0_____31292, ___0_____31293;
  wire ___0_____31294, ___0_____31295, ___0_____31296, ___0_____31297,
       ___0_____31298, ___0_____31321, ___0_____31322, ___0_____31323;
  wire ___0_____31324, ___0_____31325, ___0_____31326, ___0_____31327,
       ___0_____31328, ___0_____31331, ___0_____31332, ___0_____31333;
  wire ___0_____31334, ___0_____31335, ___0_____31336, ___0_____31337,
       ___0_____31338, ___0_____31340, ___0_____31341, ___0_____31342;
  wire ___0_____31343, ___0_____31344, ___0_____31345, ___0_____31346,
       ___0_____31349, ___0_____31350, ___0_____31351, ___0_____31352;
  wire ___0_____31353, ___0_____31354, ___0_____31355, ___0_____31356,
       ___0_____31359, ___0_____31360, ___0_____31361, ___0_____31362;
  wire ___0_____31363, ___0_____31364, ___0_____31365, ___0_____31366,
       ___0_____31369, ___0_____31370, ___0_____31371, ___0_____31372;
  wire ___0_____31373, ___0_____31374, ___0_____31375, ___0_____31376,
       ___0_____31379, ___0_____31380, ___0_____31381, ___0_____31382;
  wire ___0_____31383, ___0_____31384, ___0_____31385, ___0_____31386,
       ___0_____31389, ___0_____31390, ___0_____31391, ___0_____31392;
  wire ___0_____31393, ___0_____31394, ___0_____31395, ___0_____31396,
       ___0_____39994, ___0_____39995, ___0_____39996, ___0_____39997;
  wire ___0_____39998, ___0_____39999, ___0_____40000, ___0_____40003,
       ___0_____40004, ___0_____40005, ___0_____40006, ___0_____40007;
  wire ___0_____40008, ___0_____40009, ___0_____40010, ___0_____40013,
       ___0_____40014, ___0_____40015, ___0_____40016, ___0_____40017;
  wire ___0_____40018, ___0_____40019, ___0_____40022, ___0_____40023,
       ___0_____40024, ___0_____40025, ___0_____40026, ___0_____40027;
  wire ___0_____40028, ___0_____40030, ___0_____40031, ___0_____40032,
       ___0_____40033, ___0_____40034, ___0_____40035, ___0_____40036;
  wire ___0_____40037, ___0_____40040, ___0_____40041, ___0_____40042,
       ___0_____40043, ___0_____40044, ___0_____40045, ___0_____40046;
  wire ___0_____40047, ___0_____40050, ___0_____40051, ___0_____40052,
       ___0_____40053, ___0_____40054, ___0_____40055, ___0_____40056;
  wire ___0_____40057, ___0_____40060, ___0_____40061, ___0_____40062,
       ___0_____40063, ___0_____40064, ___0_____40065, ___0_____40066;
  wire ___0_____40067, ___0_____40090, ___0_____40091, ___0_____40092,
       ___0_____40093, ___0_____40094, ___0_____40095, ___0_____40096;
  wire ___0_____40097, ___0_____40100, ___0_____40101, ___0_____40102,
       ___0_____40103, ___0_____40104, ___0_____40105, ___0_____40106;
  wire ___0_____40107, ___0_____40110, ___0_____40111, ___0_____40112,
       ___0_____40113, ___0_____40114, ___0_____40115, ___0_____40116;
  wire ___0_____40117, ___0_____40120, ___0_____40121, ___0_____40122,
       ___0_____40123, ___0_____40124, ___0_____40125, ___0_____40126;
  wire ___0_____40127, ___0_____40130, ___0_____40131, ___0_____40132,
       ___0_____40133, ___0_____40134, ___0_____40135, ___0_____40136;
  wire ___0_____40137, ___0_____40140, ___0_____40141, ___0_____40142,
       ___0_____40143, ___0_____40144, ___0_____40145, ___0_____40146;
  wire ___0_____40147, ___0_____40150, ___0_____40151, ___0_____40152,
       ___0_____40153, ___0_____40154, ___0_____40155, ___0_____40156;
  wire ___0_____40157, ___0_____40160, ___0_____40161, ___0_____40162,
       ___0_____40163, ___0_____40164, ___0_____40165, ___0_____40166;
  wire ___0_____40188, ___0_____40189, ___0_____40190, ___0_____40191,
       ___0_____40192, ___0_____40193, ___0_____40194, ___0_____40195;
  wire ___0_____40198, ___0_____40199, ___0_____40200, ___0_____40201,
       ___0_____40202, ___0_____40203, ___0_____40204, ___0_____40205;
  wire ___0_____40207, ___0_____40208, ___0_____40209, ___0_____40210,
       ___0_____40211, ___0_____40212, ___0_____40213, ___0_____40216;
  wire ___0_____40217, ___0_____40218, ___0_____40219, ___0_____40220,
       ___0_____40221, ___0_____40222, ___0_____40224, ___0_____40225;
  wire ___0_____40226, ___0_____40227, ___0_____40228, ___0_____40229,
       ___0_____40230, ___0_____40231, ___0_____40234, ___0_____40235;
  wire ___0_____40236, ___0_____40237, ___0_____40238, ___0_____40239,
       ___0_____40240, ___0_____40241, ___0_____40244, ___0_____40245;
  wire ___0_____40246, ___0_____40247, ___0_____40248, ___0_____40249,
       ___0_____40250, ___0_____40251, ___0_____40254, ___0_____40255;
  wire ___0_____40256, ___0_____40257, ___0_____40258, ___0_____40259,
       ___0_____40260, ___0_____40261, ___0_____40284, ___0_____40285;
  wire ___0_____40286, ___0_____40287, ___0_____40288, ___0_____40289,
       ___0_____40292, ___0_____40293, ___0_____40294, ___0_____40295;
  wire ___0_____40296, ___0_____40297, ___0_____40298, ___0_____40299,
       ___0_____40302, ___0_____40303, ___0_____40304, ___0_____40305;
  wire ___0_____40306, ___0_____40307, ___0_____40308, ___0_____40310,
       ___0_____40311, ___0_____40312, ___0_____40313, ___0_____40314;
  wire ___0_____40315, ___0_____40316, ___0_____40319, ___0_____40320,
       ___0_____40321, ___0_____40322, ___0_____40323, ___0_____40324;
  wire ___0_____40326, ___0_____40327, ___0_____40328, ___0_____40329,
       ___0_____40330, ___0_____40331, ___0_____40334, ___0_____40335;
  wire ___0_____40336, ___0_____40337, ___0_____40338, ___0_____40339,
       ___0_____40340, ___0_____40341, ___0_____40344, ___0_____40345;
  wire ___0_____40346, ___0_____40347, ___0_____40348, ___0_____40349,
       ___0_____40350, ___0_____40351, ___0_____40374, ___0_____40375;
  wire ___0_____40376, ___0_____40377, ___0_____40378, ___0_____40379,
       ___0_____40380, ___0_____40381, ___0_____40384, ___0_____40385;
  wire ___0_____40386, ___0_____40387, ___0_____40388, ___0_____40389,
       ___0_____40390, ___0_____40391, ___0_____40394, ___0_____40395;
  wire ___0_____40396, ___0_____40397, ___0_____40398, ___0_____40399,
       ___0_____40400, ___0_____40401, ___0_____40404, ___0_____40405;
  wire ___0_____40406, ___0_____40407, ___0_____40408, ___0_____40409,
       ___0_____40410, ___0_____40411, ___0_____40414, ___0_____40415;
  wire ___0_____40416, ___0_____40417, ___0_____40418, ___0_____40419,
       ___0_____40422, ___0_____40423, ___0_____40424, ___0_____40425;
  wire ___0_____40426, ___0_____40427, ___0_____40428, ___0_____40429,
       ___0_____40432, ___0_____40433, ___0_____40434, ___0_____40435;
  wire ___0_____40436, ___0_____40437, ___0_____40438, ___0_____40439,
       ___0_____40442, ___0_____40443, ___0_____40444, ___0_____40445;
  wire ___0_____40446, ___0_____40447, ___0_____40448, ___0_____40449,
       ___0_____40472, ___0_____40473, ___0_____40474, ___0_____40475;
  wire ___0_____40476, ___0_____40477, ___0_____40478, ___0_____40479,
       ___0_____40482, ___0_____40483, ___0_____40484, ___0_____40485;
  wire ___0_____40486, ___0_____40487, ___0_____40488, ___0_____40489,
       ___0_____40492, ___0_____40493, ___0_____40494, ___0_____40495;
  wire ___0_____40496, ___0_____40497, ___0_____40498, ___0_____40499,
       ___0_____40502, ___0_____40503, ___0_____40504, ___0_____40505;
  wire ___0_____40506, ___0_____40507, ___0_____40508, ___0_____40509,
       ___0_____40512, ___0_____40513, ___0_____40514, ___0_____40515;
  wire ___0_____40516, ___0_____40517, ___0_____40518, ___0_____40519,
       ___0_____40522, ___0_____40523, ___0_____40524, ___0_____40525;
  wire ___0_____40526, ___0_____40527, ___0_____40528, ___0_____40529,
       ___0_____40532, ___0_____40533, ___0_____40534, ___0_____40535;
  wire ___0_____40536, ___0_____40537, ___0_____40538, ___0_____40539,
       ___0_____40542, ___0_____40543, ___0_____40544, ___0_____40545;
  wire ___0_____40546, ___0_____40547, ___0_____40548, ___0_____40549,
       ___0_____40572, ___0_____40573, ___0_____40574, ___0_____40575;
  wire ___0_____40576, ___0_____40577, ___0_____40578, ___0_____40579,
       ___0_____40582, ___0_____40583, ___0_____40584, ___0_____40585;
  wire ___0_____40586, ___0_____40587, ___0_____40588, ___0_____40589,
       ___0_____40592, ___0_____40593, ___0_____40594, ___0_____40595;
  wire ___0_____40596, ___0_____40597, ___0_____40598, ___0_____40600,
       ___0_____40601, ___0_____40602, ___0_____40603, ___0_____40604;
  wire ___0_____40605, ___0_____40606, ___0_____40607, ___0_____40610,
       ___0_____40611, ___0_____40612, ___0_____40613, ___0_____40614;
  wire ___0_____40615, ___0_____40616, ___0_____40617, ___0_____40620,
       ___0_____40621, ___0_____40622, ___0_____40623, ___0_____40624;
  wire ___0_____40625, ___0_____40626, ___0_____40627, ___0_____40630,
       ___0_____40631, ___0_____40632, ___0_____40633, ___0_____40634;
  wire ___0_____40635, ___0_____40636, ___0_____40637, ___0_____40640,
       ___0_____40641, ___0_____40642, ___0_____40643, ___0_____40644;
  wire ___0_____40646, ___0_____40647, ___0_____40649, ___0_____40650,
       ___0_____40651, ___0_____40652, ___0009__30554, ___0009__39901;
  wire ___009, ___009__23224, ___009__24177, ___009__25134,
       ___009__26059, ___009__26959, ___009__27835, ___009__28745;
  wire ___009___30633, ___009___30634, ___009___30635, ___009___30636,
       ___009___30637, ___009___30638, ___009___30639, ___009___30640;
  wire ___009___39974, ___009___39975, ___009___39976, ___009___39977,
       ___009___39978, ___009___39979, ___009___39980, ___009___39981;
  wire ___09, ___09_, ___09_0__31417, ___09_0__31427, ___09_0__31437,
       ___09_0__31447, ___09_0__31456, ___09_0__31466;
  wire ___09_0__31476, ___09_0__31486, ___09_0__40661, ___09_0__40671,
       ___09_0__40681, ___09_0__40690, ___09_0__40700, ___09_9__31426;
  wire ___09_9__31436, ___09_9__31446, ___09_9__31455, ___09_9__31465,
       ___09_9__31475, ___09_9__31485, ___09_9__31493, ___09_9__40660;
  wire ___09_9__40670, ___09_9__40680, ___09_9__40689, ___09_9__40699,
       ___09_9__40709, ___09___22354, ___09___22355, ___09___22356;
  wire ___09___22357, ___09___22358, ___09___22359, ___09___22360,
       ___09___23302, ___09___23303, ___09___23304, ___09___23305;
  wire ___09___23306, ___09___23307, ___09___23308, ___09___24258,
       ___09___24259, ___09___24260, ___09___24261, ___09___24262;
  wire ___09___24263, ___09___24264, ___09___24265, ___09___25214,
       ___09___25215, ___09___25216, ___09___25217, ___09___25218;
  wire ___09___25219, ___09___25220, ___09___26133, ___09___26134,
       ___09___26135, ___09___26136, ___09___26137, ___09___26138;
  wire ___09___27027, ___09___27028, ___09___27029, ___09___27913,
       ___09___27914, ___09___27915, ___09___27916, ___09___27917;
  wire ___09___27918, ___09___27919, ___09___27920, ___09___28825,
       ___09___28826, ___09___28827, ___09___28828, ___09___28829;
  wire ___09___28830, ___09___28831, ___09___28832, ___09____31418,
       ___09____31419, ___09____31420, ___09____31421, ___09____31422;
  wire ___09____31423, ___09____31424, ___09____31425, ___09____31428,
       ___09____31429, ___09____31430, ___09____31431, ___09____31432;
  wire ___09____31433, ___09____31434, ___09____31435, ___09____31438,
       ___09____31439, ___09____31440, ___09____31441, ___09____31442;
  wire ___09____31443, ___09____31444, ___09____31445, ___09____31448,
       ___09____31449, ___09____31450, ___09____31451, ___09____31452;
  wire ___09____31453, ___09____31454, ___09____31457, ___09____31458,
       ___09____31459, ___09____31460, ___09____31461, ___09____31462;
  wire ___09____31463, ___09____31464, ___09____31467, ___09____31468,
       ___09____31469, ___09____31470, ___09____31471, ___09____31472;
  wire ___09____31473, ___09____31474, ___09____31477, ___09____31478,
       ___09____31479, ___09____31480, ___09____31481, ___09____31482;
  wire ___09____31483, ___09____31484, ___09____31487, ___09____31488,
       ___09____31489, ___09____31490, ___09____31491, ___09____31492;
  wire ___09____40657, ___09____40658, ___09____40659, ___09____40662,
       ___09____40663, ___09____40664, ___09____40665, ___09____40666;
  wire ___09____40667, ___09____40668, ___09____40669, ___09____40672,
       ___09____40673, ___09____40674, ___09____40675, ___09____40676;
  wire ___09____40677, ___09____40678, ___09____40679, ___09____40682,
       ___09____40683, ___09____40684, ___09____40685, ___09____40686;
  wire ___09____40687, ___09____40688, ___09____40691, ___09____40692,
       ___09____40693, ___09____40694, ___09____40695, ___09____40696;
  wire ___09____40697, ___09____40698, ___09____40701, ___09____40702,
       ___09____40703, ___09____40704, ___09____40705, ___09____40706;
  wire ___09____40707, ___09____40708, ___9, ___9_, ___9_0,
       ___9_00__39071, ___9_00__39162, ___9_00__39251;
  wire ___9_00__39342, ___9_00__39433, ___9_00__39527, ___9_00__39617,
       ___9_00__39703, ___9_0__23155, ___9_0__23173, ___9_0__23182;
  wire ___9_0__23192, ___9_0__23201, ___9_0__24080, ___9_0__24090,
       ___9_0__24100, ___9_0__24109, ___9_0__24119, ___9_0__24129;
  wire ___9_0__24139, ___9_0__24149, ___9_0__25038, ___9_0__25048,
       ___9_0__25058, ___9_0__25068, ___9_0__25078, ___9_0__25087;
  wire ___9_0__25095, ___9_0__25105, ___9_0__25968, ___9_0__25978,
       ___9_0__25988, ___9_0__26004, ___9_0__26013, ___9_0__26021;
  wire ___9_0__26031, ___9_0__26873, ___9_0__26883, ___9_0__26892,
       ___9_0__26901, ___9_0__26911, ___9_0__26920, ___9_0__26930;
  wire ___9_0__26940, ___9_0__27752, ___9_0__27768, ___9_0__27777,
       ___9_0__27786, ___9_0__27795, ___9_0__27805, ___9_0__28655;
  wire ___9_0__28664, ___9_0__28673, ___9_0__28681, ___9_0__28689,
       ___9_0__28698, ___9_0__28708, ___9_0__28718, ___9_0__29570;
  wire ___9_0__29576, ___9_0__29586, ___9_0__29593, ___9_0__29602,
       ___9_0__29611, ___9_0__29620, ___9_0___39072, ___9_0___39073;
  wire ___9_0___39074, ___9_0___39075, ___9_0___39076, ___9_0___39077,
       ___9_0___39163, ___9_0___39164, ___9_0___39165, ___9_0___39166;
  wire ___9_0___39167, ___9_0___39168, ___9_0___39169, ___9_0___39170,
       ___9_0___39252, ___9_0___39253, ___9_0___39254, ___9_0___39255;
  wire ___9_0___39256, ___9_0___39257, ___9_0___39258, ___9_0___39259,
       ___9_0___39343, ___9_0___39344, ___9_0___39345, ___9_0___39346;
  wire ___9_0___39347, ___9_0___39348, ___9_0___39349, ___9_0___39350,
       ___9_0___39434, ___9_0___39435, ___9_0___39436, ___9_0___39437;
  wire ___9_0___39438, ___9_0___39439, ___9_0___39440, ___9_0___39441,
       ___9_0___39528, ___9_0___39529, ___9_0___39530, ___9_0___39531;
  wire ___9_0___39532, ___9_0___39533, ___9_0___39534, ___9_0___39618,
       ___9_0___39619, ___9_0___39620, ___9_0___39621, ___9_0___39622;
  wire ___9_0___39623, ___9_0___39624, ___9_0___39704, ___9_0___39705,
       ___9_0___39706, ___9_0___39707, ___9_0___39708, ___9_0___39709;
  wire ___9_0___39710, ___9_0___39711, ___9_09__39078, ___9_09__39171,
       ___9_09__39260, ___9_09__39351, ___9_09__39442, ___9_09__39535;
  wire ___9_09__39625, ___9_09__39712, ___9_9, ___9_9__23154,
       ___9_9__23163, ___9_9__23172, ___9_9__23181, ___9_9__23191;
  wire ___9_9__23200, ___9_9__23208, ___9_9__24089, ___9_9__24099,
       ___9_9__24108, ___9_9__24118, ___9_9__24128, ___9_9__24138;
  wire ___9_9__24148, ___9_9__24157, ___9_9__25047, ___9_9__25057,
       ___9_9__25067, ___9_9__25077, ___9_9__25094, ___9_9__25104;
  wire ___9_9__25114, ___9_9__25977, ___9_9__25987, ___9_9__25996,
       ___9_9__26003, ___9_9__26012, ___9_9__26020, ___9_9__26030;
  wire ___9_9__26040, ___9_9__26882, ___9_9__26891, ___9_9__26910,
       ___9_9__26919, ___9_9__26929, ___9_9__26939, ___9_9__26948;
  wire ___9_9__27761, ___9_9__27767, ___9_9__27776, ___9_9__27785,
       ___9_9__27794, ___9_9__27804, ___9_9__27813, ___9_9__27821;
  wire ___9_9__28663, ___9_9__28672, ___9_9__28680, ___9_9__28688,
       ___9_9__28707, ___9_9__28717, ___9_9__28727, ___9_9__29569;
  wire ___9_9__29585, ___9_9__29601, ___9_9__29610, ___9_9__29619,
       ___9_9__29627, ___9_9___39154, ___9_9___39155, ___9_9___39156;
  wire ___9_9___39157, ___9_9___39158, ___9_9___39159, ___9_9___39160,
       ___9_9___39246, ___9_9___39247, ___9_9___39248, ___9_9___39249;
  wire ___9_9___39335, ___9_9___39336, ___9_9___39337, ___9_9___39338,
       ___9_9___39339, ___9_9___39340, ___9_9___39425, ___9_9___39426;
  wire ___9_9___39427, ___9_9___39428, ___9_9___39429, ___9_9___39430,
       ___9_9___39431, ___9_9___39518, ___9_9___39519, ___9_9___39520;
  wire ___9_9___39521, ___9_9___39522, ___9_9___39523, ___9_9___39524,
       ___9_9___39525, ___9_9___39608, ___9_9___39609, ___9_9___39610;
  wire ___9_9___39611, ___9_9___39612, ___9_9___39613, ___9_9___39614,
       ___9_9___39615, ___9_9___39696, ___9_9___39697, ___9_9___39698;
  wire ___9_9___39699, ___9_9___39700, ___9_9___39701, ___9_9___39702,
       ___9_9___39788, ___9_9___39789, ___9_9___39790, ___9_9___39791;
  wire ___9_9___39792, ___9_9___39793, ___9_9___39794, ___9_9___39795,
       ___9_90__39245, ___9_90__39334, ___9_90__39424, ___9_90__39517;
  wire ___9_90__39607, ___9_90__39695, ___9_90__39787, ___9_99__39161,
       ___9_99__39250, ___9_99__39341, ___9_99__39432, ___9_99__39526;
  wire ___9_99__39616, ___9_99__39796, ___9__, ___9__0__39079,
       ___9__0__39089, ___9__0__39099, ___9__0__39108, ___9__0__39118;
  wire ___9__0__39126, ___9__0__39136, ___9__0__39146, ___9__0__39172,
       ___9__0__39182, ___9__0__39192, ___9__0__39202, ___9__0__39209;
  wire ___9__0__39228, ___9__0__39235, ___9__0__39261, ___9__0__39270,
       ___9__0__39280, ___9__0__39289, ___9__0__39299, ___9__0__39306;
  wire ___9__0__39315, ___9__0__39325, ___9__0__39352, ___9__0__39361,
       ___9__0__39370, ___9__0__39380, ___9__0__39388, ___9__0__39396;
  wire ___9__0__39406, ___9__0__39443, ___9__0__39460, ___9__0__39479,
       ___9__0__39488, ___9__0__39498, ___9__0__39507, ___9__0__39536;
  wire ___9__0__39544, ___9__0__39553, ___9__0__39561, ___9__0__39570,
       ___9__0__39578, ___9__0__39588, ___9__0__39598, ___9__0__39633;
  wire ___9__0__39643, ___9__0__39651, ___9__0__39660, ___9__0__39669,
       ___9__0__39679, ___9__0__39687, ___9__0__39713, ___9__0__39732;
  wire ___9__0__39742, ___9__0__39751, ___9__0__39760, ___9__0__39778,
       ___9__0__41371, ___9__9__39088, ___9__9__39098, ___9__9__39107;
  wire ___9__9__39117, ___9__9__39125, ___9__9__39135, ___9__9__39145,
       ___9__9__39153, ___9__9__39181, ___9__9__39191, ___9__9__39201;
  wire ___9__9__39218, ___9__9__39227, ___9__9__39234, ___9__9__39244,
       ___9__9__39279, ___9__9__39288, ___9__9__39298, ___9__9__39305;
  wire ___9__9__39314, ___9__9__39324, ___9__9__39360, ___9__9__39369,
       ___9__9__39379, ___9__9__39405, ___9__9__39415, ___9__9__39423;
  wire ___9__9__39450, ___9__9__39459, ___9__9__39469, ___9__9__39478,
       ___9__9__39487, ___9__9__39497, ___9__9__39506, ___9__9__39516;
  wire ___9__9__39543, ___9__9__39552, ___9__9__39560, ___9__9__39569,
       ___9__9__39577, ___9__9__39587, ___9__9__39597, ___9__9__39606;
  wire ___9__9__39632, ___9__9__39642, ___9__9__39650, ___9__9__39659,
       ___9__9__39668, ___9__9__39678, ___9__9__39686, ___9__9__39694;
  wire ___9__9__39722, ___9__9__39731, ___9__9__39741, ___9__9__39759,
       ___9__9__39768, ___9__9__39777, ___9__9__39786, ___9__22133;
  wire ___9__22137, ___9__22143, ___9__22156, ___9__22165,
       ___9___22190, ___9___22191, ___9___22192, ___9___22193;
  wire ___9___22194, ___9___22195, ___9___22263, ___9___22264,
       ___9___22265, ___9___22266, ___9___22267, ___9___22268;
  wire ___9___22269, ___9___22270, ___9____23140, ___9____23141,
       ___9____23142, ___9____23143, ___9____23144, ___9____23145;
  wire ___9____23146, ___9____23147, ___9____23148, ___9____23149,
       ___9____23150, ___9____23151, ___9____23152, ___9____23153;
  wire ___9____23156, ___9____23157, ___9____23158, ___9____23159,
       ___9____23160, ___9____23161, ___9____23162, ___9____23164;
  wire ___9____23165, ___9____23166, ___9____23167, ___9____23168,
       ___9____23169, ___9____23170, ___9____23171, ___9____23174;
  wire ___9____23175, ___9____23176, ___9____23177, ___9____23178,
       ___9____23179, ___9____23180, ___9____23183, ___9____23184;
  wire ___9____23185, ___9____23186, ___9____23187, ___9____23188,
       ___9____23189, ___9____23190, ___9____23193, ___9____23194;
  wire ___9____23195, ___9____23196, ___9____23197, ___9____23198,
       ___9____23199, ___9____23202, ___9____23203, ___9____23204;
  wire ___9____23205, ___9____23206, ___9____23207, ___9____24081,
       ___9____24082, ___9____24083, ___9____24084, ___9____24085;
  wire ___9____24086, ___9____24087, ___9____24088, ___9____24091,
       ___9____24092, ___9____24093, ___9____24094, ___9____24095;
  wire ___9____24096, ___9____24097, ___9____24098, ___9____24101,
       ___9____24102, ___9____24103, ___9____24104, ___9____24105;
  wire ___9____24106, ___9____24107, ___9____24110, ___9____24111,
       ___9____24112, ___9____24113, ___9____24114, ___9____24115;
  wire ___9____24116, ___9____24117, ___9____24120, ___9____24121,
       ___9____24122, ___9____24123, ___9____24124, ___9____24125;
  wire ___9____24126, ___9____24127, ___9____24130, ___9____24131,
       ___9____24132, ___9____24133, ___9____24134, ___9____24135;
  wire ___9____24136, ___9____24137, ___9____24140, ___9____24141,
       ___9____24142, ___9____24143, ___9____24144, ___9____24145;
  wire ___9____24146, ___9____24147, ___9____24150, ___9____24151,
       ___9____24152, ___9____24153, ___9____24154, ___9____24155;
  wire ___9____24156, ___9____25039, ___9____25040, ___9____25041,
       ___9____25042, ___9____25043, ___9____25044, ___9____25045;
  wire ___9____25046, ___9____25049, ___9____25050, ___9____25051,
       ___9____25052, ___9____25053, ___9____25054, ___9____25055;
  wire ___9____25056, ___9____25059, ___9____25060, ___9____25061,
       ___9____25062, ___9____25063, ___9____25064, ___9____25065;
  wire ___9____25066, ___9____25069, ___9____25070, ___9____25071,
       ___9____25072, ___9____25073, ___9____25074, ___9____25075;
  wire ___9____25076, ___9____25079, ___9____25080, ___9____25081,
       ___9____25082, ___9____25083, ___9____25084, ___9____25085;
  wire ___9____25086, ___9____25088, ___9____25089, ___9____25090,
       ___9____25091, ___9____25092, ___9____25093, ___9____25096;
  wire ___9____25097, ___9____25098, ___9____25099, ___9____25100,
       ___9____25101, ___9____25102, ___9____25103, ___9____25106;
  wire ___9____25107, ___9____25108, ___9____25109, ___9____25110,
       ___9____25111, ___9____25112, ___9____25113, ___9____25969;
  wire ___9____25970, ___9____25971, ___9____25972, ___9____25973,
       ___9____25974, ___9____25975, ___9____25976, ___9____25979;
  wire ___9____25980, ___9____25981, ___9____25982, ___9____25983,
       ___9____25984, ___9____25985, ___9____25986, ___9____25989;
  wire ___9____25990, ___9____25991, ___9____25992, ___9____25993,
       ___9____25994, ___9____25995, ___9____25997, ___9____25998;
  wire ___9____25999, ___9____26000, ___9____26001, ___9____26002,
       ___9____26005, ___9____26006, ___9____26007, ___9____26008;
  wire ___9____26009, ___9____26010, ___9____26011, ___9____26014,
       ___9____26015, ___9____26016, ___9____26017, ___9____26018;
  wire ___9____26019, ___9____26022, ___9____26023, ___9____26024,
       ___9____26025, ___9____26026, ___9____26027, ___9____26028;
  wire ___9____26029, ___9____26032, ___9____26033, ___9____26034,
       ___9____26035, ___9____26036, ___9____26037, ___9____26038;
  wire ___9____26039, ___9____26874, ___9____26875, ___9____26876,
       ___9____26877, ___9____26878, ___9____26879, ___9____26880;
  wire ___9____26881, ___9____26884, ___9____26885, ___9____26886,
       ___9____26887, ___9____26888, ___9____26889, ___9____26890;
  wire ___9____26893, ___9____26894, ___9____26895, ___9____26896,
       ___9____26897, ___9____26898, ___9____26899, ___9____26900;
  wire ___9____26902, ___9____26903, ___9____26904, ___9____26905,
       ___9____26906, ___9____26907, ___9____26908, ___9____26909;
  wire ___9____26912, ___9____26913, ___9____26914, ___9____26915,
       ___9____26916, ___9____26917, ___9____26918, ___9____26921;
  wire ___9____26922, ___9____26923, ___9____26924, ___9____26925,
       ___9____26926, ___9____26927, ___9____26928, ___9____26931;
  wire ___9____26932, ___9____26933, ___9____26934, ___9____26935,
       ___9____26936, ___9____26937, ___9____26938, ___9____26941;
  wire ___9____26942, ___9____26943, ___9____26944, ___9____26945,
       ___9____26946, ___9____26947, ___9____27753, ___9____27754;
  wire ___9____27755, ___9____27756, ___9____27757, ___9____27758,
       ___9____27759, ___9____27760, ___9____27762, ___9____27763;
  wire ___9____27764, ___9____27765, ___9____27766, ___9____27769,
       ___9____27770, ___9____27771, ___9____27772, ___9____27773;
  wire ___9____27774, ___9____27775, ___9____27778, ___9____27779,
       ___9____27780, ___9____27781, ___9____27782, ___9____27783;
  wire ___9____27784, ___9____27787, ___9____27788, ___9____27789,
       ___9____27790, ___9____27791, ___9____27792, ___9____27793;
  wire ___9____27796, ___9____27797, ___9____27798, ___9____27799,
       ___9____27800, ___9____27801, ___9____27802, ___9____27803;
  wire ___9____27806, ___9____27807, ___9____27808, ___9____27809,
       ___9____27810, ___9____27811, ___9____27812, ___9____27814;
  wire ___9____27815, ___9____27816, ___9____27817, ___9____27818,
       ___9____27819, ___9____27820, ___9____28656, ___9____28657;
  wire ___9____28658, ___9____28659, ___9____28660, ___9____28661,
       ___9____28662, ___9____28665, ___9____28666, ___9____28667;
  wire ___9____28668, ___9____28669, ___9____28670, ___9____28671,
       ___9____28674, ___9____28675, ___9____28676, ___9____28677;
  wire ___9____28678, ___9____28679, ___9____28682, ___9____28683,
       ___9____28684, ___9____28685, ___9____28686, ___9____28687;
  wire ___9____28690, ___9____28691, ___9____28692, ___9____28693,
       ___9____28694, ___9____28695, ___9____28696, ___9____28697;
  wire ___9____28699, ___9____28700, ___9____28701, ___9____28702,
       ___9____28703, ___9____28704, ___9____28705, ___9____28706;
  wire ___9____28709, ___9____28710, ___9____28711, ___9____28712,
       ___9____28713, ___9____28714, ___9____28715, ___9____28716;
  wire ___9____28719, ___9____28720, ___9____28721, ___9____28722,
       ___9____28723, ___9____28724, ___9____28725, ___9____28726;
  wire ___9____29562, ___9____29563, ___9____29564, ___9____29565,
       ___9____29566, ___9____29567, ___9____29568, ___9____29571;
  wire ___9____29572, ___9____29573, ___9____29574, ___9____29575,
       ___9____29577, ___9____29578, ___9____29579, ___9____29580;
  wire ___9____29581, ___9____29582, ___9____29583, ___9____29584,
       ___9____29587, ___9____29588, ___9____29589, ___9____29590;
  wire ___9____29591, ___9____29592, ___9____29594, ___9____29595,
       ___9____29596, ___9____29597, ___9____29598, ___9____29599;
  wire ___9____29600, ___9____29603, ___9____29604, ___9____29605,
       ___9____29606, ___9____29607, ___9____29608, ___9____29609;
  wire ___9____29612, ___9____29613, ___9____29614, ___9____29615,
       ___9____29616, ___9____29617, ___9____29618, ___9____29621;
  wire ___9____29622, ___9____29623, ___9____29624, ___9____29625,
       ___9____29626, ___9_____39080, ___9_____39081, ___9_____39082;
  wire ___9_____39083, ___9_____39084, ___9_____39085, ___9_____39086,
       ___9_____39087, ___9_____39090, ___9_____39091, ___9_____39092;
  wire ___9_____39093, ___9_____39094, ___9_____39095, ___9_____39096,
       ___9_____39097, ___9_____39100, ___9_____39101, ___9_____39102;
  wire ___9_____39103, ___9_____39104, ___9_____39105, ___9_____39106,
       ___9_____39109, ___9_____39110, ___9_____39111, ___9_____39112;
  wire ___9_____39113, ___9_____39114, ___9_____39115, ___9_____39116,
       ___9_____39119, ___9_____39120, ___9_____39121, ___9_____39122;
  wire ___9_____39123, ___9_____39124, ___9_____39127, ___9_____39128,
       ___9_____39129, ___9_____39130, ___9_____39131, ___9_____39132;
  wire ___9_____39133, ___9_____39134, ___9_____39137, ___9_____39138,
       ___9_____39139, ___9_____39140, ___9_____39141, ___9_____39142;
  wire ___9_____39143, ___9_____39144, ___9_____39147, ___9_____39148,
       ___9_____39149, ___9_____39150, ___9_____39151, ___9_____39152;
  wire ___9_____39173, ___9_____39174, ___9_____39175, ___9_____39176,
       ___9_____39177, ___9_____39178, ___9_____39179, ___9_____39180;
  wire ___9_____39183, ___9_____39184, ___9_____39185, ___9_____39186,
       ___9_____39187, ___9_____39188, ___9_____39189, ___9_____39190;
  wire ___9_____39193, ___9_____39194, ___9_____39195, ___9_____39196,
       ___9_____39197, ___9_____39198, ___9_____39199, ___9_____39200;
  wire ___9_____39203, ___9_____39204, ___9_____39205, ___9_____39206,
       ___9_____39207, ___9_____39208, ___9_____39210, ___9_____39211;
  wire ___9_____39212, ___9_____39213, ___9_____39214, ___9_____39215,
       ___9_____39216, ___9_____39217, ___9_____39219, ___9_____39220;
  wire ___9_____39221, ___9_____39222, ___9_____39223, ___9_____39224,
       ___9_____39225, ___9_____39226, ___9_____39229, ___9_____39230;
  wire ___9_____39231, ___9_____39232, ___9_____39233, ___9_____39236,
       ___9_____39237, ___9_____39238, ___9_____39239, ___9_____39240;
  wire ___9_____39241, ___9_____39242, ___9_____39243, ___9_____39262,
       ___9_____39263, ___9_____39264, ___9_____39265, ___9_____39266;
  wire ___9_____39267, ___9_____39268, ___9_____39269, ___9_____39271,
       ___9_____39272, ___9_____39273, ___9_____39274, ___9_____39275;
  wire ___9_____39276, ___9_____39277, ___9_____39278, ___9_____39281,
       ___9_____39282, ___9_____39283, ___9_____39284, ___9_____39285;
  wire ___9_____39286, ___9_____39287, ___9_____39290, ___9_____39291,
       ___9_____39292, ___9_____39293, ___9_____39294, ___9_____39295;
  wire ___9_____39296, ___9_____39297, ___9_____39300, ___9_____39301,
       ___9_____39302, ___9_____39303, ___9_____39304, ___9_____39307;
  wire ___9_____39308, ___9_____39309, ___9_____39310, ___9_____39311,
       ___9_____39312, ___9_____39313, ___9_____39316, ___9_____39317;
  wire ___9_____39318, ___9_____39319, ___9_____39320, ___9_____39321,
       ___9_____39322, ___9_____39323, ___9_____39326, ___9_____39327;
  wire ___9_____39328, ___9_____39329, ___9_____39330, ___9_____39331,
       ___9_____39332, ___9_____39333, ___9_____39353, ___9_____39354;
  wire ___9_____39355, ___9_____39356, ___9_____39357, ___9_____39358,
       ___9_____39359, ___9_____39362, ___9_____39363, ___9_____39364;
  wire ___9_____39365, ___9_____39366, ___9_____39367, ___9_____39368,
       ___9_____39371, ___9_____39372, ___9_____39373, ___9_____39374;
  wire ___9_____39375, ___9_____39376, ___9_____39377, ___9_____39378,
       ___9_____39381, ___9_____39382, ___9_____39383, ___9_____39384;
  wire ___9_____39385, ___9_____39386, ___9_____39387, ___9_____39389,
       ___9_____39390, ___9_____39391, ___9_____39392, ___9_____39393;
  wire ___9_____39394, ___9_____39395, ___9_____39397, ___9_____39398,
       ___9_____39399, ___9_____39400, ___9_____39401, ___9_____39402;
  wire ___9_____39403, ___9_____39404, ___9_____39407, ___9_____39408,
       ___9_____39409, ___9_____39410, ___9_____39411, ___9_____39412;
  wire ___9_____39413, ___9_____39414, ___9_____39416, ___9_____39417,
       ___9_____39418, ___9_____39419, ___9_____39420, ___9_____39421;
  wire ___9_____39422, ___9_____39444, ___9_____39445, ___9_____39446,
       ___9_____39447, ___9_____39448, ___9_____39449, ___9_____39451;
  wire ___9_____39452, ___9_____39453, ___9_____39454, ___9_____39455,
       ___9_____39456, ___9_____39457, ___9_____39458, ___9_____39461;
  wire ___9_____39462, ___9_____39463, ___9_____39464, ___9_____39465,
       ___9_____39466, ___9_____39467, ___9_____39468, ___9_____39470;
  wire ___9_____39471, ___9_____39472, ___9_____39473, ___9_____39474,
       ___9_____39475, ___9_____39476, ___9_____39477, ___9_____39480;
  wire ___9_____39481, ___9_____39482, ___9_____39483, ___9_____39484,
       ___9_____39485, ___9_____39486, ___9_____39489, ___9_____39490;
  wire ___9_____39491, ___9_____39492, ___9_____39493, ___9_____39494,
       ___9_____39495, ___9_____39496, ___9_____39499, ___9_____39500;
  wire ___9_____39501, ___9_____39502, ___9_____39503, ___9_____39504,
       ___9_____39505, ___9_____39508, ___9_____39509, ___9_____39510;
  wire ___9_____39511, ___9_____39512, ___9_____39513, ___9_____39514,
       ___9_____39515, ___9_____39537, ___9_____39538, ___9_____39539;
  wire ___9_____39540, ___9_____39541, ___9_____39542, ___9_____39545,
       ___9_____39546, ___9_____39547, ___9_____39548, ___9_____39549;
  wire ___9_____39550, ___9_____39551, ___9_____39554, ___9_____39555,
       ___9_____39556, ___9_____39557, ___9_____39558, ___9_____39559;
  wire ___9_____39562, ___9_____39563, ___9_____39564, ___9_____39565,
       ___9_____39566, ___9_____39567, ___9_____39568, ___9_____39571;
  wire ___9_____39572, ___9_____39573, ___9_____39574, ___9_____39575,
       ___9_____39576, ___9_____39579, ___9_____39580, ___9_____39581;
  wire ___9_____39582, ___9_____39583, ___9_____39584, ___9_____39585,
       ___9_____39586, ___9_____39589, ___9_____39590, ___9_____39591;
  wire ___9_____39592, ___9_____39593, ___9_____39594, ___9_____39595,
       ___9_____39596, ___9_____39599, ___9_____39600, ___9_____39601;
  wire ___9_____39602, ___9_____39603, ___9_____39604, ___9_____39605,
       ___9_____39626, ___9_____39627, ___9_____39628, ___9_____39629;
  wire ___9_____39630, ___9_____39631, ___9_____39634, ___9_____39635,
       ___9_____39636, ___9_____39637, ___9_____39638, ___9_____39639;
  wire ___9_____39640, ___9_____39641, ___9_____39644, ___9_____39645,
       ___9_____39646, ___9_____39647, ___9_____39648, ___9_____39649;
  wire ___9_____39652, ___9_____39653, ___9_____39654, ___9_____39655,
       ___9_____39656, ___9_____39657, ___9_____39658, ___9_____39661;
  wire ___9_____39662, ___9_____39663, ___9_____39664, ___9_____39665,
       ___9_____39666, ___9_____39667, ___9_____39670, ___9_____39671;
  wire ___9_____39672, ___9_____39673, ___9_____39674, ___9_____39675,
       ___9_____39676, ___9_____39677, ___9_____39680, ___9_____39681;
  wire ___9_____39682, ___9_____39683, ___9_____39684, ___9_____39685,
       ___9_____39688, ___9_____39689, ___9_____39690, ___9_____39691;
  wire ___9_____39692, ___9_____39693, ___9_____39714, ___9_____39715,
       ___9_____39716, ___9_____39717, ___9_____39718, ___9_____39719;
  wire ___9_____39720, ___9_____39721, ___9_____39723, ___9_____39724,
       ___9_____39725, ___9_____39726, ___9_____39727, ___9_____39728;
  wire ___9_____39729, ___9_____39730, ___9_____39733, ___9_____39734,
       ___9_____39735, ___9_____39736, ___9_____39737, ___9_____39738;
  wire ___9_____39739, ___9_____39740, ___9_____39743, ___9_____39744,
       ___9_____39745, ___9_____39746, ___9_____39747, ___9_____39748;
  wire ___9_____39749, ___9_____39750, ___9_____39752, ___9_____39753,
       ___9_____39754, ___9_____39755, ___9_____39756, ___9_____39757;
  wire ___9_____39758, ___9_____39761, ___9_____39762, ___9_____39763,
       ___9_____39764, ___9_____39765, ___9_____39766, ___9_____39767;
  wire ___9_____39769, ___9_____39770, ___9_____39771, ___9_____39772,
       ___9_____39773, ___9_____39774, ___9_____39775, ___9_____39776;
  wire ___9_____39779, ___9_____39780, ___9_____39781, ___9_____39782,
       ___9_____39783, ___9_____39784, ___9_____39785, ___0090__30632;
  wire ___0090__39973, ___090, ___090__23301, ___090__24257,
       ___090__25213, ___090__26132, ___090__27026, ___090__27912;
  wire ___090___31408, ___090___31409, ___090___31410, ___090___31411,
       ___090___31412, ___090___31413, ___090___31414, ___090___31415;
  wire ___90, ___90_, ___90_0__38988, ___90_0__38998, ___90_0__39005,
       ___90_0__39015, ___90_0__39025, ___90_0__39035;
  wire ___90_0__39044, ___90_0__39054, ___90_9__38997, ___90_9__39004,
       ___90_9__39014, ___90_9__39024, ___90_9__39034, ___90_9__39053;
  wire ___90_9__39061, ___90__22262, ___90___23134, ___90___23135,
       ___90___23136, ___90___23137, ___90___23138, ___90___23139;
  wire ___90___24071, ___90___24072, ___90___24073, ___90___24074,
       ___90___24075, ___90___24076, ___90___24077, ___90___24078;
  wire ___90___25030, ___90___25031, ___90___25032, ___90___25033,
       ___90___25034, ___90___25035, ___90___25036, ___90___25959;
  wire ___90___25960, ___90___25961, ___90___25962, ___90___25963,
       ___90___25964, ___90___25965, ___90___25966, ___90___26865;
  wire ___90___26866, ___90___26867, ___90___26868, ___90___26869,
       ___90___26870, ___90___26871, ___90___27743, ___90___27744;
  wire ___90___27745, ___90___27746, ___90___27747, ___90___27748,
       ___90___27749, ___90___27750, ___90___28647, ___90___28648;
  wire ___90___28649, ___90___28650, ___90___28651, ___90___28652,
       ___90___28653, ___90___29554, ___90___29555, ___90___29556;
  wire ___90___29557, ___90___29558, ___90___29559, ___90___29560,
       ___90____38989, ___90____38990, ___90____38991, ___90____38992;
  wire ___90____38993, ___90____38994, ___90____38995, ___90____38996,
       ___90____38999, ___90____39000, ___90____39001, ___90____39002;
  wire ___90____39003, ___90____39006, ___90____39007, ___90____39008,
       ___90____39009, ___90____39010, ___90____39011, ___90____39012;
  wire ___90____39013, ___90____39016, ___90____39017, ___90____39018,
       ___90____39019, ___90____39020, ___90____39021, ___90____39022;
  wire ___90____39023, ___90____39026, ___90____39027, ___90____39028,
       ___90____39029, ___90____39030, ___90____39031, ___90____39032;
  wire ___90____39033, ___90____39036, ___90____39037, ___90____39038,
       ___90____39039, ___90____39040, ___90____39041, ___90____39042;
  wire ___90____39043, ___90____39045, ___90____39046, ___90____39047,
       ___90____39048, ___90____39049, ___90____39050, ___90____39051;
  wire ___90____39052, ___90____39055, ___90____39056, ___90____39057,
       ___90____39058, ___90____39059, ___90____39060, ___0099__30641;
  wire ___0099__39982, ___099, ___099__23309, ___099__24266,
       ___099__25221, ___099__26139, ___099__27030, ___099__27921;
  wire ___099__28833, ___099___31495, ___099___31496, ___099___31497,
       ___099___31498, ___099___31499, ___099___31500, ___099___31501;
  wire ___099___40711, ___099___40712, ___099___40713, ___099___40714,
       ___099___40715, ___099___40716, ___099___40717, ___099___40718;
  wire ___99, ___99_, ___99_0__39807, ___99_0__39817, ___99_0__39827,
       ___99_0__39837, ___99_0__39845, ___99_0__39855;
  wire ___99_0__39864, ___99_0__39873, ___99_9__39816, ___99_9__39826,
       ___99_9__39836, ___99_9__39844, ___99_9__39854, ___99_9__39863;
  wire ___99_9__39872, ___99_9__39882, ___99__22271, ___99___23209,
       ___99___23210, ___99___23211, ___99___23212, ___99___23213;
  wire ___99___23214, ___99___23215, ___99___24159, ___99___24160,
       ___99___24161, ___99___24162, ___99___24163, ___99___24164;
  wire ___99___24165, ___99___24166, ___99___25116, ___99___25117,
       ___99___25118, ___99___25119, ___99___25120, ___99___25121;
  wire ___99___25122, ___99___25123, ___99___26042, ___99___26043,
       ___99___26044, ___99___26045, ___99___26046, ___99___26047;
  wire ___99___26048, ___99___26049, ___99___26950, ___99___26951,
       ___99___26952, ___99___26953, ___99___27823, ___99___27824;
  wire ___99___27825, ___99___27826, ___99___28729, ___99___28730,
       ___99___28731, ___99___28732, ___99___28733, ___99___28734;
  wire ___99___29629, ___99___29630, ___99___29631, ___99___29632,
       ___99___29633, ___99___29634, ___99___29635, ___99___29636;
  wire ___99____39808, ___99____39809, ___99____39810, ___99____39811,
       ___99____39812, ___99____39813, ___99____39814, ___99____39815;
  wire ___99____39818, ___99____39819, ___99____39820, ___99____39821,
       ___99____39822, ___99____39823, ___99____39824, ___99____39825;
  wire ___99____39828, ___99____39829, ___99____39830, ___99____39831,
       ___99____39832, ___99____39833, ___99____39834, ___99____39835;
  wire ___99____39838, ___99____39839, ___99____39840, ___99____39841,
       ___99____39842, ___99____39843, ___99____39846, ___99____39847;
  wire ___99____39848, ___99____39849, ___99____39850, ___99____39851,
       ___99____39852, ___99____39853, ___99____39856, ___99____39857;
  wire ___99____39858, ___99____39859, ___99____39860, ___99____39861,
       ___99____39862, ___99____39865, ___99____39866, ___99____39867;
  wire ___99____39868, ___99____39869, ___99____39870, ___99____39871,
       ___99____39874, ___99____39875, ___99____39876, ___99____39877;
  wire ___99____39878, ___99____39879, ___99____39880, ___99____39881,
       ___0900, ___900, ___900__24070, ___900__25029;
  wire ___900__25958, ___900__26864, ___900__27742, ___900__28646,
       ___900__29553, ___900___38979, ___900___38980, ___900___38981;
  wire ___900___38982, ___900___38983, ___900___38984, ___900___38985,
       ___900___38986, ___0909__31416, ___0909__40655, ___909;
  wire ___909__24079, ___909__25037, ___909__25967, ___909__26872,
       ___909__27751, ___909__28654, ___909__29561, ___909___39063;
  wire ___909___39064, ___909___39065, ___909___39066, ___909___39067,
       ___909___39068, ___909___39069, ___0990__31494, ___0990__40710;
  wire ___990, ___990__24158, ___990__25115, ___990__26041,
       ___990__26949, ___990__27822, ___990__28728, ___990__29628;
  wire ___990___39798, ___990___39799, ___990___39800, ___990___39801,
       ___990___39802, ___990___39803, ___990___39804, ___990___39805;
  wire ___0999__31502, ___0999__40719, ___999, ___999__24167,
       ___999__25124, ___999__26050, ___999__28735, ___999__29637;
  wire ___999___39884, ___999___39885, ___999___39886, ___999___39887,
       ___999___39888, ___999___39889, ___999___39890, ___9000__38978;
  wire ___9009__38987, ___9090__39062, ___9099__39070, ___9900__39797,
       ___9909__39806, ___9990__39883, ___9999__39891, ____;
  wire ____0, ____00, ____000__31503, ____000__33433, ____000__34387,
       ____000__35289, ____000__36182, ____000__37100;
  wire ____000__38038, ____000__40720, ____00__22450, ____00__22549,
       ____00__22644, ____00__22741, ____00__22839, ____00__22939;
  wire ____00__23039, ____00__23407, ____00__23502, ____00__23597,
       ____00__23692, ____00__23788, ____00__23881, ____00__23972;
  wire ____00__24267, ____00__24364, ____00__24458, ____00__24556,
       ____00__24646, ____00__24746, ____00__24839, ____00__24935;
  wire ____00__25222, ____00__25310, ____00__25407, ____00__25497,
       ____00__25586, ____00__25678, ____00__25768, ____00__25862;
  wire ____00__26140, ____00__26229, ____00__26323, ____00__26408,
       ____00__26499, ____00__26589, ____00__26775, ____00__27031;
  wire ____00__27300, ____00__27392, ____00__27480, ____00__27569,
       ____00__27654, ____00__27922, ____00__28014, ____00__28108;
  wire ____00__28200, ____00__28291, ____00__28376, ____00__28471,
       ____00__28834, ____00__28924, ____00__29009, ____00__29097;
  wire ____00__29194, ____00__29279, ____00__29369, ____00__29466,
       ____00___31504, ____00___31505, ____00___31506, ____00___31507;
  wire ____00___31508, ____00___31509, ____00___31510, ____00___31511,
       ____00___32480, ____00___32481, ____00___32482, ____00___32483;
  wire ____00___32484, ____00___32485, ____00___32486, ____00___33434,
       ____00___33435, ____00___33436, ____00___33437, ____00___33438;
  wire ____00___33439, ____00___33440, ____00___34388, ____00___34389,
       ____00___34390, ____00___34391, ____00___34392, ____00___34393;
  wire ____00___34394, ____00___35290, ____00___35291, ____00___35292,
       ____00___35293, ____00___35294, ____00___35295, ____00___35296;
  wire ____00___35297, ____00___36183, ____00___36184, ____00___36185,
       ____00___36186, ____00___36187, ____00___36188, ____00___36189;
  wire ____00___36190, ____00___37101, ____00___37102, ____00___37103,
       ____00___37104, ____00___37105, ____00___37106, ____00___37107;
  wire ____00___38039, ____00___38040, ____00___38041, ____00___38042,
       ____00___38043, ____00___38044, ____00___38045, ____00___38046;
  wire ____00___40721, ____00___40722, ____00___40723, ____00___40724,
       ____00___40725, ____00___40726, ____00___40727, ____00___40728;
  wire ____0_, ____0_0__31513, ____0_0__31523, ____0_0__31533,
       ____0_0__31543, ____0_0__31553, ____0_0__31563, ____0_0__31573;
  wire ____0_0__31583, ____0_0__32488, ____0_0__32498, ____0_0__32508,
       ____0_0__32518, ____0_0__32527, ____0_0__32537, ____0_0__32547;
  wire ____0_0__32557, ____0_0__33442, ____0_0__33452, ____0_0__33462,
       ____0_0__33471, ____0_0__33480, ____0_0__33490, ____0_0__33500;
  wire ____0_0__33510, ____0_0__34396, ____0_0__34414, ____0_0__34423,
       ____0_0__34432, ____0_0__34441, ____0_0__34451, ____0_0__34460;
  wire ____0_0__35298, ____0_0__35306, ____0_0__35315, ____0_0__35324,
       ____0_0__35334, ____0_0__35341, ____0_0__35350, ____0_0__35360;
  wire ____0_0__36192, ____0_0__36201, ____0_0__36209, ____0_0__36219,
       ____0_0__36229, ____0_0__36239, ____0_0__36249, ____0_0__36258;
  wire ____0_0__37109, ____0_0__37116, ____0_0__37124, ____0_0__37134,
       ____0_0__37144, ____0_0__37151, ____0_0__37159, ____0_0__37169;
  wire ____0_0__38056, ____0_0__38064, ____0_0__38074, ____0_0__38084,
       ____0_0__38093, ____0_0__38102, ____0_0__38112, ____0_0__40730;
  wire ____0_0__40740, ____0_0__40750, ____0_0__40760, ____0_0__40770,
       ____0_0__40780, ____0_0__40790, ____0_0__40800, ____0_9__31522;
  wire ____0_9__31532, ____0_9__31542, ____0_9__31552, ____0_9__31562,
       ____0_9__31572, ____0_9__31582, ____0_9__31592, ____0_9__32497;
  wire ____0_9__32507, ____0_9__32517, ____0_9__32526, ____0_9__32536,
       ____0_9__32546, ____0_9__32556, ____0_9__32566, ____0_9__33451;
  wire ____0_9__33461, ____0_9__33470, ____0_9__33479, ____0_9__33489,
       ____0_9__33499, ____0_9__33509, ____0_9__33519, ____0_9__34413;
  wire ____0_9__34431, ____0_9__34440, ____0_9__34450, ____0_9__34459,
       ____0_9__34469, ____0_9__35305, ____0_9__35314, ____0_9__35323;
  wire ____0_9__35333, ____0_9__35349, ____0_9__35359, ____0_9__35369,
       ____0_9__36200, ____0_9__36208, ____0_9__36218, ____0_9__36228;
  wire ____0_9__36238, ____0_9__36248, ____0_9__36257, ____0_9__36267,
       ____0_9__37123, ____0_9__37133, ____0_9__37143, ____0_9__37158;
  wire ____0_9__37168, ____0_9__37178, ____0_9__38055, ____0_9__38063,
       ____0_9__38073, ____0_9__38083, ____0_9__38101, ____0_9__38111;
  wire ____0_9__38121, ____0_9__40739, ____0_9__40749, ____0_9__40759,
       ____0_9__40769, ____0_9__40779, ____0_9__40789, ____0_9__40799;
  wire ____0_9__40809, ____0__22205, ____0__22215, ____0__22225,
       ____0__22235, ____0__22247, ____0__22281, ____0___22361;
  wire ____0___22362, ____0___22363, ____0___22364, ____0___22365,
       ____0___22366, ____0___22367, ____0___22451, ____0___22452;
  wire ____0___22453, ____0___22454, ____0___22455, ____0___22456,
       ____0___22457, ____0___22550, ____0___22551, ____0___22552;
  wire ____0___22553, ____0___22554, ____0___22555, ____0___22556,
       ____0___22557, ____0___22645, ____0___22646, ____0___22647;
  wire ____0___22648, ____0___22649, ____0___22650, ____0___22651,
       ____0___22652, ____0___22742, ____0___22743, ____0___22744;
  wire ____0___22745, ____0___22746, ____0___22747, ____0___22748,
       ____0___22749, ____0___22840, ____0___22841, ____0___22842;
  wire ____0___22843, ____0___22844, ____0___22845, ____0___22846,
       ____0___22847, ____0___22940, ____0___22941, ____0___22942;
  wire ____0___22943, ____0___22944, ____0___22945, ____0___22946,
       ____0___22947, ____0___23040, ____0___23041, ____0___23042;
  wire ____0___23043, ____0___23044, ____0___23045, ____0___23046,
       ____0___23047, ____0___23310, ____0___23311, ____0___23312;
  wire ____0___23313, ____0___23314, ____0___23315, ____0___23316,
       ____0___23317, ____0___23408, ____0___23409, ____0___23410;
  wire ____0___23411, ____0___23412, ____0___23413, ____0___23414,
       ____0___23415, ____0___23503, ____0___23504, ____0___23505;
  wire ____0___23506, ____0___23507, ____0___23508, ____0___23509,
       ____0___23598, ____0___23599, ____0___23600, ____0___23601;
  wire ____0___23602, ____0___23603, ____0___23604, ____0___23605,
       ____0___23693, ____0___23694, ____0___23695, ____0___23696;
  wire ____0___23697, ____0___23698, ____0___23699, ____0___23700,
       ____0___23789, ____0___23790, ____0___23791, ____0___23792;
  wire ____0___23793, ____0___23794, ____0___23795, ____0___23882,
       ____0___23883, ____0___23884, ____0___23885, ____0___23886;
  wire ____0___23887, ____0___23888, ____0___23889, ____0___23973,
       ____0___23974, ____0___23975, ____0___23976, ____0___23977;
  wire ____0___23978, ____0___23979, ____0___23980, ____0___24268,
       ____0___24269, ____0___24270, ____0___24271, ____0___24272;
  wire ____0___24273, ____0___24274, ____0___24275, ____0___24365,
       ____0___24366, ____0___24367, ____0___24368, ____0___24369;
  wire ____0___24370, ____0___24371, ____0___24459, ____0___24460,
       ____0___24461, ____0___24462, ____0___24463, ____0___24464;
  wire ____0___24465, ____0___24466, ____0___24557, ____0___24558,
       ____0___24559, ____0___24560, ____0___24561, ____0___24562;
  wire ____0___24563, ____0___24564, ____0___24647, ____0___24648,
       ____0___24649, ____0___24650, ____0___24651, ____0___24652;
  wire ____0___24653, ____0___24654, ____0___24747, ____0___24748,
       ____0___24749, ____0___24750, ____0___24751, ____0___24752;
  wire ____0___24753, ____0___24754, ____0___24840, ____0___24841,
       ____0___24842, ____0___24843, ____0___24844, ____0___24845;
  wire ____0___24846, ____0___24847, ____0___24936, ____0___24937,
       ____0___24938, ____0___24939, ____0___24940, ____0___24941;
  wire ____0___24942, ____0___24943, ____0___25223, ____0___25224,
       ____0___25225, ____0___25226, ____0___25227, ____0___25228;
  wire ____0___25229, ____0___25311, ____0___25312, ____0___25313,
       ____0___25314, ____0___25315, ____0___25316, ____0___25317;
  wire ____0___25408, ____0___25409, ____0___25410, ____0___25411,
       ____0___25412, ____0___25413, ____0___25414, ____0___25415;
  wire ____0___25498, ____0___25499, ____0___25500, ____0___25501,
       ____0___25502, ____0___25503, ____0___25504, ____0___25505;
  wire ____0___25587, ____0___25588, ____0___25589, ____0___25590,
       ____0___25591, ____0___25592, ____0___25593, ____0___25594;
  wire ____0___25679, ____0___25680, ____0___25681, ____0___25682,
       ____0___25683, ____0___25684, ____0___25685, ____0___25686;
  wire ____0___25769, ____0___25770, ____0___25771, ____0___25772,
       ____0___25773, ____0___25774, ____0___25775, ____0___25776;
  wire ____0___25863, ____0___25864, ____0___25865, ____0___25866,
       ____0___25867, ____0___25868, ____0___25869, ____0___25870;
  wire ____0___26141, ____0___26142, ____0___26143, ____0___26144,
       ____0___26145, ____0___26146, ____0___26147, ____0___26230;
  wire ____0___26231, ____0___26232, ____0___26233, ____0___26234,
       ____0___26235, ____0___26236, ____0___26237, ____0___26324;
  wire ____0___26325, ____0___26326, ____0___26327, ____0___26328,
       ____0___26329, ____0___26330, ____0___26409, ____0___26410;
  wire ____0___26411, ____0___26412, ____0___26413, ____0___26414,
       ____0___26415, ____0___26416, ____0___26500, ____0___26501;
  wire ____0___26502, ____0___26503, ____0___26504, ____0___26505,
       ____0___26506, ____0___26590, ____0___26591, ____0___26592;
  wire ____0___26593, ____0___26594, ____0___26595, ____0___26596,
       ____0___26597, ____0___26683, ____0___26684, ____0___26685;
  wire ____0___26686, ____0___26687, ____0___26688, ____0___26689,
       ____0___26690, ____0___26776, ____0___26777, ____0___26778;
  wire ____0___26779, ____0___26780, ____0___26781, ____0___26782,
       ____0___26783, ____0___27032, ____0___27033, ____0___27034;
  wire ____0___27035, ____0___27036, ____0___27037, ____0___27121,
       ____0___27122, ____0___27123, ____0___27124, ____0___27125;
  wire ____0___27126, ____0___27127, ____0___27209, ____0___27210,
       ____0___27211, ____0___27212, ____0___27213, ____0___27214;
  wire ____0___27301, ____0___27302, ____0___27303, ____0___27304,
       ____0___27305, ____0___27306, ____0___27393, ____0___27394;
  wire ____0___27395, ____0___27396, ____0___27397, ____0___27398,
       ____0___27399, ____0___27481, ____0___27482, ____0___27483;
  wire ____0___27484, ____0___27485, ____0___27486, ____0___27487,
       ____0___27488, ____0___27570, ____0___27571, ____0___27572;
  wire ____0___27573, ____0___27574, ____0___27575, ____0___27576,
       ____0___27655, ____0___27656, ____0___27657, ____0___27658;
  wire ____0___27923, ____0___27924, ____0___27925, ____0___27926,
       ____0___27927, ____0___27928, ____0___27929, ____0___27930;
  wire ____0___28015, ____0___28016, ____0___28017, ____0___28018,
       ____0___28019, ____0___28020, ____0___28021, ____0___28109;
  wire ____0___28110, ____0___28111, ____0___28112, ____0___28113,
       ____0___28114, ____0___28115, ____0___28116, ____0___28201;
  wire ____0___28202, ____0___28203, ____0___28204, ____0___28205,
       ____0___28206, ____0___28207, ____0___28208, ____0___28292;
  wire ____0___28293, ____0___28294, ____0___28295, ____0___28296,
       ____0___28297, ____0___28377, ____0___28378, ____0___28379;
  wire ____0___28380, ____0___28381, ____0___28382, ____0___28383,
       ____0___28472, ____0___28473, ____0___28474, ____0___28475;
  wire ____0___28476, ____0___28477, ____0___28478, ____0___28479,
       ____0___28554, ____0___28555, ____0___28556, ____0___28557;
  wire ____0___28558, ____0___28559, ____0___28560, ____0___28835,
       ____0___28836, ____0___28837, ____0___28838, ____0___28839;
  wire ____0___28840, ____0___28841, ____0___28842, ____0___28925,
       ____0___28926, ____0___28927, ____0___28928, ____0___28929;
  wire ____0___28930, ____0___29010, ____0___29011, ____0___29012,
       ____0___29013, ____0___29014, ____0___29015, ____0___29016;
  wire ____0___29017, ____0___29098, ____0___29099, ____0___29100,
       ____0___29101, ____0___29102, ____0___29103, ____0___29104;
  wire ____0___29105, ____0___29195, ____0___29196, ____0___29197,
       ____0___29198, ____0___29199, ____0___29200, ____0___29201;
  wire ____0___29202, ____0___29280, ____0___29281, ____0___29282,
       ____0___29283, ____0___29284, ____0___29285, ____0___29286;
  wire ____0___29370, ____0___29371, ____0___29372, ____0___29373,
       ____0___29374, ____0___29375, ____0___29376, ____0___29467;
  wire ____0___29468, ____0___29469, ____0___29470, ____0___29471,
       ____0___29472, ____0___29473, ____0___29474, ____0____31514;
  wire ____0____31515, ____0____31516, ____0____31517, ____0____31518,
       ____0____31519, ____0____31520, ____0____31521, ____0____31524;
  wire ____0____31525, ____0____31526, ____0____31527, ____0____31528,
       ____0____31529, ____0____31530, ____0____31531, ____0____31534;
  wire ____0____31535, ____0____31536, ____0____31537, ____0____31538,
       ____0____31539, ____0____31540, ____0____31541, ____0____31544;
  wire ____0____31545, ____0____31546, ____0____31547, ____0____31548,
       ____0____31549, ____0____31550, ____0____31551, ____0____31554;
  wire ____0____31555, ____0____31556, ____0____31557, ____0____31558,
       ____0____31559, ____0____31560, ____0____31561, ____0____31564;
  wire ____0____31565, ____0____31566, ____0____31567, ____0____31568,
       ____0____31569, ____0____31570, ____0____31571, ____0____31574;
  wire ____0____31575, ____0____31576, ____0____31577, ____0____31578,
       ____0____31579, ____0____31580, ____0____31581, ____0____31584;
  wire ____0____31585, ____0____31586, ____0____31587, ____0____31588,
       ____0____31589, ____0____31590, ____0____31591, ____0____32489;
  wire ____0____32490, ____0____32491, ____0____32492, ____0____32493,
       ____0____32494, ____0____32495, ____0____32496, ____0____32499;
  wire ____0____32500, ____0____32501, ____0____32502, ____0____32503,
       ____0____32504, ____0____32505, ____0____32506, ____0____32509;
  wire ____0____32510, ____0____32511, ____0____32512, ____0____32513,
       ____0____32514, ____0____32515, ____0____32516, ____0____32519;
  wire ____0____32520, ____0____32521, ____0____32522, ____0____32523,
       ____0____32524, ____0____32525, ____0____32528, ____0____32529;
  wire ____0____32530, ____0____32531, ____0____32532, ____0____32533,
       ____0____32534, ____0____32535, ____0____32538, ____0____32539;
  wire ____0____32540, ____0____32541, ____0____32542, ____0____32543,
       ____0____32544, ____0____32545, ____0____32548, ____0____32549;
  wire ____0____32550, ____0____32551, ____0____32552, ____0____32553,
       ____0____32554, ____0____32555, ____0____32558, ____0____32559;
  wire ____0____32560, ____0____32561, ____0____32562, ____0____32563,
       ____0____32564, ____0____32565, ____0____33443, ____0____33444;
  wire ____0____33445, ____0____33446, ____0____33447, ____0____33448,
       ____0____33449, ____0____33450, ____0____33453, ____0____33454;
  wire ____0____33455, ____0____33456, ____0____33457, ____0____33458,
       ____0____33459, ____0____33460, ____0____33463, ____0____33464;
  wire ____0____33465, ____0____33466, ____0____33467, ____0____33468,
       ____0____33469, ____0____33472, ____0____33473, ____0____33474;
  wire ____0____33475, ____0____33476, ____0____33477, ____0____33478,
       ____0____33481, ____0____33482, ____0____33483, ____0____33484;
  wire ____0____33485, ____0____33486, ____0____33487, ____0____33488,
       ____0____33491, ____0____33492, ____0____33493, ____0____33494;
  wire ____0____33495, ____0____33496, ____0____33497, ____0____33498,
       ____0____33501, ____0____33502, ____0____33503, ____0____33504;
  wire ____0____33505, ____0____33506, ____0____33507, ____0____33508,
       ____0____33511, ____0____33512, ____0____33513, ____0____33514;
  wire ____0____33515, ____0____33516, ____0____33517, ____0____33518,
       ____0____34397, ____0____34398, ____0____34399, ____0____34400;
  wire ____0____34401, ____0____34402, ____0____34403, ____0____34404,
       ____0____34405, ____0____34406, ____0____34407, ____0____34408;
  wire ____0____34409, ____0____34410, ____0____34411, ____0____34412,
       ____0____34415, ____0____34416, ____0____34417, ____0____34418;
  wire ____0____34419, ____0____34420, ____0____34421, ____0____34422,
       ____0____34424, ____0____34425, ____0____34426, ____0____34427;
  wire ____0____34428, ____0____34429, ____0____34430, ____0____34433,
       ____0____34434, ____0____34435, ____0____34436, ____0____34437;
  wire ____0____34438, ____0____34439, ____0____34442, ____0____34443,
       ____0____34444, ____0____34445, ____0____34446, ____0____34447;
  wire ____0____34448, ____0____34449, ____0____34452, ____0____34453,
       ____0____34454, ____0____34455, ____0____34456, ____0____34457;
  wire ____0____34458, ____0____34461, ____0____34462, ____0____34463,
       ____0____34464, ____0____34465, ____0____34466, ____0____34467;
  wire ____0____34468, ____0____35299, ____0____35300, ____0____35301,
       ____0____35302, ____0____35303, ____0____35304, ____0____35307;
  wire ____0____35308, ____0____35309, ____0____35310, ____0____35311,
       ____0____35312, ____0____35313, ____0____35316, ____0____35317;
  wire ____0____35318, ____0____35319, ____0____35320, ____0____35321,
       ____0____35322, ____0____35325, ____0____35326, ____0____35327;
  wire ____0____35328, ____0____35329, ____0____35330, ____0____35331,
       ____0____35332, ____0____35335, ____0____35336, ____0____35337;
  wire ____0____35338, ____0____35339, ____0____35340, ____0____35342,
       ____0____35343, ____0____35344, ____0____35345, ____0____35346;
  wire ____0____35347, ____0____35348, ____0____35351, ____0____35352,
       ____0____35353, ____0____35354, ____0____35355, ____0____35356;
  wire ____0____35357, ____0____35358, ____0____35361, ____0____35362,
       ____0____35363, ____0____35364, ____0____35365, ____0____35366;
  wire ____0____35367, ____0____35368, ____0____36193, ____0____36194,
       ____0____36195, ____0____36196, ____0____36197, ____0____36198;
  wire ____0____36199, ____0____36202, ____0____36203, ____0____36204,
       ____0____36205, ____0____36206, ____0____36207, ____0____36210;
  wire ____0____36211, ____0____36212, ____0____36213, ____0____36214,
       ____0____36215, ____0____36216, ____0____36217, ____0____36220;
  wire ____0____36221, ____0____36222, ____0____36223, ____0____36224,
       ____0____36225, ____0____36226, ____0____36227, ____0____36230;
  wire ____0____36231, ____0____36232, ____0____36233, ____0____36234,
       ____0____36235, ____0____36236, ____0____36237, ____0____36240;
  wire ____0____36241, ____0____36242, ____0____36243, ____0____36244,
       ____0____36245, ____0____36246, ____0____36247, ____0____36250;
  wire ____0____36251, ____0____36252, ____0____36253, ____0____36254,
       ____0____36255, ____0____36256, ____0____36259, ____0____36260;
  wire ____0____36261, ____0____36262, ____0____36263, ____0____36264,
       ____0____36265, ____0____36266, ____0____37110, ____0____37111;
  wire ____0____37112, ____0____37113, ____0____37114, ____0____37115,
       ____0____37117, ____0____37118, ____0____37119, ____0____37120;
  wire ____0____37121, ____0____37122, ____0____37125, ____0____37126,
       ____0____37127, ____0____37128, ____0____37129, ____0____37130;
  wire ____0____37131, ____0____37132, ____0____37135, ____0____37136,
       ____0____37137, ____0____37138, ____0____37139, ____0____37140;
  wire ____0____37141, ____0____37142, ____0____37145, ____0____37146,
       ____0____37147, ____0____37148, ____0____37149, ____0____37150;
  wire ____0____37152, ____0____37153, ____0____37154, ____0____37155,
       ____0____37156, ____0____37157, ____0____37160, ____0____37161;
  wire ____0____37162, ____0____37163, ____0____37164, ____0____37165,
       ____0____37166, ____0____37167, ____0____37170, ____0____37171;
  wire ____0____37172, ____0____37173, ____0____37174, ____0____37175,
       ____0____37176, ____0____37177, ____0____38048, ____0____38049;
  wire ____0____38050, ____0____38051, ____0____38052, ____0____38053,
       ____0____38054, ____0____38057, ____0____38058, ____0____38059;
  wire ____0____38060, ____0____38061, ____0____38062, ____0____38065,
       ____0____38066, ____0____38067, ____0____38068, ____0____38069;
  wire ____0____38070, ____0____38071, ____0____38072, ____0____38075,
       ____0____38076, ____0____38077, ____0____38078, ____0____38079;
  wire ____0____38080, ____0____38081, ____0____38082, ____0____38085,
       ____0____38086, ____0____38087, ____0____38088, ____0____38089;
  wire ____0____38090, ____0____38091, ____0____38092, ____0____38094,
       ____0____38095, ____0____38096, ____0____38097, ____0____38098;
  wire ____0____38099, ____0____38100, ____0____38103, ____0____38104,
       ____0____38105, ____0____38106, ____0____38107, ____0____38108;
  wire ____0____38109, ____0____38110, ____0____38113, ____0____38114,
       ____0____38115, ____0____38116, ____0____38117, ____0____38118;
  wire ____0____38119, ____0____38120, ____0____40731, ____0____40732,
       ____0____40733, ____0____40734, ____0____40735, ____0____40736;
  wire ____0____40737, ____0____40738, ____0____40741, ____0____40742,
       ____0____40743, ____0____40744, ____0____40745, ____0____40746;
  wire ____0____40747, ____0____40748, ____0____40751, ____0____40752,
       ____0____40753, ____0____40754, ____0____40755, ____0____40756;
  wire ____0____40757, ____0____40758, ____0____40761, ____0____40762,
       ____0____40763, ____0____40764, ____0____40765, ____0____40766;
  wire ____0____40767, ____0____40768, ____0____40771, ____0____40772,
       ____0____40773, ____0____40774, ____0____40775, ____0____40776;
  wire ____0____40777, ____0____40778, ____0____40781, ____0____40782,
       ____0____40783, ____0____40784, ____0____40785, ____0____40786;
  wire ____0____40787, ____0____40788, ____0____40791, ____0____40792,
       ____0____40793, ____0____40794, ____0____40795, ____0____40796;
  wire ____0____40797, ____0____40798, ____0____40801, ____0____40802,
       ____0____40803, ____0____40804, ____0____40805, ____0____40806;
  wire ____0____40807, ____0____40808, ____0____________0_,
       ____0____________0___21713, ____0____________9_,
       ____0____________9___21722, ____0_____________0_,
       ____0_____________0___21723;
  wire ____0______________, ____0_______________,
       ____0________________21662, ____0________________21663,
       ____0________________21664, ____0________________21665,
       ____0________________21666, ____0________________21667;
  wire ____0________________21668, ____0________________21714,
       ____0________________21715, ____0________________21716,
       ____0________________21717, ____0________________21718,
       ____0________________21719, ____0________________21720;
  wire ____0________________21721, ____0_________________21724,
       ____0_________________21725, ____0_________________21726,
       ____0_________________21727, ____009__31512, ____009__32487,
       ____009__33441;
  wire ____009__34395, ____009__36191, ____009__37108, ____009__38047,
       ____009__40729, ____09, ____09__22458, ____09__22558;
  wire ____09__22653, ____09__22750, ____09__22848, ____09__22948,
       ____09__23048, ____09__23318, ____09__23416, ____09__23510;
  wire ____09__23606, ____09__23701, ____09__23796, ____09__23890,
       ____09__23981, ____09__24276, ____09__24372, ____09__24467;
  wire ____09__24565, ____09__24655, ____09__24848, ____09__24944,
       ____09__25230, ____09__25318, ____09__25416, ____09__25506;
  wire ____09__25595, ____09__25687, ____09__25777, ____09__25871,
       ____09__26148, ____09__26238, ____09__26331, ____09__26417;
  wire ____09__26507, ____09__26598, ____09__26691, ____09__26784,
       ____09__27038, ____09__27128, ____09__27215, ____09__27307;
  wire ____09__27400, ____09__27489, ____09__27577, ____09__27659,
       ____09__27931, ____09__28022, ____09__28117, ____09__28209;
  wire ____09__28384, ____09__28480, ____09__28561, ____09__28843,
       ____09__28931, ____09__29018, ____09__29106, ____09__29203;
  wire ____09__29287, ____09__29377, ____09__29475, ____09___31594,
       ____09___31595, ____09___31596, ____09___31597, ____09___31598;
  wire ____09___31599, ____09___31600, ____09___31601, ____09___32568,
       ____09___32569, ____09___32570, ____09___32571, ____09___32572;
  wire ____09___32573, ____09___32574, ____09___33521, ____09___33522,
       ____09___33523, ____09___33524, ____09___33525, ____09___33526;
  wire ____09___33527, ____09___33528, ____09___34471, ____09___34472,
       ____09___34473, ____09___34474, ____09___34475, ____09___34476;
  wire ____09___34477, ____09___34478, ____09___35371, ____09___35372,
       ____09___35373, ____09___35374, ____09___35375, ____09___35376;
  wire ____09___35377, ____09___36269, ____09___36270, ____09___36271,
       ____09___36272, ____09___36273, ____09___36274, ____09___36275;
  wire ____09___36276, ____09___37180, ____09___37181, ____09___37182,
       ____09___37183, ____09___37184, ____09___37185, ____09___37186;
  wire ____09___37187, ____09___38123, ____09___38124, ____09___38125,
       ____09___38126, ____09___38127, ____09___38128, ____09___38129;
  wire ____09___40811, ____09___40812, ____09___40813, ____09___40814,
       ____09___40815, ____09___40816, ____09___40817, ____09___40818;
  wire ____9, ____9_, ____9_0__32391, ____9_0__32401, ____9_0__32411,
       ____9_0__32421, ____9_0__32431, ____9_0__32441;
  wire ____9_0__32451, ____9_0__32460, ____9_0__33346, ____9_0__33356,
       ____9_0__33366, ____9_0__33376, ____9_0__33385, ____9_0__33395;
  wire ____9_0__33405, ____9_0__33415, ____9_0__34297, ____9_0__34307,
       ____9_0__34317, ____9_0__34327, ____9_0__34337, ____9_0__34347;
  wire ____9_0__34357, ____9_0__34367, ____9_0__35209, ____9_0__35217,
       ____9_0__35227, ____9_0__35234, ____9_0__35243, ____9_0__35252;
  wire ____9_0__35262, ____9_0__35270, ____9_0__36107, ____9_0__36115,
       ____9_0__36122, ____9_0__36131, ____9_0__36140, ____9_0__36149;
  wire ____9_0__36162, ____9_0__37014, ____9_0__37023, ____9_0__37033,
       ____9_0__37043, ____9_0__37053, ____9_0__37060, ____9_0__37070;
  wire ____9_0__37080, ____9_0__37958, ____9_0__37968, ____9_0__37975,
       ____9_0__37985, ____9_0__37993, ____9_0__38000, ____9_0__38009;
  wire ____9_0__38019, ____9_0__38896, ____9_0__38906, ____9_0__38916,
       ____9_0__38924, ____9_0__38941, ____9_0__38951, ____9_0__38960;
  wire ____9_9__32400, ____9_9__32410, ____9_9__32420, ____9_9__32430,
       ____9_9__32440, ____9_9__32450, ____9_9__32459, ____9_9__32469;
  wire ____9_9__33355, ____9_9__33365, ____9_9__33375, ____9_9__33384,
       ____9_9__33394, ____9_9__33404, ____9_9__33414, ____9_9__33423;
  wire ____9_9__34306, ____9_9__34316, ____9_9__34326, ____9_9__34336,
       ____9_9__34346, ____9_9__34356, ____9_9__34366, ____9_9__34376;
  wire ____9_9__35216, ____9_9__35226, ____9_9__35233, ____9_9__35242,
       ____9_9__35251, ____9_9__35261, ____9_9__35269, ____9_9__35279;
  wire ____9_9__36114, ____9_9__36121, ____9_9__36130, ____9_9__36139,
       ____9_9__36148, ____9_9__36171, ____9_9__37022, ____9_9__37032;
  wire ____9_9__37042, ____9_9__37052, ____9_9__37069, ____9_9__37079,
       ____9_9__37089, ____9_9__37967, ____9_9__37974, ____9_9__37984;
  wire ____9_9__37992, ____9_9__38008, ____9_9__38018, ____9_9__38028,
       ____9_9__38905, ____9_9__38915, ____9_9__38923, ____9_9__38931;
  wire ____9_9__38940, ____9_9__38950, ____9_9__38959, ____9_9__38968,
       ____9__22189, ____9__22214, ____9__22224, ____9__22234;
  wire ____9__22246, ____9__22261, ____9___22443, ____9___22444,
       ____9___22445, ____9___22446, ____9___22447, ____9___22448;
  wire ____9___22449, ____9___22540, ____9___22541, ____9___22542,
       ____9___22543, ____9___22544, ____9___22545, ____9___22546;
  wire ____9___22547, ____9___22635, ____9___22636, ____9___22637,
       ____9___22638, ____9___22639, ____9___22640, ____9___22641;
  wire ____9___22642, ____9___22732, ____9___22733, ____9___22734,
       ____9___22735, ____9___22736, ____9___22737, ____9___22738;
  wire ____9___22739, ____9___22830, ____9___22831, ____9___22832,
       ____9___22833, ____9___22834, ____9___22835, ____9___22836;
  wire ____9___22837, ____9___22930, ____9___22931, ____9___22932,
       ____9___22933, ____9___22934, ____9___22935, ____9___22936;
  wire ____9___22937, ____9___23030, ____9___23031, ____9___23032,
       ____9___23033, ____9___23034, ____9___23035, ____9___23036;
  wire ____9___23037, ____9___23125, ____9___23126, ____9___23127,
       ____9___23128, ____9___23129, ____9___23130, ____9___23131;
  wire ____9___23132, ____9___23398, ____9___23399, ____9___23400,
       ____9___23401, ____9___23402, ____9___23403, ____9___23404;
  wire ____9___23405, ____9___23494, ____9___23495, ____9___23496,
       ____9___23497, ____9___23498, ____9___23499, ____9___23500;
  wire ____9___23588, ____9___23589, ____9___23590, ____9___23591,
       ____9___23592, ____9___23593, ____9___23594, ____9___23595;
  wire ____9___23684, ____9___23685, ____9___23686, ____9___23687,
       ____9___23688, ____9___23689, ____9___23690, ____9___23779;
  wire ____9___23780, ____9___23781, ____9___23782, ____9___23783,
       ____9___23784, ____9___23785, ____9___23786, ____9___23873;
  wire ____9___23874, ____9___23875, ____9___23876, ____9___23877,
       ____9___23878, ____9___23879, ____9___23963, ____9___23964;
  wire ____9___23965, ____9___23966, ____9___23967, ____9___23968,
       ____9___23969, ____9___23970, ____9___24061, ____9___24062;
  wire ____9___24063, ____9___24064, ____9___24065, ____9___24066,
       ____9___24067, ____9___24068, ____9___24356, ____9___24357;
  wire ____9___24358, ____9___24359, ____9___24360, ____9___24361,
       ____9___24362, ____9___24449, ____9___24450, ____9___24451;
  wire ____9___24452, ____9___24453, ____9___24454, ____9___24455,
       ____9___24456, ____9___24547, ____9___24548, ____9___24549;
  wire ____9___24550, ____9___24551, ____9___24552, ____9___24553,
       ____9___24554, ____9___24637, ____9___24638, ____9___24639;
  wire ____9___24640, ____9___24641, ____9___24642, ____9___24643,
       ____9___24644, ____9___24737, ____9___24738, ____9___24739;
  wire ____9___24740, ____9___24741, ____9___24742, ____9___24743,
       ____9___24744, ____9___24830, ____9___24831, ____9___24832;
  wire ____9___24833, ____9___24834, ____9___24835, ____9___24836,
       ____9___24837, ____9___24926, ____9___24927, ____9___24928;
  wire ____9___24929, ____9___24930, ____9___24931, ____9___24932,
       ____9___24933, ____9___25021, ____9___25022, ____9___25023;
  wire ____9___25024, ____9___25025, ____9___25026, ____9___25027,
       ____9___25301, ____9___25302, ____9___25303, ____9___25304;
  wire ____9___25305, ____9___25306, ____9___25307, ____9___25308,
       ____9___25399, ____9___25400, ____9___25401, ____9___25402;
  wire ____9___25403, ____9___25404, ____9___25405, ____9___25490,
       ____9___25491, ____9___25492, ____9___25493, ____9___25494;
  wire ____9___25495, ____9___25577, ____9___25578, ____9___25579,
       ____9___25580, ____9___25581, ____9___25582, ____9___25583;
  wire ____9___25584, ____9___25670, ____9___25671, ____9___25672,
       ____9___25673, ____9___25674, ____9___25675, ____9___25676;
  wire ____9___25759, ____9___25760, ____9___25761, ____9___25762,
       ____9___25763, ____9___25764, ____9___25765, ____9___25766;
  wire ____9___25853, ____9___25854, ____9___25855, ____9___25856,
       ____9___25857, ____9___25858, ____9___25859, ____9___25860;
  wire ____9___25949, ____9___25950, ____9___25951, ____9___25952,
       ____9___25953, ____9___25954, ____9___25955, ____9___25956;
  wire ____9___26221, ____9___26222, ____9___26223, ____9___26224,
       ____9___26225, ____9___26226, ____9___26227, ____9___26316;
  wire ____9___26317, ____9___26318, ____9___26319, ____9___26320,
       ____9___26321, ____9___26322, ____9___26401, ____9___26402;
  wire ____9___26403, ____9___26404, ____9___26405, ____9___26406,
       ____9___26491, ____9___26492, ____9___26493, ____9___26494;
  wire ____9___26495, ____9___26496, ____9___26497, ____9___26581,
       ____9___26582, ____9___26583, ____9___26584, ____9___26585;
  wire ____9___26586, ____9___26587, ____9___26674, ____9___26675,
       ____9___26676, ____9___26677, ____9___26678, ____9___26679;
  wire ____9___26680, ____9___26681, ____9___26766, ____9___26767,
       ____9___26768, ____9___26769, ____9___26770, ____9___26771;
  wire ____9___26772, ____9___26773, ____9___26858, ____9___26859,
       ____9___26860, ____9___26861, ____9___26862, ____9___27114;
  wire ____9___27115, ____9___27116, ____9___27117, ____9___27118,
       ____9___27119, ____9___27120, ____9___27205, ____9___27206;
  wire ____9___27207, ____9___27291, ____9___27292, ____9___27293,
       ____9___27294, ____9___27295, ____9___27296, ____9___27297;
  wire ____9___27298, ____9___27383, ____9___27384, ____9___27385,
       ____9___27386, ____9___27387, ____9___27388, ____9___27389;
  wire ____9___27390, ____9___27473, ____9___27474, ____9___27475,
       ____9___27476, ____9___27477, ____9___27478, ____9___27560;
  wire ____9___27561, ____9___27562, ____9___27563, ____9___27564,
       ____9___27565, ____9___27566, ____9___27567, ____9___27648;
  wire ____9___27649, ____9___27650, ____9___27651, ____9___27652,
       ____9___27733, ____9___27734, ____9___27735, ____9___27736;
  wire ____9___27737, ____9___27738, ____9___27739, ____9___27740,
       ____9___28006, ____9___28007, ____9___28008, ____9___28009;
  wire ____9___28010, ____9___28011, ____9___28012, ____9___28102,
       ____9___28103, ____9___28104, ____9___28105, ____9___28106;
  wire ____9___28192, ____9___28193, ____9___28194, ____9___28195,
       ____9___28196, ____9___28197, ____9___28198, ____9___28286;
  wire ____9___28287, ____9___28288, ____9___28289, ____9___28290,
       ____9___28370, ____9___28371, ____9___28372, ____9___28373;
  wire ____9___28374, ____9___28375, ____9___28463, ____9___28464,
       ____9___28465, ____9___28466, ____9___28467, ____9___28468;
  wire ____9___28469, ____9___28470, ____9___28547, ____9___28548,
       ____9___28549, ____9___28550, ____9___28551, ____9___28552;
  wire ____9___28553, ____9___28638, ____9___28639, ____9___28640,
       ____9___28641, ____9___28642, ____9___28643, ____9___28644;
  wire ____9___28915, ____9___28916, ____9___28917, ____9___28918,
       ____9___28919, ____9___28920, ____9___28921, ____9___28922;
  wire ____9___29000, ____9___29001, ____9___29002, ____9___29003,
       ____9___29004, ____9___29005, ____9___29006, ____9___29007;
  wire ____9___29092, ____9___29093, ____9___29094, ____9___29095,
       ____9___29186, ____9___29187, ____9___29188, ____9___29189;
  wire ____9___29190, ____9___29191, ____9___29192, ____9___29273,
       ____9___29274, ____9___29275, ____9___29276, ____9___29277;
  wire ____9___29363, ____9___29364, ____9___29365, ____9___29366,
       ____9___29367, ____9___29457, ____9___29458, ____9___29459;
  wire ____9___29460, ____9___29461, ____9___29462, ____9___29463,
       ____9___29464, ____9___29544, ____9___29545, ____9___29546;
  wire ____9___29547, ____9___29548, ____9___29549, ____9___29550,
       ____9___29551, ____9____32392, ____9____32393, ____9____32394;
  wire ____9____32395, ____9____32396, ____9____32397, ____9____32398,
       ____9____32399, ____9____32402, ____9____32403, ____9____32404;
  wire ____9____32405, ____9____32406, ____9____32407, ____9____32408,
       ____9____32409, ____9____32412, ____9____32413, ____9____32414;
  wire ____9____32415, ____9____32416, ____9____32417, ____9____32418,
       ____9____32419, ____9____32422, ____9____32423, ____9____32424;
  wire ____9____32425, ____9____32426, ____9____32427, ____9____32428,
       ____9____32429, ____9____32432, ____9____32433, ____9____32434;
  wire ____9____32435, ____9____32436, ____9____32437, ____9____32438,
       ____9____32439, ____9____32442, ____9____32443, ____9____32444;
  wire ____9____32445, ____9____32446, ____9____32447, ____9____32448,
       ____9____32449, ____9____32452, ____9____32453, ____9____32454;
  wire ____9____32455, ____9____32456, ____9____32457, ____9____32458,
       ____9____32461, ____9____32462, ____9____32463, ____9____32464;
  wire ____9____32465, ____9____32466, ____9____32467, ____9____32468,
       ____9____33347, ____9____33348, ____9____33349, ____9____33350;
  wire ____9____33351, ____9____33352, ____9____33353, ____9____33354,
       ____9____33357, ____9____33358, ____9____33359, ____9____33360;
  wire ____9____33361, ____9____33362, ____9____33363, ____9____33364,
       ____9____33367, ____9____33368, ____9____33369, ____9____33370;
  wire ____9____33371, ____9____33372, ____9____33373, ____9____33374,
       ____9____33377, ____9____33378, ____9____33379, ____9____33380;
  wire ____9____33381, ____9____33382, ____9____33383, ____9____33386,
       ____9____33387, ____9____33388, ____9____33389, ____9____33390;
  wire ____9____33391, ____9____33392, ____9____33393, ____9____33396,
       ____9____33397, ____9____33398, ____9____33399, ____9____33400;
  wire ____9____33401, ____9____33402, ____9____33403, ____9____33406,
       ____9____33407, ____9____33408, ____9____33409, ____9____33410;
  wire ____9____33411, ____9____33412, ____9____33413, ____9____33416,
       ____9____33417, ____9____33418, ____9____33419, ____9____33420;
  wire ____9____33421, ____9____33422, ____9____34298, ____9____34299,
       ____9____34300, ____9____34301, ____9____34302, ____9____34303;
  wire ____9____34304, ____9____34305, ____9____34308, ____9____34309,
       ____9____34310, ____9____34311, ____9____34312, ____9____34313;
  wire ____9____34314, ____9____34315, ____9____34318, ____9____34319,
       ____9____34320, ____9____34321, ____9____34322, ____9____34323;
  wire ____9____34324, ____9____34325, ____9____34328, ____9____34329,
       ____9____34330, ____9____34331, ____9____34332, ____9____34333;
  wire ____9____34334, ____9____34335, ____9____34338, ____9____34339,
       ____9____34340, ____9____34341, ____9____34342, ____9____34343;
  wire ____9____34344, ____9____34345, ____9____34348, ____9____34349,
       ____9____34350, ____9____34351, ____9____34352, ____9____34353;
  wire ____9____34354, ____9____34355, ____9____34358, ____9____34359,
       ____9____34360, ____9____34361, ____9____34362, ____9____34363;
  wire ____9____34364, ____9____34365, ____9____34368, ____9____34369,
       ____9____34370, ____9____34371, ____9____34372, ____9____34373;
  wire ____9____34374, ____9____34375, ____9____35210, ____9____35211,
       ____9____35212, ____9____35213, ____9____35214, ____9____35215;
  wire ____9____35218, ____9____35219, ____9____35220, ____9____35221,
       ____9____35222, ____9____35223, ____9____35224, ____9____35225;
  wire ____9____35228, ____9____35229, ____9____35230, ____9____35231,
       ____9____35232, ____9____35235, ____9____35236, ____9____35237;
  wire ____9____35238, ____9____35239, ____9____35240, ____9____35241,
       ____9____35244, ____9____35245, ____9____35246, ____9____35247;
  wire ____9____35248, ____9____35249, ____9____35250, ____9____35253,
       ____9____35254, ____9____35255, ____9____35256, ____9____35257;
  wire ____9____35258, ____9____35259, ____9____35260, ____9____35263,
       ____9____35264, ____9____35265, ____9____35266, ____9____35267;
  wire ____9____35268, ____9____35271, ____9____35272, ____9____35273,
       ____9____35274, ____9____35275, ____9____35276, ____9____35277;
  wire ____9____35278, ____9____36108, ____9____36109, ____9____36110,
       ____9____36111, ____9____36112, ____9____36113, ____9____36116;
  wire ____9____36117, ____9____36118, ____9____36119, ____9____36120,
       ____9____36123, ____9____36124, ____9____36125, ____9____36126;
  wire ____9____36127, ____9____36128, ____9____36129, ____9____36132,
       ____9____36133, ____9____36134, ____9____36135, ____9____36136;
  wire ____9____36137, ____9____36138, ____9____36141, ____9____36142,
       ____9____36143, ____9____36144, ____9____36145, ____9____36146;
  wire ____9____36147, ____9____36150, ____9____36151, ____9____36152,
       ____9____36153, ____9____36154, ____9____36155, ____9____36156;
  wire ____9____36157, ____9____36158, ____9____36159, ____9____36160,
       ____9____36161, ____9____36163, ____9____36164, ____9____36165;
  wire ____9____36166, ____9____36167, ____9____36168, ____9____36169,
       ____9____36170, ____9____37015, ____9____37016, ____9____37017;
  wire ____9____37018, ____9____37019, ____9____37020, ____9____37021,
       ____9____37024, ____9____37025, ____9____37026, ____9____37027;
  wire ____9____37028, ____9____37029, ____9____37030, ____9____37031,
       ____9____37034, ____9____37035, ____9____37036, ____9____37037;
  wire ____9____37038, ____9____37039, ____9____37040, ____9____37041,
       ____9____37044, ____9____37045, ____9____37046, ____9____37047;
  wire ____9____37048, ____9____37049, ____9____37050, ____9____37051,
       ____9____37054, ____9____37055, ____9____37056, ____9____37057;
  wire ____9____37058, ____9____37059, ____9____37061, ____9____37062,
       ____9____37063, ____9____37064, ____9____37065, ____9____37066;
  wire ____9____37067, ____9____37068, ____9____37071, ____9____37072,
       ____9____37073, ____9____37074, ____9____37075, ____9____37076;
  wire ____9____37077, ____9____37078, ____9____37081, ____9____37082,
       ____9____37083, ____9____37084, ____9____37085, ____9____37086;
  wire ____9____37087, ____9____37088, ____9____37959, ____9____37960,
       ____9____37961, ____9____37962, ____9____37963, ____9____37964;
  wire ____9____37965, ____9____37966, ____9____37969, ____9____37970,
       ____9____37971, ____9____37972, ____9____37973, ____9____37976;
  wire ____9____37977, ____9____37978, ____9____37979, ____9____37980,
       ____9____37981, ____9____37982, ____9____37983, ____9____37986;
  wire ____9____37987, ____9____37988, ____9____37989, ____9____37990,
       ____9____37991, ____9____37994, ____9____37995, ____9____37996;
  wire ____9____37997, ____9____37998, ____9____37999, ____9____38001,
       ____9____38002, ____9____38003, ____9____38004, ____9____38005;
  wire ____9____38006, ____9____38007, ____9____38010, ____9____38011,
       ____9____38012, ____9____38013, ____9____38014, ____9____38015;
  wire ____9____38016, ____9____38017, ____9____38020, ____9____38021,
       ____9____38022, ____9____38023, ____9____38024, ____9____38025;
  wire ____9____38026, ____9____38027, ____9____38897, ____9____38898,
       ____9____38899, ____9____38900, ____9____38901, ____9____38902;
  wire ____9____38903, ____9____38904, ____9____38907, ____9____38908,
       ____9____38909, ____9____38910, ____9____38911, ____9____38912;
  wire ____9____38913, ____9____38914, ____9____38917, ____9____38918,
       ____9____38919, ____9____38920, ____9____38921, ____9____38922;
  wire ____9____38925, ____9____38926, ____9____38927, ____9____38928,
       ____9____38929, ____9____38930, ____9____38932, ____9____38933;
  wire ____9____38934, ____9____38935, ____9____38936, ____9____38937,
       ____9____38938, ____9____38939, ____9____38942, ____9____38943;
  wire ____9____38944, ____9____38945, ____9____38946, ____9____38947,
       ____9____38948, ____9____38949, ____9____38952, ____9____38953;
  wire ____9____38954, ____9____38955, ____9____38956, ____9____38957,
       ____9____38958, ____9____38961, ____9____38962, ____9____38963;
  wire ____9____38964, ____9____38965, ____9____38966, ____9____38967,
       ____090__31593, ____090__32567, ____090__33520, ____090__34470;
  wire ____090__35370, ____090__36268, ____090__37179, ____090__38122,
       ____090__40810, ____90, ____90__22539, ____90__22634;
  wire ____90__22731, ____90__22829, ____90__22929, ____90__23029,
       ____90__23124, ____90__23397, ____90__23493, ____90__23587;
  wire ____90__23683, ____90__23778, ____90__23872, ____90__23962,
       ____90__24060, ____90__24355, ____90__24448, ____90__24546;
  wire ____90__24636, ____90__24736, ____90__24829, ____90__24925,
       ____90__25020, ____90__25300, ____90__25398, ____90__25489;
  wire ____90__25576, ____90__25758, ____90__25852, ____90__25948,
       ____90__26315, ____90__26400, ____90__26490, ____90__26580;
  wire ____90__26673, ____90__26857, ____90__27113, ____90__27290,
       ____90__27382, ____90__27472, ____90__27559, ____90__27647;
  wire ____90__27732, ____90__28005, ____90__28101, ____90__28191,
       ____90__28285, ____90__28369, ____90__28462, ____90__28637;
  wire ____90__28999, ____90__29185, ____90__29272, ____90__29456,
       ____90__29543, ____90___32382, ____90___32383, ____90___32384;
  wire ____90___32385, ____90___32386, ____90___32387, ____90___32388,
       ____90___32389, ____90___33338, ____90___33339, ____90___33340;
  wire ____90___33341, ____90___33342, ____90___33343, ____90___33344,
       ____90___34288, ____90___34289, ____90___34290, ____90___34291;
  wire ____90___34292, ____90___34293, ____90___34294, ____90___34295,
       ____90___35200, ____90___35201, ____90___35202, ____90___35203;
  wire ____90___35204, ____90___35205, ____90___35206, ____90___35207,
       ____90___36098, ____90___36099, ____90___36100, ____90___36101;
  wire ____90___36102, ____90___36103, ____90___36104, ____90___36105,
       ____90___37005, ____90___37006, ____90___37007, ____90___37008;
  wire ____90___37009, ____90___37010, ____90___37011, ____90___37012,
       ____90___37950, ____90___37951, ____90___37952, ____90___37953;
  wire ____90___37954, ____90___37955, ____90___37956, ____90___38889,
       ____90___38890, ____90___38891, ____90___38892, ____90___38893;
  wire ____90___38894, ____099__31602, ____099__32575, ____099__34479,
       ____099__35378, ____099__36277, ____099__37188, ____099__38130;
  wire ____099__40819, ____99, ____99__22548, ____99__22643,
       ____99__22740, ____99__22838, ____99__22938, ____99__23038;
  wire ____99__23133, ____99__23406, ____99__23501, ____99__23596,
       ____99__23691, ____99__23787, ____99__23880, ____99__23971;
  wire ____99__24069, ____99__24363, ____99__24457, ____99__24555,
       ____99__24645, ____99__24745, ____99__24838, ____99__24934;
  wire ____99__25028, ____99__25309, ____99__25406, ____99__25496,
       ____99__25585, ____99__25677, ____99__25767, ____99__25861;
  wire ____99__25957, ____99__26228, ____99__26407, ____99__26498,
       ____99__26588, ____99__26682, ____99__26774, ____99__26863;
  wire ____99__27208, ____99__27299, ____99__27391, ____99__27479,
       ____99__27568, ____99__27653, ____99__27741, ____99__28013;
  wire ____99__28107, ____99__28199, ____99__28645, ____99__28923,
       ____99__29008, ____99__29096, ____99__29193, ____99__29278;
  wire ____99__29368, ____99__29465, ____99__29552, ____99___32471,
       ____99___32472, ____99___32473, ____99___32474, ____99___32475;
  wire ____99___32476, ____99___32477, ____99___32478, ____99___33425,
       ____99___33426, ____99___33427, ____99___33428, ____99___33429;
  wire ____99___33430, ____99___33431, ____99___34378, ____99___34379,
       ____99___34380, ____99___34381, ____99___34382, ____99___34383;
  wire ____99___34384, ____99___34385, ____99___35281, ____99___35282,
       ____99___35283, ____99___35284, ____99___35285, ____99___35286;
  wire ____99___35287, ____99___36173, ____99___36174, ____99___36175,
       ____99___36176, ____99___36177, ____99___36178, ____99___36179;
  wire ____99___36180, ____99___37091, ____99___37092, ____99___37093,
       ____99___37094, ____99___37095, ____99___37096, ____99___37097;
  wire ____99___37098, ____99___38029, ____99___38030, ____99___38031,
       ____99___38032, ____99___38033, ____99___38034, ____99___38035;
  wire ____99___38036, ____99___38970, ____99___38971, ____99___38972,
       ____99___38973, ____99___38974, ____99___38975, ____99___38976;
  wire ____900__32381, ____900__33337, ____900__34287, ____900__36097,
       ____900__37004, ____900__37949, ____900__38888, ____909__32390;
  wire ____909__33345, ____909__34296, ____909__35208, ____909__36106,
       ____909__37013, ____909__37957, ____909__38895, ____990__32470;
  wire ____990__33424, ____990__34377, ____990__35280, ____990__36172,
       ____990__37090, ____990__38969, ____999__32479, ____999__33432;
  wire ____999__34386, ____999__35288, ____999__36181, ____999__37099,
       ____999__38037, ____999__38977, _____, _____0;
  wire _____00__31603, _____00__31699, _____00__31795, _____00__31894,
       _____00__31990, _____00__32186, _____00__32283, _____00__32576;
  wire _____00__32675, _____00__32872, _____00__32970, _____00__33066,
       _____00__33159, _____00__33249, _____00__33529, _____00__33622;
  wire _____00__33717, _____00__33814, _____00__33910, _____00__34004,
       _____00__34098, _____00__34191, _____00__34480, _____00__34658;
  wire _____00__34754, _____00__34847, _____00__34931, _____00__35016,
       _____00__35103, _____00__35379, _____00__35471, _____00__35565;
  wire _____00__35653, _____00__35736, _____00__35833, _____00__35923,
       _____00__36010, _____00__36278, _____00__36544, _____00__36632;
  wire _____00__36726, _____00__36823, _____00__36914, _____00__37189,
       _____00__37276, _____00__37373, _____00__37468, _____00__37566;
  wire _____00__37663, _____00__37853, _____00__38131, _____00__38227,
       _____00__38325, _____00__38419, _____00__38517, _____00__38613;
  wire _____00__38702, _____00__38800, _____00__40820, _____00__40914,
       _____00__41012, _____00__41110, _____00__41210, _____00__41309;
  wire _____0__22375, _____0__22384, _____0__22393, _____0__22403,
       _____0__22413, _____0__22423, _____0__22433, _____0__22459;
  wire _____0__22469, _____0__22479, _____0__22489, _____0__22499,
       _____0__22509, _____0__22519, _____0__22529, _____0__22559;
  wire _____0__22568, _____0__22578, _____0__22597, _____0__22605,
       _____0__22614, _____0__22624, _____0__22654, _____0__22663;
  wire _____0__22671, _____0__22681, _____0__22691, _____0__22701,
       _____0__22711, _____0__22721, _____0__22751, _____0__22761;
  wire _____0__22771, _____0__22781, _____0__22791, _____0__22801,
       _____0__22810, _____0__22849, _____0__22859, _____0__22869;
  wire _____0__22879, _____0__22889, _____0__22899, _____0__22909,
       _____0__22919, _____0__22949, _____0__22959, _____0__22969;
  wire _____0__22979, _____0__22989, _____0__22999, _____0__23009,
       _____0__23019, _____0__23049, _____0__23058, _____0__23068;
  wire _____0__23077, _____0__23086, _____0__23095, _____0__23105,
       _____0__23114, _____0__23319, _____0__23329, _____0__23339;
  wire _____0__23349, _____0__23359, _____0__23368, _____0__23377,
       _____0__23387, _____0__23417, _____0__23426, _____0__23436;
  wire _____0__23445, _____0__23454, _____0__23464, _____0__23473,
       _____0__23483, _____0__23511, _____0__23521, _____0__23530;
  wire _____0__23540, _____0__23548, _____0__23558, _____0__23568,
       _____0__23578, _____0__23607, _____0__23617, _____0__23626;
  wire _____0__23636, _____0__23646, _____0__23656, _____0__23666,
       _____0__23674, _____0__23702, _____0__23711, _____0__23728;
  wire _____0__23738, _____0__23748, _____0__23758, _____0__23768,
       _____0__23797, _____0__23807, _____0__23816, _____0__23826;
  wire _____0__23835, _____0__23843, _____0__23852, _____0__23862,
       _____0__23891, _____0__23910, _____0__23919, _____0__23929;
  wire _____0__23939, _____0__23952, _____0__23982, _____0__23992,
       _____0__24002, _____0__24012, _____0__24022, _____0__24032;
  wire _____0__24042, _____0__24277, _____0__24287, _____0__24297,
       _____0__24307, _____0__24316, _____0__24326, _____0__24336;
  wire _____0__24345, _____0__24373, _____0__24383, _____0__24393,
       _____0__24401, _____0__24411, _____0__24420, _____0__24430;
  wire _____0__24440, _____0__24468, _____0__24478, _____0__24487,
       _____0__24497, _____0__24506, _____0__24516, _____0__24526;
  wire _____0__24536, _____0__24566, _____0__24576, _____0__24585,
       _____0__24592, _____0__24601, _____0__24610, _____0__24618;
  wire _____0__24627, _____0__24656, _____0__24666, _____0__24676,
       _____0__24686, _____0__24696, _____0__24706, _____0__24716;
  wire _____0__24726, _____0__24755, _____0__24765, _____0__24775,
       _____0__24794, _____0__24803, _____0__24812, _____0__24820;
  wire _____0__24849, _____0__24867, _____0__24876, _____0__24885,
       _____0__24895, _____0__24905, _____0__24915, _____0__24945;
  wire _____0__24955, _____0__24965, _____0__24974, _____0__24991,
       _____0__25001, _____0__25010, _____0__25231, _____0__25243;
  wire _____0__25252, _____0__25262, _____0__25271, _____0__25281,
       _____0__25291, _____0__25319, _____0__25329, _____0__25339;
  wire _____0__25349, _____0__25359, _____0__25369, _____0__25379,
       _____0__25389, _____0__25417, _____0__25425, _____0__25435;
  wire _____0__25445, _____0__25453, _____0__25461, _____0__25470,
       _____0__25479, _____0__25507, _____0__25520, _____0__25528;
  wire _____0__25538, _____0__25556, _____0__25566, _____0__25596,
       _____0__25604, _____0__25614, _____0__25623, _____0__25633;
  wire _____0__25642, _____0__25651, _____0__25660, _____0__25688,
       _____0__25695, _____0__25704, _____0__25711, _____0__25721;
  wire _____0__25729, _____0__25748, _____0__25778, _____0__25786,
       _____0__25796, _____0__25806, _____0__25815, _____0__25824;
  wire _____0__25832, _____0__25842, _____0__25872, _____0__25882,
       _____0__25892, _____0__25901, _____0__25909, _____0__25918;
  wire _____0__25928, _____0__25938, _____0__26149, _____0__26159,
       _____0__26168, _____0__26177, _____0__26186, _____0__26195;
  wire _____0__26203, _____0__26211, _____0__26247, _____0__26256,
       _____0__26266, _____0__26276, _____0__26286, _____0__26295;
  wire _____0__26305, _____0__26332, _____0__26341, _____0__26349,
       _____0__26355, _____0__26363, _____0__26371, _____0__26380;
  wire _____0__26390, _____0__26418, _____0__26428, _____0__26438,
       _____0__26448, _____0__26457, _____0__26466, _____0__26474;
  wire _____0__26482, _____0__26508, _____0__26518, _____0__26528,
       _____0__26538, _____0__26547, _____0__26555, _____0__26571;
  wire _____0__26599, _____0__26608, _____0__26617, _____0__26626,
       _____0__26636, _____0__26645, _____0__26655, _____0__26665;
  wire _____0__26692, _____0__26701, _____0__26718, _____0__26728,
       _____0__26738, _____0__26748, _____0__26758, _____0__26785;
  wire _____0__26794, _____0__26804, _____0__26822, _____0__26832,
       _____0__26839, _____0__26848, _____0__27039, _____0__27047;
  wire _____0__27057, _____0__27067, _____0__27085, _____0__27093,
       _____0__27103, _____0__27129, _____0__27139, _____0__27148;
  wire _____0__27157, _____0__27167, _____0__27177, _____0__27186,
       _____0__27196, _____0__27216, _____0__27231, _____0__27241;
  wire _____0__27251, _____0__27260, _____0__27270, _____0__27280,
       _____0__27308, _____0__27317, _____0__27327, _____0__27336;
  wire _____0__27345, _____0__27354, _____0__27363, _____0__27372,
       _____0__27401, _____0__27411, _____0__27419, _____0__27427;
  wire _____0__27435, _____0__27443, _____0__27453, _____0__27463,
       _____0__27490, _____0__27499, _____0__27507, _____0__27515;
  wire _____0__27524, _____0__27543, _____0__27552, _____0__27578,
       _____0__27585, _____0__27593, _____0__27610, _____0__27620;
  wire _____0__27637, _____0__27677, _____0__27687, _____0__27696,
       _____0__27706, _____0__27714, _____0__27723, _____0__27932;
  wire _____0__27941, _____0__27950, _____0__27958, _____0__27968,
       _____0__27978, _____0__27987, _____0__28023, _____0__28032;
  wire _____0__28042, _____0__28052, _____0__28062, _____0__28072,
       _____0__28082, _____0__28118, _____0__28128, _____0__28138;
  wire _____0__28148, _____0__28158, _____0__28168, _____0__28174,
       _____0__28181, _____0__28210, _____0__28220, _____0__28229;
  wire _____0__28238, _____0__28247, _____0__28257, _____0__28276,
       _____0__28298, _____0__28306, _____0__28314, _____0__28324;
  wire _____0__28333, _____0__28342, _____0__28351, _____0__28361,
       _____0__28385, _____0__28395, _____0__28404, _____0__28414;
  wire _____0__28424, _____0__28433, _____0__28443, _____0__28453,
       _____0__28481, _____0__28502, _____0__28511, _____0__28520;
  wire _____0__28530, _____0__28538, _____0__28562, _____0__28571,
       _____0__28581, _____0__28591, _____0__28608, _____0__28618;
  wire _____0__28627, _____0__28844, _____0__28854, _____0__28863,
       _____0__28872, _____0__28881, _____0__28890, _____0__28897;
  wire _____0__28906, _____0__28932, _____0__28941, _____0__28947,
       _____0__28966, _____0__28973, _____0__28981, _____0__28990;
  wire _____0__29028, _____0__29037, _____0__29046, _____0__29055,
       _____0__29065, _____0__29075, _____0__29083, _____0__29107;
  wire _____0__29117, _____0__29127, _____0__29136, _____0__29146,
       _____0__29155, _____0__29165, _____0__29175, _____0__29204;
  wire _____0__29213, _____0__29219, _____0__29227, _____0__29235,
       _____0__29262, _____0__29288, _____0__29296, _____0__29305;
  wire _____0__29315, _____0__29325, _____0__29335, _____0__29345,
       _____0__29353, _____0__29378, _____0__29387, _____0__29397;
  wire _____0__29407, _____0__29417, _____0__29426, _____0__29436,
       _____0__29446, _____0__29476, _____0__29486, _____0__29495;
  wire _____0__29503, _____0__29510, _____0__29527, _____0__29534,
       _____0___31604, _____0___31605, _____0___31606, _____0___31607;
  wire _____0___31608, _____0___31609, _____0___31610, _____0___31611,
       _____0___31700, _____0___31701, _____0___31702, _____0___31703;
  wire _____0___31704, _____0___31705, _____0___31706, _____0___31707,
       _____0___31796, _____0___31797, _____0___31798, _____0___31799;
  wire _____0___31800, _____0___31801, _____0___31802, _____0___31803,
       _____0___31895, _____0___31896, _____0___31897, _____0___31898;
  wire _____0___31899, _____0___31900, _____0___31901, _____0___31991,
       _____0___31992, _____0___31993, _____0___31994, _____0___31995;
  wire _____0___31996, _____0___31997, _____0___31998, _____0___32090,
       _____0___32091, _____0___32092, _____0___32093, _____0___32094;
  wire _____0___32095, _____0___32096, _____0___32187, _____0___32188,
       _____0___32189, _____0___32190, _____0___32191, _____0___32192;
  wire _____0___32193, _____0___32194, _____0___32284, _____0___32285,
       _____0___32286, _____0___32287, _____0___32288, _____0___32289;
  wire _____0___32290, _____0___32291, _____0___32577, _____0___32578,
       _____0___32579, _____0___32580, _____0___32581, _____0___32582;
  wire _____0___32583, _____0___32584, _____0___32676, _____0___32677,
       _____0___32678, _____0___32679, _____0___32680, _____0___32681;
  wire _____0___32682, _____0___32683, _____0___32774, _____0___32775,
       _____0___32776, _____0___32777, _____0___32778, _____0___32779;
  wire _____0___32780, _____0___32781, _____0___32873, _____0___32874,
       _____0___32875, _____0___32876, _____0___32877, _____0___32878;
  wire _____0___32879, _____0___32880, _____0___32971, _____0___32972,
       _____0___32973, _____0___32974, _____0___32975, _____0___32976;
  wire _____0___32977, _____0___32978, _____0___33067, _____0___33068,
       _____0___33069, _____0___33070, _____0___33071, _____0___33072;
  wire _____0___33073, _____0___33160, _____0___33161, _____0___33162,
       _____0___33163, _____0___33164, _____0___33165, _____0___33166;
  wire _____0___33250, _____0___33251, _____0___33252, _____0___33253,
       _____0___33254, _____0___33255, _____0___33256, _____0___33257;
  wire _____0___33530, _____0___33531, _____0___33532, _____0___33533,
       _____0___33534, _____0___33535, _____0___33536, _____0___33623;
  wire _____0___33624, _____0___33625, _____0___33626, _____0___33627,
       _____0___33628, _____0___33629, _____0___33718, _____0___33719;
  wire _____0___33720, _____0___33721, _____0___33722, _____0___33723,
       _____0___33724, _____0___33725, _____0___33815, _____0___33816;
  wire _____0___33817, _____0___33818, _____0___33819, _____0___33820,
       _____0___33821, _____0___33822, _____0___33911, _____0___33912;
  wire _____0___33913, _____0___33914, _____0___33915, _____0___33916,
       _____0___34005, _____0___34006, _____0___34007, _____0___34008;
  wire _____0___34009, _____0___34010, _____0___34099, _____0___34100,
       _____0___34101, _____0___34102, _____0___34103, _____0___34104;
  wire _____0___34105, _____0___34106, _____0___34192, _____0___34193,
       _____0___34194, _____0___34195, _____0___34196, _____0___34197;
  wire _____0___34198, _____0___34199, _____0___34481, _____0___34482,
       _____0___34483, _____0___34484, _____0___34485, _____0___34486;
  wire _____0___34487, _____0___34569, _____0___34570, _____0___34571,
       _____0___34572, _____0___34573, _____0___34659, _____0___34660;
  wire _____0___34661, _____0___34662, _____0___34663, _____0___34664,
       _____0___34665, _____0___34666, _____0___34755, _____0___34756;
  wire _____0___34757, _____0___34758, _____0___34759, _____0___34760,
       _____0___34761, _____0___34848, _____0___34849, _____0___34850;
  wire _____0___34851, _____0___34852, _____0___34853, _____0___34932,
       _____0___34933, _____0___34934, _____0___34935, _____0___34936;
  wire _____0___34937, _____0___34938, _____0___35017, _____0___35018,
       _____0___35019, _____0___35020, _____0___35021, _____0___35022;
  wire _____0___35104, _____0___35105, _____0___35106, _____0___35107,
       _____0___35108, _____0___35109, _____0___35110, _____0___35111;
  wire _____0___35380, _____0___35381, _____0___35382, _____0___35383,
       _____0___35384, _____0___35385, _____0___35386, _____0___35472;
  wire _____0___35473, _____0___35474, _____0___35475, _____0___35476,
       _____0___35477, _____0___35478, _____0___35479, _____0___35566;
  wire _____0___35567, _____0___35568, _____0___35569, _____0___35570,
       _____0___35571, _____0___35572, _____0___35573, _____0___35654;
  wire _____0___35655, _____0___35656, _____0___35657, _____0___35658,
       _____0___35659, _____0___35660, _____0___35737, _____0___35738;
  wire _____0___35739, _____0___35740, _____0___35741, _____0___35742,
       _____0___35743, _____0___35834, _____0___35835, _____0___35836;
  wire _____0___35837, _____0___35838, _____0___35839, _____0___35840,
       _____0___35841, _____0___35924, _____0___35925, _____0___35926;
  wire _____0___35927, _____0___35928, _____0___35929, _____0___35930,
       _____0___35931, _____0___36011, _____0___36012, _____0___36013;
  wire _____0___36014, _____0___36015, _____0___36016, _____0___36279,
       _____0___36280, _____0___36281, _____0___36282, _____0___36283;
  wire _____0___36284, _____0___36285, _____0___36367, _____0___36368,
       _____0___36369, _____0___36370, _____0___36371, _____0___36372;
  wire _____0___36373, _____0___36455, _____0___36456, _____0___36457,
       _____0___36458, _____0___36459, _____0___36460, _____0___36461;
  wire _____0___36462, _____0___36545, _____0___36546, _____0___36547,
       _____0___36548, _____0___36549, _____0___36550, _____0___36633;
  wire _____0___36634, _____0___36635, _____0___36636, _____0___36637,
       _____0___36638, _____0___36639, _____0___36640, _____0___36727;
  wire _____0___36728, _____0___36729, _____0___36730, _____0___36731,
       _____0___36732, _____0___36733, _____0___36734, _____0___36824;
  wire _____0___36825, _____0___36826, _____0___36827, _____0___36828,
       _____0___36829, _____0___36830, _____0___36831, _____0___36915;
  wire _____0___36916, _____0___36917, _____0___36918, _____0___36919,
       _____0___36920, _____0___36921, _____0___36922, _____0___37190;
  wire _____0___37191, _____0___37192, _____0___37193, _____0___37194,
       _____0___37195, _____0___37196, _____0___37277, _____0___37278;
  wire _____0___37279, _____0___37280, _____0___37281, _____0___37282,
       _____0___37283, _____0___37284, _____0___37374, _____0___37375;
  wire _____0___37376, _____0___37377, _____0___37378, _____0___37379,
       _____0___37380, _____0___37469, _____0___37470, _____0___37471;
  wire _____0___37472, _____0___37473, _____0___37474, _____0___37475,
       _____0___37476, _____0___37567, _____0___37568, _____0___37569;
  wire _____0___37570, _____0___37571, _____0___37572, _____0___37664,
       _____0___37665, _____0___37666, _____0___37667, _____0___37668;
  wire _____0___37669, _____0___37670, _____0___37671, _____0___37760,
       _____0___37761, _____0___37762, _____0___37763, _____0___37764;
  wire _____0___37854, _____0___37855, _____0___37856, _____0___37857,
       _____0___37858, _____0___37859, _____0___37860, _____0___37861;
  wire _____0___38132, _____0___38133, _____0___38134, _____0___38135,
       _____0___38136, _____0___38137, _____0___38138, _____0___38139;
  wire _____0___38228, _____0___38229, _____0___38230, _____0___38231,
       _____0___38232, _____0___38233, _____0___38234, _____0___38235;
  wire _____0___38326, _____0___38327, _____0___38328, _____0___38329,
       _____0___38330, _____0___38331, _____0___38332, _____0___38333;
  wire _____0___38420, _____0___38421, _____0___38422, _____0___38423,
       _____0___38424, _____0___38425, _____0___38426, _____0___38427;
  wire _____0___38518, _____0___38519, _____0___38520, _____0___38521,
       _____0___38522, _____0___38523, _____0___38524, _____0___38525;
  wire _____0___38614, _____0___38615, _____0___38616, _____0___38617,
       _____0___38618, _____0___38619, _____0___38620, _____0___38703;
  wire _____0___38704, _____0___38705, _____0___38706, _____0___38707,
       _____0___38708, _____0___38709, _____0___38801, _____0___38802;
  wire _____0___38803, _____0___38804, _____0___38805, _____0___38806,
       _____0___38807, _____0___38808, _____0___40821, _____0___40822;
  wire _____0___40823, _____0___40824, _____0___40825, _____0___40826,
       _____0___40827, _____0___40828, _____0___40915, _____0___40916;
  wire _____0___40917, _____0___40918, _____0___40919, _____0___40920,
       _____0___40921, _____0___40922, _____0___41013, _____0___41014;
  wire _____0___41015, _____0___41016, _____0___41017, _____0___41018,
       _____0___41019, _____0___41020, _____0___41111, _____0___41112;
  wire _____0___41113, _____0___41114, _____0___41115, _____0___41116,
       _____0___41117, _____0___41118, _____0___41211, _____0___41212;
  wire _____0___41213, _____0___41214, _____0___41215, _____0___41216,
       _____0___41217, _____0___41218, _____0___41310, _____0___41311;
  wire _____0___41312, _____0___41313, _____0___41314, _____0___41315,
       _____0___41316, _____0___41317, _____09__31612, _____09__31708;
  wire _____09__31804, _____09__31902, _____09__31999, _____09__32097,
       _____09__32195, _____09__32292, _____09__32585, _____09__32684;
  wire _____09__32782, _____09__32881, _____09__32979, _____09__33074,
       _____09__33167, _____09__33258, _____09__33537, _____09__33726;
  wire _____09__33917, _____09__34011, _____09__34107, _____09__34200,
       _____09__34488, _____09__34574, _____09__34667, _____09__34854;
  wire _____09__34939, _____09__35023, _____09__35112, _____09__35387,
       _____09__35480, _____09__35574, _____09__35744, _____09__35842;
  wire _____09__35932, _____09__36017, _____09__36286, _____09__36374,
       _____09__36641, _____09__36735, _____09__36832, _____09__36923;
  wire _____09__37197, _____09__37285, _____09__37381, _____09__37477,
       _____09__37573, _____09__37672, _____09__37765, _____09__37862;
  wire _____09__38140, _____09__38236, _____09__38526, _____09__38621,
       _____09__38710, _____09__38809, _____09__40829, _____09__40923;
  wire _____09__41021, _____09__41119, _____09__41219, _____09__41318,
       _____9, _____9__22383, _____9__22392, _____9__22402;
  wire _____9__22412, _____9__22422, _____9__22432, _____9__22442,
       _____9__22468, _____9__22478, _____9__22488, _____9__22498;
  wire _____9__22508, _____9__22518, _____9__22528, _____9__22538,
       _____9__22567, _____9__22577, _____9__22587, _____9__22596;
  wire _____9__22604, _____9__22613, _____9__22623, _____9__22633,
       _____9__22662, _____9__22680, _____9__22690, _____9__22700;
  wire _____9__22710, _____9__22720, _____9__22730, _____9__22760,
       _____9__22770, _____9__22780, _____9__22790, _____9__22800;
  wire _____9__22819, _____9__22828, _____9__22858, _____9__22868,
       _____9__22878, _____9__22888, _____9__22898, _____9__22908;
  wire _____9__22918, _____9__22928, _____9__22958, _____9__22968,
       _____9__22978, _____9__22988, _____9__22998, _____9__23008;
  wire _____9__23018, _____9__23028, _____9__23057, _____9__23067,
       _____9__23076, _____9__23094, _____9__23104, _____9__23113;
  wire _____9__23123, _____9__23328, _____9__23338, _____9__23348,
       _____9__23358, _____9__23376, _____9__23386, _____9__23396;
  wire _____9__23425, _____9__23435, _____9__23444, _____9__23453,
       _____9__23463, _____9__23472, _____9__23482, _____9__23492;
  wire _____9__23520, _____9__23529, _____9__23539, _____9__23557,
       _____9__23567, _____9__23577, _____9__23586, _____9__23616;
  wire _____9__23625, _____9__23635, _____9__23645, _____9__23655,
       _____9__23665, _____9__23673, _____9__23682, _____9__23710;
  wire _____9__23718, _____9__23727, _____9__23737, _____9__23747,
       _____9__23757, _____9__23767, _____9__23777, _____9__23806;
  wire _____9__23825, _____9__23834, _____9__23842, _____9__23851,
       _____9__23861, _____9__23871, _____9__23900, _____9__23909;
  wire _____9__23918, _____9__23928, _____9__23938, _____9__23944,
       _____9__23951, _____9__23961, _____9__23991, _____9__24001;
  wire _____9__24011, _____9__24021, _____9__24031, _____9__24041,
       _____9__24051, _____9__24059, _____9__24286, _____9__24296;
  wire _____9__24306, _____9__24315, _____9__24325, _____9__24335,
       _____9__24344, _____9__24354, _____9__24382, _____9__24392;
  wire _____9__24400, _____9__24410, _____9__24419, _____9__24429,
       _____9__24439, _____9__24447, _____9__24477, _____9__24486;
  wire _____9__24496, _____9__24505, _____9__24515, _____9__24525,
       _____9__24535, _____9__24545, _____9__24575, _____9__24584;
  wire _____9__24600, _____9__24617, _____9__24635, _____9__24665,
       _____9__24675, _____9__24685, _____9__24695, _____9__24705;
  wire _____9__24715, _____9__24725, _____9__24735, _____9__24764,
       _____9__24774, _____9__24784, _____9__24793, _____9__24802;
  wire _____9__24811, _____9__24819, _____9__24828, _____9__24857,
       _____9__24866, _____9__24894, _____9__24904, _____9__24914;
  wire _____9__24924, _____9__24954, _____9__24964, _____9__24973,
       _____9__24983, _____9__24990, _____9__25000, _____9__25009;
  wire _____9__25019, _____9__25251, _____9__25261, _____9__25280,
       _____9__25290, _____9__25328, _____9__25338, _____9__25348;
  wire _____9__25358, _____9__25368, _____9__25378, _____9__25388,
       _____9__25397, _____9__25424, _____9__25434, _____9__25444;
  wire _____9__25452, _____9__25460, _____9__25469, _____9__25478,
       _____9__25488, _____9__25519, _____9__25527, _____9__25537;
  wire _____9__25546, _____9__25555, _____9__25565, _____9__25575,
       _____9__25603, _____9__25613, _____9__25622, _____9__25632;
  wire _____9__25650, _____9__25659, _____9__25669, _____9__25703,
       _____9__25710, _____9__25720, _____9__25728, _____9__25738;
  wire _____9__25747, _____9__25757, _____9__25785, _____9__25795,
       _____9__25805, _____9__25814, _____9__25823, _____9__25841;
  wire _____9__25851, _____9__25881, _____9__25891, _____9__25900,
       _____9__25908, _____9__25917, _____9__25927, _____9__25937;
  wire _____9__25947, _____9__26158, _____9__26167, _____9__26176,
       _____9__26185, _____9__26194, _____9__26202, _____9__26210;
  wire _____9__26220, _____9__26246, _____9__26255, _____9__26265,
       _____9__26275, _____9__26285, _____9__26294, _____9__26304;
  wire _____9__26314, _____9__26340, _____9__26354, _____9__26362,
       _____9__26370, _____9__26379, _____9__26389, _____9__26399;
  wire _____9__26427, _____9__26437, _____9__26447, _____9__26456,
       _____9__26465, _____9__26473, _____9__26489, _____9__26517;
  wire _____9__26527, _____9__26537, _____9__26546, _____9__26554,
       _____9__26563, _____9__26570, _____9__26616, _____9__26625;
  wire _____9__26635, _____9__26644, _____9__26654, _____9__26664,
       _____9__26672, _____9__26700, _____9__26708, _____9__26717;
  wire _____9__26727, _____9__26737, _____9__26747, _____9__26757,
       _____9__26765, _____9__26793, _____9__26803, _____9__26812;
  wire _____9__26821, _____9__26831, _____9__26838, _____9__26847,
       _____9__26856, _____9__27046, _____9__27056, _____9__27066;
  wire _____9__27075, _____9__27084, _____9__27092, _____9__27102,
       _____9__27112, _____9__27138, _____9__27147, _____9__27166;
  wire _____9__27176, _____9__27185, _____9__27195, _____9__27204,
       _____9__27222, _____9__27240, _____9__27250, _____9__27269;
  wire _____9__27279, _____9__27289, _____9__27316, _____9__27326,
       _____9__27335, _____9__27344, _____9__27362, _____9__27371;
  wire _____9__27381, _____9__27410, _____9__27426, _____9__27434,
       _____9__27442, _____9__27452, _____9__27462, _____9__27471;
  wire _____9__27498, _____9__27506, _____9__27523, _____9__27533,
       _____9__27542, _____9__27551, _____9__27558, _____9__27601;
  wire _____9__27609, _____9__27619, _____9__27628, _____9__27636,
       _____9__27646, _____9__27667, _____9__27676, _____9__27686;
  wire _____9__27695, _____9__27705, _____9__27713, _____9__27722,
       _____9__27731, _____9__27940, _____9__27949, _____9__27957;
  wire _____9__27967, _____9__27977, _____9__27986, _____9__27996,
       _____9__28004, _____9__28031, _____9__28041, _____9__28051;
  wire _____9__28061, _____9__28071, _____9__28081, _____9__28091,
       _____9__28100, _____9__28127, _____9__28137, _____9__28147;
  wire _____9__28157, _____9__28167, _____9__28173, _____9__28180,
       _____9__28190, _____9__28219, _____9__28228, _____9__28237;
  wire _____9__28246, _____9__28256, _____9__28266, _____9__28275,
       _____9__28284, _____9__28313, _____9__28323, _____9__28332;
  wire _____9__28341, _____9__28350, _____9__28360, _____9__28368,
       _____9__28394, _____9__28403, _____9__28413, _____9__28423;
  wire _____9__28432, _____9__28442, _____9__28452, _____9__28461,
       _____9__28488, _____9__28492, _____9__28501, _____9__28510;
  wire _____9__28529, _____9__28546, _____9__28570, _____9__28580,
       _____9__28590, _____9__28598, _____9__28607, _____9__28617;
  wire _____9__28626, _____9__28636, _____9__28853, _____9__28862,
       _____9__28871, _____9__28880, _____9__28896, _____9__28905;
  wire _____9__28914, _____9__28940, _____9__28946, _____9__28956,
       _____9__28965, _____9__28972, _____9__28989, _____9__28998;
  wire _____9__29027, _____9__29036, _____9__29045, _____9__29054,
       _____9__29064, _____9__29074, _____9__29082, _____9__29091;
  wire _____9__29116, _____9__29126, _____9__29135, _____9__29145,
       _____9__29164, _____9__29174, _____9__29184, _____9__29218;
  wire _____9__29234, _____9__29244, _____9__29252, _____9__29261,
       _____9__29271, _____9__29295, _____9__29304, _____9__29314;
  wire _____9__29324, _____9__29334, _____9__29344, _____9__29352,
       _____9__29362, _____9__29386, _____9__29396, _____9__29406;
  wire _____9__29416, _____9__29425, _____9__29435, _____9__29445,
       _____9__29455, _____9__29485, _____9__29502, _____9__29509;
  wire _____9__29526, _____9__29542, _____9___22049, _____9___22050,
       _____9___22051, _____9___22052, _____9___31690, _____9___31691;
  wire _____9___31692, _____9___31693, _____9___31694, _____9___31695,
       _____9___31696, _____9___31697, _____9___31786, _____9___31787;
  wire _____9___31788, _____9___31789, _____9___31790, _____9___31791,
       _____9___31792, _____9___31793, _____9___31886, _____9___31887;
  wire _____9___31888, _____9___31889, _____9___31890, _____9___31891,
       _____9___31892, _____9___31893, _____9___31981, _____9___31982;
  wire _____9___31983, _____9___31984, _____9___31985, _____9___31986,
       _____9___31987, _____9___31988, _____9___32081, _____9___32082;
  wire _____9___32083, _____9___32084, _____9___32085, _____9___32086,
       _____9___32087, _____9___32088, _____9___32177, _____9___32178;
  wire _____9___32179, _____9___32180, _____9___32181, _____9___32182,
       _____9___32183, _____9___32184, _____9___32274, _____9___32275;
  wire _____9___32276, _____9___32277, _____9___32278, _____9___32279,
       _____9___32280, _____9___32281, _____9___32372, _____9___32373;
  wire _____9___32374, _____9___32375, _____9___32376, _____9___32377,
       _____9___32378, _____9___32379, _____9___32667, _____9___32668;
  wire _____9___32669, _____9___32670, _____9___32671, _____9___32672,
       _____9___32673, _____9___32765, _____9___32766, _____9___32767;
  wire _____9___32768, _____9___32769, _____9___32770, _____9___32771,
       _____9___32772, _____9___32863, _____9___32864, _____9___32865;
  wire _____9___32866, _____9___32867, _____9___32868, _____9___32869,
       _____9___32870, _____9___32961, _____9___32962, _____9___32963;
  wire _____9___32964, _____9___32965, _____9___32966, _____9___32967,
       _____9___32968, _____9___33057, _____9___33058, _____9___33059;
  wire _____9___33060, _____9___33061, _____9___33062, _____9___33063,
       _____9___33064, _____9___33150, _____9___33151, _____9___33152;
  wire _____9___33153, _____9___33154, _____9___33155, _____9___33156,
       _____9___33157, _____9___33242, _____9___33243, _____9___33244;
  wire _____9___33245, _____9___33246, _____9___33247, _____9___33328,
       _____9___33329, _____9___33330, _____9___33331, _____9___33332;
  wire _____9___33333, _____9___33334, _____9___33335, _____9___33613,
       _____9___33614, _____9___33615, _____9___33616, _____9___33617;
  wire _____9___33618, _____9___33619, _____9___33620, _____9___33708,
       _____9___33709, _____9___33710, _____9___33711, _____9___33712;
  wire _____9___33713, _____9___33714, _____9___33715, _____9___33806,
       _____9___33807, _____9___33808, _____9___33809, _____9___33810;
  wire _____9___33811, _____9___33812, _____9___33901, _____9___33902,
       _____9___33903, _____9___33904, _____9___33905, _____9___33906;
  wire _____9___33907, _____9___33908, _____9___33995, _____9___33996,
       _____9___33997, _____9___33998, _____9___33999, _____9___34000;
  wire _____9___34001, _____9___34002, _____9___34090, _____9___34091,
       _____9___34092, _____9___34093, _____9___34094, _____9___34095;
  wire _____9___34096, _____9___34182, _____9___34183, _____9___34184,
       _____9___34185, _____9___34186, _____9___34187, _____9___34188;
  wire _____9___34189, _____9___34278, _____9___34279, _____9___34280,
       _____9___34281, _____9___34282, _____9___34283, _____9___34284;
  wire _____9___34285, _____9___34561, _____9___34562, _____9___34563,
       _____9___34564, _____9___34565, _____9___34566, _____9___34567;
  wire _____9___34650, _____9___34651, _____9___34652, _____9___34653,
       _____9___34654, _____9___34655, _____9___34656, _____9___34745;
  wire _____9___34746, _____9___34747, _____9___34748, _____9___34749,
       _____9___34750, _____9___34751, _____9___34752, _____9___34838;
  wire _____9___34839, _____9___34840, _____9___34841, _____9___34842,
       _____9___34843, _____9___34844, _____9___34845, _____9___34923;
  wire _____9___34924, _____9___34925, _____9___34926, _____9___34927,
       _____9___34928, _____9___34929, _____9___35009, _____9___35010;
  wire _____9___35011, _____9___35012, _____9___35013, _____9___35014,
       _____9___35097, _____9___35098, _____9___35099, _____9___35100;
  wire _____9___35101, _____9___35192, _____9___35193, _____9___35194,
       _____9___35195, _____9___35196, _____9___35197, _____9___35198;
  wire _____9___35462, _____9___35463, _____9___35464, _____9___35465,
       _____9___35466, _____9___35467, _____9___35468, _____9___35469;
  wire _____9___35556, _____9___35557, _____9___35558, _____9___35559,
       _____9___35560, _____9___35561, _____9___35562, _____9___35563;
  wire _____9___35645, _____9___35646, _____9___35647, _____9___35648,
       _____9___35649, _____9___35650, _____9___35651, _____9___35730;
  wire _____9___35731, _____9___35732, _____9___35733, _____9___35734,
       _____9___35824, _____9___35825, _____9___35826, _____9___35827;
  wire _____9___35828, _____9___35829, _____9___35830, _____9___35831,
       _____9___35916, _____9___35917, _____9___35918, _____9___35919;
  wire _____9___35920, _____9___35921, _____9___36001, _____9___36002,
       _____9___36003, _____9___36004, _____9___36005, _____9___36006;
  wire _____9___36007, _____9___36008, _____9___36090, _____9___36091,
       _____9___36092, _____9___36093, _____9___36094, _____9___36095;
  wire _____9___36096, _____9___36358, _____9___36359, _____9___36360,
       _____9___36361, _____9___36362, _____9___36363, _____9___36364;
  wire _____9___36365, _____9___36448, _____9___36449, _____9___36450,
       _____9___36451, _____9___36452, _____9___36453, _____9___36536;
  wire _____9___36537, _____9___36538, _____9___36539, _____9___36540,
       _____9___36541, _____9___36542, _____9___36624, _____9___36625;
  wire _____9___36626, _____9___36627, _____9___36628, _____9___36629,
       _____9___36630, _____9___36718, _____9___36719, _____9___36720;
  wire _____9___36721, _____9___36722, _____9___36723, _____9___36724,
       _____9___36725, _____9___36814, _____9___36815, _____9___36816;
  wire _____9___36817, _____9___36818, _____9___36819, _____9___36820,
       _____9___36821, _____9___36905, _____9___36906, _____9___36907;
  wire _____9___36908, _____9___36909, _____9___36910, _____9___36911,
       _____9___36912, _____9___36996, _____9___36997, _____9___36998;
  wire _____9___36999, _____9___37000, _____9___37001, _____9___37002,
       _____9___37268, _____9___37269, _____9___37270, _____9___37271;
  wire _____9___37272, _____9___37273, _____9___37274, _____9___37364,
       _____9___37365, _____9___37366, _____9___37367, _____9___37368;
  wire _____9___37369, _____9___37370, _____9___37371, _____9___37460,
       _____9___37461, _____9___37462, _____9___37463, _____9___37464;
  wire _____9___37465, _____9___37466, _____9___37557, _____9___37558,
       _____9___37559, _____9___37560, _____9___37561, _____9___37562;
  wire _____9___37563, _____9___37564, _____9___37654, _____9___37655,
       _____9___37656, _____9___37657, _____9___37658, _____9___37659;
  wire _____9___37660, _____9___37661, _____9___37752, _____9___37753,
       _____9___37754, _____9___37755, _____9___37756, _____9___37757;
  wire _____9___37758, _____9___37844, _____9___37845, _____9___37846,
       _____9___37847, _____9___37848, _____9___37849, _____9___37850;
  wire _____9___37851, _____9___37940, _____9___37941, _____9___37942,
       _____9___37943, _____9___37944, _____9___37945, _____9___37946;
  wire _____9___37947, _____9___38219, _____9___38220, _____9___38221,
       _____9___38222, _____9___38223, _____9___38224, _____9___38225;
  wire _____9___38316, _____9___38317, _____9___38318, _____9___38319,
       _____9___38320, _____9___38321, _____9___38322, _____9___38323;
  wire _____9___38410, _____9___38411, _____9___38412, _____9___38413,
       _____9___38414, _____9___38415, _____9___38416, _____9___38417;
  wire _____9___38508, _____9___38509, _____9___38510, _____9___38511,
       _____9___38512, _____9___38513, _____9___38514, _____9___38515;
  wire _____9___38604, _____9___38605, _____9___38606, _____9___38607,
       _____9___38608, _____9___38609, _____9___38610, _____9___38611;
  wire _____9___38694, _____9___38695, _____9___38696, _____9___38697,
       _____9___38698, _____9___38699, _____9___38700, _____9___38791;
  wire _____9___38792, _____9___38793, _____9___38794, _____9___38795,
       _____9___38796, _____9___38797, _____9___38798, _____9___38881;
  wire _____9___38882, _____9___38883, _____9___38884, _____9___38885,
       _____9___38886, _____9___38887, _____9___40905, _____9___40906;
  wire _____9___40907, _____9___40908, _____9___40909, _____9___40910,
       _____9___40911, _____9___40912, _____9___41003, _____9___41004;
  wire _____9___41005, _____9___41006, _____9___41007, _____9___41008,
       _____9___41009, _____9___41010, _____9___41101, _____9___41102;
  wire _____9___41103, _____9___41104, _____9___41105, _____9___41106,
       _____9___41107, _____9___41108, _____9___41201, _____9___41202;
  wire _____9___41203, _____9___41204, _____9___41205, _____9___41206,
       _____9___41207, _____9___41208, _____9___41300, _____9___41301;
  wire _____9___41302, _____9___41303, _____9___41304, _____9___41305,
       _____9___41306, _____9___41307, _____9___41369, _____9___41370;
  wire _____90__22048, _____90__31689, _____90__31785, _____90__31885,
       _____90__31980, _____90__32080, _____90__32176, _____90__32273;
  wire _____90__32371, _____90__32666, _____90__32764, _____90__32862,
       _____90__32960, _____90__33056, _____90__33149, _____90__33241;
  wire _____90__33327, _____90__33612, _____90__33707, _____90__33805,
       _____90__33900, _____90__33994, _____90__34089, _____90__34181;
  wire _____90__34277, _____90__34560, _____90__34649, _____90__34744,
       _____90__34922, _____90__35008, _____90__35096, _____90__35191;
  wire _____90__35461, _____90__35555, _____90__35644, _____90__35823,
       _____90__35915, _____90__36000, _____90__36089, _____90__36535;
  wire _____90__36623, _____90__36717, _____90__36813, _____90__36904,
       _____90__36995, _____90__37267, _____90__37363, _____90__37459;
  wire _____90__37556, _____90__37653, _____90__37751, _____90__37843,
       _____90__37939, _____90__38218, _____90__38315, _____90__38409;
  wire _____90__38507, _____90__38603, _____90__38693, _____90__38790,
       _____90__38880, _____90__40904, _____90__41002, _____90__41100;
  wire _____90__41200, _____90__41299, _____99__22053, _____99__31698,
       _____99__31794, _____99__31989, _____99__32089, _____99__32185;
  wire _____99__32282, _____99__32380, _____99__32674, _____99__32773,
       _____99__32871, _____99__32969, _____99__33065, _____99__33158;
  wire _____99__33248, _____99__33336, _____99__33621, _____99__33716,
       _____99__33813, _____99__33909, _____99__34003, _____99__34097;
  wire _____99__34190, _____99__34286, _____99__34568, _____99__34657,
       _____99__34753, _____99__34846, _____99__34930, _____99__35015;
  wire _____99__35102, _____99__35199, _____99__35470, _____99__35564,
       _____99__35652, _____99__35735, _____99__35832, _____99__35922;
  wire _____99__36009, _____99__36366, _____99__36454, _____99__36543,
       _____99__36631, _____99__36822, _____99__36913, _____99__37003;
  wire _____99__37275, _____99__37372, _____99__37467, _____99__37565,
       _____99__37662, _____99__37759, _____99__37852, _____99__37948;
  wire _____99__38226, _____99__38324, _____99__38418, _____99__38516,
       _____99__38612, _____99__38701, _____99__38799, _____99__40913;
  wire _____99__41011, _____99__41109, _____99__41209, _____99__41308,
       _____22113, _____22114, _____22115, _____22116;
  wire _____22117, _____22118, ______, ______0_, ______0__22018,
       ______0__22027, ______0__22035, ______0__22040;
  wire ______0__31613, ______0__31623, ______0__31633, ______0__31641,
       ______0__31651, ______0__31661, ______0__31671, ______0__31680;
  wire ______0__31709, ______0__31718, ______0__31728, ______0__31737,
       ______0__31747, ______0__31756, ______0__31766, ______0__31776;
  wire ______0__31805, ______0__31815, ______0__31825, ______0__31835,
       ______0__31845, ______0__31855, ______0__31865, ______0__31875;
  wire ______0__31903, ______0__31911, ______0__31921, ______0__31931,
       ______0__31940, ______0__31950, ______0__31960, ______0__31970;
  wire ______0__32000, ______0__32010, ______0__32020, ______0__32030,
       ______0__32040, ______0__32050, ______0__32060, ______0__32070;
  wire ______0__32098, ______0__32108, ______0__32118, ______0__32127,
       ______0__32137, ______0__32147, ______0__32156, ______0__32166;
  wire ______0__32196, ______0__32205, ______0__32214, ______0__32224,
       ______0__32234, ______0__32243, ______0__32253, ______0__32263;
  wire ______0__32293, ______0__32303, ______0__32313, ______0__32321,
       ______0__32331, ______0__32341, ______0__32351, ______0__32361;
  wire ______0__32586, ______0__32596, ______0__32606, ______0__32616,
       ______0__32626, ______0__32636, ______0__32646, ______0__32656;
  wire ______0__32685, ______0__32694, ______0__32704, ______0__32714,
       ______0__32724, ______0__32734, ______0__32744, ______0__32754;
  wire ______0__32783, ______0__32793, ______0__32803, ______0__32813,
       ______0__32823, ______0__32833, ______0__32843, ______0__32853;
  wire ______0__32882, ______0__32892, ______0__32902, ______0__32912,
       ______0__32930, ______0__32940, ______0__32950, ______0__32980;
  wire ______0__32990, ______0__32999, ______0__33008, ______0__33018,
       ______0__33028, ______0__33038, ______0__33046, ______0__33075;
  wire ______0__33084, ______0__33093, ______0__33103, ______0__33122,
       ______0__33132, ______0__33141, ______0__33168, ______0__33177;
  wire ______0__33186, ______0__33195, ______0__33204, ______0__33222,
       ______0__33231, ______0__33259, ______0__33268, ______0__33277;
  wire ______0__33284, ______0__33292, ______0__33302, ______0__33312,
       ______0__33538, ______0__33548, ______0__33566, ______0__33576;
  wire ______0__33585, ______0__33595, ______0__33630, ______0__33640,
       ______0__33649, ______0__33659, ______0__33669, ______0__33679;
  wire ______0__33689, ______0__33699, ______0__33727, ______0__33736,
       ______0__33746, ______0__33756, ______0__33765, ______0__33775;
  wire ______0__33785, ______0__33795, ______0__33823, ______0__33833,
       ______0__33842, ______0__33852, ______0__33861, ______0__33871;
  wire ______0__33881, ______0__33890, ______0__33918, ______0__33928,
       ______0__33937, ______0__33946, ______0__33956, ______0__33966;
  wire ______0__33984, ______0__34012, ______0__34021, ______0__34031,
       ______0__34041, ______0__34051, ______0__34060, ______0__34069;
  wire ______0__34079, ______0__34108, ______0__34117, ______0__34125,
       ______0__34134, ______0__34153, ______0__34162, ______0__34172;
  wire ______0__34201, ______0__34210, ______0__34219, ______0__34229,
       ______0__34239, ______0__34249, ______0__34259, ______0__34267;
  wire ______0__34489, ______0__34499, ______0__34508, ______0__34517,
       ______0__34524, ______0__34534, ______0__34544, ______0__34575;
  wire ______0__34585, ______0__34594, ______0__34604, ______0__34613,
       ______0__34622, ______0__34631, ______0__34639, ______0__34668;
  wire ______0__34677, ______0__34687, ______0__34697, ______0__34715,
       ______0__34725, ______0__34734, ______0__34762, ______0__34772;
  wire ______0__34780, ______0__34790, ______0__34800, ______0__34810,
       ______0__34819, ______0__34828, ______0__34855, ______0__34871;
  wire ______0__34880, ______0__34888, ______0__34897, ______0__34905,
       ______0__34915, ______0__34940, ______0__34949, ______0__34965;
  wire ______0__34975, ______0__34982, ______0__34998, ______0__35024,
       ______0__35032, ______0__35040, ______0__35050, ______0__35059;
  wire ______0__35067, ______0__35077, ______0__35087, ______0__35113,
       ______0__35122, ______0__35132, ______0__35141, ______0__35151;
  wire ______0__35161, ______0__35171, ______0__35181, ______0__35388,
       ______0__35397, ______0__35406, ______0__35416, ______0__35426;
  wire ______0__35432, ______0__35441, ______0__35451, ______0__35481,
       ______0__35489, ______0__35499, ______0__35509, ______0__35519;
  wire ______0__35528, ______0__35537, ______0__35545, ______0__35575,
       ______0__35585, ______0__35594, ______0__35603, ______0__35612;
  wire ______0__35620, ______0__35628, ______0__35636, ______0__35684,
       ______0__35694, ______0__35701, ______0__35711, ______0__35721;
  wire ______0__35745, ______0__35755, ______0__35765, ______0__35774,
       ______0__35784, ______0__35793, ______0__35803, ______0__35813;
  wire ______0__35843, ______0__35853, ______0__35863, ______0__35871,
       ______0__35880, ______0__35889, ______0__35897, ______0__35933;
  wire ______0__35942, ______0__35948, ______0__35957, ______0__35965,
       ______0__35975, ______0__35983, ______0__35993, ______0__36018;
  wire ______0__36028, ______0__36038, ______0__36047, ______0__36056,
       ______0__36065, ______0__36081, ______0__36287, ______0__36302;
  wire ______0__36309, ______0__36319, ______0__36329, ______0__36338,
       ______0__36348, ______0__36375, ______0__36385, ______0__36394;
  wire ______0__36404, ______0__36410, ______0__36428, ______0__36438,
       ______0__36463, ______0__36473, ______0__36481, ______0__36491;
  wire ______0__36499, ______0__36508, ______0__36516, ______0__36526,
       ______0__36551, ______0__36561, ______0__36570, ______0__36580;
  wire ______0__36589, ______0__36598, ______0__36604, ______0__36614,
       ______0__36642, ______0__36651, ______0__36660, ______0__36669;
  wire ______0__36677, ______0__36687, ______0__36697, ______0__36707,
       ______0__36736, ______0__36746, ______0__36756, ______0__36766;
  wire ______0__36775, ______0__36784, ______0__36793, ______0__36803,
       ______0__36833, ______0__36842, ______0__36851, ______0__36860;
  wire ______0__36869, ______0__36879, ______0__36889, ______0__36897,
       ______0__36924, ______0__36932, ______0__36942, ______0__36951;
  wire ______0__36961, ______0__36970, ______0__36978, ______0__36985,
       ______0__37198, ______0__37205, ______0__37222, ______0__37232;
  wire ______0__37248, ______0__37257, ______0__37286, ______0__37295,
       ______0__37305, ______0__37315, ______0__37325, ______0__37335;
  wire ______0__37345, ______0__37354, ______0__37382, ______0__37391,
       ______0__37401, ______0__37411, ______0__37420, ______0__37430;
  wire ______0__37440, ______0__37450, ______0__37478, ______0__37488,
       ______0__37498, ______0__37507, ______0__37516, ______0__37526;
  wire ______0__37536, ______0__37546, ______0__37574, ______0__37584,
       ______0__37594, ______0__37604, ______0__37613, ______0__37623;
  wire ______0__37633, ______0__37643, ______0__37673, ______0__37683,
       ______0__37693, ______0__37702, ______0__37711, ______0__37721;
  wire ______0__37731, ______0__37741, ______0__37766, ______0__37776,
       ______0__37786, ______0__37796, ______0__37805, ______0__37814;
  wire ______0__37824, ______0__37833, ______0__37863, ______0__37872,
       ______0__37882, ______0__37892, ______0__37901, ______0__37910;
  wire ______0__37920, ______0__37929, ______0__38141, ______0__38151,
       ______0__38161, ______0__38170, ______0__38179, ______0__38189;
  wire ______0__38199, ______0__38209, ______0__38237, ______0__38246,
       ______0__38256, ______0__38266, ______0__38276, ______0__38286;
  wire ______0__38295, ______0__38305, ______0__38334, ______0__38343,
       ______0__38352, ______0__38362, ______0__38371, ______0__38381;
  wire ______0__38391, ______0__38401, ______0__38428, ______0__38438,
       ______0__38448, ______0__38458, ______0__38467, ______0__38477;
  wire ______0__38487, ______0__38497, ______0__38527, ______0__38537,
       ______0__38546, ______0__38555, ______0__38565, ______0__38575;
  wire ______0__38585, ______0__38594, ______0__38622, ______0__38631,
       ______0__38640, ______0__38648, ______0__38656, ______0__38664;
  wire ______0__38673, ______0__38683, ______0__38711, ______0__38721,
       ______0__38731, ______0__38740, ______0__38750, ______0__38760;
  wire ______0__38770, ______0__38780, ______0__38810, ______0__38820,
       ______0__38827, ______0__38837, ______0__38845, ______0__38855;
  wire ______0__38865, ______0__38873, ______0__40830, ______0__40840,
       ______0__40850, ______0__40860, ______0__40884, ______0__40894;
  wire ______0__40924, ______0__40934, ______0__40944, ______0__40953,
       ______0__40963, ______0__40973, ______0__40983, ______0__40992;
  wire ______0__41022, ______0__41032, ______0__41042, ______0__41052,
       ______0__41062, ______0__41072, ______0__41082, ______0__41092;
  wire ______0__41120, ______0__41130, ______0__41140, ______0__41150,
       ______0__41160, ______0__41170, ______0__41180, ______0__41190;
  wire ______0__41220, ______0__41230, ______0__41240, ______0__41250,
       ______0__41260, ______0__41270, ______0__41279, ______0__41289;
  wire ______0__41319, ______0__41329, ______0__41339, ______0__41349,
       ______0__41359, ______0__41366, ______0___22054, ______0___22055;
  wire ______0___22056, ______0___22057, ______0___22058, ______09,
       ______9__22017, ______9__22026, ______9__22030, ______9__22034;
  wire ______9__31622, ______9__31632, ______9__31640, ______9__31650,
       ______9__31660, ______9__31670, ______9__31679, ______9__31688;
  wire ______9__31717, ______9__31727, ______9__31736, ______9__31746,
       ______9__31755, ______9__31765, ______9__31775, ______9__31814;
  wire ______9__31824, ______9__31834, ______9__31844, ______9__31854,
       ______9__31864, ______9__31874, ______9__31884, ______9__31910;
  wire ______9__31920, ______9__31930, ______9__31939, ______9__31949,
       ______9__31959, ______9__31969, ______9__31979, ______9__32009;
  wire ______9__32019, ______9__32029, ______9__32039, ______9__32049,
       ______9__32059, ______9__32069, ______9__32079, ______9__32107;
  wire ______9__32117, ______9__32126, ______9__32136, ______9__32146,
       ______9__32155, ______9__32165, ______9__32175, ______9__32204;
  wire ______9__32213, ______9__32223, ______9__32233, ______9__32242,
       ______9__32252, ______9__32262, ______9__32272, ______9__32302;
  wire ______9__32312, ______9__32320, ______9__32330, ______9__32340,
       ______9__32350, ______9__32360, ______9__32370, ______9__32595;
  wire ______9__32605, ______9__32615, ______9__32625, ______9__32635,
       ______9__32645, ______9__32655, ______9__32665, ______9__32693;
  wire ______9__32703, ______9__32713, ______9__32723, ______9__32733,
       ______9__32743, ______9__32753, ______9__32763, ______9__32792;
  wire ______9__32802, ______9__32812, ______9__32822, ______9__32832,
       ______9__32842, ______9__32852, ______9__32861, ______9__32891;
  wire ______9__32901, ______9__32911, ______9__32921, ______9__32929,
       ______9__32939, ______9__32949, ______9__32959, ______9__32989;
  wire ______9__32998, ______9__33007, ______9__33017, ______9__33027,
       ______9__33037, ______9__33045, ______9__33055, ______9__33083;
  wire ______9__33092, ______9__33102, ______9__33112, ______9__33121,
       ______9__33131, ______9__33140, ______9__33148, ______9__33176;
  wire ______9__33185, ______9__33194, ______9__33203, ______9__33213,
       ______9__33221, ______9__33230, ______9__33240, ______9__33267;
  wire ______9__33276, ______9__33283, ______9__33301, ______9__33311,
       ______9__33326, ______9__33547, ______9__33556, ______9__33565;
  wire ______9__33575, ______9__33584, ______9__33594, ______9__33604,
       ______9__33639, ______9__33648, ______9__33658, ______9__33668;
  wire ______9__33678, ______9__33688, ______9__33698, ______9__33706,
       ______9__33735, ______9__33745, ______9__33755, ______9__33764;
  wire ______9__33774, ______9__33784, ______9__33794, ______9__33804,
       ______9__33832, ______9__33841, ______9__33851, ______9__33860;
  wire ______9__33870, ______9__33880, ______9__33889, ______9__33899,
       ______9__33927, ______9__33936, ______9__33945, ______9__33955;
  wire ______9__33965, ______9__33975, ______9__33983, ______9__33993,
       ______9__34020, ______9__34030, ______9__34040, ______9__34050;
  wire ______9__34059, ______9__34068, ______9__34078, ______9__34088,
       ______9__34116, ______9__34124, ______9__34133, ______9__34143;
  wire ______9__34152, ______9__34161, ______9__34171, ______9__34180,
       ______9__34209, ______9__34218, ______9__34228, ______9__34238;
  wire ______9__34248, ______9__34258, ______9__34266, ______9__34276,
       ______9__34498, ______9__34507, ______9__34516, ______9__34523;
  wire ______9__34533, ______9__34543, ______9__34553, ______9__34584,
       ______9__34593, ______9__34603, ______9__34612, ______9__34621;
  wire ______9__34630, ______9__34638, ______9__34648, ______9__34676,
       ______9__34686, ______9__34696, ______9__34705, ______9__34714;
  wire ______9__34724, ______9__34743, ______9__34771, ______9__34779,
       ______9__34789, ______9__34799, ______9__34809, ______9__34818;
  wire ______9__34827, ______9__34837, ______9__34863, ______9__34870,
       ______9__34887, ______9__34896, ______9__34904, ______9__34914;
  wire ______9__34948, ______9__34964, ______9__34974, ______9__34981,
       ______9__34997, ______9__35007, ______9__35039, ______9__35049;
  wire ______9__35066, ______9__35076, ______9__35086, ______9__35095,
       ______9__35121, ______9__35131, ______9__35140, ______9__35150;
  wire ______9__35160, ______9__35170, ______9__35180, ______9__35190,
       ______9__35396, ______9__35405, ______9__35415, ______9__35425;
  wire ______9__35431, ______9__35440, ______9__35450, ______9__35460,
       ______9__35498, ______9__35508, ______9__35518, ______9__35527;
  wire ______9__35536, ______9__35544, ______9__35554, ______9__35584,
       ______9__35593, ______9__35602, ______9__35619, ______9__35627;
  wire ______9__35643, ______9__35667, ______9__35675, ______9__35683,
       ______9__35693, ______9__35710, ______9__35720, ______9__35754;
  wire ______9__35764, ______9__35773, ______9__35783, ______9__35792,
       ______9__35802, ______9__35812, ______9__35822, ______9__35852;
  wire ______9__35862, ______9__35870, ______9__35879, ______9__35888,
       ______9__35896, ______9__35906, ______9__35941, ______9__35947;
  wire ______9__35956, ______9__35964, ______9__35974, ______9__35982,
       ______9__35992, ______9__35999, ______9__36027, ______9__36037;
  wire ______9__36055, ______9__36064, ______9__36072, ______9__36080,
       ______9__36088, ______9__36295, ______9__36308, ______9__36318;
  wire ______9__36328, ______9__36337, ______9__36347, ______9__36357,
       ______9__36384, ______9__36403, ______9__36419, ______9__36427;
  wire ______9__36437, ______9__36447, ______9__36472, ______9__36490,
       ______9__36498, ______9__36507, ______9__36515, ______9__36525;
  wire ______9__36534, ______9__36560, ______9__36569, ______9__36579,
       ______9__36588, ______9__36597, ______9__36603, ______9__36613;
  wire ______9__36622, ______9__36659, ______9__36668, ______9__36676,
       ______9__36686, ______9__36696, ______9__36706, ______9__36716;
  wire ______9__36745, ______9__36755, ______9__36765, ______9__36774,
       ______9__36783, ______9__36792, ______9__36802, ______9__36812;
  wire ______9__36841, ______9__36850, ______9__36859, ______9__36868,
       ______9__36878, ______9__36888, ______9__36896, ______9__36903;
  wire ______9__36931, ______9__36941, ______9__36950, ______9__36960,
       ______9__36969, ______9__36977, ______9__36984, ______9__36994;
  wire ______9__37214, ______9__37231, ______9__37240, ______9__37247,
       ______9__37256, ______9__37266, ______9__37294, ______9__37304;
  wire ______9__37314, ______9__37324, ______9__37334, ______9__37344,
       ______9__37353, ______9__37362, ______9__37390, ______9__37400;
  wire ______9__37410, ______9__37419, ______9__37429, ______9__37439,
       ______9__37449, ______9__37458, ______9__37487, ______9__37497;
  wire ______9__37506, ______9__37515, ______9__37525, ______9__37535,
       ______9__37545, ______9__37555, ______9__37583, ______9__37593;
  wire ______9__37603, ______9__37622, ______9__37632, ______9__37642,
       ______9__37652, ______9__37682, ______9__37692, ______9__37701;
  wire ______9__37710, ______9__37720, ______9__37730, ______9__37740,
       ______9__37750, ______9__37775, ______9__37785, ______9__37795;
  wire ______9__37804, ______9__37813, ______9__37823, ______9__37832,
       ______9__37842, ______9__37871, ______9__37881, ______9__37891;
  wire ______9__37900, ______9__37909, ______9__37919, ______9__37928,
       ______9__37938, ______9__38150, ______9__38160, ______9__38169;
  wire ______9__38188, ______9__38198, ______9__38208, ______9__38217,
       ______9__38245, ______9__38255, ______9__38265, ______9__38275;
  wire ______9__38285, ______9__38294, ______9__38304, ______9__38314,
       ______9__38342, ______9__38351, ______9__38361, ______9__38370;
  wire ______9__38380, ______9__38390, ______9__38400, ______9__38408,
       ______9__38437, ______9__38447, ______9__38457, ______9__38466;
  wire ______9__38476, ______9__38486, ______9__38496, ______9__38506,
       ______9__38536, ______9__38545, ______9__38554, ______9__38564;
  wire ______9__38574, ______9__38584, ______9__38593, ______9__38602,
       ______9__38630, ______9__38639, ______9__38647, ______9__38655;
  wire ______9__38672, ______9__38682, ______9__38692, ______9__38720,
       ______9__38730, ______9__38739, ______9__38749, ______9__38759;
  wire ______9__38769, ______9__38779, ______9__38789, ______9__38819,
       ______9__38826, ______9__38836, ______9__38844, ______9__38854;
  wire ______9__38864, ______9__38879, ______9__40839, ______9__40849,
       ______9__40859, ______9__40883, ______9__40893, ______9__40903;
  wire ______9__40933, ______9__40943, ______9__40952, ______9__40962,
       ______9__40972, ______9__40982, ______9__40991, ______9__41001;
  wire ______9__41031, ______9__41041, ______9__41051, ______9__41061,
       ______9__41071, ______9__41081, ______9__41091, ______9__41099;
  wire ______9__41129, ______9__41139, ______9__41149, ______9__41159,
       ______9__41169, ______9__41179, ______9__41189, ______9__41199;
  wire ______9__41229, ______9__41239, ______9__41249, ______9__41259,
       ______9__41269, ______9__41278, ______9__41288, ______9__41298;
  wire ______9__41328, ______9__41338, ______9__41348, ______9__41358,
       ______22119, ______22120, ______22121, ______22122;
  wire ______22123, ______22124, ______22125, ______22126, ______22127,
       ______22128, ______22129, ______22130;
  wire ______22131, ______22132, ______22135, ______22136, ______22138,
       ______22139, ______22140, ______22141;
  wire ______22142, ______22144, ______22145, ______22146, ______22147,
       ______22148, ______22150, ______22151;
  wire ______22152, ______22153, ______22154, ______22155, ______22158,
       ______22159, ______22160, ______22161;
  wire ______22162, ______22163, ______22164, _______22172,
       _______22173, _______22174, _______22175, _______22176;
  wire _______22177, _______22178, _______22179, _______22180,
       _______22181, _______22182, _______22183, _______22184;
  wire _______22185, _______22186, _______22187, _______22188,
       _______22206, _______22207, _______22208, _______22209;
  wire _______22210, _______22211, _______22212, _______22213,
       _______22216, _______22217, _______22218, _______22219;
  wire _______22220, _______22221, _______22222, _______22223,
       _______22226, _______22227, _______22228, _______22229;
  wire _______22230, _______22231, _______22232, _______22233,
       _______22236, _______22237, _______22238, _______22239;
  wire _______22240, _______22241, _______22242, _______22243,
       _______22244, _______22245, _______22248, _______22249;
  wire _______22250, _______22251, _______22252, _______22253,
       _______22254, _______22255, _______22256, _______22257;
  wire _______22258, _______22259, _______22260, _______22277,
       _______22278, _______22279, _______22280, _______22282;
  wire _______22283, _______22284, _______22285, _______22286,
       ________, ________22013, ________22368, ________22369;
  wire ________22370, ________22371, ________22372, ________22373,
       ________22374, ________22376, ________22377, ________22378;
  wire ________22379, ________22380, ________22381, ________22382,
       ________22385, ________22386, ________22387, ________22388;
  wire ________22389, ________22390, ________22391, ________22394,
       ________22395, ________22396, ________22397, ________22398;
  wire ________22399, ________22400, ________22401, ________22404,
       ________22405, ________22406, ________22407, ________22408;
  wire ________22409, ________22410, ________22411, ________22414,
       ________22415, ________22416, ________22417, ________22418;
  wire ________22419, ________22420, ________22421, ________22424,
       ________22425, ________22426, ________22427, ________22428;
  wire ________22429, ________22430, ________22431, ________22434,
       ________22435, ________22436, ________22437, ________22438;
  wire ________22439, ________22440, ________22441, ________22460,
       ________22461, ________22462, ________22463, ________22464;
  wire ________22465, ________22466, ________22467, ________22470,
       ________22471, ________22472, ________22473, ________22474;
  wire ________22475, ________22476, ________22477, ________22480,
       ________22481, ________22482, ________22483, ________22484;
  wire ________22485, ________22486, ________22487, ________22490,
       ________22491, ________22492, ________22493, ________22494;
  wire ________22495, ________22496, ________22497, ________22500,
       ________22501, ________22502, ________22503, ________22504;
  wire ________22505, ________22506, ________22507, ________22510,
       ________22511, ________22512, ________22513, ________22514;
  wire ________22515, ________22516, ________22517, ________22520,
       ________22521, ________22522, ________22523, ________22524;
  wire ________22525, ________22526, ________22527, ________22530,
       ________22531, ________22532, ________22533, ________22534;
  wire ________22535, ________22536, ________22537, ________22560,
       ________22561, ________22562, ________22563, ________22564;
  wire ________22565, ________22566, ________22569, ________22570,
       ________22571, ________22572, ________22573, ________22574;
  wire ________22575, ________22576, ________22579, ________22580,
       ________22581, ________22582, ________22583, ________22584;
  wire ________22585, ________22586, ________22588, ________22589,
       ________22590, ________22591, ________22592, ________22593;
  wire ________22594, ________22595, ________22598, ________22599,
       ________22600, ________22601, ________22602, ________22603;
  wire ________22606, ________22607, ________22608, ________22609,
       ________22610, ________22611, ________22612, ________22615;
  wire ________22616, ________22617, ________22618, ________22619,
       ________22620, ________22621, ________22622, ________22625;
  wire ________22626, ________22627, ________22628, ________22629,
       ________22630, ________22631, ________22632, ________22655;
  wire ________22656, ________22657, ________22658, ________22659,
       ________22660, ________22661, ________22664, ________22665;
  wire ________22666, ________22667, ________22668, ________22669,
       ________22670, ________22672, ________22673, ________22674;
  wire ________22675, ________22676, ________22677, ________22678,
       ________22679, ________22682, ________22683, ________22684;
  wire ________22685, ________22686, ________22687, ________22688,
       ________22689, ________22692, ________22693, ________22694;
  wire ________22695, ________22696, ________22697, ________22698,
       ________22699, ________22702, ________22703, ________22704;
  wire ________22705, ________22706, ________22707, ________22708,
       ________22709, ________22712, ________22713, ________22714;
  wire ________22715, ________22716, ________22717, ________22718,
       ________22719, ________22722, ________22723, ________22724;
  wire ________22725, ________22726, ________22727, ________22728,
       ________22729, ________22752, ________22753, ________22754;
  wire ________22755, ________22756, ________22757, ________22758,
       ________22759, ________22762, ________22763, ________22764;
  wire ________22765, ________22766, ________22767, ________22768,
       ________22769, ________22772, ________22773, ________22774;
  wire ________22775, ________22776, ________22777, ________22778,
       ________22779, ________22782, ________22783, ________22784;
  wire ________22785, ________22786, ________22787, ________22788,
       ________22789, ________22792, ________22793, ________22794;
  wire ________22795, ________22796, ________22797, ________22798,
       ________22799, ________22802, ________22803, ________22804;
  wire ________22805, ________22806, ________22807, ________22808,
       ________22809, ________22811, ________22812, ________22813;
  wire ________22814, ________22815, ________22816, ________22817,
       ________22818, ________22820, ________22821, ________22822;
  wire ________22823, ________22824, ________22825, ________22826,
       ________22827, ________22850, ________22851, ________22852;
  wire ________22853, ________22854, ________22855, ________22856,
       ________22857, ________22860, ________22861, ________22862;
  wire ________22863, ________22864, ________22865, ________22866,
       ________22867, ________22870, ________22871, ________22872;
  wire ________22873, ________22874, ________22875, ________22876,
       ________22877, ________22880, ________22881, ________22882;
  wire ________22883, ________22884, ________22885, ________22886,
       ________22887, ________22890, ________22891, ________22892;
  wire ________22893, ________22894, ________22895, ________22896,
       ________22897, ________22900, ________22901, ________22902;
  wire ________22903, ________22904, ________22905, ________22906,
       ________22907, ________22910, ________22911, ________22912;
  wire ________22913, ________22914, ________22915, ________22916,
       ________22917, ________22920, ________22921, ________22922;
  wire ________22923, ________22924, ________22925, ________22926,
       ________22927, ________22950, ________22951, ________22952;
  wire ________22953, ________22954, ________22955, ________22956,
       ________22957, ________22960, ________22961, ________22962;
  wire ________22963, ________22964, ________22965, ________22966,
       ________22967, ________22970, ________22971, ________22972;
  wire ________22973, ________22974, ________22975, ________22976,
       ________22977, ________22980, ________22981, ________22982;
  wire ________22983, ________22984, ________22985, ________22986,
       ________22987, ________22990, ________22991, ________22992;
  wire ________22993, ________22994, ________22995, ________22996,
       ________22997, ________23000, ________23001, ________23002;
  wire ________23003, ________23004, ________23005, ________23006,
       ________23007, ________23010, ________23011, ________23012;
  wire ________23013, ________23014, ________23015, ________23016,
       ________23017, ________23020, ________23021, ________23022;
  wire ________23023, ________23024, ________23025, ________23026,
       ________23027, ________23050, ________23051, ________23052;
  wire ________23053, ________23054, ________23055, ________23056,
       ________23059, ________23060, ________23061, ________23062;
  wire ________23063, ________23064, ________23065, ________23066,
       ________23069, ________23070, ________23071, ________23072;
  wire ________23073, ________23074, ________23075, ________23078,
       ________23079, ________23080, ________23081, ________23082;
  wire ________23083, ________23084, ________23085, ________23087,
       ________23088, ________23089, ________23090, ________23091;
  wire ________23092, ________23093, ________23096, ________23097,
       ________23098, ________23099, ________23100, ________23101;
  wire ________23102, ________23103, ________23106, ________23107,
       ________23108, ________23109, ________23110, ________23111;
  wire ________23112, ________23115, ________23116, ________23117,
       ________23118, ________23119, ________23120, ________23121;
  wire ________23122, ________23320, ________23321, ________23322,
       ________23323, ________23324, ________23325, ________23326;
  wire ________23327, ________23330, ________23331, ________23332,
       ________23333, ________23334, ________23335, ________23336;
  wire ________23337, ________23340, ________23341, ________23342,
       ________23343, ________23344, ________23345, ________23346;
  wire ________23347, ________23350, ________23351, ________23352,
       ________23353, ________23354, ________23355, ________23356;
  wire ________23357, ________23360, ________23361, ________23362,
       ________23363, ________23364, ________23365, ________23366;
  wire ________23367, ________23369, ________23370, ________23371,
       ________23372, ________23373, ________23374, ________23375;
  wire ________23378, ________23379, ________23380, ________23381,
       ________23382, ________23383, ________23384, ________23385;
  wire ________23388, ________23389, ________23390, ________23391,
       ________23392, ________23393, ________23394, ________23395;
  wire ________23418, ________23419, ________23420, ________23421,
       ________23422, ________23423, ________23424, ________23427;
  wire ________23428, ________23429, ________23430, ________23431,
       ________23432, ________23433, ________23434, ________23437;
  wire ________23438, ________23439, ________23440, ________23441,
       ________23442, ________23443, ________23446, ________23447;
  wire ________23448, ________23449, ________23450, ________23451,
       ________23452, ________23455, ________23456, ________23457;
  wire ________23458, ________23459, ________23460, ________23461,
       ________23462, ________23465, ________23466, ________23467;
  wire ________23468, ________23469, ________23470, ________23471,
       ________23474, ________23475, ________23476, ________23477;
  wire ________23478, ________23479, ________23480, ________23481,
       ________23484, ________23485, ________23486, ________23487;
  wire ________23488, ________23489, ________23490, ________23491,
       ________23512, ________23513, ________23514, ________23515;
  wire ________23516, ________23517, ________23518, ________23519,
       ________23522, ________23523, ________23524, ________23525;
  wire ________23526, ________23527, ________23528, ________23531,
       ________23532, ________23533, ________23534, ________23535;
  wire ________23536, ________23537, ________23538, ________23541,
       ________23542, ________23543, ________23544, ________23545;
  wire ________23546, ________23547, ________23549, ________23550,
       ________23551, ________23552, ________23553, ________23554;
  wire ________23555, ________23556, ________23559, ________23560,
       ________23561, ________23562, ________23563, ________23564;
  wire ________23565, ________23566, ________23569, ________23570,
       ________23571, ________23572, ________23573, ________23574;
  wire ________23575, ________23576, ________23579, ________23580,
       ________23581, ________23582, ________23583, ________23584;
  wire ________23585, ________23608, ________23609, ________23610,
       ________23611, ________23612, ________23613, ________23614;
  wire ________23615, ________23618, ________23619, ________23620,
       ________23621, ________23622, ________23623, ________23624;
  wire ________23627, ________23628, ________23629, ________23630,
       ________23631, ________23632, ________23633, ________23634;
  wire ________23637, ________23638, ________23639, ________23640,
       ________23641, ________23642, ________23643, ________23644;
  wire ________23647, ________23648, ________23649, ________23650,
       ________23651, ________23652, ________23653, ________23654;
  wire ________23657, ________23658, ________23659, ________23660,
       ________23661, ________23662, ________23663, ________23664;
  wire ________23667, ________23668, ________23669, ________23670,
       ________23671, ________23672, ________23675, ________23676;
  wire ________23677, ________23678, ________23679, ________23680,
       ________23681, ________23703, ________23704, ________23705;
  wire ________23706, ________23707, ________23708, ________23709,
       ________23712, ________23713, ________23714, ________23715;
  wire ________23716, ________23717, ________23719, ________23720,
       ________23721, ________23722, ________23723, ________23724;
  wire ________23725, ________23726, ________23729, ________23730,
       ________23731, ________23732, ________23733, ________23734;
  wire ________23735, ________23736, ________23739, ________23740,
       ________23741, ________23742, ________23743, ________23744;
  wire ________23745, ________23746, ________23749, ________23750,
       ________23751, ________23752, ________23753, ________23754;
  wire ________23755, ________23756, ________23759, ________23760,
       ________23761, ________23762, ________23763, ________23764;
  wire ________23765, ________23766, ________23769, ________23770,
       ________23771, ________23772, ________23773, ________23774;
  wire ________23775, ________23776, ________23798, ________23799,
       ________23800, ________23801, ________23802, ________23803;
  wire ________23804, ________23805, ________23808, ________23809,
       ________23810, ________23811, ________23812, ________23813;
  wire ________23814, ________23815, ________23817, ________23818,
       ________23819, ________23820, ________23821, ________23822;
  wire ________23823, ________23824, ________23827, ________23828,
       ________23829, ________23830, ________23831, ________23832;
  wire ________23833, ________23836, ________23837, ________23838,
       ________23839, ________23840, ________23841, ________23844;
  wire ________23845, ________23846, ________23847, ________23848,
       ________23849, ________23850, ________23853, ________23854;
  wire ________23855, ________23856, ________23857, ________23858,
       ________23859, ________23860, ________23863, ________23864;
  wire ________23865, ________23866, ________23867, ________23868,
       ________23869, ________23870, ________23892, ________23893;
  wire ________23894, ________23895, ________23896, ________23897,
       ________23898, ________23899, ________23901, ________23902;
  wire ________23903, ________23904, ________23905, ________23906,
       ________23907, ________23908, ________23911, ________23912;
  wire ________23913, ________23914, ________23915, ________23916,
       ________23917, ________23920, ________23921, ________23922;
  wire ________23923, ________23924, ________23925, ________23926,
       ________23927, ________23930, ________23931, ________23932;
  wire ________23933, ________23934, ________23935, ________23936,
       ________23937, ________23940, ________23941, ________23942;
  wire ________23943, ________23945, ________23946, ________23947,
       ________23948, ________23949, ________23950, ________23953;
  wire ________23954, ________23955, ________23956, ________23957,
       ________23958, ________23959, ________23960, ________23983;
  wire ________23984, ________23985, ________23986, ________23987,
       ________23988, ________23989, ________23990, ________23993;
  wire ________23994, ________23995, ________23996, ________23997,
       ________23998, ________23999, ________24000, ________24003;
  wire ________24004, ________24005, ________24006, ________24007,
       ________24008, ________24009, ________24010, ________24013;
  wire ________24014, ________24015, ________24016, ________24017,
       ________24018, ________24019, ________24020, ________24023;
  wire ________24024, ________24025, ________24026, ________24027,
       ________24028, ________24029, ________24030, ________24033;
  wire ________24034, ________24035, ________24036, ________24037,
       ________24038, ________24039, ________24040, ________24043;
  wire ________24044, ________24045, ________24046, ________24047,
       ________24048, ________24049, ________24050, ________24052;
  wire ________24053, ________24054, ________24055, ________24056,
       ________24057, ________24058, ________24278, ________24279;
  wire ________24280, ________24281, ________24282, ________24283,
       ________24284, ________24285, ________24288, ________24289;
  wire ________24290, ________24291, ________24292, ________24293,
       ________24294, ________24295, ________24298, ________24299;
  wire ________24300, ________24301, ________24302, ________24303,
       ________24304, ________24305, ________24308, ________24309;
  wire ________24310, ________24311, ________24312, ________24313,
       ________24314, ________24317, ________24318, ________24319;
  wire ________24320, ________24321, ________24322, ________24323,
       ________24324, ________24327, ________24328, ________24329;
  wire ________24330, ________24331, ________24332, ________24333,
       ________24334, ________24337, ________24338, ________24339;
  wire ________24340, ________24341, ________24342, ________24343,
       ________24346, ________24347, ________24348, ________24349;
  wire ________24350, ________24351, ________24352, ________24353,
       ________24374, ________24375, ________24376, ________24377;
  wire ________24378, ________24379, ________24380, ________24381,
       ________24384, ________24385, ________24386, ________24387;
  wire ________24388, ________24389, ________24390, ________24391,
       ________24394, ________24395, ________24396, ________24397;
  wire ________24398, ________24399, ________24402, ________24403,
       ________24404, ________24405, ________24406, ________24407;
  wire ________24408, ________24409, ________24412, ________24413,
       ________24414, ________24415, ________24416, ________24417;
  wire ________24418, ________24421, ________24422, ________24423,
       ________24424, ________24425, ________24426, ________24427;
  wire ________24428, ________24431, ________24432, ________24433,
       ________24434, ________24435, ________24436, ________24437;
  wire ________24438, ________24441, ________24442, ________24443,
       ________24444, ________24445, ________24446, ________24469;
  wire ________24470, ________24471, ________24472, ________24473,
       ________24474, ________24475, ________24476, ________24479;
  wire ________24480, ________24481, ________24482, ________24483,
       ________24484, ________24485, ________24488, ________24489;
  wire ________24490, ________24491, ________24492, ________24493,
       ________24494, ________24495, ________24498, ________24499;
  wire ________24500, ________24501, ________24502, ________24503,
       ________24504, ________24507, ________24508, ________24509;
  wire ________24510, ________24511, ________24512, ________24513,
       ________24514, ________24517, ________24518, ________24519;
  wire ________24520, ________24521, ________24522, ________24523,
       ________24524, ________24527, ________24528, ________24529;
  wire ________24530, ________24531, ________24532, ________24533,
       ________24534, ________24537, ________24538, ________24539;
  wire ________24540, ________24541, ________24542, ________24543,
       ________24544, ________24567, ________24568, ________24569;
  wire ________24570, ________24571, ________24572, ________24573,
       ________24574, ________24577, ________24578, ________24579;
  wire ________24580, ________24581, ________24582, ________24583,
       ________24586, ________24587, ________24588, ________24589;
  wire ________24590, ________24591, ________24593, ________24594,
       ________24595, ________24596, ________24597, ________24598;
  wire ________24599, ________24602, ________24603, ________24604,
       ________24605, ________24606, ________24607, ________24608;
  wire ________24609, ________24611, ________24612, ________24613,
       ________24614, ________24615, ________24616, ________24619;
  wire ________24620, ________24621, ________24622, ________24623,
       ________24624, ________24625, ________24626, ________24628;
  wire ________24629, ________24630, ________24631, ________24632,
       ________24633, ________24634, ________24657, ________24658;
  wire ________24659, ________24660, ________24661, ________24662,
       ________24663, ________24664, ________24667, ________24668;
  wire ________24669, ________24670, ________24671, ________24672,
       ________24673, ________24674, ________24677, ________24678;
  wire ________24679, ________24680, ________24681, ________24682,
       ________24683, ________24684, ________24687, ________24688;
  wire ________24689, ________24690, ________24691, ________24692,
       ________24693, ________24694, ________24697, ________24698;
  wire ________24699, ________24700, ________24701, ________24702,
       ________24703, ________24704, ________24707, ________24708;
  wire ________24709, ________24710, ________24711, ________24712,
       ________24713, ________24714, ________24717, ________24718;
  wire ________24719, ________24720, ________24721, ________24722,
       ________24723, ________24724, ________24727, ________24728;
  wire ________24729, ________24730, ________24731, ________24732,
       ________24733, ________24734, ________24756, ________24757;
  wire ________24758, ________24759, ________24760, ________24761,
       ________24762, ________24763, ________24766, ________24767;
  wire ________24768, ________24769, ________24770, ________24771,
       ________24772, ________24773, ________24776, ________24777;
  wire ________24778, ________24779, ________24780, ________24781,
       ________24782, ________24783, ________24785, ________24786;
  wire ________24787, ________24788, ________24789, ________24790,
       ________24791, ________24792, ________24795, ________24796;
  wire ________24797, ________24798, ________24799, ________24800,
       ________24801, ________24804, ________24805, ________24806;
  wire ________24807, ________24808, ________24809, ________24810,
       ________24813, ________24814, ________24815, ________24816;
  wire ________24817, ________24818, ________24821, ________24822,
       ________24823, ________24824, ________24825, ________24826;
  wire ________24827, ________24850, ________24851, ________24852,
       ________24853, ________24854, ________24855, ________24856;
  wire ________24858, ________24859, ________24860, ________24861,
       ________24862, ________24863, ________24864, ________24865;
  wire ________24868, ________24869, ________24870, ________24871,
       ________24872, ________24873, ________24874, ________24875;
  wire ________24877, ________24878, ________24879, ________24880,
       ________24881, ________24882, ________24883, ________24884;
  wire ________24886, ________24887, ________24888, ________24889,
       ________24890, ________24891, ________24892, ________24893;
  wire ________24896, ________24897, ________24898, ________24899,
       ________24900, ________24901, ________24902, ________24903;
  wire ________24906, ________24907, ________24908, ________24909,
       ________24910, ________24911, ________24912, ________24913;
  wire ________24916, ________24917, ________24918, ________24919,
       ________24920, ________24921, ________24922, ________24923;
  wire ________24946, ________24947, ________24948, ________24949,
       ________24950, ________24951, ________24952, ________24953;
  wire ________24956, ________24957, ________24958, ________24959,
       ________24960, ________24961, ________24962, ________24963;
  wire ________24966, ________24967, ________24968, ________24969,
       ________24970, ________24971, ________24972, ________24975;
  wire ________24976, ________24977, ________24978, ________24979,
       ________24980, ________24981, ________24982, ________24984;
  wire ________24985, ________24986, ________24987, ________24988,
       ________24989, ________24992, ________24993, ________24994;
  wire ________24995, ________24996, ________24997, ________24998,
       ________24999, ________25002, ________25003, ________25004;
  wire ________25005, ________25006, ________25007, ________25008,
       ________25011, ________25012, ________25013, ________25014;
  wire ________25015, ________25016, ________25017, ________25018,
       ________25232, ________25233, ________25234, ________25235;
  wire ________25236, ________25237, ________25238, ________25239,
       ________25240, ________25241, ________25242, ________25244;
  wire ________25245, ________25246, ________25247, ________25248,
       ________25249, ________25250, ________25253, ________25254;
  wire ________25255, ________25256, ________25257, ________25258,
       ________25259, ________25260, ________25263, ________25264;
  wire ________25265, ________25266, ________25267, ________25268,
       ________25269, ________25270, ________25272, ________25273;
  wire ________25274, ________25275, ________25276, ________25277,
       ________25278, ________25279, ________25282, ________25283;
  wire ________25284, ________25285, ________25286, ________25287,
       ________25288, ________25289, ________25292, ________25293;
  wire ________25294, ________25295, ________25296, ________25297,
       ________25298, ________25299, ________25320, ________25321;
  wire ________25322, ________25323, ________25324, ________25325,
       ________25326, ________25327, ________25330, ________25331;
  wire ________25332, ________25333, ________25334, ________25335,
       ________25336, ________25337, ________25340, ________25341;
  wire ________25342, ________25343, ________25344, ________25345,
       ________25346, ________25347, ________25350, ________25351;
  wire ________25352, ________25353, ________25354, ________25355,
       ________25356, ________25357, ________25360, ________25361;
  wire ________25362, ________25363, ________25364, ________25365,
       ________25366, ________25367, ________25370, ________25371;
  wire ________25372, ________25373, ________25374, ________25375,
       ________25376, ________25377, ________25380, ________25381;
  wire ________25382, ________25383, ________25384, ________25385,
       ________25386, ________25387, ________25390, ________25391;
  wire ________25392, ________25393, ________25394, ________25395,
       ________25396, ________25418, ________25419, ________25420;
  wire ________25421, ________25422, ________25423, ________25426,
       ________25427, ________25428, ________25429, ________25430;
  wire ________25431, ________25432, ________25433, ________25436,
       ________25437, ________25438, ________25439, ________25440;
  wire ________25441, ________25442, ________25443, ________25446,
       ________25447, ________25448, ________25449, ________25450;
  wire ________25451, ________25454, ________25455, ________25456,
       ________25457, ________25458, ________25459, ________25462;
  wire ________25463, ________25464, ________25465, ________25466,
       ________25467, ________25468, ________25471, ________25472;
  wire ________25473, ________25474, ________25475, ________25476,
       ________25477, ________25480, ________25481, ________25482;
  wire ________25483, ________25484, ________25485, ________25486,
       ________25487, ________25508, ________25509, ________25510;
  wire ________25511, ________25512, ________25513, ________25514,
       ________25515, ________25516, ________25517, ________25518;
  wire ________25521, ________25522, ________25523, ________25524,
       ________25525, ________25526, ________25529, ________25530;
  wire ________25531, ________25532, ________25533, ________25534,
       ________25535, ________25536, ________25539, ________25540;
  wire ________25541, ________25542, ________25543, ________25544,
       ________25545, ________25547, ________25548, ________25549;
  wire ________25550, ________25551, ________25552, ________25553,
       ________25554, ________25557, ________25558, ________25559;
  wire ________25560, ________25561, ________25562, ________25563,
       ________25564, ________25567, ________25568, ________25569;
  wire ________25570, ________25571, ________25572, ________25573,
       ________25574, ________25597, ________25598, ________25599;
  wire ________25600, ________25601, ________25602, ________25605,
       ________25606, ________25607, ________25608, ________25609;
  wire ________25610, ________25611, ________25612, ________25615,
       ________25616, ________25617, ________25618, ________25619;
  wire ________25620, ________25621, ________25624, ________25625,
       ________25626, ________25627, ________25628, ________25629;
  wire ________25630, ________25631, ________25634, ________25635,
       ________25636, ________25637, ________25638, ________25639;
  wire ________25640, ________25641, ________25643, ________25644,
       ________25645, ________25646, ________25647, ________25648;
  wire ________25649, ________25652, ________25653, ________25654,
       ________25655, ________25656, ________25657, ________25658;
  wire ________25661, ________25662, ________25663, ________25664,
       ________25665, ________25666, ________25667, ________25668;
  wire ________25689, ________25690, ________25691, ________25692,
       ________25693, ________25694, ________25696, ________25697;
  wire ________25698, ________25699, ________25700, ________25701,
       ________25702, ________25705, ________25706, ________25707;
  wire ________25708, ________25709, ________25712, ________25713,
       ________25714, ________25715, ________25716, ________25717;
  wire ________25718, ________25719, ________25722, ________25723,
       ________25724, ________25725, ________25726, ________25727;
  wire ________25730, ________25731, ________25732, ________25733,
       ________25734, ________25735, ________25736, ________25737;
  wire ________25739, ________25740, ________25741, ________25742,
       ________25743, ________25744, ________25745, ________25746;
  wire ________25749, ________25750, ________25751, ________25752,
       ________25753, ________25754, ________25755, ________25756;
  wire ________25779, ________25780, ________25781, ________25782,
       ________25783, ________25784, ________25787, ________25788;
  wire ________25789, ________25790, ________25791, ________25792,
       ________25793, ________25794, ________25797, ________25798;
  wire ________25799, ________25800, ________25801, ________25802,
       ________25803, ________25804, ________25807, ________25808;
  wire ________25809, ________25810, ________25811, ________25812,
       ________25813, ________25816, ________25817, ________25818;
  wire ________25819, ________25820, ________25821, ________25822,
       ________25825, ________25826, ________25827, ________25828;
  wire ________25829, ________25830, ________25831, ________25833,
       ________25834, ________25835, ________25836, ________25837;
  wire ________25838, ________25839, ________25840, ________25843,
       ________25844, ________25845, ________25846, ________25847;
  wire ________25848, ________25849, ________25850, ________25873,
       ________25874, ________25875, ________25876, ________25877;
  wire ________25878, ________25879, ________25880, ________25883,
       ________25884, ________25885, ________25886, ________25887;
  wire ________25888, ________25889, ________25890, ________25893,
       ________25894, ________25895, ________25896, ________25897;
  wire ________25898, ________25899, ________25902, ________25903,
       ________25904, ________25905, ________25906, ________25907;
  wire ________25910, ________25911, ________25912, ________25913,
       ________25914, ________25915, ________25916, ________25919;
  wire ________25920, ________25921, ________25922, ________25923,
       ________25924, ________25925, ________25926, ________25929;
  wire ________25930, ________25931, ________25932, ________25933,
       ________25934, ________25935, ________25936, ________25939;
  wire ________25940, ________25941, ________25942, ________25943,
       ________25944, ________25945, ________25946, ________26150;
  wire ________26151, ________26152, ________26153, ________26154,
       ________26155, ________26156, ________26157, ________26160;
  wire ________26161, ________26162, ________26163, ________26164,
       ________26165, ________26166, ________26169, ________26170;
  wire ________26171, ________26172, ________26173, ________26174,
       ________26175, ________26178, ________26179, ________26180;
  wire ________26181, ________26182, ________26183, ________26184,
       ________26187, ________26188, ________26189, ________26190;
  wire ________26191, ________26192, ________26193, ________26196,
       ________26197, ________26198, ________26199, ________26200;
  wire ________26201, ________26204, ________26205, ________26206,
       ________26207, ________26208, ________26209, ________26212;
  wire ________26213, ________26214, ________26215, ________26216,
       ________26217, ________26218, ________26219, ________26239;
  wire ________26240, ________26241, ________26242, ________26243,
       ________26244, ________26245, ________26248, ________26249;
  wire ________26250, ________26251, ________26252, ________26253,
       ________26254, ________26257, ________26258, ________26259;
  wire ________26260, ________26261, ________26262, ________26263,
       ________26264, ________26267, ________26268, ________26269;
  wire ________26270, ________26271, ________26272, ________26273,
       ________26274, ________26277, ________26278, ________26279;
  wire ________26280, ________26281, ________26282, ________26283,
       ________26284, ________26287, ________26288, ________26289;
  wire ________26290, ________26291, ________26292, ________26293,
       ________26296, ________26297, ________26298, ________26299;
  wire ________26300, ________26301, ________26302, ________26303,
       ________26306, ________26307, ________26308, ________26309;
  wire ________26310, ________26311, ________26312, ________26313,
       ________26333, ________26334, ________26335, ________26336;
  wire ________26337, ________26338, ________26339, ________26342,
       ________26343, ________26344, ________26345, ________26346;
  wire ________26347, ________26348, ________26350, ________26351,
       ________26352, ________26353, ________26356, ________26357;
  wire ________26358, ________26359, ________26360, ________26361,
       ________26364, ________26365, ________26366, ________26367;
  wire ________26368, ________26369, ________26372, ________26373,
       ________26374, ________26375, ________26376, ________26377;
  wire ________26378, ________26381, ________26382, ________26383,
       ________26384, ________26385, ________26386, ________26387;
  wire ________26388, ________26391, ________26392, ________26393,
       ________26394, ________26395, ________26396, ________26397;
  wire ________26398, ________26419, ________26420, ________26421,
       ________26422, ________26423, ________26424, ________26425;
  wire ________26426, ________26429, ________26430, ________26431,
       ________26432, ________26433, ________26434, ________26435;
  wire ________26436, ________26439, ________26440, ________26441,
       ________26442, ________26443, ________26444, ________26445;
  wire ________26446, ________26449, ________26450, ________26451,
       ________26452, ________26453, ________26454, ________26455;
  wire ________26458, ________26459, ________26460, ________26461,
       ________26462, ________26463, ________26464, ________26467;
  wire ________26468, ________26469, ________26470, ________26471,
       ________26472, ________26475, ________26476, ________26477;
  wire ________26478, ________26479, ________26480, ________26481,
       ________26483, ________26484, ________26485, ________26486;
  wire ________26487, ________26488, ________26509, ________26510,
       ________26511, ________26512, ________26513, ________26514;
  wire ________26515, ________26516, ________26519, ________26520,
       ________26521, ________26522, ________26523, ________26524;
  wire ________26525, ________26526, ________26529, ________26530,
       ________26531, ________26532, ________26533, ________26534;
  wire ________26535, ________26536, ________26539, ________26540,
       ________26541, ________26542, ________26543, ________26544;
  wire ________26545, ________26548, ________26549, ________26550,
       ________26551, ________26552, ________26553, ________26556;
  wire ________26557, ________26558, ________26559, ________26560,
       ________26561, ________26562, ________26564, ________26565;
  wire ________26566, ________26567, ________26568, ________26569,
       ________26572, ________26573, ________26574, ________26575;
  wire ________26576, ________26577, ________26578, ________26579,
       ________26600, ________26601, ________26602, ________26603;
  wire ________26604, ________26605, ________26606, ________26607,
       ________26609, ________26610, ________26611, ________26612;
  wire ________26613, ________26614, ________26615, ________26618,
       ________26619, ________26620, ________26621, ________26622;
  wire ________26623, ________26624, ________26627, ________26628,
       ________26629, ________26630, ________26631, ________26632;
  wire ________26633, ________26634, ________26637, ________26638,
       ________26639, ________26640, ________26641, ________26642;
  wire ________26643, ________26646, ________26647, ________26648,
       ________26649, ________26650, ________26651, ________26652;
  wire ________26653, ________26656, ________26657, ________26658,
       ________26659, ________26660, ________26661, ________26662;
  wire ________26663, ________26666, ________26667, ________26668,
       ________26669, ________26670, ________26671, ________26693;
  wire ________26694, ________26695, ________26696, ________26697,
       ________26698, ________26699, ________26702, ________26703;
  wire ________26704, ________26705, ________26706, ________26707,
       ________26709, ________26710, ________26711, ________26712;
  wire ________26713, ________26714, ________26715, ________26716,
       ________26719, ________26720, ________26721, ________26722;
  wire ________26723, ________26724, ________26725, ________26726,
       ________26729, ________26730, ________26731, ________26732;
  wire ________26733, ________26734, ________26735, ________26736,
       ________26739, ________26740, ________26741, ________26742;
  wire ________26743, ________26744, ________26745, ________26746,
       ________26749, ________26750, ________26751, ________26752;
  wire ________26753, ________26754, ________26755, ________26756,
       ________26759, ________26760, ________26761, ________26762;
  wire ________26763, ________26764, ________26786, ________26787,
       ________26788, ________26789, ________26790, ________26791;
  wire ________26792, ________26795, ________26796, ________26797,
       ________26798, ________26799, ________26800, ________26801;
  wire ________26802, ________26805, ________26806, ________26807,
       ________26808, ________26809, ________26810, ________26811;
  wire ________26813, ________26814, ________26815, ________26816,
       ________26817, ________26818, ________26819, ________26820;
  wire ________26823, ________26824, ________26825, ________26826,
       ________26827, ________26828, ________26829, ________26830;
  wire ________26833, ________26834, ________26835, ________26836,
       ________26837, ________26840, ________26841, ________26842;
  wire ________26843, ________26844, ________26845, ________26846,
       ________26849, ________26850, ________26851, ________26852;
  wire ________26853, ________26854, ________26855, ________27040,
       ________27041, ________27042, ________27043, ________27044;
  wire ________27045, ________27048, ________27049, ________27050,
       ________27051, ________27052, ________27053, ________27054;
  wire ________27055, ________27058, ________27059, ________27060,
       ________27061, ________27062, ________27063, ________27064;
  wire ________27065, ________27068, ________27069, ________27070,
       ________27071, ________27072, ________27073, ________27074;
  wire ________27076, ________27077, ________27078, ________27079,
       ________27080, ________27081, ________27082, ________27083;
  wire ________27086, ________27087, ________27088, ________27089,
       ________27090, ________27091, ________27094, ________27095;
  wire ________27096, ________27097, ________27098, ________27099,
       ________27100, ________27101, ________27104, ________27105;
  wire ________27106, ________27107, ________27108, ________27109,
       ________27110, ________27111, ________27130, ________27131;
  wire ________27132, ________27133, ________27134, ________27135,
       ________27136, ________27137, ________27140, ________27141;
  wire ________27142, ________27143, ________27144, ________27145,
       ________27146, ________27149, ________27150, ________27151;
  wire ________27152, ________27153, ________27154, ________27155,
       ________27156, ________27158, ________27159, ________27160;
  wire ________27161, ________27162, ________27163, ________27164,
       ________27165, ________27168, ________27169, ________27170;
  wire ________27171, ________27172, ________27173, ________27174,
       ________27175, ________27178, ________27179, ________27180;
  wire ________27181, ________27182, ________27183, ________27184,
       ________27187, ________27188, ________27189, ________27190;
  wire ________27191, ________27192, ________27193, ________27194,
       ________27197, ________27198, ________27199, ________27200;
  wire ________27201, ________27202, ________27203, ________27217,
       ________27218, ________27219, ________27220, ________27221;
  wire ________27223, ________27224, ________27225, ________27226,
       ________27227, ________27228, ________27229, ________27230;
  wire ________27232, ________27233, ________27234, ________27235,
       ________27236, ________27237, ________27238, ________27239;
  wire ________27242, ________27243, ________27244, ________27245,
       ________27246, ________27247, ________27248, ________27249;
  wire ________27252, ________27253, ________27254, ________27255,
       ________27256, ________27257, ________27258, ________27259;
  wire ________27261, ________27262, ________27263, ________27264,
       ________27265, ________27266, ________27267, ________27268;
  wire ________27271, ________27272, ________27273, ________27274,
       ________27275, ________27276, ________27277, ________27278;
  wire ________27281, ________27282, ________27283, ________27284,
       ________27285, ________27286, ________27287, ________27288;
  wire ________27309, ________27310, ________27311, ________27312,
       ________27313, ________27314, ________27315, ________27318;
  wire ________27319, ________27320, ________27321, ________27322,
       ________27323, ________27324, ________27325, ________27328;
  wire ________27329, ________27330, ________27331, ________27332,
       ________27333, ________27334, ________27337, ________27338;
  wire ________27339, ________27340, ________27341, ________27342,
       ________27343, ________27346, ________27347, ________27348;
  wire ________27349, ________27350, ________27351, ________27352,
       ________27353, ________27355, ________27356, ________27357;
  wire ________27358, ________27359, ________27360, ________27361,
       ________27364, ________27365, ________27366, ________27367;
  wire ________27368, ________27369, ________27370, ________27373,
       ________27374, ________27375, ________27376, ________27377;
  wire ________27378, ________27379, ________27380, ________27402,
       ________27403, ________27404, ________27405, ________27406;
  wire ________27407, ________27408, ________27409, ________27412,
       ________27413, ________27414, ________27415, ________27416;
  wire ________27417, ________27418, ________27420, ________27421,
       ________27422, ________27423, ________27424, ________27425;
  wire ________27428, ________27429, ________27430, ________27431,
       ________27432, ________27433, ________27436, ________27437;
  wire ________27438, ________27439, ________27440, ________27441,
       ________27444, ________27445, ________27446, ________27447;
  wire ________27448, ________27449, ________27450, ________27451,
       ________27454, ________27455, ________27456, ________27457;
  wire ________27458, ________27459, ________27460, ________27461,
       ________27464, ________27465, ________27466, ________27467;
  wire ________27468, ________27469, ________27470, ________27491,
       ________27492, ________27493, ________27494, ________27495;
  wire ________27496, ________27497, ________27500, ________27501,
       ________27502, ________27503, ________27504, ________27505;
  wire ________27508, ________27509, ________27510, ________27511,
       ________27512, ________27513, ________27514, ________27516;
  wire ________27517, ________27518, ________27519, ________27520,
       ________27521, ________27522, ________27525, ________27526;
  wire ________27527, ________27528, ________27529, ________27530,
       ________27531, ________27532, ________27534, ________27535;
  wire ________27536, ________27537, ________27538, ________27539,
       ________27540, ________27541, ________27544, ________27545;
  wire ________27546, ________27547, ________27548, ________27549,
       ________27550, ________27553, ________27554, ________27555;
  wire ________27556, ________27557, ________27579, ________27580,
       ________27581, ________27582, ________27583, ________27584;
  wire ________27586, ________27587, ________27588, ________27589,
       ________27590, ________27591, ________27592, ________27594;
  wire ________27595, ________27596, ________27597, ________27598,
       ________27599, ________27600, ________27602, ________27603;
  wire ________27604, ________27605, ________27606, ________27607,
       ________27608, ________27611, ________27612, ________27613;
  wire ________27614, ________27615, ________27616, ________27617,
       ________27618, ________27621, ________27622, ________27623;
  wire ________27624, ________27625, ________27626, ________27627,
       ________27629, ________27630, ________27631, ________27632;
  wire ________27633, ________27634, ________27635, ________27638,
       ________27639, ________27640, ________27641, ________27642;
  wire ________27643, ________27644, ________27645, ________27660,
       ________27661, ________27662, ________27663, ________27664;
  wire ________27665, ________27666, ________27668, ________27669,
       ________27670, ________27671, ________27672, ________27673;
  wire ________27674, ________27675, ________27678, ________27679,
       ________27680, ________27681, ________27682, ________27683;
  wire ________27684, ________27685, ________27688, ________27689,
       ________27690, ________27691, ________27692, ________27693;
  wire ________27694, ________27697, ________27698, ________27699,
       ________27700, ________27701, ________27702, ________27703;
  wire ________27704, ________27707, ________27708, ________27709,
       ________27710, ________27711, ________27712, ________27715;
  wire ________27716, ________27717, ________27718, ________27719,
       ________27720, ________27721, ________27724, ________27725;
  wire ________27726, ________27727, ________27728, ________27729,
       ________27730, ________27933, ________27934, ________27935;
  wire ________27936, ________27937, ________27938, ________27939,
       ________27942, ________27943, ________27944, ________27945;
  wire ________27946, ________27947, ________27948, ________27951,
       ________27952, ________27953, ________27954, ________27955;
  wire ________27956, ________27959, ________27960, ________27961,
       ________27962, ________27963, ________27964, ________27965;
  wire ________27966, ________27969, ________27970, ________27971,
       ________27972, ________27973, ________27974, ________27975;
  wire ________27976, ________27979, ________27980, ________27981,
       ________27982, ________27983, ________27984, ________27985;
  wire ________27988, ________27989, ________27990, ________27991,
       ________27992, ________27993, ________27994, ________27995;
  wire ________27997, ________27998, ________27999, ________28000,
       ________28001, ________28002, ________28003, ________28024;
  wire ________28025, ________28026, ________28027, ________28028,
       ________28029, ________28030, ________28033, ________28034;
  wire ________28035, ________28036, ________28037, ________28038,
       ________28039, ________28040, ________28043, ________28044;
  wire ________28045, ________28046, ________28047, ________28048,
       ________28049, ________28050, ________28053, ________28054;
  wire ________28055, ________28056, ________28057, ________28058,
       ________28059, ________28060, ________28063, ________28064;
  wire ________28065, ________28066, ________28067, ________28068,
       ________28069, ________28070, ________28073, ________28074;
  wire ________28075, ________28076, ________28077, ________28078,
       ________28079, ________28080, ________28083, ________28084;
  wire ________28085, ________28086, ________28087, ________28088,
       ________28089, ________28090, ________28092, ________28093;
  wire ________28094, ________28095, ________28096, ________28097,
       ________28098, ________28099, ________28119, ________28120;
  wire ________28121, ________28122, ________28123, ________28124,
       ________28125, ________28126, ________28129, ________28130;
  wire ________28131, ________28132, ________28133, ________28134,
       ________28135, ________28136, ________28139, ________28140;
  wire ________28141, ________28142, ________28143, ________28144,
       ________28145, ________28146, ________28149, ________28150;
  wire ________28151, ________28152, ________28153, ________28154,
       ________28155, ________28156, ________28159, ________28160;
  wire ________28161, ________28162, ________28163, ________28164,
       ________28165, ________28166, ________28169, ________28170;
  wire ________28171, ________28172, ________28175, ________28176,
       ________28177, ________28178, ________28179, ________28182;
  wire ________28183, ________28184, ________28185, ________28186,
       ________28187, ________28188, ________28189, ________28211;
  wire ________28212, ________28213, ________28214, ________28215,
       ________28216, ________28217, ________28218, ________28221;
  wire ________28222, ________28223, ________28224, ________28225,
       ________28226, ________28227, ________28230, ________28231;
  wire ________28232, ________28233, ________28234, ________28235,
       ________28236, ________28239, ________28240, ________28241;
  wire ________28242, ________28243, ________28244, ________28245,
       ________28248, ________28249, ________28250, ________28251;
  wire ________28252, ________28253, ________28254, ________28255,
       ________28258, ________28259, ________28260, ________28261;
  wire ________28262, ________28263, ________28264, ________28265,
       ________28267, ________28268, ________28269, ________28270;
  wire ________28271, ________28272, ________28273, ________28274,
       ________28277, ________28278, ________28279, ________28280;
  wire ________28281, ________28282, ________28283, ________28299,
       ________28300, ________28301, ________28302, ________28303;
  wire ________28304, ________28305, ________28307, ________28308,
       ________28309, ________28310, ________28311, ________28312;
  wire ________28315, ________28316, ________28317, ________28318,
       ________28319, ________28320, ________28321, ________28322;
  wire ________28325, ________28326, ________28327, ________28328,
       ________28329, ________28330, ________28331, ________28334;
  wire ________28335, ________28336, ________28337, ________28338,
       ________28339, ________28340, ________28343, ________28344;
  wire ________28345, ________28346, ________28347, ________28348,
       ________28349, ________28352, ________28353, ________28354;
  wire ________28355, ________28356, ________28357, ________28358,
       ________28359, ________28362, ________28363, ________28364;
  wire ________28365, ________28366, ________28367, ________28386,
       ________28387, ________28388, ________28389, ________28390;
  wire ________28391, ________28392, ________28393, ________28396,
       ________28397, ________28398, ________28399, ________28400;
  wire ________28401, ________28402, ________28405, ________28406,
       ________28407, ________28408, ________28409, ________28410;
  wire ________28411, ________28412, ________28415, ________28416,
       ________28417, ________28418, ________28419, ________28420;
  wire ________28421, ________28422, ________28425, ________28426,
       ________28427, ________28428, ________28429, ________28430;
  wire ________28431, ________28434, ________28435, ________28436,
       ________28437, ________28438, ________28439, ________28440;
  wire ________28441, ________28444, ________28445, ________28446,
       ________28447, ________28448, ________28449, ________28450;
  wire ________28451, ________28454, ________28455, ________28456,
       ________28457, ________28458, ________28459, ________28460;
  wire ________28482, ________28483, ________28484, ________28485,
       ________28486, ________28487, ________28489, ________28490;
  wire ________28491, ________28493, ________28494, ________28495,
       ________28496, ________28497, ________28498, ________28499;
  wire ________28500, ________28503, ________28504, ________28505,
       ________28506, ________28507, ________28508, ________28509;
  wire ________28512, ________28513, ________28514, ________28515,
       ________28516, ________28517, ________28518, ________28519;
  wire ________28521, ________28522, ________28523, ________28524,
       ________28525, ________28526, ________28527, ________28528;
  wire ________28531, ________28532, ________28533, ________28534,
       ________28535, ________28536, ________28537, ________28539;
  wire ________28540, ________28541, ________28542, ________28543,
       ________28544, ________28545, ________28563, ________28564;
  wire ________28565, ________28566, ________28567, ________28568,
       ________28569, ________28572, ________28573, ________28574;
  wire ________28575, ________28576, ________28577, ________28578,
       ________28579, ________28582, ________28583, ________28584;
  wire ________28585, ________28586, ________28587, ________28588,
       ________28589, ________28592, ________28593, ________28594;
  wire ________28595, ________28596, ________28597, ________28599,
       ________28600, ________28601, ________28602, ________28603;
  wire ________28604, ________28605, ________28606, ________28609,
       ________28610, ________28611, ________28612, ________28613;
  wire ________28614, ________28615, ________28616, ________28619,
       ________28620, ________28621, ________28622, ________28623;
  wire ________28624, ________28625, ________28628, ________28629,
       ________28630, ________28631, ________28632, ________28633;
  wire ________28634, ________28635, ________28845, ________28846,
       ________28847, ________28848, ________28849, ________28850;
  wire ________28851, ________28852, ________28855, ________28856,
       ________28857, ________28858, ________28859, ________28860;
  wire ________28861, ________28864, ________28865, ________28866,
       ________28867, ________28868, ________28869, ________28870;
  wire ________28873, ________28874, ________28875, ________28876,
       ________28877, ________28878, ________28879, ________28882;
  wire ________28883, ________28884, ________28885, ________28886,
       ________28887, ________28888, ________28889, ________28891;
  wire ________28892, ________28893, ________28894, ________28895,
       ________28898, ________28899, ________28900, ________28901;
  wire ________28902, ________28903, ________28904, ________28907,
       ________28908, ________28909, ________28910, ________28911;
  wire ________28912, ________28913, ________28933, ________28934,
       ________28935, ________28936, ________28937, ________28938;
  wire ________28939, ________28942, ________28943, ________28944,
       ________28945, ________28948, ________28949, ________28950;
  wire ________28951, ________28952, ________28953, ________28954,
       ________28955, ________28957, ________28958, ________28959;
  wire ________28960, ________28961, ________28962, ________28963,
       ________28964, ________28967, ________28968, ________28969;
  wire ________28970, ________28971, ________28974, ________28975,
       ________28976, ________28977, ________28978, ________28979;
  wire ________28980, ________28982, ________28983, ________28984,
       ________28985, ________28986, ________28987, ________28988;
  wire ________28991, ________28992, ________28993, ________28994,
       ________28995, ________28996, ________28997, ________29019;
  wire ________29020, ________29021, ________29022, ________29023,
       ________29024, ________29025, ________29026, ________29029;
  wire ________29030, ________29031, ________29032, ________29033,
       ________29034, ________29035, ________29038, ________29039;
  wire ________29040, ________29041, ________29042, ________29043,
       ________29044, ________29047, ________29048, ________29049;
  wire ________29050, ________29051, ________29052, ________29053,
       ________29056, ________29057, ________29058, ________29059;
  wire ________29060, ________29061, ________29062, ________29063,
       ________29066, ________29067, ________29068, ________29069;
  wire ________29070, ________29071, ________29072, ________29073,
       ________29076, ________29077, ________29078, ________29079;
  wire ________29080, ________29081, ________29084, ________29085,
       ________29086, ________29087, ________29088, ________29089;
  wire ________29090, ________29108, ________29109, ________29110,
       ________29111, ________29112, ________29113, ________29114;
  wire ________29115, ________29118, ________29119, ________29120,
       ________29121, ________29122, ________29123, ________29124;
  wire ________29125, ________29128, ________29129, ________29130,
       ________29131, ________29132, ________29133, ________29134;
  wire ________29137, ________29138, ________29139, ________29140,
       ________29141, ________29142, ________29143, ________29144;
  wire ________29147, ________29148, ________29149, ________29150,
       ________29151, ________29152, ________29153, ________29154;
  wire ________29156, ________29157, ________29158, ________29159,
       ________29160, ________29161, ________29162, ________29163;
  wire ________29166, ________29167, ________29168, ________29169,
       ________29170, ________29171, ________29172, ________29173;
  wire ________29176, ________29177, ________29178, ________29179,
       ________29180, ________29181, ________29182, ________29183;
  wire ________29205, ________29206, ________29207, ________29208,
       ________29209, ________29210, ________29211, ________29212;
  wire ________29214, ________29215, ________29216, ________29217,
       ________29220, ________29221, ________29222, ________29223;
  wire ________29224, ________29225, ________29226, ________29228,
       ________29229, ________29230, ________29231, ________29232;
  wire ________29233, ________29236, ________29237, ________29238,
       ________29239, ________29240, ________29241, ________29242;
  wire ________29243, ________29245, ________29246, ________29247,
       ________29248, ________29249, ________29250, ________29251;
  wire ________29253, ________29254, ________29255, ________29256,
       ________29257, ________29258, ________29259, ________29260;
  wire ________29263, ________29264, ________29265, ________29266,
       ________29267, ________29268, ________29269, ________29270;
  wire ________29289, ________29290, ________29291, ________29292,
       ________29293, ________29294, ________29297, ________29298;
  wire ________29299, ________29300, ________29301, ________29302,
       ________29303, ________29306, ________29307, ________29308;
  wire ________29309, ________29310, ________29311, ________29312,
       ________29313, ________29316, ________29317, ________29318;
  wire ________29319, ________29320, ________29321, ________29322,
       ________29323, ________29326, ________29327, ________29328;
  wire ________29329, ________29330, ________29331, ________29332,
       ________29333, ________29336, ________29337, ________29338;
  wire ________29339, ________29340, ________29341, ________29342,
       ________29343, ________29346, ________29347, ________29348;
  wire ________29349, ________29350, ________29351, ________29354,
       ________29355, ________29356, ________29357, ________29358;
  wire ________29359, ________29360, ________29361, ________29379,
       ________29380, ________29381, ________29382, ________29383;
  wire ________29384, ________29385, ________29388, ________29389,
       ________29390, ________29391, ________29392, ________29393;
  wire ________29394, ________29395, ________29398, ________29399,
       ________29400, ________29401, ________29402, ________29403;
  wire ________29404, ________29405, ________29408, ________29409,
       ________29410, ________29411, ________29412, ________29413;
  wire ________29414, ________29415, ________29418, ________29419,
       ________29420, ________29421, ________29422, ________29423;
  wire ________29424, ________29427, ________29428, ________29429,
       ________29430, ________29431, ________29432, ________29433;
  wire ________29434, ________29437, ________29438, ________29439,
       ________29440, ________29441, ________29442, ________29443;
  wire ________29444, ________29447, ________29448, ________29449,
       ________29450, ________29451, ________29452, ________29453;
  wire ________29454, ________29477, ________29478, ________29479,
       ________29480, ________29481, ________29482, ________29483;
  wire ________29484, ________29487, ________29488, ________29489,
       ________29490, ________29491, ________29492, ________29493;
  wire ________29494, ________29496, ________29497, ________29498,
       ________29499, ________29500, ________29501, ________29504;
  wire ________29505, ________29506, ________29507, ________29508,
       ________29511, ________29512, ________29513, ________29514;
  wire ________29515, ________29516, ________29517, ________29518,
       ________29519, ________29520, ________29521, ________29522;
  wire ________29523, ________29524, ________29525, ________29528,
       ________29529, ________29530, ________29531, ________29532;
  wire ________29533, ________29535, ________29536, ________29537,
       ________29538, ________29539, ________29540, ________29541;
  wire _________0_, _________9_, _________22014, _________22015,
       _________22016, _________22019, _________22020, _________22021;
  wire _________22022, _________22023, _________22024, _________22025,
       _________22028, _________22029, _________22031, _________22032;
  wire _________22033, _________22036, _________22037, _________22038,
       _________22039, _________22041, _________22042, _________22043;
  wire _________22044, _________22045, _________22046, _________22047,
       _________31614, _________31615, _________31616, _________31617;
  wire _________31618, _________31619, _________31620, _________31621,
       _________31624, _________31625, _________31626, _________31627;
  wire _________31628, _________31629, _________31630, _________31631,
       _________31634, _________31635, _________31636, _________31637;
  wire _________31638, _________31639, _________31642, _________31643,
       _________31644, _________31645, _________31646, _________31647;
  wire _________31648, _________31649, _________31652, _________31653,
       _________31654, _________31655, _________31656, _________31657;
  wire _________31658, _________31659, _________31662, _________31663,
       _________31664, _________31665, _________31666, _________31667;
  wire _________31668, _________31669, _________31672, _________31673,
       _________31674, _________31675, _________31676, _________31677;
  wire _________31678, _________31681, _________31682, _________31683,
       _________31684, _________31685, _________31686, _________31687;
  wire _________31710, _________31711, _________31712, _________31713,
       _________31714, _________31715, _________31716, _________31719;
  wire _________31720, _________31721, _________31722, _________31723,
       _________31724, _________31725, _________31726, _________31729;
  wire _________31730, _________31731, _________31732, _________31733,
       _________31734, _________31735, _________31738, _________31739;
  wire _________31740, _________31741, _________31742, _________31743,
       _________31744, _________31745, _________31748, _________31749;
  wire _________31750, _________31751, _________31752, _________31753,
       _________31754, _________31757, _________31758, _________31759;
  wire _________31760, _________31761, _________31762, _________31763,
       _________31764, _________31767, _________31768, _________31769;
  wire _________31770, _________31771, _________31772, _________31773,
       _________31774, _________31777, _________31778, _________31779;
  wire _________31780, _________31781, _________31782, _________31783,
       _________31784, _________31806, _________31807, _________31808;
  wire _________31809, _________31810, _________31811, _________31812,
       _________31813, _________31816, _________31817, _________31818;
  wire _________31819, _________31820, _________31821, _________31822,
       _________31823, _________31826, _________31827, _________31828;
  wire _________31829, _________31830, _________31831, _________31832,
       _________31833, _________31836, _________31837, _________31838;
  wire _________31839, _________31840, _________31841, _________31842,
       _________31843, _________31846, _________31847, _________31848;
  wire _________31849, _________31850, _________31851, _________31852,
       _________31853, _________31856, _________31857, _________31858;
  wire _________31859, _________31860, _________31861, _________31862,
       _________31863, _________31866, _________31867, _________31868;
  wire _________31869, _________31870, _________31871, _________31872,
       _________31873, _________31876, _________31877, _________31878;
  wire _________31879, _________31880, _________31881, _________31882,
       _________31883, _________31904, _________31905, _________31906;
  wire _________31907, _________31908, _________31909, _________31912,
       _________31913, _________31914, _________31915, _________31916;
  wire _________31917, _________31918, _________31919, _________31922,
       _________31923, _________31924, _________31925, _________31926;
  wire _________31927, _________31928, _________31929, _________31932,
       _________31933, _________31934, _________31935, _________31936;
  wire _________31937, _________31938, _________31941, _________31942,
       _________31943, _________31944, _________31945, _________31946;
  wire _________31947, _________31948, _________31951, _________31952,
       _________31953, _________31954, _________31955, _________31956;
  wire _________31957, _________31958, _________31961, _________31962,
       _________31963, _________31964, _________31965, _________31966;
  wire _________31967, _________31968, _________31971, _________31972,
       _________31973, _________31974, _________31975, _________31976;
  wire _________31977, _________31978, _________32001, _________32002,
       _________32003, _________32004, _________32005, _________32006;
  wire _________32007, _________32008, _________32011, _________32012,
       _________32013, _________32014, _________32015, _________32016;
  wire _________32017, _________32018, _________32021, _________32022,
       _________32023, _________32024, _________32025, _________32026;
  wire _________32027, _________32028, _________32031, _________32032,
       _________32033, _________32034, _________32035, _________32036;
  wire _________32037, _________32038, _________32041, _________32042,
       _________32043, _________32044, _________32045, _________32046;
  wire _________32047, _________32048, _________32051, _________32052,
       _________32053, _________32054, _________32055, _________32056;
  wire _________32057, _________32058, _________32061, _________32062,
       _________32063, _________32064, _________32065, _________32066;
  wire _________32067, _________32068, _________32071, _________32072,
       _________32073, _________32074, _________32075, _________32076;
  wire _________32077, _________32078, _________32099, _________32100,
       _________32101, _________32102, _________32103, _________32104;
  wire _________32105, _________32106, _________32109, _________32110,
       _________32111, _________32112, _________32113, _________32114;
  wire _________32115, _________32116, _________32119, _________32120,
       _________32121, _________32122, _________32123, _________32124;
  wire _________32125, _________32128, _________32129, _________32130,
       _________32131, _________32132, _________32133, _________32134;
  wire _________32135, _________32138, _________32139, _________32140,
       _________32141, _________32142, _________32143, _________32144;
  wire _________32145, _________32148, _________32149, _________32150,
       _________32151, _________32152, _________32153, _________32154;
  wire _________32157, _________32158, _________32159, _________32160,
       _________32161, _________32162, _________32163, _________32164;
  wire _________32167, _________32168, _________32169, _________32170,
       _________32171, _________32172, _________32173, _________32174;
  wire _________32197, _________32198, _________32199, _________32200,
       _________32201, _________32202, _________32203, _________32206;
  wire _________32207, _________32208, _________32209, _________32210,
       _________32211, _________32212, _________32215, _________32216;
  wire _________32217, _________32218, _________32219, _________32220,
       _________32221, _________32222, _________32225, _________32226;
  wire _________32227, _________32228, _________32229, _________32230,
       _________32231, _________32232, _________32235, _________32236;
  wire _________32237, _________32238, _________32239, _________32240,
       _________32241, _________32244, _________32245, _________32246;
  wire _________32247, _________32248, _________32249, _________32250,
       _________32251, _________32254, _________32255, _________32256;
  wire _________32257, _________32258, _________32259, _________32260,
       _________32261, _________32264, _________32265, _________32266;
  wire _________32267, _________32268, _________32269, _________32270,
       _________32271, _________32294, _________32295, _________32296;
  wire _________32297, _________32298, _________32299, _________32300,
       _________32301, _________32304, _________32305, _________32306;
  wire _________32307, _________32308, _________32309, _________32310,
       _________32311, _________32314, _________32315, _________32316;
  wire _________32317, _________32318, _________32319, _________32322,
       _________32323, _________32324, _________32325, _________32326;
  wire _________32327, _________32328, _________32329, _________32332,
       _________32333, _________32334, _________32335, _________32336;
  wire _________32337, _________32338, _________32339, _________32342,
       _________32343, _________32344, _________32345, _________32346;
  wire _________32347, _________32348, _________32349, _________32352,
       _________32353, _________32354, _________32355, _________32356;
  wire _________32357, _________32358, _________32359, _________32362,
       _________32363, _________32364, _________32365, _________32366;
  wire _________32367, _________32368, _________32369, _________32587,
       _________32588, _________32589, _________32590, _________32591;
  wire _________32592, _________32593, _________32594, _________32597,
       _________32598, _________32599, _________32600, _________32601;
  wire _________32602, _________32603, _________32604, _________32607,
       _________32608, _________32609, _________32610, _________32611;
  wire _________32612, _________32613, _________32614, _________32617,
       _________32618, _________32619, _________32620, _________32621;
  wire _________32622, _________32623, _________32624, _________32627,
       _________32628, _________32629, _________32630, _________32631;
  wire _________32632, _________32633, _________32634, _________32637,
       _________32638, _________32639, _________32640, _________32641;
  wire _________32642, _________32643, _________32644, _________32647,
       _________32648, _________32649, _________32650, _________32651;
  wire _________32652, _________32653, _________32654, _________32657,
       _________32658, _________32659, _________32660, _________32661;
  wire _________32662, _________32663, _________32664, _________32686,
       _________32687, _________32688, _________32689, _________32690;
  wire _________32691, _________32692, _________32695, _________32696,
       _________32697, _________32698, _________32699, _________32700;
  wire _________32701, _________32702, _________32705, _________32706,
       _________32707, _________32708, _________32709, _________32710;
  wire _________32711, _________32712, _________32715, _________32716,
       _________32717, _________32718, _________32719, _________32720;
  wire _________32721, _________32722, _________32725, _________32726,
       _________32727, _________32728, _________32729, _________32730;
  wire _________32731, _________32732, _________32735, _________32736,
       _________32737, _________32738, _________32739, _________32740;
  wire _________32741, _________32742, _________32745, _________32746,
       _________32747, _________32748, _________32749, _________32750;
  wire _________32751, _________32752, _________32755, _________32756,
       _________32757, _________32758, _________32759, _________32760;
  wire _________32761, _________32762, _________32784, _________32785,
       _________32786, _________32787, _________32788, _________32789;
  wire _________32790, _________32791, _________32794, _________32795,
       _________32796, _________32797, _________32798, _________32799;
  wire _________32800, _________32801, _________32804, _________32805,
       _________32806, _________32807, _________32808, _________32809;
  wire _________32810, _________32811, _________32814, _________32815,
       _________32816, _________32817, _________32818, _________32819;
  wire _________32820, _________32821, _________32824, _________32825,
       _________32826, _________32827, _________32828, _________32829;
  wire _________32830, _________32831, _________32834, _________32835,
       _________32836, _________32837, _________32838, _________32839;
  wire _________32840, _________32841, _________32844, _________32845,
       _________32846, _________32847, _________32848, _________32849;
  wire _________32850, _________32851, _________32854, _________32855,
       _________32856, _________32857, _________32858, _________32859;
  wire _________32860, _________32883, _________32884, _________32885,
       _________32886, _________32887, _________32888, _________32889;
  wire _________32890, _________32893, _________32894, _________32895,
       _________32896, _________32897, _________32898, _________32899;
  wire _________32900, _________32903, _________32904, _________32905,
       _________32906, _________32907, _________32908, _________32909;
  wire _________32910, _________32913, _________32914, _________32915,
       _________32916, _________32917, _________32918, _________32919;
  wire _________32920, _________32922, _________32923, _________32924,
       _________32925, _________32926, _________32927, _________32928;
  wire _________32931, _________32932, _________32933, _________32934,
       _________32935, _________32936, _________32937, _________32938;
  wire _________32941, _________32942, _________32943, _________32944,
       _________32945, _________32946, _________32947, _________32948;
  wire _________32951, _________32952, _________32953, _________32954,
       _________32955, _________32956, _________32957, _________32958;
  wire _________32981, _________32982, _________32983, _________32984,
       _________32985, _________32986, _________32987, _________32988;
  wire _________32991, _________32992, _________32993, _________32994,
       _________32995, _________32996, _________32997, _________33000;
  wire _________33001, _________33002, _________33003, _________33004,
       _________33005, _________33006, _________33009, _________33010;
  wire _________33011, _________33012, _________33013, _________33014,
       _________33015, _________33016, _________33019, _________33020;
  wire _________33021, _________33022, _________33023, _________33024,
       _________33025, _________33026, _________33029, _________33030;
  wire _________33031, _________33032, _________33033, _________33034,
       _________33035, _________33036, _________33039, _________33040;
  wire _________33041, _________33042, _________33043, _________33044,
       _________33047, _________33048, _________33049, _________33050;
  wire _________33051, _________33052, _________33053, _________33054,
       _________33076, _________33077, _________33078, _________33079;
  wire _________33080, _________33081, _________33082, _________33085,
       _________33086, _________33087, _________33088, _________33089;
  wire _________33090, _________33091, _________33094, _________33095,
       _________33096, _________33097, _________33098, _________33099;
  wire _________33100, _________33101, _________33104, _________33105,
       _________33106, _________33107, _________33108, _________33109;
  wire _________33110, _________33111, _________33113, _________33114,
       _________33115, _________33116, _________33117, _________33118;
  wire _________33119, _________33120, _________33123, _________33124,
       _________33125, _________33126, _________33127, _________33128;
  wire _________33129, _________33130, _________33133, _________33134,
       _________33135, _________33136, _________33137, _________33138;
  wire _________33139, _________33142, _________33143, _________33144,
       _________33145, _________33146, _________33147, _________33169;
  wire _________33170, _________33171, _________33172, _________33173,
       _________33174, _________33175, _________33178, _________33179;
  wire _________33180, _________33181, _________33182, _________33183,
       _________33184, _________33187, _________33188, _________33189;
  wire _________33190, _________33191, _________33192, _________33193,
       _________33196, _________33197, _________33198, _________33199;
  wire _________33200, _________33201, _________33202, _________33205,
       _________33206, _________33207, _________33208, _________33209;
  wire _________33210, _________33211, _________33212, _________33214,
       _________33215, _________33216, _________33217, _________33218;
  wire _________33219, _________33220, _________33223, _________33224,
       _________33225, _________33226, _________33227, _________33228;
  wire _________33229, _________33232, _________33233, _________33234,
       _________33235, _________33236, _________33237, _________33238;
  wire _________33239, _________33260, _________33261, _________33262,
       _________33263, _________33264, _________33265, _________33266;
  wire _________33269, _________33270, _________33271, _________33272,
       _________33273, _________33274, _________33275, _________33278;
  wire _________33279, _________33280, _________33281, _________33282,
       _________33285, _________33286, _________33287, _________33288;
  wire _________33289, _________33290, _________33291, _________33293,
       _________33294, _________33295, _________33296, _________33297;
  wire _________33298, _________33299, _________33300, _________33303,
       _________33304, _________33305, _________33306, _________33307;
  wire _________33308, _________33309, _________33310, _________33313,
       _________33314, _________33315, _________33316, _________33317;
  wire _________33318, _________33319, _________33320, _________33321,
       _________33322, _________33323, _________33324, _________33325;
  wire _________33539, _________33540, _________33541, _________33542,
       _________33543, _________33544, _________33545, _________33546;
  wire _________33549, _________33550, _________33551, _________33552,
       _________33553, _________33554, _________33555, _________33557;
  wire _________33558, _________33559, _________33560, _________33561,
       _________33562, _________33563, _________33564, _________33567;
  wire _________33568, _________33569, _________33570, _________33571,
       _________33572, _________33573, _________33574, _________33577;
  wire _________33578, _________33579, _________33580, _________33581,
       _________33582, _________33583, _________33586, _________33587;
  wire _________33588, _________33589, _________33590, _________33591,
       _________33592, _________33593, _________33596, _________33597;
  wire _________33598, _________33599, _________33600, _________33601,
       _________33602, _________33603, _________33605, _________33606;
  wire _________33607, _________33608, _________33609, _________33610,
       _________33611, _________33631, _________33632, _________33633;
  wire _________33634, _________33635, _________33636, _________33637,
       _________33638, _________33641, _________33642, _________33643;
  wire _________33644, _________33645, _________33646, _________33647,
       _________33650, _________33651, _________33652, _________33653;
  wire _________33654, _________33655, _________33656, _________33657,
       _________33660, _________33661, _________33662, _________33663;
  wire _________33664, _________33665, _________33666, _________33667,
       _________33670, _________33671, _________33672, _________33673;
  wire _________33674, _________33675, _________33676, _________33677,
       _________33680, _________33681, _________33682, _________33683;
  wire _________33684, _________33685, _________33686, _________33687,
       _________33690, _________33691, _________33692, _________33693;
  wire _________33694, _________33695, _________33696, _________33697,
       _________33700, _________33701, _________33702, _________33703;
  wire _________33704, _________33705, _________33728, _________33729,
       _________33730, _________33731, _________33732, _________33733;
  wire _________33734, _________33737, _________33738, _________33739,
       _________33740, _________33741, _________33742, _________33743;
  wire _________33744, _________33747, _________33748, _________33749,
       _________33750, _________33751, _________33752, _________33753;
  wire _________33754, _________33757, _________33758, _________33759,
       _________33760, _________33761, _________33762, _________33763;
  wire _________33766, _________33767, _________33768, _________33769,
       _________33770, _________33771, _________33772, _________33773;
  wire _________33776, _________33777, _________33778, _________33779,
       _________33780, _________33781, _________33782, _________33783;
  wire _________33786, _________33787, _________33788, _________33789,
       _________33790, _________33791, _________33792, _________33793;
  wire _________33796, _________33797, _________33798, _________33799,
       _________33800, _________33801, _________33802, _________33803;
  wire _________33824, _________33825, _________33826, _________33827,
       _________33828, _________33829, _________33830, _________33831;
  wire _________33834, _________33835, _________33836, _________33837,
       _________33838, _________33839, _________33840, _________33843;
  wire _________33844, _________33845, _________33846, _________33847,
       _________33848, _________33849, _________33850, _________33853;
  wire _________33854, _________33855, _________33856, _________33857,
       _________33858, _________33859, _________33862, _________33863;
  wire _________33864, _________33865, _________33866, _________33867,
       _________33868, _________33869, _________33872, _________33873;
  wire _________33874, _________33875, _________33876, _________33877,
       _________33878, _________33879, _________33882, _________33883;
  wire _________33884, _________33885, _________33886, _________33887,
       _________33888, _________33891, _________33892, _________33893;
  wire _________33894, _________33895, _________33896, _________33897,
       _________33898, _________33919, _________33920, _________33921;
  wire _________33922, _________33923, _________33924, _________33925,
       _________33926, _________33929, _________33930, _________33931;
  wire _________33932, _________33933, _________33934, _________33935,
       _________33938, _________33939, _________33940, _________33941;
  wire _________33942, _________33943, _________33944, _________33947,
       _________33948, _________33949, _________33950, _________33951;
  wire _________33952, _________33953, _________33954, _________33957,
       _________33958, _________33959, _________33960, _________33961;
  wire _________33962, _________33963, _________33964, _________33967,
       _________33968, _________33969, _________33970, _________33971;
  wire _________33972, _________33973, _________33974, _________33976,
       _________33977, _________33978, _________33979, _________33980;
  wire _________33981, _________33982, _________33985, _________33986,
       _________33987, _________33988, _________33989, _________33990;
  wire _________33991, _________33992, _________34013, _________34014,
       _________34015, _________34016, _________34017, _________34018;
  wire _________34019, _________34022, _________34023, _________34024,
       _________34025, _________34026, _________34027, _________34028;
  wire _________34029, _________34032, _________34033, _________34034,
       _________34035, _________34036, _________34037, _________34038;
  wire _________34039, _________34042, _________34043, _________34044,
       _________34045, _________34046, _________34047, _________34048;
  wire _________34049, _________34052, _________34053, _________34054,
       _________34055, _________34056, _________34057, _________34058;
  wire _________34061, _________34062, _________34063, _________34064,
       _________34065, _________34066, _________34067, _________34070;
  wire _________34071, _________34072, _________34073, _________34074,
       _________34075, _________34076, _________34077, _________34080;
  wire _________34081, _________34082, _________34083, _________34084,
       _________34085, _________34086, _________34087, _________34109;
  wire _________34110, _________34111, _________34112, _________34113,
       _________34114, _________34115, _________34118, _________34119;
  wire _________34120, _________34121, _________34122, _________34123,
       _________34126, _________34127, _________34128, _________34129;
  wire _________34130, _________34131, _________34132, _________34135,
       _________34136, _________34137, _________34138, _________34139;
  wire _________34140, _________34141, _________34142, _________34144,
       _________34145, _________34146, _________34147, _________34148;
  wire _________34149, _________34150, _________34151, _________34154,
       _________34155, _________34156, _________34157, _________34158;
  wire _________34159, _________34160, _________34163, _________34164,
       _________34165, _________34166, _________34167, _________34168;
  wire _________34169, _________34170, _________34173, _________34174,
       _________34175, _________34176, _________34177, _________34178;
  wire _________34179, _________34202, _________34203, _________34204,
       _________34205, _________34206, _________34207, _________34208;
  wire _________34211, _________34212, _________34213, _________34214,
       _________34215, _________34216, _________34217, _________34220;
  wire _________34221, _________34222, _________34223, _________34224,
       _________34225, _________34226, _________34227, _________34230;
  wire _________34231, _________34232, _________34233, _________34234,
       _________34235, _________34236, _________34237, _________34240;
  wire _________34241, _________34242, _________34243, _________34244,
       _________34245, _________34246, _________34247, _________34250;
  wire _________34251, _________34252, _________34253, _________34254,
       _________34255, _________34256, _________34257, _________34260;
  wire _________34261, _________34262, _________34263, _________34264,
       _________34265, _________34268, _________34269, _________34270;
  wire _________34271, _________34272, _________34273, _________34274,
       _________34275, _________34490, _________34491, _________34492;
  wire _________34493, _________34494, _________34495, _________34496,
       _________34497, _________34500, _________34501, _________34502;
  wire _________34503, _________34504, _________34505, _________34506,
       _________34509, _________34510, _________34511, _________34512;
  wire _________34513, _________34514, _________34515, _________34518,
       _________34519, _________34520, _________34521, _________34522;
  wire _________34525, _________34526, _________34527, _________34528,
       _________34529, _________34530, _________34531, _________34532;
  wire _________34535, _________34536, _________34537, _________34538,
       _________34539, _________34540, _________34541, _________34542;
  wire _________34545, _________34546, _________34547, _________34548,
       _________34549, _________34550, _________34551, _________34552;
  wire _________34554, _________34555, _________34556, _________34557,
       _________34558, _________34559, _________34576, _________34577;
  wire _________34578, _________34579, _________34580, _________34581,
       _________34582, _________34583, _________34586, _________34587;
  wire _________34588, _________34589, _________34590, _________34591,
       _________34592, _________34595, _________34596, _________34597;
  wire _________34598, _________34599, _________34600, _________34601,
       _________34602, _________34605, _________34606, _________34607;
  wire _________34608, _________34609, _________34610, _________34611,
       _________34614, _________34615, _________34616, _________34617;
  wire _________34618, _________34619, _________34620, _________34623,
       _________34624, _________34625, _________34626, _________34627;
  wire _________34628, _________34629, _________34632, _________34633,
       _________34634, _________34635, _________34636, _________34637;
  wire _________34640, _________34641, _________34642, _________34643,
       _________34644, _________34645, _________34646, _________34647;
  wire _________34669, _________34670, _________34671, _________34672,
       _________34673, _________34674, _________34675, _________34678;
  wire _________34679, _________34680, _________34681, _________34682,
       _________34683, _________34684, _________34685, _________34688;
  wire _________34689, _________34690, _________34691, _________34692,
       _________34693, _________34694, _________34695, _________34698;
  wire _________34699, _________34700, _________34701, _________34702,
       _________34703, _________34704, _________34706, _________34707;
  wire _________34708, _________34709, _________34710, _________34711,
       _________34712, _________34713, _________34716, _________34717;
  wire _________34718, _________34719, _________34720, _________34721,
       _________34722, _________34723, _________34726, _________34727;
  wire _________34728, _________34729, _________34730, _________34731,
       _________34732, _________34733, _________34735, _________34736;
  wire _________34737, _________34738, _________34739, _________34740,
       _________34741, _________34742, _________34763, _________34764;
  wire _________34765, _________34766, _________34767, _________34768,
       _________34769, _________34770, _________34773, _________34774;
  wire _________34775, _________34776, _________34777, _________34778,
       _________34781, _________34782, _________34783, _________34784;
  wire _________34785, _________34786, _________34787, _________34788,
       _________34791, _________34792, _________34793, _________34794;
  wire _________34795, _________34796, _________34797, _________34798,
       _________34801, _________34802, _________34803, _________34804;
  wire _________34805, _________34806, _________34807, _________34808,
       _________34811, _________34812, _________34813, _________34814;
  wire _________34815, _________34816, _________34817, _________34820,
       _________34821, _________34822, _________34823, _________34824;
  wire _________34825, _________34826, _________34829, _________34830,
       _________34831, _________34832, _________34833, _________34834;
  wire _________34835, _________34836, _________34856, _________34857,
       _________34858, _________34859, _________34860, _________34861;
  wire _________34862, _________34864, _________34865, _________34866,
       _________34867, _________34868, _________34869, _________34872;
  wire _________34873, _________34874, _________34875, _________34876,
       _________34877, _________34878, _________34879, _________34881;
  wire _________34882, _________34883, _________34884, _________34885,
       _________34886, _________34889, _________34890, _________34891;
  wire _________34892, _________34893, _________34894, _________34895,
       _________34898, _________34899, _________34900, _________34901;
  wire _________34902, _________34903, _________34906, _________34907,
       _________34908, _________34909, _________34910, _________34911;
  wire _________34912, _________34913, _________34916, _________34917,
       _________34918, _________34919, _________34920, _________34921;
  wire _________34941, _________34942, _________34943, _________34944,
       _________34945, _________34946, _________34947, _________34950;
  wire _________34951, _________34952, _________34953, _________34954,
       _________34955, _________34956, _________34957, _________34958;
  wire _________34959, _________34960, _________34961, _________34962,
       _________34963, _________34966, _________34967, _________34968;
  wire _________34969, _________34970, _________34971, _________34972,
       _________34973, _________34976, _________34977, _________34978;
  wire _________34979, _________34980, _________34983, _________34984,
       _________34985, _________34986, _________34987, _________34988;
  wire _________34989, _________34990, _________34991, _________34992,
       _________34993, _________34994, _________34995, _________34996;
  wire _________34999, _________35000, _________35001, _________35002,
       _________35003, _________35004, _________35005, _________35006;
  wire _________35025, _________35026, _________35027, _________35028,
       _________35029, _________35030, _________35031, _________35033;
  wire _________35034, _________35035, _________35036, _________35037,
       _________35038, _________35041, _________35042, _________35043;
  wire _________35044, _________35045, _________35046, _________35047,
       _________35048, _________35051, _________35052, _________35053;
  wire _________35054, _________35055, _________35056, _________35057,
       _________35058, _________35060, _________35061, _________35062;
  wire _________35063, _________35064, _________35065, _________35068,
       _________35069, _________35070, _________35071, _________35072;
  wire _________35073, _________35074, _________35075, _________35078,
       _________35079, _________35080, _________35081, _________35082;
  wire _________35083, _________35084, _________35085, _________35088,
       _________35089, _________35090, _________35091, _________35092;
  wire _________35093, _________35094, _________35114, _________35115,
       _________35116, _________35117, _________35118, _________35119;
  wire _________35120, _________35123, _________35124, _________35125,
       _________35126, _________35127, _________35128, _________35129;
  wire _________35130, _________35133, _________35134, _________35135,
       _________35136, _________35137, _________35138, _________35139;
  wire _________35142, _________35143, _________35144, _________35145,
       _________35146, _________35147, _________35148, _________35149;
  wire _________35152, _________35153, _________35154, _________35155,
       _________35156, _________35157, _________35158, _________35159;
  wire _________35162, _________35163, _________35164, _________35165,
       _________35166, _________35167, _________35168, _________35169;
  wire _________35172, _________35173, _________35174, _________35175,
       _________35176, _________35177, _________35178, _________35179;
  wire _________35182, _________35183, _________35184, _________35185,
       _________35186, _________35187, _________35188, _________35189;
  wire _________35389, _________35390, _________35391, _________35392,
       _________35393, _________35394, _________35395, _________35398;
  wire _________35399, _________35400, _________35401, _________35402,
       _________35403, _________35404, _________35407, _________35408;
  wire _________35409, _________35410, _________35411, _________35412,
       _________35413, _________35414, _________35417, _________35418;
  wire _________35419, _________35420, _________35421, _________35422,
       _________35423, _________35424, _________35427, _________35428;
  wire _________35429, _________35430, _________35433, _________35434,
       _________35435, _________35436, _________35437, _________35438;
  wire _________35439, _________35442, _________35443, _________35444,
       _________35445, _________35446, _________35447, _________35448;
  wire _________35449, _________35452, _________35453, _________35454,
       _________35455, _________35456, _________35457, _________35458;
  wire _________35459, _________35482, _________35483, _________35484,
       _________35485, _________35486, _________35487, _________35488;
  wire _________35490, _________35491, _________35492, _________35493,
       _________35494, _________35495, _________35496, _________35497;
  wire _________35500, _________35501, _________35502, _________35503,
       _________35504, _________35505, _________35506, _________35507;
  wire _________35510, _________35511, _________35512, _________35513,
       _________35514, _________35515, _________35516, _________35517;
  wire _________35520, _________35521, _________35522, _________35523,
       _________35524, _________35525, _________35526, _________35529;
  wire _________35530, _________35531, _________35532, _________35533,
       _________35534, _________35535, _________35538, _________35539;
  wire _________35540, _________35541, _________35542, _________35543,
       _________35546, _________35547, _________35548, _________35549;
  wire _________35550, _________35551, _________35552, _________35553,
       _________35576, _________35577, _________35578, _________35579;
  wire _________35580, _________35581, _________35582, _________35583,
       _________35586, _________35587, _________35588, _________35589;
  wire _________35590, _________35591, _________35592, _________35595,
       _________35596, _________35597, _________35598, _________35599;
  wire _________35600, _________35601, _________35604, _________35605,
       _________35606, _________35607, _________35608, _________35609;
  wire _________35610, _________35611, _________35613, _________35614,
       _________35615, _________35616, _________35617, _________35618;
  wire _________35621, _________35622, _________35623, _________35624,
       _________35625, _________35626, _________35629, _________35630;
  wire _________35631, _________35632, _________35633, _________35634,
       _________35635, _________35637, _________35638, _________35639;
  wire _________35640, _________35641, _________35642, _________35661,
       _________35662, _________35663, _________35664, _________35665;
  wire _________35666, _________35668, _________35669, _________35670,
       _________35671, _________35672, _________35673, _________35674;
  wire _________35676, _________35677, _________35678, _________35679,
       _________35680, _________35681, _________35682, _________35685;
  wire _________35686, _________35687, _________35688, _________35689,
       _________35690, _________35691, _________35692, _________35695;
  wire _________35696, _________35697, _________35698, _________35699,
       _________35700, _________35702, _________35703, _________35704;
  wire _________35705, _________35706, _________35707, _________35708,
       _________35709, _________35712, _________35713, _________35714;
  wire _________35715, _________35716, _________35717, _________35718,
       _________35719, _________35722, _________35723, _________35724;
  wire _________35725, _________35726, _________35727, _________35728,
       _________35729, _________35746, _________35747, _________35748;
  wire _________35749, _________35750, _________35751, _________35752,
       _________35753, _________35756, _________35757, _________35758;
  wire _________35759, _________35760, _________35761, _________35762,
       _________35763, _________35766, _________35767, _________35768;
  wire _________35769, _________35770, _________35771, _________35772,
       _________35775, _________35776, _________35777, _________35778;
  wire _________35779, _________35780, _________35781, _________35782,
       _________35785, _________35786, _________35787, _________35788;
  wire _________35789, _________35790, _________35791, _________35794,
       _________35795, _________35796, _________35797, _________35798;
  wire _________35799, _________35800, _________35801, _________35804,
       _________35805, _________35806, _________35807, _________35808;
  wire _________35809, _________35810, _________35811, _________35814,
       _________35815, _________35816, _________35817, _________35818;
  wire _________35819, _________35820, _________35821, _________35844,
       _________35845, _________35846, _________35847, _________35848;
  wire _________35849, _________35850, _________35851, _________35854,
       _________35855, _________35856, _________35857, _________35858;
  wire _________35859, _________35860, _________35861, _________35864,
       _________35865, _________35866, _________35867, _________35868;
  wire _________35869, _________35872, _________35873, _________35874,
       _________35875, _________35876, _________35877, _________35878;
  wire _________35881, _________35882, _________35883, _________35884,
       _________35885, _________35886, _________35887, _________35890;
  wire _________35891, _________35892, _________35893, _________35894,
       _________35895, _________35898, _________35899, _________35900;
  wire _________35901, _________35902, _________35903, _________35904,
       _________35905, _________35907, _________35908, _________35909;
  wire _________35910, _________35911, _________35912, _________35913,
       _________35914, _________35934, _________35935, _________35936;
  wire _________35937, _________35938, _________35939, _________35940,
       _________35943, _________35944, _________35945, _________35946;
  wire _________35949, _________35950, _________35951, _________35952,
       _________35953, _________35954, _________35955, _________35958;
  wire _________35959, _________35960, _________35961, _________35962,
       _________35963, _________35966, _________35967, _________35968;
  wire _________35969, _________35970, _________35971, _________35972,
       _________35973, _________35976, _________35977, _________35978;
  wire _________35979, _________35980, _________35981, _________35984,
       _________35985, _________35986, _________35987, _________35988;
  wire _________35989, _________35990, _________35991, _________35994,
       _________35995, _________35996, _________35997, _________35998;
  wire _________36019, _________36020, _________36021, _________36022,
       _________36023, _________36024, _________36025, _________36026;
  wire _________36029, _________36030, _________36031, _________36032,
       _________36033, _________36034, _________36035, _________36036;
  wire _________36039, _________36040, _________36041, _________36042,
       _________36043, _________36044, _________36045, _________36046;
  wire _________36048, _________36049, _________36050, _________36051,
       _________36052, _________36053, _________36054, _________36057;
  wire _________36058, _________36059, _________36060, _________36061,
       _________36062, _________36063, _________36066, _________36067;
  wire _________36068, _________36069, _________36070, _________36071,
       _________36073, _________36074, _________36075, _________36076;
  wire _________36077, _________36078, _________36079, _________36082,
       _________36083, _________36084, _________36085, _________36086;
  wire _________36087, _________36288, _________36289, _________36290,
       _________36291, _________36292, _________36293, _________36294;
  wire _________36296, _________36297, _________36298, _________36299,
       _________36300, _________36301, _________36303, _________36304;
  wire _________36305, _________36306, _________36307, _________36310,
       _________36311, _________36312, _________36313, _________36314;
  wire _________36315, _________36316, _________36317, _________36320,
       _________36321, _________36322, _________36323, _________36324;
  wire _________36325, _________36326, _________36327, _________36330,
       _________36331, _________36332, _________36333, _________36334;
  wire _________36335, _________36336, _________36339, _________36340,
       _________36341, _________36342, _________36343, _________36344;
  wire _________36345, _________36346, _________36349, _________36350,
       _________36351, _________36352, _________36353, _________36354;
  wire _________36355, _________36356, _________36376, _________36377,
       _________36378, _________36379, _________36380, _________36381;
  wire _________36382, _________36383, _________36386, _________36387,
       _________36388, _________36389, _________36390, _________36391;
  wire _________36392, _________36393, _________36395, _________36396,
       _________36397, _________36398, _________36399, _________36400;
  wire _________36401, _________36402, _________36405, _________36406,
       _________36407, _________36408, _________36409, _________36411;
  wire _________36412, _________36413, _________36414, _________36415,
       _________36416, _________36417, _________36418, _________36420;
  wire _________36421, _________36422, _________36423, _________36424,
       _________36425, _________36426, _________36429, _________36430;
  wire _________36431, _________36432, _________36433, _________36434,
       _________36435, _________36436, _________36439, _________36440;
  wire _________36441, _________36442, _________36443, _________36444,
       _________36445, _________36446, _________36464, _________36465;
  wire _________36466, _________36467, _________36468, _________36469,
       _________36470, _________36471, _________36474, _________36475;
  wire _________36476, _________36477, _________36478, _________36479,
       _________36480, _________36482, _________36483, _________36484;
  wire _________36485, _________36486, _________36487, _________36488,
       _________36489, _________36492, _________36493, _________36494;
  wire _________36495, _________36496, _________36497, _________36500,
       _________36501, _________36502, _________36503, _________36504;
  wire _________36505, _________36506, _________36509, _________36510,
       _________36511, _________36512, _________36513, _________36514;
  wire _________36517, _________36518, _________36519, _________36520,
       _________36521, _________36522, _________36523, _________36524;
  wire _________36527, _________36528, _________36529, _________36530,
       _________36531, _________36532, _________36533, _________36552;
  wire _________36553, _________36554, _________36555, _________36556,
       _________36557, _________36558, _________36559, _________36562;
  wire _________36563, _________36564, _________36565, _________36566,
       _________36567, _________36568, _________36571, _________36572;
  wire _________36573, _________36574, _________36575, _________36576,
       _________36577, _________36578, _________36581, _________36582;
  wire _________36583, _________36584, _________36585, _________36586,
       _________36587, _________36590, _________36591, _________36592;
  wire _________36593, _________36594, _________36595, _________36596,
       _________36599, _________36600, _________36601, _________36602;
  wire _________36605, _________36606, _________36607, _________36608,
       _________36609, _________36610, _________36611, _________36612;
  wire _________36615, _________36616, _________36617, _________36618,
       _________36619, _________36620, _________36621, _________36643;
  wire _________36644, _________36645, _________36646, _________36647,
       _________36648, _________36649, _________36650, _________36652;
  wire _________36653, _________36654, _________36655, _________36656,
       _________36657, _________36658, _________36661, _________36662;
  wire _________36663, _________36664, _________36665, _________36666,
       _________36667, _________36670, _________36671, _________36672;
  wire _________36673, _________36674, _________36675, _________36678,
       _________36679, _________36680, _________36681, _________36682;
  wire _________36683, _________36684, _________36685, _________36688,
       _________36689, _________36690, _________36691, _________36692;
  wire _________36693, _________36694, _________36695, _________36698,
       _________36699, _________36700, _________36701, _________36702;
  wire _________36703, _________36704, _________36705, _________36708,
       _________36709, _________36710, _________36711, _________36712;
  wire _________36713, _________36714, _________36715, _________36737,
       _________36738, _________36739, _________36740, _________36741;
  wire _________36742, _________36743, _________36744, _________36747,
       _________36748, _________36749, _________36750, _________36751;
  wire _________36752, _________36753, _________36754, _________36757,
       _________36758, _________36759, _________36760, _________36761;
  wire _________36762, _________36763, _________36764, _________36767,
       _________36768, _________36769, _________36770, _________36771;
  wire _________36772, _________36773, _________36776, _________36777,
       _________36778, _________36779, _________36780, _________36781;
  wire _________36782, _________36785, _________36786, _________36787,
       _________36788, _________36789, _________36790, _________36791;
  wire _________36794, _________36795, _________36796, _________36797,
       _________36798, _________36799, _________36800, _________36801;
  wire _________36804, _________36805, _________36806, _________36807,
       _________36808, _________36809, _________36810, _________36811;
  wire _________36834, _________36835, _________36836, _________36837,
       _________36838, _________36839, _________36840, _________36843;
  wire _________36844, _________36845, _________36846, _________36847,
       _________36848, _________36849, _________36852, _________36853;
  wire _________36854, _________36855, _________36856, _________36857,
       _________36858, _________36861, _________36862, _________36863;
  wire _________36864, _________36865, _________36866, _________36867,
       _________36870, _________36871, _________36872, _________36873;
  wire _________36874, _________36875, _________36876, _________36877,
       _________36880, _________36881, _________36882, _________36883;
  wire _________36884, _________36885, _________36886, _________36887,
       _________36890, _________36891, _________36892, _________36893;
  wire _________36894, _________36895, _________36898, _________36899,
       _________36900, _________36901, _________36902, _________36925;
  wire _________36926, _________36927, _________36928, _________36929,
       _________36930, _________36933, _________36934, _________36935;
  wire _________36936, _________36937, _________36938, _________36939,
       _________36940, _________36943, _________36944, _________36945;
  wire _________36946, _________36947, _________36948, _________36949,
       _________36952, _________36953, _________36954, _________36955;
  wire _________36956, _________36957, _________36958, _________36959,
       _________36962, _________36963, _________36964, _________36965;
  wire _________36966, _________36967, _________36968, _________36971,
       _________36972, _________36973, _________36974, _________36975;
  wire _________36976, _________36979, _________36980, _________36981,
       _________36982, _________36983, _________36986, _________36987;
  wire _________36988, _________36989, _________36990, _________36991,
       _________36992, _________36993, _________37199, _________37200;
  wire _________37201, _________37202, _________37203, _________37204,
       _________37206, _________37207, _________37208, _________37209;
  wire _________37210, _________37211, _________37212, _________37213,
       _________37215, _________37216, _________37217, _________37218;
  wire _________37219, _________37220, _________37221, _________37223,
       _________37224, _________37225, _________37226, _________37227;
  wire _________37228, _________37229, _________37230, _________37233,
       _________37234, _________37235, _________37236, _________37237;
  wire _________37238, _________37239, _________37241, _________37242,
       _________37243, _________37244, _________37245, _________37246;
  wire _________37249, _________37250, _________37251, _________37252,
       _________37253, _________37254, _________37255, _________37258;
  wire _________37259, _________37260, _________37261, _________37262,
       _________37263, _________37264, _________37265, _________37287;
  wire _________37288, _________37289, _________37290, _________37291,
       _________37292, _________37293, _________37296, _________37297;
  wire _________37298, _________37299, _________37300, _________37301,
       _________37302, _________37303, _________37306, _________37307;
  wire _________37308, _________37309, _________37310, _________37311,
       _________37312, _________37313, _________37316, _________37317;
  wire _________37318, _________37319, _________37320, _________37321,
       _________37322, _________37323, _________37326, _________37327;
  wire _________37328, _________37329, _________37330, _________37331,
       _________37332, _________37333, _________37336, _________37337;
  wire _________37338, _________37339, _________37340, _________37341,
       _________37342, _________37343, _________37346, _________37347;
  wire _________37348, _________37349, _________37350, _________37351,
       _________37352, _________37355, _________37356, _________37357;
  wire _________37358, _________37359, _________37360, _________37361,
       _________37383, _________37384, _________37385, _________37386;
  wire _________37387, _________37388, _________37389, _________37392,
       _________37393, _________37394, _________37395, _________37396;
  wire _________37397, _________37398, _________37399, _________37402,
       _________37403, _________37404, _________37405, _________37406;
  wire _________37407, _________37408, _________37409, _________37412,
       _________37413, _________37414, _________37415, _________37416;
  wire _________37417, _________37418, _________37421, _________37422,
       _________37423, _________37424, _________37425, _________37426;
  wire _________37427, _________37428, _________37431, _________37432,
       _________37433, _________37434, _________37435, _________37436;
  wire _________37437, _________37438, _________37441, _________37442,
       _________37443, _________37444, _________37445, _________37446;
  wire _________37447, _________37448, _________37451, _________37452,
       _________37453, _________37454, _________37455, _________37456;
  wire _________37457, _________37479, _________37480, _________37481,
       _________37482, _________37483, _________37484, _________37485;
  wire _________37486, _________37489, _________37490, _________37491,
       _________37492, _________37493, _________37494, _________37495;
  wire _________37496, _________37499, _________37500, _________37501,
       _________37502, _________37503, _________37504, _________37505;
  wire _________37508, _________37509, _________37510, _________37511,
       _________37512, _________37513, _________37514, _________37517;
  wire _________37518, _________37519, _________37520, _________37521,
       _________37522, _________37523, _________37524, _________37527;
  wire _________37528, _________37529, _________37530, _________37531,
       _________37532, _________37533, _________37534, _________37537;
  wire _________37538, _________37539, _________37540, _________37541,
       _________37542, _________37543, _________37544, _________37547;
  wire _________37548, _________37549, _________37550, _________37551,
       _________37552, _________37553, _________37554, _________37575;
  wire _________37576, _________37577, _________37578, _________37579,
       _________37580, _________37581, _________37582, _________37585;
  wire _________37586, _________37587, _________37588, _________37589,
       _________37590, _________37591, _________37592, _________37595;
  wire _________37596, _________37597, _________37598, _________37599,
       _________37600, _________37601, _________37602, _________37605;
  wire _________37606, _________37607, _________37608, _________37609,
       _________37610, _________37611, _________37612, _________37614;
  wire _________37615, _________37616, _________37617, _________37618,
       _________37619, _________37620, _________37621, _________37624;
  wire _________37625, _________37626, _________37627, _________37628,
       _________37629, _________37630, _________37631, _________37634;
  wire _________37635, _________37636, _________37637, _________37638,
       _________37639, _________37640, _________37641, _________37644;
  wire _________37645, _________37646, _________37647, _________37648,
       _________37649, _________37650, _________37651, _________37674;
  wire _________37675, _________37676, _________37677, _________37678,
       _________37679, _________37680, _________37681, _________37684;
  wire _________37685, _________37686, _________37687, _________37688,
       _________37689, _________37690, _________37691, _________37694;
  wire _________37695, _________37696, _________37697, _________37698,
       _________37699, _________37700, _________37703, _________37704;
  wire _________37705, _________37706, _________37707, _________37708,
       _________37709, _________37712, _________37713, _________37714;
  wire _________37715, _________37716, _________37717, _________37718,
       _________37719, _________37722, _________37723, _________37724;
  wire _________37725, _________37726, _________37727, _________37728,
       _________37729, _________37732, _________37733, _________37734;
  wire _________37735, _________37736, _________37737, _________37738,
       _________37739, _________37742, _________37743, _________37744;
  wire _________37745, _________37746, _________37747, _________37748,
       _________37749, _________37767, _________37768, _________37769;
  wire _________37770, _________37771, _________37772, _________37773,
       _________37774, _________37777, _________37778, _________37779;
  wire _________37780, _________37781, _________37782, _________37783,
       _________37784, _________37787, _________37788, _________37789;
  wire _________37790, _________37791, _________37792, _________37793,
       _________37794, _________37797, _________37798, _________37799;
  wire _________37800, _________37801, _________37802, _________37803,
       _________37806, _________37807, _________37808, _________37809;
  wire _________37810, _________37811, _________37812, _________37815,
       _________37816, _________37817, _________37818, _________37819;
  wire _________37820, _________37821, _________37822, _________37825,
       _________37826, _________37827, _________37828, _________37829;
  wire _________37830, _________37831, _________37834, _________37835,
       _________37836, _________37837, _________37838, _________37839;
  wire _________37840, _________37841, _________37864, _________37865,
       _________37866, _________37867, _________37868, _________37869;
  wire _________37870, _________37873, _________37874, _________37875,
       _________37876, _________37877, _________37878, _________37879;
  wire _________37880, _________37883, _________37884, _________37885,
       _________37886, _________37887, _________37888, _________37889;
  wire _________37890, _________37893, _________37894, _________37895,
       _________37896, _________37897, _________37898, _________37899;
  wire _________37902, _________37903, _________37904, _________37905,
       _________37906, _________37907, _________37908, _________37911;
  wire _________37912, _________37913, _________37914, _________37915,
       _________37916, _________37917, _________37918, _________37921;
  wire _________37922, _________37923, _________37924, _________37925,
       _________37926, _________37927, _________37930, _________37931;
  wire _________37932, _________37933, _________37934, _________37935,
       _________37936, _________37937, _________38142, _________38143;
  wire _________38144, _________38145, _________38146, _________38147,
       _________38148, _________38149, _________38152, _________38153;
  wire _________38154, _________38155, _________38156, _________38157,
       _________38158, _________38159, _________38162, _________38163;
  wire _________38164, _________38165, _________38166, _________38167,
       _________38168, _________38171, _________38172, _________38173;
  wire _________38174, _________38175, _________38176, _________38177,
       _________38178, _________38180, _________38181, _________38182;
  wire _________38183, _________38184, _________38185, _________38186,
       _________38187, _________38190, _________38191, _________38192;
  wire _________38193, _________38194, _________38195, _________38196,
       _________38197, _________38200, _________38201, _________38202;
  wire _________38203, _________38204, _________38205, _________38206,
       _________38207, _________38210, _________38211, _________38212;
  wire _________38213, _________38214, _________38215, _________38216,
       _________38238, _________38239, _________38240, _________38241;
  wire _________38242, _________38243, _________38244, _________38247,
       _________38248, _________38249, _________38250, _________38251;
  wire _________38252, _________38253, _________38254, _________38257,
       _________38258, _________38259, _________38260, _________38261;
  wire _________38262, _________38263, _________38264, _________38267,
       _________38268, _________38269, _________38270, _________38271;
  wire _________38272, _________38273, _________38274, _________38277,
       _________38278, _________38279, _________38280, _________38281;
  wire _________38282, _________38283, _________38284, _________38287,
       _________38288, _________38289, _________38290, _________38291;
  wire _________38292, _________38293, _________38296, _________38297,
       _________38298, _________38299, _________38300, _________38301;
  wire _________38302, _________38303, _________38306, _________38307,
       _________38308, _________38309, _________38310, _________38311;
  wire _________38312, _________38313, _________38335, _________38336,
       _________38337, _________38338, _________38339, _________38340;
  wire _________38341, _________38344, _________38345, _________38346,
       _________38347, _________38348, _________38349, _________38350;
  wire _________38353, _________38354, _________38355, _________38356,
       _________38357, _________38358, _________38359, _________38360;
  wire _________38363, _________38364, _________38365, _________38366,
       _________38367, _________38368, _________38369, _________38372;
  wire _________38373, _________38374, _________38375, _________38376,
       _________38377, _________38378, _________38379, _________38382;
  wire _________38383, _________38384, _________38385, _________38386,
       _________38387, _________38388, _________38389, _________38392;
  wire _________38393, _________38394, _________38395, _________38396,
       _________38397, _________38398, _________38399, _________38402;
  wire _________38403, _________38404, _________38405, _________38406,
       _________38407, _________38429, _________38430, _________38431;
  wire _________38432, _________38433, _________38434, _________38435,
       _________38436, _________38439, _________38440, _________38441;
  wire _________38442, _________38443, _________38444, _________38445,
       _________38446, _________38449, _________38450, _________38451;
  wire _________38452, _________38453, _________38454, _________38455,
       _________38456, _________38459, _________38460, _________38461;
  wire _________38462, _________38463, _________38464, _________38465,
       _________38468, _________38469, _________38470, _________38471;
  wire _________38472, _________38473, _________38474, _________38475,
       _________38478, _________38479, _________38480, _________38481;
  wire _________38482, _________38483, _________38484, _________38485,
       _________38488, _________38489, _________38490, _________38491;
  wire _________38492, _________38493, _________38494, _________38495,
       _________38498, _________38499, _________38500, _________38501;
  wire _________38502, _________38503, _________38504, _________38505,
       _________38528, _________38529, _________38530, _________38531;
  wire _________38532, _________38533, _________38534, _________38535,
       _________38538, _________38539, _________38540, _________38541;
  wire _________38542, _________38543, _________38544, _________38547,
       _________38548, _________38549, _________38550, _________38551;
  wire _________38552, _________38553, _________38556, _________38557,
       _________38558, _________38559, _________38560, _________38561;
  wire _________38562, _________38563, _________38566, _________38567,
       _________38568, _________38569, _________38570, _________38571;
  wire _________38572, _________38573, _________38576, _________38577,
       _________38578, _________38579, _________38580, _________38581;
  wire _________38582, _________38583, _________38586, _________38587,
       _________38588, _________38589, _________38590, _________38591;
  wire _________38592, _________38595, _________38596, _________38597,
       _________38598, _________38599, _________38600, _________38601;
  wire _________38623, _________38624, _________38625, _________38626,
       _________38627, _________38628, _________38629, _________38632;
  wire _________38633, _________38634, _________38635, _________38636,
       _________38637, _________38638, _________38641, _________38642;
  wire _________38643, _________38644, _________38645, _________38646,
       _________38649, _________38650, _________38651, _________38652;
  wire _________38653, _________38654, _________38657, _________38658,
       _________38659, _________38660, _________38661, _________38662;
  wire _________38663, _________38665, _________38666, _________38667,
       _________38668, _________38669, _________38670, _________38671;
  wire _________38674, _________38675, _________38676, _________38677,
       _________38678, _________38679, _________38680, _________38681;
  wire _________38684, _________38685, _________38686, _________38687,
       _________38688, _________38689, _________38690, _________38691;
  wire _________38712, _________38713, _________38714, _________38715,
       _________38716, _________38717, _________38718, _________38719;
  wire _________38722, _________38723, _________38724, _________38725,
       _________38726, _________38727, _________38728, _________38729;
  wire _________38732, _________38733, _________38734, _________38735,
       _________38736, _________38737, _________38738, _________38741;
  wire _________38742, _________38743, _________38744, _________38745,
       _________38746, _________38747, _________38748, _________38751;
  wire _________38752, _________38753, _________38754, _________38755,
       _________38756, _________38757, _________38758, _________38761;
  wire _________38762, _________38763, _________38764, _________38765,
       _________38766, _________38767, _________38768, _________38771;
  wire _________38772, _________38773, _________38774, _________38775,
       _________38776, _________38777, _________38778, _________38781;
  wire _________38782, _________38783, _________38784, _________38785,
       _________38786, _________38787, _________38788, _________38811;
  wire _________38812, _________38813, _________38814, _________38815,
       _________38816, _________38817, _________38818, _________38821;
  wire _________38822, _________38823, _________38824, _________38825,
       _________38828, _________38829, _________38830, _________38831;
  wire _________38832, _________38833, _________38834, _________38835,
       _________38838, _________38839, _________38840, _________38841;
  wire _________38842, _________38843, _________38846, _________38847,
       _________38848, _________38849, _________38850, _________38851;
  wire _________38852, _________38853, _________38856, _________38857,
       _________38858, _________38859, _________38860, _________38861;
  wire _________38862, _________38863, _________38866, _________38867,
       _________38868, _________38869, _________38870, _________38871;
  wire _________38872, _________38874, _________38875, _________38876,
       _________38877, _________38878, _________40656, _________40831;
  wire _________40832, _________40833, _________40834, _________40835,
       _________40836, _________40837, _________40838, _________40841;
  wire _________40842, _________40843, _________40844, _________40845,
       _________40846, _________40847, _________40848, _________40851;
  wire _________40852, _________40853, _________40854, _________40855,
       _________40856, _________40857, _________40858, _________40861;
  wire _________40862, _________40863, _________40864, _________40865,
       _________40866, _________40867, _________40868, _________40869;
  wire _________40870, _________40871, _________40872, _________40873,
       _________40874, _________40875, _________40876, _________40877;
  wire _________40878, _________40879, _________40880, _________40881,
       _________40882, _________40885, _________40886, _________40887;
  wire _________40888, _________40889, _________40890, _________40891,
       _________40892, _________40895, _________40896, _________40897;
  wire _________40898, _________40899, _________40900, _________40901,
       _________40902, _________40925, _________40926, _________40927;
  wire _________40928, _________40929, _________40930, _________40931,
       _________40932, _________40935, _________40936, _________40937;
  wire _________40938, _________40939, _________40940, _________40941,
       _________40942, _________40945, _________40946, _________40947;
  wire _________40948, _________40949, _________40950, _________40951,
       _________40954, _________40955, _________40956, _________40957;
  wire _________40958, _________40959, _________40960, _________40961,
       _________40964, _________40965, _________40966, _________40967;
  wire _________40968, _________40969, _________40970, _________40971,
       _________40974, _________40975, _________40976, _________40977;
  wire _________40978, _________40979, _________40980, _________40981,
       _________40984, _________40985, _________40986, _________40987;
  wire _________40988, _________40989, _________40990, _________40993,
       _________40994, _________40995, _________40996, _________40997;
  wire _________40998, _________40999, _________41000, _________41023,
       _________41024, _________41025, _________41026, _________41027;
  wire _________41028, _________41029, _________41030, _________41033,
       _________41034, _________41035, _________41036, _________41037;
  wire _________41038, _________41039, _________41040, _________41043,
       _________41044, _________41045, _________41046, _________41047;
  wire _________41048, _________41049, _________41050, _________41053,
       _________41054, _________41055, _________41056, _________41057;
  wire _________41058, _________41059, _________41060, _________41063,
       _________41064, _________41065, _________41066, _________41067;
  wire _________41068, _________41069, _________41070, _________41073,
       _________41074, _________41075, _________41076, _________41077;
  wire _________41078, _________41079, _________41080, _________41083,
       _________41084, _________41085, _________41086, _________41087;
  wire _________41088, _________41089, _________41090, _________41093,
       _________41094, _________41095, _________41096, _________41097;
  wire _________41098, _________41121, _________41122, _________41123,
       _________41124, _________41125, _________41126, _________41127;
  wire _________41128, _________41131, _________41132, _________41133,
       _________41134, _________41135, _________41136, _________41137;
  wire _________41138, _________41141, _________41142, _________41143,
       _________41144, _________41145, _________41146, _________41147;
  wire _________41148, _________41151, _________41152, _________41153,
       _________41154, _________41155, _________41156, _________41157;
  wire _________41158, _________41161, _________41162, _________41163,
       _________41164, _________41165, _________41166, _________41167;
  wire _________41168, _________41171, _________41172, _________41173,
       _________41174, _________41175, _________41176, _________41177;
  wire _________41178, _________41181, _________41182, _________41183,
       _________41184, _________41185, _________41186, _________41187;
  wire _________41188, _________41191, _________41192, _________41193,
       _________41194, _________41195, _________41196, _________41197;
  wire _________41198, _________41221, _________41222, _________41223,
       _________41224, _________41225, _________41226, _________41227;
  wire _________41228, _________41231, _________41232, _________41233,
       _________41234, _________41235, _________41236, _________41237;
  wire _________41238, _________41241, _________41242, _________41243,
       _________41244, _________41245, _________41246, _________41247;
  wire _________41248, _________41251, _________41252, _________41253,
       _________41254, _________41255, _________41256, _________41257;
  wire _________41258, _________41261, _________41262, _________41263,
       _________41264, _________41265, _________41266, _________41267;
  wire _________41268, _________41271, _________41272, _________41273,
       _________41274, _________41275, _________41276, _________41277;
  wire _________41280, _________41281, _________41282, _________41283,
       _________41284, _________41285, _________41286, _________41287;
  wire _________41290, _________41291, _________41292, _________41293,
       _________41294, _________41295, _________41296, _________41297;
  wire _________41320, _________41321, _________41322, _________41323,
       _________41324, _________41325, _________41326, _________41327;
  wire _________41330, _________41331, _________41332, _________41333,
       _________41334, _________41335, _________41336, _________41337;
  wire _________41340, _________41341, _________41342, _________41343,
       _________41344, _________41345, _________41346, _________41347;
  wire _________41350, _________41351, _________41352, _________41353,
       _________41354, _________41355, _________41356, _________41357;
  wire _________41360, _________41361, _________41362, _________41363,
       _________41364, _________41365, _________41367, _________41372;
  wire __________, __________0_, __________9_, __________9___22107,
       __________22059, __________22060, __________22061,
       __________22062;
  wire __________22063, ___________, ___________9___22071,
       ____________, ____________22078, _____________22079,
       _____________22080, _____________22081;
  wire _____________22082, _____________22083, _____________22084,
       _____________22085, _____________22086, _____________22087,
       _____________22088, _____________22097;
  wire _____________22098, _____________22099, _____________22100,
       _____________22101, _____________22102, ______________22064,
       ______________22065, ______________22066;
  wire ______________22067, ______________22068, ______________22103,
       ______________22104, ______________22105, ______________22106,
       ______________22108, ______________22109;
  wire ______________22110, ______________22111, ______________22112,
       _______________0, _______________22069, _______________22070,
       _______________22072, _______________22073;
  wire _______________22074, _______________22075,
       _______________22076, _______________22077, _________________0_,
       _________________0___21676, _________________0___21687,
       _________________0___21702;
  wire _________________0___21728, _________________0___21740,
       _________________9_, _________________9___21685,
       _________________9___21696, _________________9___21711,
       _________________9___21737, _________________9___21749;
  wire __________________0_, __________________0___21686,
       __________________0___21697, __________________0___21712,
       __________________0___21738, __________________0___21750,
       ___________________, ____________________;
  wire _____________________21669, _____________________21670,
       _____________________21671, _____________________21672,
       _____________________21673, _____________________21674,
       _____________________21675, _____________________21677;
  wire _____________________21678, _____________________21679,
       _____________________21680, _____________________21681,
       _____________________21682, _____________________21683,
       _____________________21684, _____________________21688;
  wire _____________________21689, _____________________21690,
       _____________________21691, _____________________21692,
       _____________________21693, _____________________21694,
       _____________________21695, _____________________21703;
  wire _____________________21704, _____________________21705,
       _____________________21706, _____________________21707,
       _____________________21708, _____________________21709,
       _____________________21710, _____________________21729;
  wire _____________________21730, _____________________21731,
       _____________________21732, _____________________21733,
       _____________________21734, _____________________21735,
       _____________________21736, _____________________21741;
  wire _____________________21742, _____________________21743,
       _____________________21744, _____________________21745,
       _____________________21746, _____________________21747,
       _____________________21748, ______________________21698;
  wire ______________________21699, ______________________21700,
       ______________________21701, ______________________21739,
       ______________________21751, ______________________21752,
       ______________________21753,
       __________________________________9__________;
  wire _____________________________________0___0_,
       _____________________________________0___0___21760,
       _____________________________________0____,
       _____________________________________0_____,
       _____________________________________0______21754,
       _____________________________________0______21755,
       _____________________________________0______21756,
       _____________________________________0______21757;
  wire _____________________________________0_______21758,
       _____________________________________0_______21759,
       _____________________________________9___0_,
       _____________________________________9___0___21880,
       _____________________________________9____,
       _____________________________________9_____,
       _____________________________________9______21876,
       _____________________________________9______21877;
  wire _____________________________________9_______21878,
       _____________________________________9_______21879,
       _____________________________________9_______21881,
       _____________________________________9_______21882,
       _____________________________________9_______21883,
       _____________________________________9_______21884,
       ______________________________________0__0_,
       ______________________________________0___0_;
  wire ______________________________________0___9_,
       ______________________________________0____,
       ______________________________________0_____,
       ______________________________________0______21885,
       ______________________________________0______21886,
       ______________________________________0______21887,
       ______________________________________0_______21888,
       ______________________________________0_______21889;
  wire ______________________________________0_______21890,
       ______________________________________0_______21891,
       ______________________________________0_______21892,
       ______________________________________0_______21893,
       ______________________________________0_______21894,
       ________________________________________0_,
       ________________________________________0___21771,
       ________________________________________0___21788;
  wire ________________________________________0___21816,
       ________________________________________0___21829,
       ________________________________________0___21863,
       ________________________________________9_,
       _________________________________________0_,
       _________________________________________0___21786,
       _________________________________________0___21794,
       _________________________________________0___21798;
  wire _________________________________________0___21814,
       _________________________________________0___21821,
       _________________________________________0___21824,
       _________________________________________0___21840,
       _________________________________________0___21856,
       _________________________________________0___21862,
       _________________________________________0___21895,
       _________________________________________0___21939;
  wire _________________________________________0___21952,
       _________________________________________0___21968,
       _________________________________________9_,
       _________________________________________9___21779,
       _________________________________________9___21803,
       _________________________________________9___21855,
       _________________________________________9___21861,
       _________________________________________9___21874;
  wire _________________________________________9___21901,
       _________________________________________9___21929,
       _________________________________________9___21943,
       __________________________________________,
       __________________________________________0_,
       __________________________________________0___21919,
       __________________________________________0___21935,
       __________________________________________0___21944;
  wire __________________________________________0___21959,
       __________________________________________0___21981,
       __________________________________________9_,
       __________________________________________9___21918,
       __________________________________________9___21923,
       __________________________________________9___21934,
       __________________________________________9___21947,
       __________________________________________9___21951;
  wire __________________________________________9___21966,
       __________________________________________9___21977,
       ___________________________________________,
       ____________________________________________,
       ____________________________________________21761,
       ____________________________________________21762,
       ____________________________________________21763,
       ____________________________________________21764;
  wire ____________________________________________21772,
       ____________________________________________21773,
       ____________________________________________21774,
       ____________________________________________21789,
       ____________________________________________21790,
       ____________________________________________21791,
       ____________________________________________21792,
       ____________________________________________21793;
  wire ____________________________________________21804,
       ____________________________________________21805,
       ____________________________________________21806,
       ____________________________________________21807,
       ____________________________________________21817,
       ____________________________________________21818,
       ____________________________________________21819,
       ____________________________________________21820;
  wire ____________________________________________21830,
       ____________________________________________21831,
       ____________________________________________21832,
       ____________________________________________21833,
       ____________________________________________21834,
       ____________________________________________21846,
       ____________________________________________21847,
       ____________________________________________21848;
  wire ____________________________________________21849,
       ____________________________________________21850,
       ____________________________________________21851,
       ____________________________________________21864,
       ____________________________________________21865,
       ____________________________________________21866,
       ____________________________________________21867,
       ____________________________________________21868;
  wire _____________________________________________21765,
       _____________________________________________21766,
       _____________________________________________21767,
       _____________________________________________21768,
       _____________________________________________21769,
       _____________________________________________21770,
       _____________________________________________21775,
       _____________________________________________21776;
  wire _____________________________________________21777,
       _____________________________________________21778,
       _____________________________________________21780,
       _____________________________________________21781,
       _____________________________________________21782,
       _____________________________________________21783,
       _____________________________________________21784,
       _____________________________________________21785;
  wire _____________________________________________21787,
       _____________________________________________21795,
       _____________________________________________21796,
       _____________________________________________21797,
       _____________________________________________21799,
       _____________________________________________21800,
       _____________________________________________21801,
       _____________________________________________21802;
  wire _____________________________________________21808,
       _____________________________________________21809,
       _____________________________________________21810,
       _____________________________________________21811,
       _____________________________________________21812,
       _____________________________________________21813,
       _____________________________________________21815,
       _____________________________________________21822;
  wire _____________________________________________21823,
       _____________________________________________21825,
       _____________________________________________21826,
       _____________________________________________21827,
       _____________________________________________21828,
       _____________________________________________21835,
       _____________________________________________21836,
       _____________________________________________21837;
  wire _____________________________________________21838,
       _____________________________________________21839,
       _____________________________________________21841,
       _____________________________________________21842,
       _____________________________________________21843,
       _____________________________________________21844,
       _____________________________________________21845,
       _____________________________________________21852;
  wire _____________________________________________21853,
       _____________________________________________21854,
       _____________________________________________21857,
       _____________________________________________21858,
       _____________________________________________21859,
       _____________________________________________21860,
       _____________________________________________21869,
       _____________________________________________21870;
  wire _____________________________________________21871,
       _____________________________________________21872,
       _____________________________________________21873,
       _____________________________________________21875,
       _____________________________________________21896,
       _____________________________________________21897,
       _____________________________________________21898,
       _____________________________________________21899;
  wire _____________________________________________21900,
       _____________________________________________21907,
       _____________________________________________21908,
       _____________________________________________21909,
       _____________________________________________21910,
       _____________________________________________21924,
       _____________________________________________21925,
       _____________________________________________21926;
  wire _____________________________________________21927,
       _____________________________________________21928,
       _____________________________________________21940,
       _____________________________________________21941,
       _____________________________________________21942,
       _____________________________________________21953,
       _____________________________________________21954,
       _____________________________________________21969;
  wire _____________________________________________21970,
       _____________________________________________21971,
       _____________________________________________21972,
       _____________________________________________21973,
       _____________________________________________21974,
       ______________________________________________21902,
       ______________________________________________21903,
       ______________________________________________21904;
  wire ______________________________________________21905,
       ______________________________________________21906,
       ______________________________________________21911,
       ______________________________________________21912,
       ______________________________________________21913,
       ______________________________________________21914,
       ______________________________________________21915,
       ______________________________________________21916;
  wire ______________________________________________21917,
       ______________________________________________21920,
       ______________________________________________21921,
       ______________________________________________21922,
       ______________________________________________21930,
       ______________________________________________21931,
       ______________________________________________21932,
       ______________________________________________21933;
  wire ______________________________________________21936,
       ______________________________________________21937,
       ______________________________________________21938,
       ______________________________________________21945,
       ______________________________________________21946,
       ______________________________________________21948,
       ______________________________________________21949,
       ______________________________________________21950;
  wire ______________________________________________21955,
       ______________________________________________21956,
       ______________________________________________21957,
       ______________________________________________21958,
       ______________________________________________21960,
       ______________________________________________21961,
       ______________________________________________21962,
       ______________________________________________21963;
  wire ______________________________________________21964,
       ______________________________________________21965,
       ______________________________________________21967,
       ______________________________________________21975,
       ______________________________________________21976,
       ______________________________________________21978,
       ______________________________________________21979,
       ______________________________________________21980;
  wire ______________________________________________21982,
       _______________________________________________________________,
       _______________________________________________________________0,
       _______________________________________________________________0__21998,
       _______________________________________________________________0__22006,
       _______________________________________________________________0__22010,
       _______________________________________________________________9,
       _______________________________________________________________9__21995;
  wire ________________________________________________________________,
       _________________________________________________________________21991,
       _________________________________________________________________22000,
       _________________________________________________________________22001,
       __________________________________________________________________21983,
       __________________________________________________________________21984,
       __________________________________________________________________21985,
       __________________________________________________________________21986;
  wire __________________________________________________________________21987,
       __________________________________________________________________21988,
       __________________________________________________________________21989,
       __________________________________________________________________21990,
       __________________________________________________________________21992,
       __________________________________________________________________21993,
       __________________________________________________________________21994,
       __________________________________________________________________21996;
  wire __________________________________________________________________21997,
       __________________________________________________________________21999,
       __________________________________________________________________22002,
       __________________________________________________________________22003,
       __________________________________________________________________22004,
       __________________________________________________________________22005,
       __________________________________________________________________22007,
       __________________________________________________________________22008;
  wire __________________________________________________________________22009,
       __________________________________________________________________22011,
       __________________________________________________________________22012,
       ______________________________________________________________________________________0,
       ______________________________________________________________________________________0__22093,
       ______________________________________________________________________________________0__22096,
       _______________________________________________________________________________________,
       _________________________________________________________________________________________22089;
  wire _________________________________________________________________________________________22090,
       _________________________________________________________________________________________22091,
       _________________________________________________________________________________________22092,
       _________________________________________________________________________________________22094,
       _________________________________________________________________________________________22095;
  dffacs1 ________________________________________________(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40410), .Q
       (______________________________________________21982));
  nnd2s1 ____0_______0(.DIN1 (___0_____40409), .DIN2 (___0__0__40403),
       .Q (___0_____40410));
  nnd2s1 ____0______9_(.DIN1 (___0_____40407), .DIN2 (___0_____40400),
       .Q (___0_____40409));
  dffacs1 ________________________________________________495156(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40408), .Q (___0_____40414));
  dffacs1 ______________________________________________0_(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40406), .Q
       (__________________________________________0___21981));
  dffacs1 _______________________________________(.CLRB (reset), .CLK
       (clk), .DIN (___0_____40405), .QN (___0_____40447));
  nnd2s1 ____0_0______(.DIN1 (___0__9__40402), .DIN2 (___0_9___40358),
       .Q (___0_____40408));
  xor2s1 ____0________(.DIN1 (___0_____40398), .DIN2 (___00____39971),
       .Q (___0_____40407));
  nnd2s1 ____0_9______(.DIN1 (___0_____40401), .DIN2 (__90____29694),
       .Q (___0_____40406));
  dffacs1 ______________________________________________9_(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40404), .Q (___0_____40607));
  nnd2s1 ____0____9___(.DIN1 (___0_____40399), .DIN2 (___0__9__40392),
       .Q (___0_____40405));
  nnd2s1 ____0________495157(.DIN1 (___0_____40397), .DIN2
       (___0_____40376), .Q (___0_____40404));
  nnd2s1 ____0______09(.DIN1 (___0_____40386), .DIN2 (___0_____40394),
       .Q (___0__0__40403));
  nor2s1 ____0________495158(.DIN1 (___0_____40395), .DIN2
       (___0_9___40355), .Q (___0__9__40402));
  nnd2s1 ____0_____900(.DIN1 (___0_____40396), .DIN2 (___0_____40400),
       .Q (___0_____40401));
  dffacs1 ________________________________________________495159(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40391), .Q
       (______________________________________________21980));
  dffacs1 _______________________________________495160(.CLRB (reset),
       .CLK (clk), .DIN (___0__0__40393), .QN (___0_____40448));
  nor2s1 ____0_9____9_(.DIN1 (______9__38730), .DIN2 (___0_____40388),
       .Q (___0_____40399));
  nor2s1 ____0________495161(.DIN1 (___00____39937), .DIN2
       (___0_____40390), .Q (___0_____40398));
  nor2s1 ____0_0______495162(.DIN1 (________29138), .DIN2
       (___0_____40384), .Q (___0_____40397));
  xor2s1 ____0________495163(.DIN1 (___00____39938), .DIN2
       (___0_____40389), .Q (___0_____40396));
  nor2s1 ____0________495164(.DIN1 (___0_____40385), .DIN2
       (___0_9___40354), .Q (___0_____40395));
  xor2s1 ____0_____9__(.DIN1 (_________22031), .DIN2 (________23117),
       .Q (___0_____40394));
  nnd2s1 ____0______0_(.DIN1 (___0__0__40383), .DIN2 (___0__9__40392),
       .Q (___0__0__40393));
  nnd2s1 ____0________495165(.DIN1 (___0_9___40360), .DIN2
       (___0_____40387), .Q (___0_____40391));
  nor2s1 ____0________495166(.DIN1 (___00____39936), .DIN2
       (___0_____40389), .Q (___0_____40390));
  nor2s1 ____0_0_____0(.DIN1 (_________22031), .DIN2 (___0_____40380),
       .Q (___0_____40388));
  nnd2s1 ____0_____0__(.DIN1 (___0_____40386), .DIN2 (___0_____40379),
       .Q (___0_____40387));
  nor2s1 ____0_9____0_(.DIN1 (____9____38963), .DIN2 (___0_____40378),
       .Q (___0_____40385));
  and2s1 ____0______9_495167(.DIN1 (___0__9__40382), .DIN2
       (___0_____40400), .Q (___0_____40384));
  nor2s1 ____0________495168(.DIN1 (_____9__26399), .DIN2
       (___0_____40381), .Q (___0__0__40383));
  dffacs1 ________________________________________________495169(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40377), .QN
       (_________22031));
  nor2s1 ____0_______495170(.DIN1 (___00____39919), .DIN2
       (___0_____40375), .Q (___0_____40389));
  xor2s1 ____0_____0_9(.DIN1 (___00____39920), .DIN2 (___0_____40374),
       .Q (___0__9__40382));
  nor2s1 ____0_9______495171(.DIN1 (___0__0__40373), .DIN2
       (___0_____40380), .Q (___0_____40381));
  xor2s1 ____0____990_(.DIN1 (_______22237), .DIN2 (___0_____40604), .Q
       (___0_____40379));
  xor2s1 ____0_______495172(.DIN1
       (______________________________________________21979), .DIN2
       (___0_____40604), .Q (___0_____40378));
  nnd2s1 ____0______9_495173(.DIN1 (___0_09__40372), .DIN2
       (___0_____40376), .Q (___0_____40377));
  and2s1 ____0_0______495174(.DIN1 (___0_____40374), .DIN2
       (___00____39907), .Q (___0_____40375));
  hi1s1 ____0__(.DIN (___0_____40604), .Q (___0__0__40373));
  dffacs1 ________________________________________________495175(.CLRB
       (reset), .CLK (clk), .DIN (___0_0___40371), .Q (___0_____40604));
  nor2s1 ____0________495176(.DIN1 (________29128), .DIN2
       (___0_0___40370), .Q (___0_09__40372));
  xor2s1 ____0________495177(.DIN1 (___0_0___40369), .DIN2
       (_________37547), .Q (___0_____40374));
  nnd2s1 ____0____9___495178(.DIN1 (___0_0___40368), .DIN2
       (___0_____40376), .Q (___0_0___40371));
  and2s1 ____0________495179(.DIN1 (___0_0___40367), .DIN2
       (___0_____40400), .Q (___0_0___40370));
  nnd2s1 ____0______495180(.DIN1 (___0_0___40366), .DIN2
       (___0_____40103), .Q (___0_0___40369));
  nor2s1 ____0________495181(.DIN1 (_____0__29146), .DIN2
       (___0_0___40364), .Q (___0_0___40368));
  xor2s1 ____0_9___900(.DIN1 (___0_____40111), .DIN2 (___0_0___40365),
       .Q (___0_0___40367));
  nnd2s1 ____0_0____9_(.DIN1 (___0_0___40365), .DIN2 (___0_____40102),
       .Q (___0_0___40366));
  and2s1 ____0________495182(.DIN1 (___0_00__40363), .DIN2
       (___0_____40400), .Q (___0_0___40364));
  nor2s1 ____0________495183(.DIN1 (___0__0__40119), .DIN2
       (___0_99__40362), .Q (___0_0___40365));
  xor2s1 ____0________495184(.DIN1 (___0_____40120), .DIN2
       (___0_9___40361), .Q (___0_00__40363));
  nor2s1 ____0________495185(.DIN1 (___0__9__40118), .DIN2
       (___0_9___40361), .Q (___0_99__40362));
  dffacs1 ________________________________________________495186(.CLRB
       (reset), .CLK (clk), .DIN (___0_9___40359), .Q (___0_____40415));
  nnd2s1 ____0_____9__495187(.DIN1 (___0_9___40356), .DIN2
       (___0_____40400), .Q (___0_9___40360));
  dffacs1 ________________________________________________495188(.CLRB
       (reset), .CLK (clk), .DIN (___0_9___40357), .Q
       (______________________________________________21979));
  nnd2s1 ____0______0_495189(.DIN1 (___0_90__40353), .DIN2
       (___0_9___40358), .Q (___0_9___40359));
  nnd2s1 ____09_______(.DIN1 (___0__9__40352), .DIN2 (___0_9___40077),
       .Q (___0_9___40361));
  nnd2s1 ____0_9______495190(.DIN1 (___0_____40350), .DIN2
       (___9____29614), .Q (___0_9___40357));
  xor2s1 ____09______0(.DIN1 (___0_0___40086), .DIN2 (___0_____40351),
       .Q (___0_9___40356));
  and2s1 ____090___0__(.DIN1 (___0_____40349), .DIN2 (___0_9___40354),
       .Q (___0_9___40355));
  and2s1 ____09_____0_(.DIN1 (___0_____40348), .DIN2 (___0_____40347),
       .Q (___0_90__40353));
  nnd2s1 ____09_____9_(.DIN1 (___0_____40351), .DIN2 (___0_00__40079),
       .Q (___0__9__40352));
  nnd2s1 ____09_______495191(.DIN1 (___0_____40345), .DIN2
       (___0_9___40354), .Q (___0_____40350));
  dffacs1 _______________________________________495192(.CLRB (reset),
       .CLK (clk), .DIN (___0_____40346), .QN (______________22109));
  xor2s1 ____09______495193(.DIN1 (___0_____40339), .DIN2
       (___909___39065), .Q (___0_____40349));
  nor2s1 _____00___0_9(.DIN1 (___0_____40344), .DIN2 (___0_____40327),
       .Q (___0_____40348));
  nnd2s1 ____099______(.DIN1 (___0__0__40343), .DIN2 (___9_____39764),
       .Q (___0_____40351));
  nnd2s1 ____09___990_(.DIN1 (___0_____40326), .DIN2 (___0_____40341),
       .Q (___0_____40347));
  nnd2s1 _____0______0(.DIN1 (___09___26133), .DIN2 (___0_____40340),
       .Q (___0_____40346));
  xor2s1 _____0_____9_(.DIN1 (___0__9__40342), .DIN2 (___990___39805),
       .Q (___0_____40345));
  nor2s1 _____0_______(.DIN1 (___0_____40338), .DIN2 (___0_____40320),
       .Q (___0_____40344));
  nnd2s1 _____0_______495194(.DIN1 (___0__9__40342), .DIN2
       (___9_____39765), .Q (___0__0__40343));
  nor2s1 _____0_______495195(.DIN1
       (______________________________________________21978), .DIN2
       (________28146), .Q (___0_____40341));
  nnd2s1 _____0___9___(.DIN1 (_________32712), .DIN2
       (______________________________________________21978), .Q
       (___0_____40340));
  xor2s1 _____0_______495196(.DIN1 (___0_____40337), .DIN2
       (___0__0__40333), .Q (___0_____40339));
  hi1s1 _____0_(.DIN
       (______________________________________________21978), .Q
       (___0_____40338));
  nnd2s1 ______0____09(.DIN1 (___0_____40335), .DIN2 (___0_____40336),
       .Q (___0__9__40342));
  dffacs1 ________________________________________________495197(.CLRB
       (reset), .CLK (clk), .DIN (___0__9__40332), .Q
       (______________________________________________21978));
  and2s1 _____________(.DIN1 (___0_____40336), .DIN2 (___0_____40334),
       .Q (___0_____40337));
  nnd2s1 __________900(.DIN1 (___0_____40334), .DIN2 (___0__0__40333),
       .Q (___0_____40335));
  nnd2s1 ___________9_(.DIN1 (___0_____40330), .DIN2 (__9_____30213),
       .Q (___0__9__40332));
  or2s1 _____________495198(.DIN1
       (______________________________________________21963), .DIN2
       (___0_____40331), .Q (___0_____40336));
  nnd2s1 _____________495199(.DIN1 (___0_____40331), .DIN2
       (______________________________________________21963), .Q
       (___0_____40334));
  nnd2s1 _____________495200(.DIN1 (___0_____40329), .DIN2
       (___0_9___40354), .Q (___0_____40330));
  nnd2s1 _____________495201(.DIN1 (___0_____40328), .DIN2
       (___0_____40036), .Q (___0_____40331));
  xor2s1 __________9__(.DIN1 (___0__0__40039), .DIN2 (___09____40692),
       .Q (___0_____40329));
  nnd2s1 ______9____0_(.DIN1 (___09____40692), .DIN2 (___0_____40037),
       .Q (___0_____40328));
  dffacs1 ______________________________________________0_495202(.CLRB
       (reset), .CLK (clk), .DIN (___0__0__40325), .Q (______9__22030));
  nor2s1 ____________0(.DIN1 (___0_____40326), .DIN2 (___0_____40322),
       .Q (___0_____40327));
  nnd2s1 __________0__(.DIN1 (___0_____40321), .DIN2 (___0_9___40358),
       .Q (___0__0__40325));
  xor2s1 _____________495203(.DIN1 (___9_____39547), .DIN2
       (___09____40694), .Q (___0_____40322));
  dffacs1 ________________________________________________495204(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40319), .Q (___0_____40602));
  and2s1 ____________495205(.DIN1 (___0__9__40317), .DIN2
       (___0_____40320), .Q (___0_____40321));
  nor2s1 __________0_9(.DIN1 (___9_____39514), .DIN2 (___09____40694),
       .Q (___0_____40324));
  dffacs1 ______________________________________________9_495206(.CLRB
       (reset), .CLK (clk), .DIN (___0__0__40318), .Q
       (__________________________________________9___21977));
  nnd2s1 _____________495207(.DIN1 (___0_____40315), .DIN2
       (___0_9___40358), .Q (___0_____40319));
  dffacs1 ________________________________________________495208(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40316), .Q (_________22029));
  nnd2s1 ______9__990_(.DIN1 (___0_____40285), .DIN2 (___0_____40314),
       .Q (___0__0__40318));
  and2s1 ____________495209(.DIN1 (___0_____40313), .DIN2
       (____9___29276), .Q (___0__9__40317));
  nnd2s1 _____________495210(.DIN1 (___0_____40312), .DIN2
       (___0_0___40281), .Q (___0_____40316));
  and2s1 _____________495211(.DIN1 (___0_____40311), .DIN2
       (____9___28548), .Q (___0_____40315));
  nnd2s1 _____________495212(.DIN1 (___0_____40310), .DIN2
       (inData[18]), .Q (___0_____40314));
  nnd2s1 _________9___(.DIN1 (___0__0__40309), .DIN2 (___0_9___40354),
       .Q (___0_____40313));
  nor2s1 ___________09(.DIN1 (___0_____40306), .DIN2 (___0_____40251),
       .Q (___0_____40312));
  nnd2s1 _____________495213(.DIN1 (___0_____40305), .DIN2
       (___0_9___40354), .Q (___0_____40311));
  nor2s1 ______0___900(.DIN1 (___0_____40304), .DIN2 (___0_____40294),
       .Q (___0_____40310));
  xor2s1 ___________9_495214(.DIN1 (___0__0__40301), .DIN2
       (___9_0___39166), .Q (___0__0__40309));
  nor2s1 _____________495215(.DIN1 (___0_____40302), .DIN2
       (___0_____40284), .Q (___0_____40306));
  xor2s1 _____________495216(.DIN1 (___9_____39458), .DIN2
       (___0_____40303), .Q (___0_____40305));
  xor2s1 __________9__495217(.DIN1 (___0_____40296), .DIN2
       (_______22233), .Q (___0_____40304));
  nor2s1 ___________0_(.DIN1 (___9_____39457), .DIN2 (___0_____40303),
       .Q (___0_____40307));
  dffacs1 ________________________________________________495218(.CLRB
       (reset), .CLK (clk), .DIN (___0__9__40300), .Q
       (______________________________________________21976));
  dffacs1 _______________________________________495219(.CLRB (reset),
       .CLK (clk), .DIN (___0_____40299), .QN (___0_90__40451));
  nor2s1 _____________495220(.DIN1 (___99____39814), .DIN2
       (___0_____40297), .Q (___0_____40302));
  xor2s1 _____________495221(.DIN1 (___0__9__40290), .DIN2
       (___0__0__40291), .Q (___0__0__40301));
  dffacs1 ________________________________________________495222(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40298), .Q (___0_____40416));
  nnd2s1 ____________495223(.DIN1 (___0_____40259), .DIN2
       (___0_____40295), .Q (___0__9__40300));
  nnd2s1 __________0__495224(.DIN1 (___0_0___30836), .DIN2
       (___0_____40293), .Q (___0_____40299));
  nor2s1 ___________0_495225(.DIN1 (___0_____40289), .DIN2
       (___0_____40292), .Q (___0_____40303));
  nnd2s1 ___________9_495226(.DIN1 (___0_____40288), .DIN2
       (___0__9__40232), .Q (___0_____40298));
  xor2s1 ______0______(.DIN1
       (______________________________________________21976), .DIN2
       (___0_____40600), .Q (___0_____40297));
  xor2s1 ____________495227(.DIN1 (_________22029), .DIN2
       (___0_____40600), .Q (___0_____40296));
  or2s1 __________0_495228(.DIN1 (___0_____40600), .DIN2
       (___0_____40294), .Q (___0_____40295));
  nnd2s1 _____________495229(.DIN1 (___0_9___40270), .DIN2
       (___0_____40600), .Q (___0_____40293));
  nor2s1 _________990_(.DIN1 (___0__0__40291), .DIN2 (___09____40658),
       .Q (___0_____40292));
  nor2s1 ____________495230(.DIN1 (___0_____40289), .DIN2
       (___09____40658), .Q (___0__9__40290));
  nor2s1 ___________9_495231(.DIN1 (___0_____40287), .DIN2
       (___0__9__40223), .Q (___0_____40288));
  dffacs1 ________________________________________________495232(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40286), .Q
       (______________________________________________21975));
  dffacs1 ________________________________________________495233(.CLRB
       (reset), .CLK (clk), .DIN (___0_09__40282), .Q (___0_____40600));
  nor2s1 _____________495234(.DIN1 (___0_0___40278), .DIN2
       (___0_____40188), .Q (___0_____40287));
  nor2s1 _____________495235(.DIN1
       (__________________________________________0___21959), .DIN2
       (___0__0__40283), .Q (___0_____40289));
  nnd2s1 _________9___495236(.DIN1 (___0_____40234), .DIN2
       (___0_0___40279), .Q (___0_____40286));
  dffacs1 _______________________________________495237(.CLRB (reset),
       .CLK (clk), .DIN (___0_0___40280), .QN (_________22016));
  dffacs1 _____________________0_(.CLRB (reset), .CLK (clk), .DIN
       (___0_0___40277), .Q (_________________0___21676));
  nnd2s1 ______9______(.DIN1 (___0_0___40275), .DIN2 (___0_____40284),
       .Q (___0_____40285));
  nnd2s1 ___________495238(.DIN1 (___0_0___40276), .DIN2
       (___0_0___40281), .Q (___0_09__40282));
  nnd2s1 _____________495239(.DIN1 (___0_9___40271), .DIN2
       (_____9__28452), .Q (___0_0___40280));
  nnd2s1 ______9___900(.DIN1 (___0_9___40269), .DIN2 (___990___39803),
       .Q (___0__0__40283));
  or2s1 ___________9_495240(.DIN1 (___0_00__40273), .DIN2
       (___0_____40294), .Q (___0_0___40279));
  nor2s1 _____________495241(.DIN1 (_____00__34847), .DIN2
       (___0_0___40274), .Q (___0_0___40278));
  or2s1 _____________495242(.DIN1 (________29152), .DIN2
       (___0_99__40272), .Q (___0_0___40277));
  nor2s1 _____________495243(.DIN1 (___0____27002), .DIN2
       (___0_9___40267), .Q (___0_0___40276));
  xor2s1 _____________495244(.DIN1 (___99____39813), .DIN2
       (___0_9___40268), .Q (___0_0___40275));
  xor2s1 ______0___9__(.DIN1 (___0_____40605), .DIN2 (___0__9__40608),
       .Q (___0_0___40274));
  xor2s1 ___________0_495245(.DIN1 (___0_____40605), .DIN2
       (___0__9__40242), .Q (___0_00__40273));
  nnd2s1 _____________495246(.DIN1 (___0_____31066), .DIN2
       (___0_9___40265), .Q (___0_99__40272));
  nnd2s1 _____________495247(.DIN1 (___0_9___40270), .DIN2
       (___0_9___40266), .Q (___0_9___40271));
  nnd2s1 _____9______0(.DIN1 (___0_9___40268), .DIN2 (___990___39804),
       .Q (___0_9___40269));
  and2s1 _____9____0__(.DIN1 (___0_9___40264), .DIN2 (___0_____40284),
       .Q (___0_9___40267));
  hi1s1 _____90(.DIN (___0_____40605), .Q (___0_9___40266));
  nnd2s1 _____9_____0_(.DIN1 (___0_90__40263), .DIN2 (_________31715),
       .Q (___0_9___40265));
  nor2s1 _____9_____9_(.DIN1 (___99____39881), .DIN2 (___0__9__40262),
       .Q (___0_9___40268));
  dffacs1 ________________________________________________495248(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40260), .QN
       (___0_____40605));
  xor2s1 _____9_______(.DIN1 (___99_9__39882), .DIN2 (___0_____40261),
       .Q (___0_9___40264));
  nnd2s1 _____9______495249(.DIN1 (___0_____40258), .DIN2
       (___0_____30684), .Q (___0_90__40263));
  and2s1 _____0____0_9(.DIN1 (___0_____40261), .DIN2 (___99____39865),
       .Q (___0__9__40262));
  nnd2s1 _____9_______495250(.DIN1 (___0_____40257), .DIN2
       (___0_0___40281), .Q (___0_____40260));
  nnd2s1 _____0___990_(.DIN1 (___0_____40256), .DIN2 (___0_____40284),
       .Q (___0_____40259));
  nor2s1 _____99_____0(.DIN1 (_____9___31789), .DIN2 (___0_____40255),
       .Q (___0_____40258));
  nor2s1 _____0_____9_495251(.DIN1 (___9_0___39163), .DIN2
       (___0_____40254), .Q (___0_____40261));
  nor2s1 _____00______(.DIN1 (___0__9__40252), .DIN2 (___0_____40241),
       .Q (___0_____40257));
  xor2s1 _____0_______495252(.DIN1 (___9_0___39169), .DIN2
       (___0__0__40253), .Q (___0_____40256));
  nnd2s1 _____0_______495253(.DIN1 (___0_____40250), .DIN2
       (________27660), .Q (___0_____40255));
  and2s1 _________9___495254(.DIN1 (___0__0__40253), .DIN2
       (___9_99__39161), .Q (___0_____40254));
  nor2s1 _____0_______495255(.DIN1 (___0_____40249), .DIN2
       (___0_____40284), .Q (___0__9__40252));
  and2s1 ______0____495256(.DIN1 (___0_____40248), .DIN2
       (___0_____40284), .Q (___0_____40251));
  nor2s1 _____0_______495257(.DIN1 (____9___25856), .DIN2
       (___0_____40247), .Q (___0_____40250));
  nor2s1 __________495258(.DIN1 (___9__9__39181), .DIN2
       (___0_____40245), .Q (___0__0__40253));
  dffacs1 _______________________________________495259(.CLRB (reset),
       .CLK (clk), .DIN (___0_____40246), .QN (_________22015));
  nor2s1 _____09____9_(.DIN1 (___9____25102), .DIN2 (___0__0__40243),
       .Q (___0_____40249));
  xor2s1 _____________495260(.DIN1 (___9__0__39182), .DIN2
       (___0_____40244), .Q (___0_____40248));
  nnd2s1 _____________495261(.DIN1 (_____0___35657), .DIN2
       (___0_____40240), .Q (___0_____40247));
  nnd2s1 _____________495262(.DIN1 (________28616), .DIN2
       (___0_____40239), .Q (___0_____40246));
  nor2s1 _____________495263(.DIN1 (___9_____39180), .DIN2
       (___0_____40244), .Q (___0_____40245));
  xnr2s1 __________9__495264(.DIN1 (___0__9__40608), .DIN2
       (___0_____40416), .Q (___0__0__40243));
  nnd2s1 ___________0_495265(.DIN1 (___0_____40238), .DIN2
       (______________________________________________21975), .Q
       (___0__9__40242));
  and2s1 ______0______495266(.DIN1 (___0_____40237), .DIN2
       (___0_____40284), .Q (___0_____40241));
  or2s1 _____________495267(.DIN1 (___0__9__40608), .DIN2
       (_________32260), .Q (___0_____40240));
  nnd2s1 ______9_____0(.DIN1 (________23538), .DIN2 (___0__9__40608),
       .Q (___0_____40239));
  nor2s1 __________0__495268(.DIN1 (____9____38936), .DIN2
       (___0_____40236), .Q (___0_____40244));
  hi1s1 _______(.DIN (___0__9__40608), .Q (___0_____40238));
  xor2s1 ___________0_495269(.DIN1 (___90____39011), .DIN2
       (___0_____40235), .Q (___0_____40237));
  dffacs1 ________________________________________________495270(.CLRB
       (reset), .CLK (clk), .DIN (___0__0__40233), .Q (___0__9__40608));
  and2s1 ___________9_495271(.DIN1 (___0_____40235), .DIN2
       (___90____39010), .Q (___0_____40236));
  nnd2s1 _____________495272(.DIN1 (___0_____40231), .DIN2
       (___0_____40284), .Q (___0_____40234));
  nnd2s1 ____________495273(.DIN1 (___0_____40230), .DIN2
       (___0__9__40232), .Q (___0__0__40233));
  nor2s1 __________0_495274(.DIN1 (_____9___38792), .DIN2
       (___0_____40229), .Q (___0_____40235));
  xor2s1 ______0______495275(.DIN1 (_________38866), .DIN2
       (___0_____40228), .Q (___0_____40231));
  nor2s1 ______9__990_495276(.DIN1 (________27358), .DIN2
       (___0_____40227), .Q (___0_____40230));
  nor2s1 ____________495277(.DIN1 (_____90__38790), .DIN2
       (___0_____40228), .Q (___0_____40229));
  nor2s1 ___________9_495278(.DIN1 (___0_____40222), .DIN2
       (___0_____40226), .Q (___0_____40227));
  nor2s1 _____________495279(.DIN1 (___0_____40225), .DIN2
       (___09____40696), .Q (___0_____40228));
  xor2s1 _____________495280(.DIN1 (___0_____40221), .DIN2
       (_________38395), .Q (___0_____40226));
  nor2s1 _____________495281(.DIN1 (___0__9__40158), .DIN2
       (___0_____40224), .Q (___0_____40225));
  nnd2s1 _________9___495282(.DIN1 (___0_____40220), .DIN2
       (___9_____39537), .Q (___0_____40224));
  nor2s1 ______9____09(.DIN1 (___0_____40222), .DIN2 (___0_____40218),
       .Q (___0__9__40223));
  xor2s1 ______0______495283(.DIN1 (___9__0__39561), .DIN2
       (___0_____40219), .Q (___0_____40221));
  nnd2s1 __________495284(.DIN1 (___099___40718), .DIN2
       (___0_____40219), .Q (___0_____40220));
  xor2s1 _____________495285(.DIN1 (___0_____40216), .DIN2
       (______________________________________________21955), .Q
       (___0_____40218));
  dffacs1 ________________________________________________495286(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40217), .Q (___0_____40611));
  nor2s1 _____________495287(.DIN1 (___0__0__40215), .DIN2
       (___0_____40213), .Q (___0_____40219));
  dffacs1 ______________________________________________0_495288(.CLRB
       (reset), .CLK (clk), .DIN (___0__9__40214), .QN
       (___0_____40417));
  nnd2s1 _____________495289(.DIN1 (___0_____40211), .DIN2
       (___0__9__40232), .Q (___0_____40217));
  nor2s1 _____________495290(.DIN1 (___0__0__40215), .DIN2
       (___0_____40212), .Q (___0_____40216));
  nnd2s1 __________9__495291(.DIN1 (___0_____40210), .DIN2
       (___0__9__40232), .Q (___0__9__40214));
  nor2s1 ______9____0_495292(.DIN1
       (______________________________________________21955), .DIN2
       (___0_____40212), .Q (___0_____40213));
  nor2s1 ______0______495293(.DIN1 (________27132), .DIN2
       (___0_____40209), .Q (___0_____40211));
  nor2s1 _____________495294(.DIN1 (___0_____40208), .DIN2
       (_________38578), .Q (___0__0__40215));
  nor2s1 ____________495295(.DIN1 (________27111), .DIN2
       (___0_____40207), .Q (___0_____40210));
  nor2s1 __________0__495296(.DIN1 (___09____40698), .DIN2
       (_____0___38523), .Q (___0_____40212));
  nor2s1 ___________0_495297(.DIN1 (___0_____40222), .DIN2
       (___0__0__40206), .Q (___0_____40209));
  hi1s1 _______495298(.DIN (___09____40698), .Q (___0_____40208));
  nor2s1 ___________9_495299(.DIN1 (___0_____40222), .DIN2
       (___0_____40204), .Q (___0_____40207));
  xor2s1 ____________495300(.DIN1 (___0_____40205), .DIN2
       (___9_____39666), .Q (___0__0__40206));
  xor2s1 _____________495301(.DIN1 (___0_____40203), .DIN2
       (_________36349), .Q (___0_____40204));
  xor2s1 _________990_495302(.DIN1 (___0_____40201), .DIN2
       (____9____37036), .Q (___0_____40205));
  xor2s1 ____________495303(.DIN1
       (__________________________________________________________________22009),
       .DIN2 (___0_____40199), .Q (___0_____40203));
  dffacs1 _______________________________________________(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40202), .Q
       (_____________________________________________21973));
  dffacs1 _____________________________________________9_(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40200), .Q (___0_____40418));
  nnd2s1 ___________9_495304(.DIN1 (___0_9___40170), .DIN2
       (___0__0__40197), .Q (___0_____40202));
  nor2s1 _____________495305(.DIN1 (___0_____40198), .DIN2
       (___0__9__40196), .Q (___0_____40201));
  nnd2s1 ______0______495306(.DIN1 (___0_____40195), .DIN2
       (___0__9__40232), .Q (___0_____40200));
  nor2s1 _____________495307(.DIN1 (___0_____40198), .DIN2
       (___0_____40194), .Q (___0_____40199));
  nnd2s1 _________9___495308(.DIN1 (___0_____40192), .DIN2
       (inData[14]), .Q (___0__0__40197));
  and2s1 _____________495309(.DIN1 (___0_____40193), .DIN2
       (__________________________________________________________________22009),
       .Q (___0__9__40196));
  nor2s1 ___________495310(.DIN1 (_____9__27112), .DIN2
       (___0_____40189), .Q (___0_____40195));
  hi1s1 _______495311(.DIN (___0_____40193), .Q (___0_____40194));
  nor2s1 ______9______495312(.DIN1 (___0__0__40187), .DIN2
       (___0_____40166), .Q (___0_____40192));
  nor2s1 __________495313(.DIN1 (___0_____40190), .DIN2
       (___0_____40191), .Q (___0_____40198));
  dffacs1 ______________________________________(.CLRB (reset), .CLK
       (clk), .DIN (___0_09__40186), .Q (___0_9___40453));
  nnd2s1 ___________9_495314(.DIN1 (___0_____40191), .DIN2
       (___0_____40190), .Q (___0_____40193));
  and2s1 ______9______495315(.DIN1 (___0_0___40185), .DIN2
       (___0_____40188), .Q (___0_____40189));
  xor2s1 _____________495316(.DIN1 (___0_0___40182), .DIN2
       (___0_____40160), .Q (___0__0__40187));
  nnd2s1 ______0______495317(.DIN1 (___0_90__40168), .DIN2
       (___0_0___40184), .Q (___0_09__40186));
  nor2s1 _____________495318(.DIN1 (_________37876), .DIN2
       (___0_0___40183), .Q (___0_____40190));
  nnd2s1 __________9__495319(.DIN1 (___0_00__40177), .DIN2
       (___0_0___40181), .Q (___0_0___40185));
  nor2s1 ___________0_495320(.DIN1 (___0_0___40178), .DIN2
       (________24008), .Q (___0_0___40184));
  xor2s1 _____________495321(.DIN1 (___0_0___40180), .DIN2
       (_________38675), .Q (___0_0___40183));
  dffacs1 _______________________________________________495322(.CLRB
       (reset), .CLK (clk), .DIN (___0_0___40179), .Q
       (_____________________________________________21974));
  xor2s1 _____________495323(.DIN1
       (_____________________________________________21971), .DIN2
       (___0_____40419), .Q (___0_0___40182));
  nnd2s1 ______9_____495324(.DIN1 (___0_0___40180), .DIN2
       (_________37836), .Q (___0_0___40181));
  nnd2s1 __________0__495325(.DIN1 (___0_9___40175), .DIN2
       (________28405), .Q (___0_0___40179));
  and2s1 ___________0_495326(.DIN1 (___9_____39746), .DIN2
       (_____________________________________________21971), .Q
       (___0_0___40178));
  nnd2s1 _____90____9_(.DIN1 (_________37878), .DIN2 (___0_99__40176),
       .Q (___0_00__40177));
  nor2s1 _____9_______495327(.DIN1 (_________37877), .DIN2
       (___0_99__40176), .Q (___0_0___40180));
  dffacs1 _______________________________________________495328(.CLRB
       (reset), .CLK (clk), .DIN (___0_9___40174), .QN
       (_____________________________________________21971));
  nnd2s1 _____9______495329(.DIN1 (___0_9___40173), .DIN2
       (___0_____40188), .Q (___0_9___40175));
  nor2s1 _____9____0_9(.DIN1 (______9__37813), .DIN2 (___0_9___40172),
       .Q (___0_99__40176));
  nnd2s1 _____9_______495330(.DIN1 (___0__0__40149), .DIN2
       (___0_9___40171), .Q (___0_9___40174));
  xor2s1 _____9___990_(.DIN1 (______0__37814), .DIN2 (___09_0__40700),
       .Q (___0_9___40173));
  and2s1 _____9______495331(.DIN1 (___09_0__40700), .DIN2
       (_________37726), .Q (___0_9___40172));
  dffacs1 ______________________________________495332(.CLRB (reset),
       .CLK (clk), .DIN (___0_9___40169), .QN (_________22014));
  nnd2s1 _____99____9_(.DIN1 (___0__9__40167), .DIN2 (inData[28]), .Q
       (___0_9___40171));
  nnd2s1 _____00______495333(.DIN1 (___0_____40165), .DIN2
       (___0_____40156), .Q (___0_9___40170));
  nnd2s1 _____0_______495334(.DIN1 (___0_90__40168), .DIN2
       (___0_____40164), .Q (___0_9___40169));
  nor2s1 _____0___9___495335(.DIN1 (___0_____40162), .DIN2
       (___0_____40166), .Q (___0__9__40167));
  xor2s1 _____0_______495336(.DIN1 (___0_____40163), .DIN2
       (_________38451), .Q (___0_____40165));
  nor2s1 _____0_____09(.DIN1 (___0__0__40159), .DIN2 (_____9__24665),
       .Q (___0_____40164));
  dffacs1 _______________________________________________495337(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40161), .Q (___0_____40419));
  xor2s1 _____0____900(.DIN1 (___0_____40419), .DIN2
       (_____________________________________________21972), .Q
       (___0_____40162));
  nnd2s1 _____09____9_495338(.DIN1 (___0_____40157), .DIN2
       (__9_____29815), .Q (___0_____40161));
  nnd2s1 ______0______495339(.DIN1
       (_____________________________________________21972), .DIN2
       (_____________________________________________21973), .Q
       (___0_____40160));
  nor2s1 _____________495340(.DIN1
       (_____________________________________________21972), .DIN2
       (____0___23882), .Q (___0__0__40159));
  xor2s1 _____________495341(.DIN1 (___0_____40155), .DIN2
       (___0__9__40158), .Q (___0_____40163));
  dffacs1 _______________________________________________495342(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40154), .Q
       (_____________________________________________21972));
  nnd2s1 _____________495343(.DIN1 (___0_____40153), .DIN2
       (___0_____40156), .Q (___0_____40157));
  nnd2s1 __________9__495344(.DIN1 (___0_____40152), .DIN2
       (_________37347), .Q (___0_____40155));
  nnd2s1 ___________0_495345(.DIN1 (___0_____40150), .DIN2
       (__9_____29938), .Q (___0_____40154));
  xor2s1 _____________495346(.DIN1 (_____9___37371), .DIN2
       (___0_____40151), .Q (___0_____40153));
  nnd2s1 _____________495347(.DIN1 (___0_____40151), .DIN2
       (_________37351), .Q (___0_____40152));
  nnd2s1 ______9_____495348(.DIN1 (___0__9__40148), .DIN2
       (___0_____40156), .Q (___0_____40150));
  nnd2s1 ______0___0__(.DIN1 (___0_____40147), .DIN2 (____90___37012),
       .Q (___0_____40151));
  nnd2s1 ___________0_495349(.DIN1 (___0_____40145), .DIN2
       (___0_____40156), .Q (___0__0__40149));
  xor2s1 ___________9_495350(.DIN1 (____9_0__37033), .DIN2
       (___0_____40146), .Q (___0__9__40148));
  nnd2s1 _____________495351(.DIN1 (___0_____40146), .DIN2
       (____90___37006), .Q (___0_____40147));
  xor2s1 ____________495352(.DIN1 (___0_____40143), .DIN2
       (___0_____40423), .Q (___0_____40145));
  nnd2s1 __________0_495353(.DIN1 (___0_____40144), .DIN2
       (___0_____40142), .Q (___0_____40146));
  nnd2s1 _____________495354(.DIN1 (___0_____40141), .DIN2
       (___0_____40423), .Q (___0_____40144));
  nnd2s1 _________990_495355(.DIN1 (___0_____40142), .DIN2
       (___0_____40141), .Q (___0_____40143));
  dffacs1 _______________________________________________495356(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40140), .Q
       (_____________________________________________21970));
  nnd2s1 ____________495357(.DIN1 (___0__0__40139), .DIN2
       (_________36964), .Q (___0_____40141));
  nnd2s1 ___________9_495358(.DIN1 (___0__9__40138), .DIN2
       (_________36946), .Q (___0_____40142));
  nnd2s1 ______9______495359(.DIN1 (___0_____40136), .DIN2
       (_________36607), .Q (___0_____40140));
  dffacs1 ______________________________________________9_495360(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40137), .Q
       (__________________________________________9___21951));
  hi1s1 _______495361(.DIN (___0__9__40138), .Q (___0__0__40139));
  nnd2s1 _____________495362(.DIN1 (___0_9___40072), .DIN2
       (___0_____40135), .Q (___0_____40137));
  nnd2s1 _____________495363(.DIN1 (___0_____40134), .DIN2
       (___0_____40156), .Q (___0_____40136));
  xor2s1 _________9___495364(.DIN1 (___0_____40133), .DIN2
       (___9_____39784), .Q (___0__9__40138));
  nnd2s1 _____________495365(.DIN1 (___0_____40115), .DIN2
       (___0_____40132), .Q (___0_____40135));
  xor2s1 ___________495366(.DIN1 (___0__0__40129), .DIN2
       (___0_____40130), .Q (___0_____40134));
  nnd2s1 ______0______495367(.DIN1 (___0_____40131), .DIN2
       (___0__9__40128), .Q (___0_____40133));
  nor2s1 ______9___495368(.DIN1 (___0_____40126), .DIN2
       (___90___28648), .Q (___0_____40132));
  nnd2s1 ___________9_495369(.DIN1 (___0_____40130), .DIN2
       (___0_____40127), .Q (___0_____40131));
  and2s1 _____________495370(.DIN1 (___0__9__40128), .DIN2
       (___0_____40127), .Q (___0__0__40129));
  xor2s1 _____________495371(.DIN1
       (__________________________________________________________________22003),
       .DIN2 (___0__9__40108), .Q (___0_____40126));
  dffacs1 ________________________________________________495372(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40124), .Q
       (______________________________________________21967));
  or2s1 _____________495373(.DIN1
       (__________________________________________________________________22003),
       .DIN2 (___0_____40125), .Q (___0_____40127));
  nnd2s1 _____________495374(.DIN1 (___0_____40125), .DIN2
       (__________________________________________________________________22003),
       .Q (___0__9__40128));
  nnd2s1 __________9__495375(.DIN1 (___999___39889), .DIN2
       (___0_____40123), .Q (___0_____40124));
  dffacs1 _______________________________________________495376(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40122), .QN
       (__________________________________________________________________22003));
  nnd2s1 ______9____0_495377(.DIN1 (___0_____40100), .DIN2
       (___0_____40424), .Q (___0_____40123));
  nnd2s1 _____________495378(.DIN1 (___0_____40121), .DIN2
       (___9_____39494), .Q (___0_____40122));
  dffacs1 ________________________________________________495379(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40117), .QN
       (___0_____40424));
  nor2s1 _____________495380(.DIN1 (___0_____40116), .DIN2
       (____00__28834), .Q (___0_____40121));
  or2s1 ____________495381(.DIN1 (___0__0__40119), .DIN2
       (___0__9__40118), .Q (___0_____40120));
  nnd2s1 __________0__495382(.DIN1 (___0_____40114), .DIN2
       (___0_90__40168), .Q (___0_____40117));
  and2s1 ___________0_495383(.DIN1 (___0_____40115), .DIN2
       (___0_____40113), .Q (___0_____40116));
  nor2s1 ______9____9_(.DIN1 (___0_____40112), .DIN2 (___9_9___39792),
       .Q (___0__0__40119));
  xor2s1 _____________495384(.DIN1 (________25522), .DIN2
       (___0_____40107), .Q (___0_____40114));
  nor2s1 ______0_____0(.DIN1
       (______________________________________________21965), .DIN2
       (___99____39809), .Q (___0__9__40118));
  dffacs1 ______________________________________________0_495385(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40110), .QN
       (___0__0__40421));
  nnd2s1 __________0_495386(.DIN1 (___0__0__40109), .DIN2 (inData[20]),
       .Q (___0_____40113));
  hi1s1 _______495387(.DIN
       (______________________________________________21965), .Q
       (___0_____40112));
  xor2s1 _____________495388(.DIN1 (___0_____40104), .DIN2
       (___9_____39582), .Q (___0_____40111));
  nnd2s1 _________990_495389(.DIN1 (___0_____40106), .DIN2
       (___9909__39806), .Q (___0_____40110));
  dffacs1 ________________________________________________495390(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40105), .QN
       (______________________________________________21965));
  xor2s1 ____________495391(.DIN1
       (______________________________________________21949), .DIN2
       (___0__9__40108), .Q (___0__0__40109));
  xor2s1 ___________9_495392(.DIN1 (___0__0__40099), .DIN2
       (___0_9___40645), .Q (___0_____40107));
  and2s1 _____________495393(.DIN1 (________28514), .DIN2
       (___0_____40101), .Q (___0_____40106));
  nor2s1 _____________495394(.DIN1
       (______________________________________________21949), .DIN2
       (___0__0__39993), .Q (___0_____40105));
  nnd2s1 ______9______495395(.DIN1 (___0_____40103), .DIN2
       (___0_____40102), .Q (___0_____40104));
  nnd2s1 ______0__9___(.DIN1 (___0_____40100), .DIN2 (________22013),
       .Q (___0_____40101));
  xor2s1 _____________495396(.DIN1 (___0_____40096), .DIN2
       (___0_9___40073), .Q (___0__0__40099));
  dffacs1 ________________________________________________495397(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40097), .QN
       (______________________________________________21949));
  xor2s1 ___________495398(.DIN1 (___0_____40093), .DIN2
       (___0__9__40098), .Q (___0_____40103));
  dffacs1 ______________________________________________0_495399(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40094), .Q (________22013));
  nnd2s1 _____________495400(.DIN1 (___0__0__40089), .DIN2
       (___0_____40095), .Q (___0_____40097));
  xor2s1 ______0___495401(.DIN1 (___0_0___40087), .DIN2
       (___0__0__40648), .Q (___0_____40096));
  dffacs1 ________________________________________________495402(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40091), .Q (___0_____40425));
  nnd2s1 ___________9_495403(.DIN1 (___0_9___40070), .DIN2
       (___0_____40090), .Q (___0_____40095));
  nnd2s1 _____________495404(.DIN1 (___0_09__40088), .DIN2
       (___0_90__40168), .Q (___0_____40094));
  nor2s1 ______9______495405(.DIN1
       (__________________________________________________________________22008),
       .DIN2 (___0_____40092), .Q (___0_____40093));
  nnd2s1 _____________495406(.DIN1 (___0_____40092), .DIN2
       (__________________________________________________________________22008),
       .Q (___0_____40102));
  nnd2s1 _____________495407(.DIN1 (___0_0___40085), .DIN2
       (___0__9__40048), .Q (___0_____40091));
  nor2s1 __________9__495408(.DIN1
       (__________________________________________9___21951), .DIN2
       (___0_0___40084), .Q (___0_____40090));
  dffacs1 ________________________________________________495409(.CLRB
       (reset), .CLK (clk), .DIN (___0_0___40082), .Q
       (__________________________________________________________________22008));
  and2s1 ___________0_495410(.DIN1 (___0_____40053), .DIN2
       (___0_0___40083), .Q (___0__0__40089));
  xor2s1 _____________495411(.DIN1 (___0_9___40075), .DIN2
       (___0_0___40080), .Q (___0_09__40088));
  nor2s1 _____9_______495412(.DIN1 (___0_____40067), .DIN2
       (___0_0___40081), .Q (___0_0___40087));
  xor2s1 _____90_____0(.DIN1
       (__________________________________________________________________22012),
       .DIN2 (___0_99__40078), .Q (___0_0___40086));
  and2s1 _____9____0__495413(.DIN1 (___0_9___40074), .DIN2
       (___0_9___40071), .Q (___0_0___40085));
  nnd2s1 _____9_____0_495414(.DIN1 (___0_9___40076), .DIN2
       (__________________________________________9___21951), .Q
       (___0__9__40108));
  or2s1 ___________9_495415(.DIN1
       (______________________________________________21950), .DIN2
       (________26731), .Q (___0_0___40084));
  nnd2s1 _____________495416(.DIN1 (___0_____40063), .DIN2
       (______________________________________________21950), .Q
       (___0_0___40083));
  or2s1 ______9_____495417(.DIN1
       (______________________________________________21950), .DIN2
       (___99_0__39817), .Q (___0_0___40082));
  and2s1 _____9____0_495418(.DIN1 (___0_90__40069), .DIN2
       (___0_0___40080), .Q (___0_0___40081));
  or2s1 _____9_______495419(.DIN1
       (__________________________________________________________________22012),
       .DIN2 (___0_99__40078), .Q (___0_00__40079));
  nnd2s1 _____9___990_495420(.DIN1 (___0_99__40078), .DIN2
       (__________________________________________________________________22012),
       .Q (___0_9___40077));
  hi1s1 _____9_(.DIN
       (______________________________________________21950), .Q
       (___0_9___40076));
  xor2s1 _____00_____0(.DIN1 (___0__9__40068), .DIN2 (___0_____40045),
       .Q (___0_9___40075));
  nor2s1 _____0_____9_495421(.DIN1 (___0_____40066), .DIN2
       (___0_0___39989), .Q (___0_9___40074));
  nnd2s1 _____0_______495422(.DIN1 (___0_____40065), .DIN2
       (___009___39981), .Q (___0_9___40073));
  nnd2s1 _____99______(.DIN1 (___0_____40062), .DIN2 (___9_____39219),
       .Q (___0_9___40072));
  nnd2s1 _____0_______495423(.DIN1 (___0_9___40070), .DIN2
       (___0_____40061), .Q (___0_9___40071));
  dffacs1 ________________________________________________495424(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40064), .QN
       (______________________________________________21950));
  nnd2s1 _____0___9___495425(.DIN1 (___0__9__40068), .DIN2
       (__________________________________________________________________21993),
       .Q (___0_90__40069));
  nor2s1 _____0_______495426(.DIN1
       (__________________________________________________________________21993),
       .DIN2 (___0__9__40068), .Q (___0_____40067));
  dffacs1 ________________________________________________495427(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40060), .QN
       (__________________________________________________________________22012));
  nor2s1 _____09____09(.DIN1 (___0__0__40059), .DIN2 (___0__0__40021),
       .Q (___0_____40066));
  nor2s1 ______0______495428(.DIN1 (___009___39980), .DIN2
       (___0_____40056), .Q (___0_____40065));
  nnd2s1 __________495429(.DIN1 (___0__9__40058), .DIN2
       (___0_____40047), .Q (___0_0___40080));
  or2s1 _____0_____9_495430(.DIN1 (___0_____40063), .DIN2
       (___0_____40054), .Q (___0_____40064));
  xor2s1 _____0_______495431(.DIN1 (___0_____40052), .DIN2
       (___0_____40057), .Q (___0_____40062));
  nor2s1 _____________495432(.DIN1 (_________22028), .DIN2
       (___0_____40026), .Q (___0_____40061));
  nnd2s1 _____________495433(.DIN1 (________23899), .DIN2
       (_________22028), .Q (___0_____40060));
  xor2s1 _____________495434(.DIN1 (___009___39977), .DIN2
       (___0_____40055), .Q (___0__9__40068));
  hi1s1 _______495435(.DIN (_________22028), .Q (___0__0__40059));
  nnd2s1 __________9__495436(.DIN1 (___0_____40057), .DIN2
       (___0_____40044), .Q (___0__9__40058));
  and2s1 ______9____0_495437(.DIN1 (___0_____40055), .DIN2
       (___0_0___39985), .Q (___0_____40056));
  nor2s1 _____________495438(.DIN1 (___0_9___40070), .DIN2
       (___0_____40050), .Q (___0_____40054));
  nnd2s1 _____________495439(.DIN1 (___0_____40051), .DIN2
       (___0____26076), .Q (___0_____40053));
  dffacs1 ________________________________________________495440(.CLRB
       (reset), .CLK (clk), .DIN (___0__0__40049), .QN
       (_________22028));
  xor2s1 ____________495441(.DIN1
       (__________________________________________________________________21993),
       .DIN2 (___0_____40046), .Q (___0_____40052));
  nor2s1 __________0__495442(.DIN1 (___0_____40015), .DIN2
       (___0_____40042), .Q (___0_____40057));
  nor2s1 ______9____0_495443(.DIN1 (___0_____40040), .DIN2
       (___0_____40043), .Q (___0_____40055));
  xor2s1 ___________9_495444(.DIN1 (___0_____40034), .DIN2
       (___0_____40027), .Q (___0_____40051));
  xor2s1 _____________495445(.DIN1 (___0_____40030), .DIN2
       (___0_____40041), .Q (___0_____40050));
  nnd2s1 ____________495446(.DIN1 (___0__9__40038), .DIN2
       (___0__9__40048), .Q (___0__0__40049));
  nnd2s1 __________0_495447(.DIN1 (___0_____40046), .DIN2
       (___0_____40045), .Q (___0_____40047));
  or2s1 _____________495448(.DIN1 (___0_____40045), .DIN2
       (___0_____40046), .Q (___0_____40044));
  nor2s1 ______0__990_(.DIN1 (___00_9__39911), .DIN2 (___0_____40031),
       .Q (___0_____40043));
  nor2s1 ____________495449(.DIN1 (___0_____40019), .DIN2
       (___0_____40041), .Q (___0_____40042));
  nor2s1 ___________9_495450(.DIN1 (___00____39967), .DIN2
       (___0_____40033), .Q (___0_____40040));
  xor2s1 _____________495451(.DIN1
       (______________________________________________21962), .DIN2
       (___9__9__39606), .Q (___0__0__40039));
  and2s1 _____________495452(.DIN1 (___0__9__40029), .DIN2
       (___09____40702), .Q (___0__9__40038));
  xor2s1 _____________495453(.DIN1 (___00____39933), .DIN2
       (___0_____40032), .Q (___0_____40046));
  or2s1 _________9___495454(.DIN1
       (______________________________________________21962), .DIN2
       (___0_____40035), .Q (___0_____40037));
  nnd2s1 _____________495455(.DIN1 (___0_____40035), .DIN2
       (______________________________________________21962), .Q
       (___0_____40036));
  xor2s1 ___________495456(.DIN1 (___0_____40024), .DIN2
       (___9_0___39709), .Q (___0_____40034));
  and2s1 _____________495457(.DIN1 (___0_____40032), .DIN2
       (___00_0__39912), .Q (___0_____40033));
  and2s1 __________495458(.DIN1 (___0_____40032), .DIN2
       (___00_0__39930), .Q (___0_____40031));
  xor2s1 ___________9_495459(.DIN1 (___0_____40025), .DIN2
       (______________________________________________21938), .Q
       (___0_____40030));
  nor2s1 _____________495460(.DIN1 (___0_____40023), .DIN2
       (___0_____40028), .Q (___0_____40041));
  nor2s1 ______0______495461(.DIN1 (___0_____40022), .DIN2
       (___0_____40014), .Q (___0__9__40029));
  dffacs1 ________________________________________________495462(.CLRB
       (reset), .CLK (clk), .DIN (___0__9__40020), .QN
       (______________________________________________21962));
  and2s1 ______9______495463(.DIN1 (___0_____40017), .DIN2
       (___0_____40027), .Q (___0_____40028));
  xor2s1 __________9__495464(.DIN1 (___0_____40013), .DIN2
       (___9_____39312), .Q (___0_____40032));
  xor2s1 ______0______495465(.DIN1 (___0_____40018), .DIN2
       (_________41343), .Q (___0_____40025));
  or2s1 _____________495466(.DIN1 (___0_____40023), .DIN2
       (___0_____40016), .Q (___0_____40024));
  nor2s1 ____________495467(.DIN1 (______0__22027), .DIN2
       (___0__0__40021), .Q (___0_____40022));
  nor2s1 __________0__495468(.DIN1 (______0__22027), .DIN2
       (___9_____39575), .Q (___0__9__40020));
  nor2s1 ___________0_495469(.DIN1
       (______________________________________________21938), .DIN2
       (___0_____40018), .Q (___0_____40019));
  hi1s1 _______495470(.DIN (___0_____40016), .Q (___0_____40017));
  and2s1 ___________9_495471(.DIN1 (___0_____40018), .DIN2
       (______________________________________________21938), .Q
       (___0_____40015));
  nor2s1 _____________495472(.DIN1 (___0_9___40070), .DIN2
       (___0__0__40012), .Q (___0_____40014));
  nnd2s1 ____________495473(.DIN1 (___0__9__40011), .DIN2
       (___0009__39901), .Q (___0_____40013));
  xor2s1 ______9___0_9(.DIN1 (___0_____40008), .DIN2 (___99_0__39864),
       .Q (___0_____40016));
  dffacs1 ________________________________________________495474(.CLRB
       (reset), .CLK (clk), .DIN (___0_____40009), .Q (______0__22027));
  xor2s1 _____________495475(.DIN1 (___00____39909), .DIN2
       (___0_____40010), .Q (___0_____40018));
  xor2s1 _________990_495476(.DIN1 (___0_____40005), .DIN2
       (___0_0___39987), .Q (___0__0__40012));
  nnd2s1 ____________495477(.DIN1 (___0_____40010), .DIN2
       (___000___39899), .Q (___0__9__40011));
  nnd2s1 ______0____9_(.DIN1 (___0_____40006), .DIN2 (___0__9__40048),
       .Q (___0_____40009));
  nor2s1 _____________495478(.DIN1
       (__________________________________________________________________21997),
       .DIN2 (___0_____40007), .Q (___0_____40008));
  and2s1 _____________495479(.DIN1 (___0_____40007), .DIN2
       (__________________________________________________________________21997),
       .Q (___0_____40023));
  xnr2s1 ______0______495480(.DIN1 (_____9___36721), .DIN2
       (___0_____40003), .Q (___0_____40010));
  and2s1 _________9___495481(.DIN1 (___0_____40004), .DIN2
       (___0__0__40021), .Q (___0_____40006));
  xor2s1 _____________495482(.DIN1 (________23476), .DIN2
       (___0__0__40002), .Q (___0_____40005));
  xor2s1 ______9____495483(.DIN1 (___0__9__40001), .DIN2
       (___99____39870), .Q (___0_____40007));
  nor2s1 _____________495484(.DIN1 (___0_____40000), .DIN2
       (___00____39943), .Q (___0_____40004));
  nnd2s1 ______0___495485(.DIN1 (___0_____39997), .DIN2
       (___99____39877), .Q (___0_____40003));
  nnd2s1 ___________9_495486(.DIN1 (___0_____39999), .DIN2
       (___0_0___39988), .Q (___0_____40027));
  xor2s1 _____________495487(.DIN1 (___0_____39998), .DIN2
       (_________36301), .Q (___0__0__40002));
  xor2s1 _____________495488(.DIN1 (___0_____39996), .DIN2
       (___0_____40092), .Q (___0__9__40001));
  nor2s1 _____________495489(.DIN1 (___0_____39995), .DIN2
       (___0____26076), .Q (___0_____40000));
  dffacs1 ________________________________________________495490(.CLRB
       (reset), .CLK (clk), .DIN (___0_____39994), .QN
       (______________________________________________21963));
  or2s1 _____________495491(.DIN1 (___0_____39998), .DIN2
       (___0_0___39986), .Q (___0_____39999));
  nnd2s1 __________9__495492(.DIN1 (___0_____39996), .DIN2
       (___000___39897), .Q (___0_____39997));
  nnd2s1 ___________0_495493(.DIN1 (___0_9___40070), .DIN2
       (___0_____40026), .Q (___0__0__40021));
  nnd2s1 _____________495494(.DIN1 (___0_____40426), .DIN2
       (___0_____40425), .Q (___0_____39995));
  nor2s1 _____________495495(.DIN1 (___0_____40425), .DIN2
       (___0_____40426), .Q (___0_____40026));
  nor2s1 ______9_____495496(.DIN1 (___0_____40426), .DIN2
       (___0__0__39993), .Q (___0_____39994));
  xor2s1 __________0__495497(.DIN1 (___0_0___39991), .DIN2
       (___0_____40323), .Q (___0_____39996));
  xor2s1 ___________0_495498(.DIN1 (___0_09__39992), .DIN2
       (___0_00__39983), .Q (___0_____39998));
  dffacs1 ________________________________________________495499(.CLRB
       (reset), .CLK (clk), .DIN (___0_0___39990), .Q (___0_____40426));
  xor2s1 _____9_____9_495500(.DIN1 (___009___39975), .DIN2
       (___0_____40308), .Q (___0_09__39992));
  nnd2s1 _____9_______495501(.DIN1 (___0_0___39984), .DIN2
       (___009___39974), .Q (___0_0___39991));
  nnd2s1 ____________495502(.DIN1 (___0099__39982), .DIN2
       (___0__9__40048), .Q (___0_0___39990));
  dffacs1 ________________________________________________495503(.CLRB
       (reset), .CLK (clk), .DIN (___0090__39973), .QN
       (______________________________________________21937));
  nor2s1 __________0_495504(.DIN1 (___0_9___40070), .DIN2
       (___00_9__39972), .Q (___0_0___39989));
  or2s1 ______9______495505(.DIN1
       (______________________________________________21937), .DIN2
       (___0_0___39987), .Q (___0_0___39988));
  and2s1 _____90__990_(.DIN1 (___0_0___39987), .DIN2
       (______________________________________________21937), .Q
       (___0_0___39986));
  xor2s1 _____9______495506(.DIN1 (___009___39976), .DIN2
       (___00____41368), .Q (___0_0___39985));
  or2s1 _____0_____9_495507(.DIN1 (___0_00__39983), .DIN2
       (___00____39969), .Q (___0_0___39984));
  nor2s1 _____________495508(.DIN1 (________26829), .DIN2
       (___00____39968), .Q (___0099__39982));
  nnd2s1 _____9_______495509(.DIN1 (___009___39978), .DIN2
       (___009___39979), .Q (___009___39981));
  nor2s1 _____9_______495510(.DIN1 (___009___39979), .DIN2
       (___009___39978), .Q (___009___39980));
  nnd2s1 _____99__9___(.DIN1 (___009___39976), .DIN2 (___009___39978),
       .Q (___009___39977));
  and2s1 _____0_______495511(.DIN1 (___009___39974), .DIN2
       (___09____40659), .Q (___009___39975));
  nnd2s1 ___________495512(.DIN1 (___00____39966), .DIN2
       (___9_9___39793), .Q (___0090__39973));
  xor2s1 _____9_______495513(.DIN1 (___09_0__40690), .DIN2
       (___00_0__39964), .Q (___00_9__39972));
  nor2s1 _____9____900(.DIN1 (___00____39958), .DIN2 (___00____39965),
       .Q (___0_0___39987));
  xnr2s1 _____00____9_(.DIN1
       (______________________________________________21967), .DIN2
       (___00____39970), .Q (___00____39971));
  hi1s1 _______495514(.DIN (___09____40659), .Q (___00____39969));
  nor2s1 _____9_______495515(.DIN1 (___0_9___40070), .DIN2
       (___00_9__39963), .Q (___00____39968));
  nnd2s1 _____0_______495516(.DIN1 (___0__0__40648), .DIN2
       (___00____39967), .Q (___009___39976));
  or2s1 _____0_______495517(.DIN1 (___00____39967), .DIN2
       (___00____39970), .Q (___009___39978));
  nnd2s1 _____________495518(.DIN1 (________27077), .DIN2
       (__________________________________________________________________21997),
       .Q (___00____39966));
  dffacs1 _____________________________________________9_495519(.CLRB
       (reset), .CLK (clk), .DIN (___00____39961), .QN
       (_________________________________________9___21943));
  nor2s1 _____0_____0_(.DIN1 (___00____39960), .DIN2 (___00_0__39964),
       .Q (___00____39965));
  nnd2s1 _____________495520(.DIN1 (___00____39962), .DIN2
       (___99____39866), .Q (___009___39974));
  dffacs1 ______________________________________________9_495521(.CLRB
       (reset), .CLK (clk), .DIN (___00____39957), .QN
       (__________________________________________________________________21993));
  xor2s1 _____0_______495522(.DIN1 (___00____39954), .DIN2
       (______________________________________________21936), .Q
       (___00_9__39963));
  xor2s1 __________0__495523(.DIN1 (___00____39952), .DIN2
       (___9_9___39790), .Q (___00____39970));
  nnd2s1 ___________0_495524(.DIN1 (_____9___38698), .DIN2
       (___00_9__39955), .Q (___00____39961));
  dffacs1 ________________________________________________495525(.CLRB
       (reset), .CLK (clk), .DIN (___00_0__39956), .QN
       (__________________________________________________________________21997));
  nor2s1 _____0_____9_495526(.DIN1
       (__________________________________________________________________21996),
       .DIN2 (___00____39959), .Q (___00____39960));
  and2s1 _____09______(.DIN1 (___00____39959), .DIN2
       (__________________________________________________________________21996),
       .Q (___00____39958));
  or2s1 ____________495527(.DIN1 (___00____39951), .DIN2
       (_________37837), .Q (___00____39957));
  xnr2s1 __________0_495528(.DIN1 (_________38650), .DIN2
       (___09____40704), .Q (___00____39962));
  nor2s1 _____________495529(.DIN1 (___00____39953), .DIN2
       (___00____39950), .Q (___00_0__39964));
  nnd2s1 _________990_495530(.DIN1 (________27640), .DIN2
       (___00_0__39949), .Q (___00_0__39956));
  nnd2s1 ____________495531(.DIN1 (___00___24169), .DIN2
       (___00_9__39948), .Q (___00_9__39955));
  nor2s1 ___________9_495532(.DIN1 (___00____39953), .DIN2
       (___00____39947), .Q (___00____39954));
  xor2s1 _____________495533(.DIN1 (___00____39942), .DIN2
       (___00____41368), .Q (___00____39959));
  xor2s1 _____________495534(.DIN1 (___00_0__39939), .DIN2
       (___0_9___40645), .Q (___00____39952));
  nnd2s1 _____________495535(.DIN1 (_____9__25881), .DIN2
       (___00____39944), .Q (___00____39951));
  dffacs1 ________________________________________________495536(.CLRB
       (reset), .CLK (clk), .DIN (___00____39945), .QN
       (___0_____40432));
  and2s1 _________9___495537(.DIN1 (___00____39946), .DIN2
       (______________________________________________21936), .Q
       (___00____39950));
  nor2s1 ______0____495538(.DIN1 (___99____39857), .DIN2
       (___00____39935), .Q (___00_0__39949));
  xor2s1 _____________495539(.DIN1
       (_____________________________________________21941), .DIN2
       (__________________________________________9___21923), .Q
       (___00_9__39948));
  dffacs1 ________________________________________________495540(.CLRB
       (reset), .CLK (clk), .DIN (___00____39934), .Q
       (______________________________________________21938));
  hi1s1 _______495541(.DIN (___00____39946), .Q (___00____39947));
  nnd2s1 __________495542(.DIN1 (___00____39932), .DIN2
       (___9_____39644), .Q (___00____39945));
  or2s1 ______0____9_495543(.DIN1
       (__________________________________________9___21923), .DIN2
       (______9__37419), .Q (___00____39944));
  nor2s1 ______0______495544(.DIN1 (___0_9___40070), .DIN2
       (___00____39931), .Q (___00____39943));
  xor2s1 _____________495545(.DIN1 (___00____39924), .DIN2
       (___99____39846), .Q (___00____39942));
  nor2s1 _____________495546(.DIN1 (___00____39940), .DIN2
       (___00____39941), .Q (___00____39953));
  nnd2s1 _____________495547(.DIN1 (___00____39941), .DIN2
       (___00____39940), .Q (___00____39946));
  xor2s1 __________9__495548(.DIN1 (___9_90__39607), .DIN2
       (___00____39923), .Q (___00_0__39939));
  nor2s1 _____________495549(.DIN1 (___00____39937), .DIN2
       (___00____39936), .Q (___00____39938));
  nor2s1 ______9______495550(.DIN1 (___00____39927), .DIN2
       (___00____39925), .Q (___00____39935));
  nnd2s1 ____________495551(.DIN1 (________27642), .DIN2
       (___00____39926), .Q (___00____39934));
  xor2s1 __________0__495552(.DIN1 (___00____39908), .DIN2
       (___00____39967), .Q (___00____39933));
  nor2s1 ___________0_495553(.DIN1 (___00_0__39922), .DIN2
       (___00____39903), .Q (___00____39932));
  dffacs1 ______________________________________________9_495554(.CLRB
       (reset), .CLK (clk), .DIN (___00_9__39921), .Q
       (__________________________________________9___21923));
  xor2s1 ______0____9_495555(.DIN1 (___00____39915), .DIN2
       (_________38155), .Q (___00____39931));
  xor2s1 _____________495556(.DIN1 (___00____39913), .DIN2
       (___9_____39542), .Q (___00____39941));
  and2s1 ____________495557(.DIN1 (___00____39967), .DIN2
       (___0__0__40421), .Q (___00____39936));
  nor2s1 __________0_495558(.DIN1 (___0__0__40421), .DIN2
       (___00____39967), .Q (___00____39937));
  nnd2s1 _____________495559(.DIN1 (___00____39967), .DIN2
       (___00____39910), .Q (___00_0__39930));
  nor2s1 _____00____9_495560(.DIN1 (____0_0__38093), .DIN2
       (___00____39917), .Q (___00____39927));
  nnd2s1 _____0_______495561(.DIN1 (___00____39925), .DIN2
       (___0_____40434), .Q (___00____39926));
  xor2s1 _____________495562(.DIN1 (___99____39847), .DIN2
       (___00____39918), .Q (___00____39924));
  dffacs1 ________________________________________________495563(.CLRB
       (reset), .CLK (clk), .DIN (___00____39916), .Q (______9__22026));
  nor2s1 _____________495564(.DIN1 (___9_0___39621), .DIN2
       (___00____39905), .Q (___00____39923));
  nor2s1 _____9___9___(.DIN1
       (______________________________________________21921), .DIN2
       (___00_0__39902), .Q (___00_0__39922));
  nnd2s1 _____________495565(.DIN1 (___00____39914), .DIN2
       (___00___24170), .Q (___00_9__39921));
  nor2s1 ______0____495566(.DIN1 (___00____39919), .DIN2
       (___00____39906), .Q (___00____39920));
  xor2s1 _____________495567(.DIN1 (___99____39811), .DIN2
       (___999___39887), .Q (___00____39940));
  or2s1 __________495568(.DIN1 (___99____39848), .DIN2
       (___00____39918), .Q (___00____39928));
  dffacs1 ________________________________________________495569(.CLRB
       (reset), .CLK (clk), .DIN (___000___39896), .QN
       (___0_____40434));
  nnd2s1 ___________9_495570(.DIN1 (___000___39895), .DIN2
       (___000___39900), .Q (___00____39917));
  xor2s1 _____________495571(.DIN1 (___9_0___39623), .DIN2
       (___00____39904), .Q (___00____39967));
  nnd2s1 ______9______495572(.DIN1 (___999___39888), .DIN2
       (___99____39861), .Q (___00____39916));
  xor2s1 _____________495573(.DIN1 (___09____40706), .DIN2
       (___999___39886), .Q (___00____39915));
  nnd2s1 _____________495574(.DIN1 (___9999__39891), .DIN2
       (___9__9__39659), .Q (___00____39914));
  nor2s1 __________9__495575(.DIN1 (___999___39885), .DIN2
       (___999___39890), .Q (___00____39913));
  xor2s1 ______9____0_495576(.DIN1 (___00_9__39911), .DIN2
       (___00____39910), .Q (___00_0__39912));
  xor2s1 _____________495577(.DIN1 (___99____39880), .DIN2
       (___00_9__39911), .Q (___00____39909));
  xor2s1 _____________495578(.DIN1 (_________37687), .DIN2
       (___00_9__39911), .Q (___00____39908));
  hi1s1 _______495579(.DIN (___00____39906), .Q (___00____39907));
  nor2s1 ____________495580(.DIN1 (___9_0___39622), .DIN2
       (___00____39904), .Q (___00____39905));
  dffacs1 ________________________________________________495581(.CLRB
       (reset), .CLK (clk), .DIN (___0000__39892), .Q
       (______________________________________________21921));
  and2s1 ______0___0__495582(.DIN1 (___00_0__39902), .DIN2
       (___000___39894), .Q (___00____39903));
  nnd2s1 ___________0_495583(.DIN1 (___00_9__39911), .DIN2
       (___000___39898), .Q (___0009__39901));
  nnd2s1 ___________9_495584(.DIN1 (___9990__39883), .DIN2
       (___9_____39773), .Q (___000___39900));
  or2s1 _____________495585(.DIN1 (___000___39898), .DIN2
       (___00_9__39911), .Q (___000___39899));
  nor2s1 ____________495586(.DIN1 (___990___39800), .DIN2
       (___99____39879), .Q (___00____39918));
  xor2s1 _____90___0_9(.DIN1 (___99____39871), .DIN2 (_________36854),
       .Q (___000___39897));
  nnd2s1 _____________495587(.DIN1 (___999___39884), .DIN2 (___9_9), .Q
       (___000___39896));
  and2s1 _____9___990_495588(.DIN1 (___00_9__39911), .DIN2
       (__________________________________________9___21966), .Q
       (___00____39919));
  nor2s1 _____9______495589(.DIN1
       (__________________________________________9___21966), .DIN2
       (___00_9__39911), .Q (___00____39906));
  nnd2s1 ___________9_495590(.DIN1 (___000___39893), .DIN2
       (___99____39875), .Q (___000___39895));
  xnr2s1 _____________495591(.DIN1
       (______________________________________________21936), .DIN2
       (___000___39893), .Q (___000___39894));
  nnd2s1 _____________495592(.DIN1 (___9_____39484), .DIN2
       (___99____39876), .Q (___0000__39892));
  xnr2s1 _____________495593(.DIN1 (___9_____39231), .DIN2
       (___99____39868), .Q (___9999__39891));
  and2s1 _________9___495594(.DIN1 (___09____40706), .DIN2
       (___99____39851), .Q (___999___39890));
  nnd2s1 _____________495595(.DIN1 (________29086), .DIN2
       (___99____39869), .Q (___999___39889));
  nor2s1 ___________495596(.DIN1 (___99____39820), .DIN2
       (___99____39874), .Q (___999___39888));
  xor2s1 _____9_______495597(.DIN1 (___99____39878), .DIN2
       (_____9___38512), .Q (___999___39887));
  nor2s1 ______0___495598(.DIN1 (___9_____39600), .DIN2
       (___99_0__39873), .Q (___00____39904));
  nor2s1 ___________9_495599(.DIN1 (___99____39850), .DIN2
       (___999___39885), .Q (___999___39886));
  xor2s1 _____________495600(.DIN1 (___99____39856), .DIN2
       (___9_9___39696), .Q (___999___39884));
  or2s1 _____________495601(.DIN1
       (______________________________________________21936), .DIN2
       (______________________________________________21937), .Q
       (___9990__39883));
  or2s1 _____________495602(.DIN1 (___99_9__39863), .DIN2
       (___99____39881), .Q (___99_9__39882));
  dffacs1 ________________________________________________495603(.CLRB
       (reset), .CLK (clk), .DIN (___99____39860), .QN
       (______________________________________________21960));
  xor2s1 _____09______495604(.DIN1 (___0_____40092), .DIN2
       (_________38372), .Q (___99____39880));
  nor2s1 _____0____9__(.DIN1 (___9_9___39795), .DIN2 (___99____39878),
       .Q (___99____39879));
  nnd2s1 ______9____0_495605(.DIN1 (___0_____40092), .DIN2
       (___99____39867), .Q (___99____39877));
  dffacs1 ______________________________________________0_495606(.CLRB
       (reset), .CLK (clk), .DIN (___99____39862), .QN
       (___0_____40427));
  xnr2s1 _____________495607(.DIN1 (___99_9__39872), .DIN2
       (___9_____39601), .Q (___00_9__39911));
  nnd2s1 _____________495608(.DIN1 (___99____39859), .DIN2 (inData[4]),
       .Q (___99____39876));
  hi1s1 ______0(.DIN
       (______________________________________________21936), .Q
       (___99____39875));
  nor2s1 ______9_____495609(.DIN1 (___9_____39743), .DIN2
       (___99____39858), .Q (___99____39874));
  nor2s1 __________0__495610(.DIN1 (___9_____39599), .DIN2
       (___99_9__39872), .Q (___99_0__39873));
  or2s1 ___________0_495611(.DIN1 (___99____39870), .DIN2
       (___0_____40092), .Q (___99____39871));
  xor2s1 ___________9_495612(.DIN1 (___99_9__39844), .DIN2
       (___9___22267), .Q (___99____39869));
  nnd2s1 _____9______495613(.DIN1 (___99_9__39854), .DIN2
       (___9_____39538), .Q (___99____39868));
  and2s1 ______9___0_495614(.DIN1 (___99____39870), .DIN2
       (___900___38985), .Q (___99____39867));
  nor2s1 _____________495615(.DIN1 (____9___26770), .DIN2
       (___99_0__39855), .Q (___999___39885));
  dffacs1 ________________________________________________495616(.CLRB
       (reset), .CLK (clk), .DIN (___99____39852), .Q
       (______________________________________________21936));
  xnr2s1 ______9__990_495617(.DIN1 (___99_0__39864), .DIN2
       (___99_9__39863), .Q (___99____39865));
  nnd2s1 ____________495618(.DIN1 (___99____39849), .DIN2
       (___99____39861), .Q (___99____39862));
  nnd2s1 ___________9_495619(.DIN1 (________29087), .DIN2
       (___99_0__39845), .Q (___99____39860));
  xor2s1 ______0______495620(.DIN1 (___99____39840), .DIN2
       (___0_____40650), .Q (___99____39878));
  xor2s1 _____9_______495621(.DIN1 (___99____39835), .DIN2
       (_____9___37654), .Q (___99____39881));
  nor2s1 _____________495622(.DIN1 (___99____39838), .DIN2
       (___9_9___39610), .Q (___99____39859));
  xor2s1 _________9___495623(.DIN1 (___99____39832), .DIN2
       (___9_____39752), .Q (___99____39866));
  nor2s1 ______0______495624(.DIN1 (___9_90__39517), .DIN2
       (___99____39842), .Q (___99_9__39872));
  hi1s1 _______495625(.DIN (___000___39898), .Q (___0_____40092));
  xor2s1 _____9_____09(.DIN1 (___9_____39783), .DIN2 (___99____39825),
       .Q (___99____39858));
  nor2s1 _____________495626(.DIN1 (___0_____40603), .DIN2
       (________26254), .Q (___99____39857));
  xor2s1 _____99___900(.DIN1 (___99____39853), .DIN2 (___99____39808),
       .Q (___99____39856));
  nor2s1 _____________495627(.DIN1 (___9_____39779), .DIN2
       (___99____39839), .Q (___0_00__39983));
  xor2s1 _____9_______495628(.DIN1 (___99____39833), .DIN2
       (___9__9__39731), .Q (___99_0__39855));
  nnd2s1 _____0_______495629(.DIN1 (___99____39853), .DIN2
       (___9_9___39522), .Q (___99_9__39854));
  nnd2s1 _____________495630(.DIN1 (___99____39828), .DIN2
       (________23478), .Q (___99____39852));
  hi1s1 _____9_495631(.DIN (___99____39850), .Q (___99____39851));
  xor2s1 __________9__495632(.DIN1 (___9_____39584), .DIN2
       (___99____39841), .Q (___000___39898));
  nnd2s1 ______0____0_(.DIN1 (___99____39830), .DIN2 (___99____39831),
       .Q (___99____39870));
  nor2s1 _____99______495633(.DIN1 (___99____39824), .DIN2
       (___9_____39744), .Q (___99____39849));
  and2s1 _____________495634(.DIN1 (___99____39847), .DIN2
       (___99____39846), .Q (___99____39848));
  nnd2s1 _____0______495635(.DIN1 (___0_____40100), .DIN2
       (______________________________________________21948), .Q
       (___99_0__39845));
  xor2s1 _____0____0__(.DIN1 (___0__0__40421), .DIN2
       (__________________________________________________________________22011),
       .Q (___99_9__39844));
  nor2s1 ___________0_495636(.DIN1 (___99____39846), .DIN2
       (___99____39847), .Q (___99____39843));
  dffacs1 ________________________________________________495637(.CLRB
       (reset), .CLK (clk), .DIN (___99_9__39826), .Q
       (______________________________________________21946));
  and2s1 ___________9_495638(.DIN1 (___99____39841), .DIN2
       (___9_9___39519), .Q (___99____39842));
  nnd2s1 _____________495639(.DIN1 (___99____39823), .DIN2
       (___9__0__39742), .Q (___99____39840));
  xor2s1 ____________495640(.DIN1 (___99____39812), .DIN2
       (____90___36104), .Q (___99____39839));
  xor2s1 _____9____0_495641(.DIN1 (___0_____40435), .DIN2
       (___0_____40610), .Q (___99____39838));
  dffacs1 ________________________________________________495642(.CLRB
       (reset), .CLK (clk), .DIN (___99____39821), .QN
       (___0_____40603));
  or2s1 ____________495643(.DIN1
       (__________________________________________________________________22011),
       .DIN2 (___99____39834), .Q (___99____39835));
  and2s1 ___________9_495644(.DIN1 (___99____39834), .DIN2
       (__________________________________________________________________22011),
       .Q (___99_9__39863));
  nor2s1 _____0_______495645(.DIN1
       (_________________________________________________________________21991),
       .DIN2 (___99____39833), .Q (___99____39850));
  and2s1 _____________495646(.DIN1 (___99____39831), .DIN2
       (___99____39829), .Q (___99____39832));
  nnd2s1 _____________495647(.DIN1 (___99____39829), .DIN2
       (___99_0__39827), .Q (___99____39830));
  nnd2s1 _____0___9___495648(.DIN1 (________26568), .DIN2
       (___0_____40435), .Q (___99____39828));
  xor2s1 _____________495649(.DIN1 (___990___39801), .DIN2
       (___99_0__39827), .Q (___99____39847));
  nnd2s1 ___________495650(.DIN1 (___9_9___39614), .DIN2
       (___99_9__39816), .Q (___99_9__39826));
  dffacs1 ________________________________________________495651(.CLRB
       (reset), .CLK (clk), .DIN (___99____39818), .Q
       (______________________________________________21948));
  xor2s1 _____________495652(.DIN1 (___99____39822), .DIN2
       (___0_____40308), .Q (___99____39825));
  nor2s1 __________495653(.DIN1 (___99____39815), .DIN2
       (___99____39819), .Q (___99____39824));
  nnd2s1 ___________9_495654(.DIN1 (___99____39810), .DIN2
       (___9_____39781), .Q (___99____39853));
  nor2s1 _____________495655(.DIN1 (___9_____39739), .DIN2
       (___9900__39797), .Q (___99____39823));
  or2s1 ______0______495656(.DIN1 (___9_____39775), .DIN2
       (___99____39822), .Q (___99_0__39837));
  dffacs1 ________________________________________________495657(.CLRB
       (reset), .CLK (clk), .DIN (___99_0__39807), .Q
       (__________________________________________________________________22011));
  nnd2s1 _____________495658(.DIN1 (___9_9___39794), .DIN2 (___9_9), .Q
       (___99____39821));
  xor2s1 _____________495659(.DIN1 (___09____40708), .DIN2
       (___090__23301), .Q (___99____39841));
  xor2s1 ______9___9__(.DIN1 (___9_____39785), .DIN2 (___9_99__39796),
       .Q (___99____39833));
  nor2s1 ___________0_495660(.DIN1 (___9_90__39787), .DIN2
       (___99____39819), .Q (___99____39820));
  nor2s1 _____________495661(.DIN1 (___99_0__39817), .DIN2
       (___9_9___39788), .Q (___99____39818));
  nnd2s1 _____________495662(.DIN1 (___9_____39782), .DIN2
       (inData[28]), .Q (___99_9__39816));
  nor2s1 ____________495663(.DIN1 (___99____39814), .DIN2
       (___9_9___39789), .Q (___99____39815));
  xor2s1 ______9___0__(.DIN1
       (__________________________________________________________________22007),
       .DIN2 (___9_____39276), .Q (___99____39813));
  nor2s1 ___________0_495664(.DIN1 (___9_____39767), .DIN2
       (___9_9___39791), .Q (___99____39812));
  xor2s1 ______0____9_495665(.DIN1 (___990___39799), .DIN2
       (___990___39798), .Q (___99____39811));
  nnd2s1 _____________495666(.DIN1 (___9_____39776), .DIN2
       (___9_____39539), .Q (___99____39810));
  dffacs1 ________________________________________________495667(.CLRB
       (reset), .CLK (clk), .DIN (___9__9__39777), .QN
       (___0_____40435));
  nnd2s1 _____0______495668(.DIN1 (___99____39809), .DIN2
       (___99____39808), .Q (___99____39829));
  dffacs1 ________________________________________________495669(.CLRB
       (reset), .CLK (clk), .DIN (___9__0__39778), .QN
       (__________________________________________________________________21996));
  nnd2s1 __________0_495670(.DIN1 (___9_____39772), .DIN2
       (___9909__39806), .Q (___99_0__39807));
  xnr2s1 _____________495671(.DIN1 (___99_9__39836), .DIN2
       (___9_____39766), .Q (___990___39805));
  or2s1 _________990_495672(.DIN1
       (__________________________________________________________________22007),
       .DIN2 (___990___39802), .Q (___990___39804));
  nnd2s1 ____________495673(.DIN1 (___990___39802), .DIN2
       (__________________________________________________________________22007),
       .Q (___990___39803));
  xor2s1 ___________9_495674(.DIN1 (___9__9__39768), .DIN2
       (____9____38909), .Q (___990___39801));
  nor2s1 ______9______495675(.DIN1 (___9_____39734), .DIN2
       (___9_____39771), .Q (___99____39822));
  and2s1 _____________495676(.DIN1 (___990___39799), .DIN2
       (___990___39798), .Q (___990___39800));
  nor2s1 _____90______(.DIN1 (___9_____39719), .DIN2 (___9_99__39796),
       .Q (___9900__39797));
  nor2s1 _____9___9___495677(.DIN1 (___990___39798), .DIN2
       (___990___39799), .Q (___9_9___39795));
  nor2s1 ______0______495678(.DIN1 (___09_9__40660), .DIN2
       (___9_____39780), .Q (___9_9___39794));
  nnd2s1 ___________495679(.DIN1 (___00____39925), .DIN2
       (_________22022), .Q (___9_9___39793));
  nnd2s1 _____0_______495680(.DIN1 (___9_9___39792), .DIN2
       (___9_00__39527), .Q (___99____39831));
  xor2s1 _____9____495681(.DIN1 (___9_____39753), .DIN2
       (___9_9___39790), .Q (___9_9___39791));
  xor2s1 ___________9_495682(.DIN1 (______9__22026), .DIN2
       (___9__9__39786), .Q (___9_9___39789));
  xor2s1 _____________495683(.DIN1 (___9_____39770), .DIN2
       (___9_____39735), .Q (___9_9___39788));
  xor2s1 _____________495684(.DIN1
       (______________________________________________21946), .DIN2
       (___9__9__39786), .Q (___9_90__39787));
  xor2s1 ______9______495685(.DIN1 (___9_____39755), .DIN2
       (___9_____39784), .Q (___9_____39785));
  xor2s1 _____________495686(.DIN1 (________26155), .DIN2
       (___9_____39774), .Q (___9_____39783));
  nor2s1 __________9__495687(.DIN1 (___9_____39763), .DIN2
       (___9_____39657), .Q (___9_____39782));
  nnd2s1 ___________0_495688(.DIN1 (___9_____39780), .DIN2
       (___9__9__39569), .Q (___9_____39781));
  xor2s1 _____9_______495689(.DIN1 (___9__0__39751), .DIN2
       (_____9___36360), .Q (___9_____39779));
  nnd2s1 ____________495690(.DIN1 (___0_90__40168), .DIN2
       (___9__9__39759), .Q (___9__0__39778));
  nnd2s1 ______9___0__495691(.DIN1 (___9__9__39668), .DIN2
       (___9__0__39760), .Q (___9__9__39777));
  nnd2s1 ___________0_495692(.DIN1 (___9_____39761), .DIN2
       (___9__0__39306), .Q (___9_____39776));
  hi1s1 ______495693(.DIN (___9_9___39792), .Q (___99____39809));
  and2s1 ___________9_495694(.DIN1 (___9_____39774), .DIN2
       (___9_____39773), .Q (___9_____39775));
  nor2s1 _____________495695(.DIN1 (________28259), .DIN2
       (___9_____39756), .Q (___9_____39772));
  nor2s1 ____________495696(.DIN1 (___9_____39733), .DIN2
       (___9_____39770), .Q (___9_____39771));
  nor2s1 ______9___0_495697(.DIN1 (___9_____39773), .DIN2
       (___9_____39774), .Q (___9_____39769));
  dffacs1 ______________________________________________9_495698(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39757), .Q
       (__________________________________________________________________22007));
  dffacs1 ________________________________________________495699(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39754), .QN
       (_________22022));
  xor2s1 _________990_495700(.DIN1 (___9_____39750), .DIN2
       (_________38463), .Q (___9_99__39796));
  xor2s1 ____________495701(.DIN1 (___9_____39740), .DIN2
       (___9_____39749), .Q (___990___39799));
  xor2s1 ___________9_495702(.DIN1 (___9_____39565), .DIN2
       (___9_____39762), .Q (___9_9___39792));
  xnr2s1 _____________495703(.DIN1 (___9_____39767), .DIN2
       (___0_99__40078), .Q (___9__9__39768));
  nnd2s1 _____0_______495704(.DIN1 (___9_____39765), .DIN2
       (___9_____39764), .Q (___9_____39766));
  xor2s1 ______9______495705(.DIN1 (___0_____40427), .DIN2
       (__________________________________________9___21947), .Q
       (___9_____39763));
  nnd2s1 _____________495706(.DIN1 (___9_____39758), .DIN2
       (___9__0__39315), .Q (___9_____39761));
  nnd2s1 ___________495707(.DIN1 (___9_____39667), .DIN2
       (___9_____39745), .Q (___9__0__39760));
  nor2s1 _____________495708(.DIN1 (___9_____39747), .DIN2
       (________23527), .Q (___9__9__39759));
  nor2s1 __________495709(.DIN1 (___09____40657), .DIN2
       (___9_____39758), .Q (___9_____39780));
  or2s1 _____9_____9_495710(.DIN1
       (__________________________________________9___21947), .DIN2
       (___0__0__39993), .Q (___9_____39757));
  and2s1 _____9_______495711(.DIN1 (___0_____40100), .DIN2
       (___0_____40601), .Q (___9_____39756));
  xor2s1 _____00______495712(.DIN1 (___9__0__39732), .DIN2
       (___9_____39718), .Q (___9_____39755));
  nor2s1 _____9_______495713(.DIN1 (________26698), .DIN2
       (__________________________________________9___21947), .Q
       (___9__9__39786));
  xor2s1 _____0_______495714(.DIN1 (___9_____39730), .DIN2
       (_________35523), .Q (___9_____39770));
  nnd2s1 __________9__495715(.DIN1 (___9_____39736), .DIN2 (___9_9), .Q
       (___9_____39754));
  nnd2s1 ___________0_495716(.DIN1 (___0_99__40078), .DIN2
       (___9_____39752), .Q (___9_____39753));
  nor2s1 ______0______495717(.DIN1 (___9_____39752), .DIN2
       (___0_99__40078), .Q (___9__0__39751));
  xor2s1 _____________495718(.DIN1 (___9_____39729), .DIN2
       (___9_9___39700), .Q (___9_____39774));
  nor2s1 ____________495719(.DIN1 (___9_____39748), .DIN2
       (___9__9__39741), .Q (___99____39846));
  nor2s1 ______0___0__495720(.DIN1 (___9__0__39713), .DIN2
       (___9_____39728), .Q (___9_____39750));
  nor2s1 ___________0_495721(.DIN1 (___9_____39725), .DIN2
       (___9_____39748), .Q (___9_____39749));
  xor2s1 ___________9_495722(.DIN1 (___9_____39716), .DIN2
       (_________38680), .Q (___9_____39765));
  and2s1 _____________495723(.DIN1 (___9_____39746), .DIN2
       (___0_____40610), .Q (___9_____39747));
  or2s1 ____________495724(.DIN1 (___0_____40610), .DIN2
       (_____9__25927), .Q (___9_____39745));
  nor2s1 ______9___0_495725(.DIN1 (___9_0___39534), .DIN2
       (___9_____39727), .Q (___9_____39762));
  nor2s1 ______9______495726(.DIN1 (___9_____39354), .DIN2
       (___9_____39723), .Q (___9_____39758));
  nor2s1 _____0___990_495727(.DIN1 (___9_____39743), .DIN2
       (___9__9__39722), .Q (___9_____39744));
  dffacs1 ________________________________________________495728(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39721), .Q (___0_____40601));
  nnd2s1 ______9_____495729(.DIN1 (___9_____39737), .DIN2
       (___9_____39738), .Q (___9__0__39742));
  dffacs1 ______________________________________________9_495730(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39720), .QN
       (__________________________________________9___21947));
  and2s1 ___________9_495731(.DIN1 (___9_____39724), .DIN2
       (___9_____39740), .Q (___9__9__39741));
  nor2s1 _____________495732(.DIN1 (___9_____39738), .DIN2
       (___9_____39737), .Q (___9_____39739));
  xor2s1 _____9_______495733(.DIN1 (___9_____39367), .DIN2
       (___0990__40710), .Q (___9_____39736));
  xnr2s1 ______0______495734(.DIN1 (___9_____39726), .DIN2
       (___9_____39583), .Q (___0_99__40078));
  nor2s1 _________9___495735(.DIN1 (___9_____39734), .DIN2
       (___9_____39733), .Q (___9_____39735));
  xor2s1 ______9______495736(.DIN1 (___9_____39717), .DIN2
       (___9__9__39731), .Q (___9__0__39732));
  nor2s1 ___________495737(.DIN1 (___9__9__39632), .DIN2
       (___9_0___39711), .Q (___9_____39730));
  xor2s1 _____________495738(.DIN1 (___09_0__40661), .DIN2
       (___9_____39627), .Q (___9_____39729));
  nnd2s1 __________495739(.DIN1 (___9_09__39712), .DIN2
       (___9_0___39707), .Q (___9_____39728));
  nor2s1 ___________9_495740(.DIN1 (___9_0___39530), .DIN2
       (___9_____39726), .Q (___9_____39727));
  hi1s1 ______9(.DIN (___9_____39724), .Q (___9_____39725));
  nor2s1 _____99______495741(.DIN1 (___9_____39355), .DIN2
       (___0990__40710), .Q (___9_____39723));
  dffacs1 ________________________________________________495742(.CLRB
       (reset), .CLK (clk), .DIN (___9_0___39708), .Q (___0_____40610));
  xor2s1 _____________495743(.DIN1 (___9_____39654), .DIN2
       (___9_0___39710), .Q (___9__9__39722));
  nnd2s1 _____________495744(.DIN1 (___9_00__39703), .DIN2
       (___0_90__40168), .Q (___9_____39721));
  nnd2s1 _____________495745(.DIN1 (___9_0___39704), .DIN2
       (________27201), .Q (___9_____39720));
  nor2s1 __________9__495746(.DIN1 (___9_____39718), .DIN2
       (___9_____39717), .Q (___9_____39719));
  nor2s1 ___________0_495747(.DIN1
       (______________________________________________21964), .DIN2
       (___9_____39715), .Q (___9_____39716));
  nnd2s1 _____________495748(.DIN1 (___9_____39715), .DIN2
       (___9_____39714), .Q (___9_____39724));
  nor2s1 _____________495749(.DIN1 (___9_____39714), .DIN2
       (___9_____39715), .Q (___9_____39748));
  nnd2s1 ____________495750(.DIN1 (___9_____39717), .DIN2
       (___9_____39718), .Q (___9_____39737));
  nnd2s1 __________0__495751(.DIN1 (___9_____39715), .DIN2
       (______________________________________________21964), .Q
       (___9_____39764));
  nor2s1 ______9____0_495752(.DIN1 (___9_0___39705), .DIN2
       (___9_0___39706), .Q (___9__0__39713));
  nnd2s1 ___________9_495753(.DIN1 (___9_____39685), .DIN2
       (___9_9___39702), .Q (___9_09__39712));
  and2s1 _____________495754(.DIN1 (___9_0___39710), .DIN2
       (___9_____39638), .Q (___9_0___39711));
  xor2s1 ____________495755(.DIN1 (___9__9__39694), .DIN2
       (___9_0___39709), .Q (___9_____39733));
  nnd2s1 _____00___0_495756(.DIN1 (___9_9___39697), .DIN2 (___9_9), .Q
       (___9_0___39708));
  nnd2s1 ______9______495757(.DIN1 (___9_0___39706), .DIN2
       (___9_0___39705), .Q (___9_0___39707));
  nor2s1 ____________495758(.DIN1 (___9_____39580), .DIN2
       (___9_9___39699), .Q (___9_____39726));
  nnd2s1 ___________9_495759(.DIN1 (___9_90__39695), .DIN2
       (___99____39819), .Q (___9_0___39704));
  xor2s1 _____________495760(.DIN1 (___9_____39691), .DIN2
       (___9_____39319), .Q (___9_00__39703));
  xor2s1 _____________495761(.DIN1 (___9_____39692), .DIN2
       (___9_____39399), .Q (___9_____39717));
  xor2s1 _________9___495762(.DIN1 (___9_9___39608), .DIN2
       (___9_9___39698), .Q (___9_____39715));
  nnd2s1 _____9_______495763(.DIN1 (___9_9___39701), .DIN2
       (___9_9___39700), .Q (___9_9___39702));
  and2s1 _____9_____495764(.DIN1 (___9_9___39698), .DIN2
       (___9__0__39578), .Q (___9_9___39699));
  nor2s1 _____________495765(.DIN1 (___9_____39596), .DIN2
       (___9_____39690), .Q (___9_0___39710));
  xor2s1 __________495766(.DIN1 (___9_____39684), .DIN2
       (___9_9___39696), .Q (___9_9___39697));
  nor2s1 _____9_______495767(.DIN1 (___9_9___39700), .DIN2
       (___9_9___39701), .Q (___9_0___39706));
  xor2s1 _____________495768(.DIN1 (___9_____39639), .DIN2
       (___9_____39689), .Q (___9_90__39695));
  nor2s1 _____________495769(.DIN1
       (__________________________________________________________________21994),
       .DIN2 (___9_____39693), .Q (___9_____39734));
  nnd2s1 _____________495770(.DIN1 (___9_____39693), .DIN2
       (__________________________________________________________________21994),
       .Q (___9__9__39694));
  nor2s1 _____9____9__(.DIN1 (___9_____39393), .DIN2 (___9__9__39686),
       .Q (___990___39798));
  xor2s1 _____9_____0_495771(.DIN1 (___9_____39398), .DIN2
       (___0__0__40333), .Q (___9_____39692));
  xor2s1 _____________495772(.DIN1 (___9_____39681), .DIN2
       (__________________________________________________________________21999),
       .Q (___9_____39691));
  nor2s1 _____________495773(.DIN1 (___9_____39594), .DIN2
       (___9_____39689), .Q (___9_____39690));
  nnd2s1 _____0______495774(.DIN1 (___9_____39682), .DIN2
       (___9_____39655), .Q (___9_9___39698));
  dffacs1 ________________________________________________495775(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39683), .Q
       (______________________________________________21945));
  xor2s1 _____0_____9_495776(.DIN1 (___9__0__39679), .DIN2
       (____9____38944), .Q (___9_9___39701));
  and2s1 _____0_______495777(.DIN1 (___0__0__40333), .DIN2
       (___9_____39400), .Q (___9__9__39686));
  xor2s1 _____0______495778(.DIN1 (___9_____39671), .DIN2
       (___9_____39675), .Q (___9_____39693));
  xor2s1 __________0_495779(.DIN1 (___9__0__41371), .DIN2
       (___099___40714), .Q (___9_____39684));
  dffacs1 ________________________________________________495780(.CLRB
       (reset), .CLK (clk), .DIN (___9__9__39678), .QN
       (______________________________________________21922));
  xnr2s1 _____________495781(.DIN1 (_________41252), .DIN2
       (___099___40712), .Q (___9_9___39700));
  dffacs1 ______________________________________________9_495782(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39677), .Q
       (__________________________________________9___21918));
  nnd2s1 ______0__990_495783(.DIN1 (___9_____39447), .DIN2
       (___9_____39672), .Q (___9_____39683));
  nor2s1 ____________495784(.DIN1 (___9_____39680), .DIN2
       (___9_____39674), .Q (___9_____39689));
  xor2s1 ___________9_495785(.DIN1 (___9_____39664), .DIN2
       (___9_____39397), .Q (___9_____39682));
  nnd2s1 _____________495786(.DIN1 (___9_____39676), .DIN2
       (___9_____39670), .Q (___9_____39685));
  nor2s1 _____________495787(.DIN1 (___9_____39144), .DIN2
       (___099___40714), .Q (___9__0__39687));
  or2s1 _____0_______495788(.DIN1 (___9_____39680), .DIN2
       (___9_____39673), .Q (___9_____39681));
  xor2s1 ______9__9___(.DIN1 (___9_____39649), .DIN2 (___9__9__39650),
       .Q (___9__0__39679));
  xor2s1 _____________495789(.DIN1 (___9_____39656), .DIN2
       (___9_____39663), .Q (___0__0__40333));
  nnd2s1 ___________495790(.DIN1 (___9__0__39660), .DIN2
       (________25464), .Q (___9__9__39678));
  nnd2s1 _____________495791(.DIN1 (___9_____39661), .DIN2
       (___9_____39630), .Q (___9_____39677));
  dffacs1 ________________________________________________495792(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39662), .Q
       (______________________________________________21915));
  nnd2s1 ______9___495793(.DIN1 (___9__0__39669), .DIN2
       (___9_____39675), .Q (___9_____39676));
  nor2s1 _____9_____9_495794(.DIN1
       (__________________________________________________________________21999),
       .DIN2 (___9_____39673), .Q (___9_____39674));
  nnd2s1 _____________495795(.DIN1 (___9_____39658), .DIN2
       (inData[30]), .Q (___9_____39672));
  and2s1 ______0______495796(.DIN1 (___9_____39670), .DIN2
       (___9__0__39669), .Q (___9_____39671));
  or2s1 _____________495797(.DIN1 (___9_____39667), .DIN2
       (___9_____39646), .Q (___9__9__39668));
  nor2s1 ___________0_495798(.DIN1 (___9_____39647), .DIN2
       (___9__0__39651), .Q (___9_____39718));
  dffacs1 ________________________________________________495799(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39645), .Q
       (__________________________________________________________________21994));
  nor2s1 _____0_______495800(.DIN1 (___9__0__39643), .DIN2
       (___9_____39665), .Q (___9_____39666));
  or2s1 _____________495801(.DIN1 (___9_____39635), .DIN2
       (___9_____39663), .Q (___9_____39664));
  nor2s1 _____09_____0(.DIN1 (___9_____39466), .DIN2 (___9__9__39642),
       .Q (___9_____39680));
  nnd2s1 ______0___0__495802(.DIN1 (___9_____39631), .DIN2
       (___9_____39628), .Q (___9_____39662));
  nor2s1 ___________0_495803(.DIN1 (___9_____39629), .DIN2
       (___9_____39636), .Q (___9_____39661));
  nnd2s1 ______9____9_495804(.DIN1 (___9__0__39633), .DIN2
       (___9__9__39659), .Q (___9__0__39660));
  dffacs1 __________________________________________0_____(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39640), .Q (___0__9__40440));
  nor2s1 _____9_______495805(.DIN1 (___9_____39626), .DIN2
       (___9_____39657), .Q (___9_____39658));
  and2s1 ____________495806(.DIN1 (___9_____39634), .DIN2
       (___9_____39655), .Q (___9_____39656));
  xor2s1 __________0_495807(.DIN1 (________22470), .DIN2
       (___9_____39637), .Q (___9_____39654));
  nnd2s1 _____________495808(.DIN1 (___9_____39652), .DIN2
       (___9_____39653), .Q (___9_____39670));
  or2s1 _________990_495809(.DIN1 (___9_____39653), .DIN2
       (___9_____39652), .Q (___9__0__39669));
  nor2s1 _____0______495810(.DIN1 (___9_____39467), .DIN2
       (___9_____39641), .Q (___9_____39673));
  nor2s1 _____________495811(.DIN1 (___9__9__39650), .DIN2
       (___9_____39648), .Q (___9__0__39651));
  nor2s1 _____________495812(.DIN1 (___9_____39648), .DIN2
       (___9_____39647), .Q (___9_____39649));
  xor2s1 ______0______495813(.DIN1 (___9_9___39612), .DIN2
       (______________________________________________21905), .Q
       (___9_____39646));
  nnd2s1 _____9_______495814(.DIN1 (___9_0___39618), .DIN2
       (___9_____39644), .Q (___9_____39645));
  hi1s1 _______495815(.DIN (___9_____39641), .Q (___9__9__39642));
  nnd2s1 ___________495816(.DIN1 (___9_99__39616), .DIN2
       (___9_____39548), .Q (___9_____39640));
  xor2s1 _____________495817(.DIN1 (___9_9___39609), .DIN2
       (_________38860), .Q (___9_____39639));
  or2s1 __________495818(.DIN1
       (__________________________________________0___21935), .DIN2
       (___9_____39637), .Q (___9_____39638));
  nor2s1 ___________9_495819(.DIN1 (___9_9___39615), .DIN2
       (_____99__38418), .Q (___9_____39665));
  nnd2s1 _____9_______495820(.DIN1 (___9__0__39352), .DIN2
       (___9_9___39613), .Q (___9_____39636));
  hi1s1 _______495821(.DIN (___9_____39634), .Q (___9_____39635));
  xor2s1 ______9______495822(.DIN1 (___9_____39605), .DIN2
       (___99_9__39836), .Q (___9__0__39633));
  and2s1 _____________495823(.DIN1 (___9_____39637), .DIN2
       (__________________________________________0___21935), .Q
       (___9__9__39632));
  and2s1 _____9_______495824(.DIN1 (___909___39064), .DIN2
       (___9_____39630), .Q (___9_____39631));
  nor2s1 _____9____9__495825(.DIN1 (______22125), .DIN2
       (___9_____39628), .Q (___9_____39629));
  xor2s1 ______9____0_495826(.DIN1 (___099___40716), .DIN2
       (___9_____39627), .Q (___9_____39663));
  xor2s1 _____________495827(.DIN1 (___9__0__39598), .DIN2
       (___9_9___39425), .Q (___9_____39626));
  xnr2s1 ______0_____495828(.DIN1 (_________38666), .DIN2
       (___9__9__39597), .Q (___9_____39641));
  xor2s1 __________0__495829(.DIN1 (___9_____39589), .DIN2
       (___9__9__39125), .Q (___9_____39653));
  xor2s1 ___________0_495830(.DIN1 (___9_____39590), .DIN2
       (___9_____39461), .Q (___9_____39634));
  nor2s1 ___________9_495831(.DIN1 (___0_____40422), .DIN2
       (_____9___38413), .Q (___9__0__39643));
  nor2s1 __________0_495832(.DIN1 (___9_0___39622), .DIN2
       (___9_0___39621), .Q (___9_0___39623));
  nor2s1 ____9____990_(.DIN1 (_____0__26195), .DIN2 (___9_____39604),
       .Q (___9_0___39618));
  and2s1 ____________495833(.DIN1 (___0_____40035), .DIN2
       (___9_00__39617), .Q (___9_____39648));
  nor2s1 ___________9_495834(.DIN1 (___9_00__39617), .DIN2
       (___0_____40035), .Q (___9_____39647));
  and2s1 ______0______495835(.DIN1 (___9_____39593), .DIN2
       (________25662), .Q (___9_99__39616));
  hi1s1 _______495836(.DIN (___0_____40422), .Q (___9_9___39615));
  nnd2s1 _____________495837(.DIN1 (___9_____39592), .DIN2
       (___99____39819), .Q (___9_9___39614));
  xor2s1 _____________495838(.DIN1 (___9_____39585), .DIN2
       (___9__0__39507), .Q (___9_____39637));
  nnd2s1 ____9_9__9___(.DIN1 (___9_9___39611), .DIN2 (___9__0__39588),
       .Q (___9_9___39613));
  xor2s1 ____9________(.DIN1 (___9_____39602), .DIN2 (___9_0___39349),
       .Q (___9_9___39612));
  nnd2s1 ___________495839(.DIN1 (___9_____39591), .DIN2
       (___9_____39551), .Q (___9_____39652));
  nnd2s1 ____9________495840(.DIN1 (___9_9___39611), .DIN2
       (___9__9__39587), .Q (___9_____39630));
  or2s1 ____9_____900(.DIN1 (___9_____39586), .DIN2 (___9_9___39610),
       .Q (___9_____39628));
  xor2s1 ______0____9_495841(.DIN1 (___9_____39595), .DIN2
       (________23832), .Q (___9_9___39609));
  xor2s1 _____________495842(.DIN1 (___9_90__39607), .DIN2
       (___9_____39579), .Q (___9_9___39608));
  dffacs1 ________________________________________________495843(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39576), .QN
       (___0_____40422));
  nnd2s1 ____90_______(.DIN1 (___9_____39603), .DIN2 (___90____39028),
       .Q (___9_____39655));
  nor2s1 ____90_______495844(.DIN1 (___9_____39557), .DIN2
       (___9_____39574), .Q (___9_09__39625));
  hi1s1 ____90_(.DIN (___9__9__39606), .Q (___0_____40035));
  xor2s1 ____9_____9__(.DIN1 (___9_____39568), .DIN2 (___9__9__39218),
       .Q (___9_____39605));
  nor2s1 ____9______0_(.DIN1 (___9_____39573), .DIN2 (___00_0__39902),
       .Q (___9_____39604));
  nor2s1 ____90_______495845(.DIN1 (___99____39808), .DIN2
       (___9_____39603), .Q (___9_0___39621));
  nor2s1 ____9________495846(.DIN1 (___9_____39097), .DIN2
       (___9_____39602), .Q (___9_0___39620));
  dffacs1 __________________________________________0_____495847(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39581), .QN
       (______________________________________0_______21894));
  nor2s1 ____________495848(.DIN1 (___9_____39600), .DIN2
       (___9_____39599), .Q (___9_____39601));
  xor2s1 __________0__495849(.DIN1 (___0_____40428), .DIN2
       (_________22025), .Q (___9__0__39598));
  nor2s1 ___________0_495850(.DIN1 (___9_____39504), .DIN2
       (___9_____39571), .Q (___9__9__39597));
  nor2s1 ___________9_495851(.DIN1
       (__________________________________________9___21934), .DIN2
       (___9_____39595), .Q (___9_____39596));
  and2s1 ______9______495852(.DIN1 (___9_____39595), .DIN2
       (__________________________________________9___21934), .Q
       (___9_____39594));
  nor2s1 ____________495853(.DIN1 (________27070), .DIN2
       (___9__0__39570), .Q (___9_____39593));
  xor2s1 ______0___0_9(.DIN1 (___9_9___39524), .DIN2 (___9__9__39560),
       .Q (___9_____39592));
  nor2s1 _____9_______495854(.DIN1 (___9__9__39552), .DIN2
       (___9_____39567), .Q (___9_____39591));
  nnd2s1 ____90___990_(.DIN1 (___9_____39572), .DIN2 (___900___38981),
       .Q (___9_____39590));
  xor2s1 ____90______0(.DIN1 (___9_____39558), .DIN2 (___9_09__39535),
       .Q (___9_____39589));
  nor2s1 ____9______9_(.DIN1
       (__________________________________________9___21918), .DIN2
       (______________________________________________21920), .Q
       (___9__0__39588));
  nor2s1 ____9_0______(.DIN1
       (______________________________________________21917), .DIN2
       (______________________________________________21920), .Q
       (___9__9__39587));
  nnd2s1 ____9________495855(.DIN1
       (______________________________________________21920), .DIN2
       (______________________________________________21917), .Q
       (___9_____39586));
  or2s1 _____9_______495856(.DIN1 (___9_0___39532), .DIN2
       (___9_____39767), .Q (___9_____39740));
  xor2s1 ____9____9___(.DIN1 (___9_____39562), .DIN2 (_________37452),
       .Q (___9__9__39606));
  xor2s1 ____9_0______495857(.DIN1 (___9__0__39498), .DIN2
       (___9_____39566), .Q (___9_____39585));
  xor2s1 ___________495858(.DIN1 (___9_____39540), .DIN2
       (___9_9___39518), .Q (___9_____39584));
  xor2s1 _____________495859(.DIN1 (___9_____39541), .DIN2
       (___9_____39582), .Q (___9_____39583));
  nnd2s1 _____9____495860(.DIN1 (___9_____39559), .DIN2
       (_____0__25688), .Q (___9_____39581));
  nor2s1 ____90_____9_(.DIN1 (___9_____39579), .DIN2 (___9__9__39577),
       .Q (___9_____39580));
  nnd2s1 ____90_______495861(.DIN1 (___9__9__39577), .DIN2
       (___9_____39579), .Q (___9__0__39578));
  or2s1 _____________495862(.DIN1 (_________22025), .DIN2
       (___9_____39575), .Q (___9_____39576));
  xor2s1 ____9________495863(.DIN1 (___9_0___39529), .DIN2
       (____9____38944), .Q (___9_____39574));
  hi1s1 ____9_9(.DIN
       (______________________________________________21920), .Q
       (___9_____39573));
  hi1s1 ____9__(.DIN (___9_____39572), .Q (___9_____39603));
  nor2s1 ____9_____9__495864(.DIN1 (____99___38976), .DIN2
       (___9_____39556), .Q (___9_____39602));
  xor2s1 ____9______0_495865(.DIN1 (___9_____39563), .DIN2
       (_____0___38422), .Q (___9_0___39622));
  dffacs1 __________________________________________0_____495866(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39549), .QN
       (___0_____40617));
  xor2s1 _____________495867(.DIN1 (___9_9___39525), .DIN2
       (_____00__35736), .Q (___9_____39571));
  nor2s1 ____900______(.DIN1 (____0___25683), .DIN2 (___9__0__39544),
       .Q (___9__0__39570));
  xor2s1 ____9_______0(.DIN1 (___9__9__39516), .DIN2 (___9__9__39569),
       .Q (___9_____39600));
  xor2s1 ____9_____0__(.DIN1 (___9_____39510), .DIN2 (_____9___38611),
       .Q (___9_____39599));
  xor2s1 ____9______0_495868(.DIN1 (___9_____39475), .DIN2
       (___9_____39512), .Q (___9_____39595));
  nor2s1 ____9______9_495869(.DIN1 (___9__9__39324), .DIN2
       (___9__9__39543), .Q (___9_____39767));
  xor2s1 ____00_______(.DIN1 (___9_____39555), .DIN2
       (_______________________________________________________________9),
       .Q (___9_____39568));
  nor2s1 ____9_______495870(.DIN1 (___9_____39499), .DIN2
       (___9_____39566), .Q (___9_____39567));
  nor2s1 ____9_____0_9(.DIN1 (___9_____39564), .DIN2 (___9_____39545),
       .Q (___9_____39565));
  nor2s1 ____9_0______495871(.DIN1 (___9_9___39523), .DIN2
       (___9_____39563), .Q (___9_____39572));
  hi1s1 ____9_495872(.DIN (___9__9__39577), .Q (___9_90__39607));
  nor2s1 ____9____990_495873(.DIN1 (___9_09__39442), .DIN2
       (___9_0___39531), .Q (___9_____39675));
  dffacs1 ________________________________________________495874(.CLRB
       (reset), .CLK (clk), .DIN (___9_0___39528), .QN
       (______________________________________________21920));
  xor2s1 ____9_______495875(.DIN1 (___9_____39496), .DIN2
       (___9__9__39506), .Q (___9_____39562));
  xnr2s1 ___________9_495876(.DIN1 (____9_9__38931), .DIN2
       (___9_____39505), .Q (___9__9__39560));
  nor2s1 ____9________495877(.DIN1 (________25529), .DIN2
       (___9_9___39521), .Q (___9_____39559));
  xor2s1 ____9________495878(.DIN1 (___9_____39557), .DIN2
       (___9_____39546), .Q (___9_____39558));
  dffacs1 ________________________________________________495879(.CLRB
       (reset), .CLK (clk), .DIN (___9_99__39526), .Q (_________22025));
  nnd2s1 ____9________495880(.DIN1 (___9_9___39520), .DIN2
       (___9_____39383), .Q (___9__9__39577));
  and2s1 ____00___9___(.DIN1 (___9_____39555), .DIN2 (___9000__38978),
       .Q (___9_____39556));
  nor2s1 ____99_______(.DIN1 (___9_9___39790), .DIN2 (___9_____39550),
       .Q (___9__9__39552));
  nnd2s1 ____99____900(.DIN1 (___9_____39550), .DIN2 (___9_9___39790),
       .Q (___9_____39551));
  nnd2s1 ____00_____9_(.DIN1 (___9_____39508), .DIN2 (___9_____39548),
       .Q (___9_____39549));
  xor2s1 ____9________495881(.DIN1 (___9_____39546), .DIN2
       (______________________________________________21961), .Q
       (___9_____39547));
  xor2s1 ____9_0______495882(.DIN1 (___9_____39472), .DIN2
       (___0_9___40645), .Q (___9__0__39544));
  xor2s1 ____9________495883(.DIN1 (___0_9___40645), .DIN2
       (___9_____39542), .Q (___9__9__39543));
  xor2s1 ____9________495884(.DIN1 (___9_0___39533), .DIN2
       (___0_9___40645), .Q (___9_____39541));
  xor2s1 ____9_9___9__(.DIN1 (___9_____39539), .DIN2 (___0_9___40645),
       .Q (___9_____39540));
  nnd2s1 ____9______0_495885(.DIN1 (___9_00__39527), .DIN2
       (___9_9___39696), .Q (___9_____39538));
  nor2s1 ____9________495886(.DIN1 (___9_____39474), .DIN2
       (___9_____39502), .Q (___9_____39566));
  nnd2s1 _____90______495887(.DIN1 (___9_____39537), .DIN2
       (___099___40718), .Q (___9__0__39561));
  nor2s1 ____9_______495888(.DIN1 (___9_00__39527), .DIN2
       (___9_____39454), .Q (___9_____39563));
  nnd2s1 ____00____0__(.DIN1 (___9_____39546), .DIN2 (___9_09__39535),
       .Q (___9__0__39536));
  and2s1 ____9______0_495889(.DIN1 (___9_00__39527), .DIN2
       (___9_0___39533), .Q (___9_0___39534));
  nor2s1 ____9______9_495890(.DIN1 (___9__9__39305), .DIN2
       (___9_00__39527), .Q (___9_0___39532));
  nor2s1 ____999______(.DIN1 (___9_____39511), .DIN2 (___9__9__39497),
       .Q (___9_0___39531));
  nor2s1 ____9_______495891(.DIN1 (___9_0___39533), .DIN2
       (___9_00__39527), .Q (___9_0___39530));
  or2s1 ____00____0_9(.DIN1 (___9_09__39535), .DIN2 (___9_____39546),
       .Q (___9_0___39529));
  nnd2s1 ____00_______495892(.DIN1 (___9_____39500), .DIN2
       (___9_____39329), .Q (___9_0___39528));
  nor2s1 ____9____990_495893(.DIN1 (___9_____39278), .DIN2
       (___9_00__39527), .Q (___9_____39564));
  dffacs1 _________________________________________9_____(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39503), .QN
       (_____________________________________9_______21884));
  nnd2s1 _____99_____495894(.DIN1 (___9_____39491), .DIN2 (___9_9), .Q
       (___9_99__39526));
  dffacs1 ________________(.CLRB (reset), .CLK (clk), .DIN
       (___9_____39490), .Q (outData[31]));
  nnd2s1 ____9______9_495895(.DIN1 (___9_____39493), .DIN2
       (___9_9___39524), .Q (___9_9___39525));
  nor2s1 ____9________495896(.DIN1 (___99____39808), .DIN2
       (___9_____39453), .Q (___9_9___39523));
  nnd2s1 ____9________495897(.DIN1 (___0_9___40645), .DIN2
       (______________________________________________21906), .Q
       (___9_9___39522));
  nor2s1 ____9_9______(.DIN1 (___99____39808), .DIN2 (___9__0__39460),
       .Q (___9_9___39521));
  nnd2s1 ____9____9___495898(.DIN1 (___9_____39381), .DIN2
       (___0_9___40645), .Q (___9_9___39520));
  nnd2s1 ____9________495899(.DIN1 (___9_9___39518), .DIN2
       (___0_9___40645), .Q (___9_9___39519));
  nor2s1 ____9______09(.DIN1 (___0_9___40645), .DIN2 (___9_9___39518),
       .Q (___9_90__39517));
  nor2s1 ____9________495900(.DIN1 (___99____39808), .DIN2
       (___9_____39509), .Q (___9__9__39516));
  nnd2s1 ____9_____495901(.DIN1 (___9_____39513), .DIN2
       (______________________________________________21961), .Q
       (___9_____39515));
  nor2s1 ____9______9_495902(.DIN1
       (______________________________________________21961), .DIN2
       (___9_____39513), .Q (___9_____39514));
  xnr2s1 ____9________495903(.DIN1 (___9_____39511), .DIN2
       (___9_____39501), .Q (___9_____39512));
  nnd2s1 ____9_9______495904(.DIN1 (___9_____39509), .DIN2
       (___99____39808), .Q (___9_____39510));
  and2s1 ____0_9______495905(.DIN1 (___9_____39483), .DIN2
       (____0___25682), .Q (___9_____39508));
  nor2s1 ____9________495906(.DIN1 (___9_0___39256), .DIN2
       (___99____39808), .Q (___9_____39545));
  nor2s1 ____0_____9__495907(.DIN1 (___9_____39463), .DIN2
       (___9__0__39507), .Q (___9_____39550));
  nnd2s1 ____0______0_495908(.DIN1 (___9__9__39506), .DIN2
       (___9__0__39488), .Q (___9__0__39553));
  nnd2s1 ____0________495909(.DIN1 (___9_____39489), .DIN2
       (____9_9__38968), .Q (___9_____39555));
  dffacs1 __________________________________________0_____495910(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39485), .Q (___0_____40616));
  dffacs1 ________________________________________________495911(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39495), .Q
       (__________________________________________________________________22002));
  nor2s1 ____9________495912(.DIN1 (___9_____39504), .DIN2
       (___9_____39492), .Q (___9_____39505));
  nnd2s1 ____9_______495913(.DIN1 (___9_____39184), .DIN2
       (___9_____39482), .Q (___9_____39503));
  xor2s1 ____909___0__(.DIN1 (___9__9__39478), .DIN2 (_________38869),
       .Q (___9_____39537));
  hi1s1 ____99_(.DIN (___9_____39490), .Q (___9_00__39527));
  nor2s1 ____99_____0_(.DIN1 (___9_____39476), .DIN2 (___9_____39501),
       .Q (___9_____39502));
  or2s1 ____0______9_495914(.DIN1 (___9_____39667), .DIN2
       (___9_____39480), .Q (___9_____39500));
  nor2s1 ____0________495915(.DIN1 (___9__0__39498), .DIN2
       (___09____40662), .Q (___9_____39499));
  nnd2s1 ____0_______495916(.DIN1 (___9_____39481), .DIN2
       (___9__0__39443), .Q (___9__9__39497));
  xor2s1 ____0_____0_495917(.DIN1 (___9_____39509), .DIN2
       (___9__9__39487), .Q (___9_____39496));
  hi1s1 ____0__495918(.DIN (___9_____39513), .Q (___9_____39546));
  nnd2s1 ____9________495919(.DIN1 (___9__0__39479), .DIN2
       (___9_____39494), .Q (___9_____39495));
  hi1s1 ____9_495920(.DIN (___9_____39492), .Q (___9_____39493));
  nor2s1 ____9____990_495921(.DIN1 (___9_____39477), .DIN2
       (____99___38974), .Q (___9_____39491));
  xor2s1 ____0_______495922(.DIN1 (___9_9___39429), .DIN2
       (___9_____39462), .Q (___9_____39513));
  nb1s1 ____990(.DIN (___9_____39490), .Q (___99____39808));
  xor2s1 ____0_9____9_495923(.DIN1 (___9_____39456), .DIN2
       (____9____38944), .Q (___9_____39489));
  or2s1 ____0________495924(.DIN1 (___9__9__39487), .DIN2
       (___9_____39509), .Q (___9__0__39488));
  and2s1 ____0________495925(.DIN1 (___9_____39509), .DIN2
       (___9__9__39487), .Q (___9_____39486));
  nnd2s1 ____0________495926(.DIN1 (___9_____39471), .DIN2
       (___9____25086), .Q (___9_____39485));
  or2s1 ____0____9___495927(.DIN1 (___9_____39667), .DIN2
       (___9_____39470), .Q (___9_____39484));
  nnd2s1 ____0________495928(.DIN1 (___9_____39473), .DIN2
       (___9_90__39245), .Q (___9_____39483));
  hi1s1 ____0__495929(.DIN (___09____40662), .Q (___9__0__39507));
  nnd2s1 ____00_____09(.DIN1 (___9_____39468), .DIN2 (___9____24154),
       .Q (___9_____39482));
  xor2s1 ____9________495930(.DIN1 (___9_____39449), .DIN2
       (___9_9___39790), .Q (___9_____39492));
  xor2s1 ____00_____9_495931(.DIN1 (___9__9__39450), .DIN2
       (___9_____39295), .Q (___9_____39490));
  nnd2s1 ____0________495932(.DIN1 (___9_____39465), .DIN2
       (_________41264), .Q (___9_____39481));
  xor2s1 ____0_0______495933(.DIN1 (___9_0___39437), .DIN2
       (___9_0___39170), .Q (___9_____39480));
  nor2s1 ____0________495934(.DIN1 (___9_____39375), .DIN2
       (___9__9__39469), .Q (___9_____39501));
  nor2s1 ____99____9__(.DIN1 (________28415), .DIN2 (___9_____39448),
       .Q (___9__0__39479));
  nnd2s1 ____9______0_495935(.DIN1 (_________38733), .DIN2
       (__________________________________________________________________22004),
       .Q (___9__9__39478));
  nor2s1 ____9________495936(.DIN1 (___09____40663), .DIN2
       (_________38838), .Q (___9_____39477));
  xor2s1 ____0_9______495937(.DIN1 (___9_____39451), .DIN2
       (___9_0___39624), .Q (___9_____39476));
  nor2s1 ____0_0_____495938(.DIN1 (___9_____39474), .DIN2
       (___9_____39452), .Q (___9_____39475));
  nnd2s1 ____0_____0__495939(.DIN1 (___9_____39472), .DIN2
       (___9_0___39439), .Q (___9_____39473));
  nnd2s1 ____0______0_495940(.DIN1 (___9_0___39440), .DIN2
       (___9__9__39459), .Q (___9_____39471));
  xor2s1 ____0______9_495941(.DIN1 (___90_0__39005), .DIN2
       (___9_____39455), .Q (___9_____39470));
  dffacs1 ________________495942(.CLRB (reset), .CLK (clk), .DIN
       (___9_0___39441), .Q (outData[17]));
  xor2s1 ____0________495943(.DIN1 (____000__40720), .DIN2
       (___99_0__39827), .Q (___9_____39509));
  nnd2s1 ____0_______495944(.DIN1 (___9_0___39435), .DIN2
       (___9_____39374), .Q (___9__9__39469));
  nnd2s1 ____0_____0_495945(.DIN1 (___9_00__39433), .DIN2
       (___9_0___39436), .Q (___9_____39468));
  hi1s1 ____0__495946(.DIN (___9_____39466), .Q (___9_____39467));
  nor2s1 ____0________495947(.DIN1 (___9_____39464), .DIN2
       (___9_____39444), .Q (___9_____39465));
  hi1s1 ____0__495948(.DIN (___9_____39463), .Q (___9__0__39498));
  xor2s1 ____0____990_495949(.DIN1 (___9__9__39423), .DIN2
       (___9_____39461), .Q (___9_____39462));
  nnd2s1 ____0_______495950(.DIN1 (___9_____39472), .DIN2
       (___9__9__39459), .Q (___9__0__39460));
  nor2s1 ____0______9_495951(.DIN1 (___9_____39457), .DIN2
       (___9_____39445), .Q (___9_____39458));
  nor2s1 ______0______495952(.DIN1 (___90_9__39004), .DIN2
       (___9_____39455), .Q (___9_____39456));
  hi1s1 ____0__495953(.DIN (___9_____39453), .Q (___9_____39454));
  nnd2s1 ____0________495954(.DIN1 (___9_9___39430), .DIN2
       (___9_____39413), .Q (___9__9__39506));
  hi1s1 ____0__495955(.DIN (___9_____39451), .Q (___9_____39452));
  xor2s1 ____0____9___495956(.DIN1 (_________22037), .DIN2
       (___0_____40445), .Q (___9__9__39450));
  nnd2s1 ____0_0______495957(.DIN1 (___9_____39446), .DIN2
       (_________22023), .Q (___9_____39449));
  nor2s1 ____0______495958(.DIN1 (___0_____40606), .DIN2
       (___0_____40115), .Q (___9_____39448));
  nnd2s1 ____0_0______495959(.DIN1 (___9_9___39426), .DIN2
       (___99____39819), .Q (___9_____39447));
  xor2s1 ____0_____495960(.DIN1 (___9__9__39405), .DIN2
       (___9_0___39434), .Q (___9_____39466));
  dffacs1 ________________________________________________495961(.CLRB
       (reset), .CLK (clk), .DIN (___9_9___39427), .QN
       (__________________________________________________________________22004));
  nor2s1 ____009____9_(.DIN1 (_________22023), .DIN2 (___9_____39446),
       .Q (___9_____39504));
  nor2s1 ____0________495962(.DIN1 (___9_____39204), .DIN2
       (___9_____39419), .Q (___9__0__39443));
  and2s1 ____0________495963(.DIN1 (___9_____39421), .DIN2
       (___9_____39511), .Q (___9_09__39442));
  nnd2s1 ____0________495964(.DIN1 (_________37595), .DIN2
       (___9_9___39428), .Q (___9_0___39441));
  nnd2s1 _____0_______495965(.DIN1 (___9_0___39438), .DIN2
       (___9_09__39351), .Q (___9_0___39440));
  nnd2s1 _____0____9__495966(.DIN1 (___9_0___39438), .DIN2
       (___99_0__39827), .Q (___9_0___39439));
  xor2s1 ___________0_495967(.DIN1 (___9_____39411), .DIN2
       (___9_____39414), .Q (___9_0___39437));
  nnd2s1 ____0________495968(.DIN1 (___9_90__39424), .DIN2
       (___90____39042), .Q (___9_____39463));
  nnd2s1 ____0_9______495969(.DIN1 (___9_____39422), .DIN2
       (___9_____39394), .Q (___9_____39453));
  or2s1 ____0_______495970(.DIN1 (_________22037), .DIN2
       (___9_____39283), .Q (___9_0___39436));
  nnd2s1 ____0_____0__495971(.DIN1 (___9_0___39434), .DIN2
       (___9_0___39343), .Q (___9_0___39435));
  nnd2s1 ____0______0_495972(.DIN1 (________25395), .DIN2
       (_________22037), .Q (___9_00__39433));
  nnd2s1 ____0______9_495973(.DIN1 (___9_____39417), .DIN2
       (___9_____39365), .Q (___9_9___39524));
  nor2s1 ____0________495974(.DIN1 (___9_9___39431), .DIN2
       (___9_99__39432), .Q (___9_____39474));
  nnd2s1 ____0_______495975(.DIN1 (___9_99__39432), .DIN2
       (___9_9___39431), .Q (___9_____39451));
  nnd2s1 ____09____0_9(.DIN1 (___9_9___39429), .DIN2 (___9_____39402),
       .Q (___9_9___39430));
  nor2s1 _____00__990_(.DIN1
       (______________________________________________21960), .DIN2
       (___9_____39412), .Q (___9_____39445));
  xor2s1 ____090_____0(.DIN1 (___9_____39420), .DIN2 (___9_____39207),
       .Q (___9_____39444));
  nor2s1 ___________9_495976(.DIN1 (___9_____39409), .DIN2
       (___9__9__39415), .Q (___9_____39455));
  nnd2s1 _____________495977(.DIN1 (___9_____39418), .DIN2
       (___9_____39752), .Q (___9_____39472));
  nnd2s1 ____09_______495978(.DIN1 (___9_9___39339), .DIN2
       (___9_____39408), .Q (___9_9___39428));
  nnd2s1 ____0________495979(.DIN1 (______9__38496), .DIN2
       (___0__0__40609), .Q (___9_9___39427));
  dffacs1 ________________________________________________495980(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39407), .QN
       (___0_____40606));
  xor2s1 ____0_9__9___(.DIN1 (___9_____39376), .DIN2 (___9_____39416),
       .Q (___9_9___39426));
  nnd2s1 ____0________495981(.DIN1 (___0__0__40609), .DIN2
       (______________________________________________21945), .Q
       (___9_9___39425));
  nor2s1 ____0_0____09(.DIN1 (___9_____39356), .DIN2 (___9_____39404),
       .Q (___9_90__39424));
  xor2s1 ____0________495982(.DIN1 (___9_____39391), .DIN2
       (___9_0___39619), .Q (___9_____39446));
  xor2s1 __________495983(.DIN1 (___9_9___39518), .DIN2
       (___9_____39401), .Q (___9__9__39423));
  nnd2s1 _____0_____9_495984(.DIN1 (___9__0__39396), .DIN2
       (___99_0__39827), .Q (___9_____39422));
  nor2s1 _____0_______495985(.DIN1 (___9_____39188), .DIN2
       (___9_____39420), .Q (___9_____39421));
  nor2s1 _____0_______495986(.DIN1 (___9_____39208), .DIN2
       (___9_____39420), .Q (___9_____39419));
  nor2s1 _____0_______495987(.DIN1 (_____9__22577), .DIN2
       (___9_____39420), .Q (___9_____39457));
  hi1s1 _______495988(.DIN (___9_____39418), .Q (___9_0___39438));
  dffacs1 ______________________________________________0_495989(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39395), .Q
       (__________________________________________0___21919));
  dffacs1 ________________________________________________495990(.CLRB
       (reset), .CLK (clk), .DIN (___9__0__39406), .Q (___0_____40428));
  or2s1 ____0_9______495991(.DIN1 (___9_____39416), .DIN2
       (___9_____39363), .Q (___9_____39417));
  xor2s1 ____0______0_495992(.DIN1 (___9_____39403), .DIN2
       (___90____39057), .Q (___9_99__39432));
  nnd2s1 ____0________495993(.DIN1 (___9_____39389), .DIN2
       (___9_____39318), .Q (___9_0___39434));
  dffacs1 ______________________________________495994(.CLRB (reset),
       .CLK (clk), .DIN (___9_____39390), .QN (_________22037));
  nor2s1 _____________495995(.DIN1 (___9_____39414), .DIN2
       (___9_____39410), .Q (___9__9__39415));
  nnd2s1 ____________495996(.DIN1 (___9_9___39518), .DIN2
       (____9____38947), .Q (___9_____39413));
  hi1s1 _______495997(.DIN (___9_____39420), .Q (___9_____39412));
  nor2s1 ______0___0__495998(.DIN1 (___9_____39410), .DIN2
       (___9_____39409), .Q (___9_____39411));
  nnd2s1 ___________0_495999(.DIN1 (___9__0__39388), .DIN2
       (___9_9___39336), .Q (___9_9___39429));
  nor2s1 ___________9_496000(.DIN1 (___9_____39127), .DIN2
       (___9_____39387), .Q (___9_____39418));
  xor2s1 ______0______496001(.DIN1 (___9__9__39244), .DIN2
       (outData[24]), .Q (___9_____39408));
  nnd2s1 ____0_______496002(.DIN1 (___9_____39377), .DIN2
       (___0_90__40168), .Q (___9_____39407));
  nnd2s1 ____0_0___0_9(.DIN1 (___9_____39378), .DIN2 (___99____39861),
       .Q (___9__0__39406));
  xor2s1 ____0________496003(.DIN1 (___9_____39357), .DIN2
       (_________34647), .Q (___9__9__39405));
  nor2s1 _____09__990_(.DIN1 (___90_0__39025), .DIN2 (___9_____39403),
       .Q (___9_____39404));
  nnd2s1 ____________496004(.DIN1 (___9__9__39379), .DIN2
       (___9_____39401), .Q (___9_____39402));
  dffacs1 ________________________________________________496005(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39371), .QN
       (___0__0__40609));
  or2s1 ___________9_496006(.DIN1 (___9_____39392), .DIN2
       (___9_____39399), .Q (___9_____39400));
  xor2s1 _____________496007(.DIN1 (___9_____39397), .DIN2
       (___9_____39386), .Q (___9_____39398));
  xor2s1 _____________496008(.DIN1 (___9_____39382), .DIN2
       (_________41343), .Q (___9__0__39396));
  nnd2s1 _____________496009(.DIN1 (___9__0__39370), .DIN2
       (___9____24142), .Q (___9_____39395));
  nnd2s1 _________9___496010(.DIN1 (___9__9__39369), .DIN2
       (___9_____39752), .Q (___9_____39394));
  and2s1 _____________496011(.DIN1 (___9_____39399), .DIN2
       (___9_____39392), .Q (___9_____39393));
  xor2s1 ___________496012(.DIN1 (___9_9___39337), .DIN2
       (____00___40722), .Q (___9_____39420));
  xor2s1 ____0_____496013(.DIN1 (___9_0___39346), .DIN2
       (___9_____39359), .Q (___9_____39391));
  or2s1 ____09_____9_496014(.DIN1 (___9_0___39344), .DIN2
       (___9_____39366), .Q (___9_____39390));
  nor2s1 _____0_______496015(.DIN1 (___9_____39320), .DIN2
       (___9__9__39360), .Q (___9_____39389));
  nnd2s1 ______9______496016(.DIN1 (____00___40722), .DIN2
       (___9_9___39335), .Q (___9__0__39388));
  nnd2s1 _____________496017(.DIN1 (___9_____39386), .DIN2
       (___9_____39082), .Q (___9_____39387));
  nor2s1 ____0________496018(.DIN1 (___9_____39291), .DIN2
       (___9_____39362), .Q (___9_____39416));
  or2s1 ___________0_496019(.DIN1 (___9_____39752), .DIN2
       (___9_____39382), .Q (___9_____39383));
  nnd2s1 _____________496020(.DIN1 (___9_____39368), .DIN2
       (___9_____39752), .Q (___9_____39381));
  nor2s1 _____________496021(.DIN1
       (__________________________________________________________________21985),
       .DIN2 (___9__0__39380), .Q (___9_____39409));
  nor2s1 ____________496022(.DIN1 (___9_____39353), .DIN2
       (___9_____39386), .Q (___9_00__39617));
  and2s1 __________0__496023(.DIN1 (___9__0__39380), .DIN2
       (__________________________________________________________________21985),
       .Q (___9_____39410));
  hi1s1 _______496024(.DIN (___9__9__39379), .Q (___9_9___39518));
  nor2s1 ____0______0_496025(.DIN1 (_____0__25660), .DIN2
       (___9_0___39347), .Q (___9_____39378));
  xor2s1 ____0_0____9_496026(.DIN1 (___9_____39292), .DIN2
       (___9__0__39361), .Q (___9_____39377));
  xor2s1 ____0________496027(.DIN1 (________22772), .DIN2
       (___9_____39364), .Q (___9_____39376));
  nor2s1 ____________496028(.DIN1 (___9_____39372), .DIN2
       (___9_____39373), .Q (___9_____39375));
  nnd2s1 ______9___0_496029(.DIN1 (___9_____39373), .DIN2
       (___9_____39372), .Q (___9_____39374));
  nnd2s1 ____0________496030(.DIN1 (___9_0___39348), .DIN2 (___9_9), .Q
       (___9_____39371));
  xor2s1 _________990_496031(.DIN1 (___90____39026), .DIN2
       (___0__0__40291), .Q (___9_____39403));
  nnd2s1 ____________496032(.DIN1 (___9_90__39334), .DIN2
       (___9__9__39659), .Q (___9__0__39370));
  dffacs1 ______________0_(.CLRB (reset), .CLK (clk), .DIN
       (___9_9___39340), .Q (outData[30]));
  hi1s1 _______496033(.DIN (___9_____39368), .Q (___9__9__39369));
  xor2s1 ______0____9_496034(.DIN1
       (______________________________________________21906), .DIN2
       (___9__9__39324), .Q (___9_____39367));
  hi1s1 _______496035(.DIN (___9_____39386), .Q (___9_____39392));
  xor2s1 _____________496036(.DIN1 (____00___40724), .DIN2
       (___9_____39358), .Q (___9__9__39379));
  dffacs1 ________________________________________________496037(.CLRB
       (reset), .CLK (clk), .DIN (___9_9___39338), .Q
       (__________________________________________________________________21999));
  dffacs1 ____________________________________0_(.CLRB (reset), .CLK
       (clk), .DIN (___9_0___39345), .QN (___0_____40582));
  nnd2s1 _____________496038(.DIN1 (___9_____39331), .DIN2
       (___9_____39311), .Q (___9_____39366));
  or2s1 ____09_______496039(.DIN1
       (______________________________________________21933), .DIN2
       (___9_____39364), .Q (___9_____39365));
  and2s1 ____09___9___(.DIN1 (___9_____39364), .DIN2
       (______________________________________________21933), .Q
       (___9_____39363));
  nor2s1 ____09_______496040(.DIN1 (___9_____39290), .DIN2
       (___9__0__39361), .Q (___9_____39362));
  nor2s1 ___________496041(.DIN1 (___9_____39330), .DIN2
       (___9_____39359), .Q (___9__9__39360));
  dffacs1 ______________9_(.CLRB (reset), .CLK (clk), .DIN
       (___9_____39358), .Q (outData[29]));
  xor2s1 _____________496042(.DIN1 (___9__0__39280), .DIN2
       (___9_00__39342), .Q (___9_____39357));
  nor2s1 __________496043(.DIN1 (___90____39058), .DIN2
       (___0__0__40291), .Q (___9_____39356));
  nor2s1 ___________9_496044(.DIN1 (___9_9___39696), .DIN2
       (___9__9__39324), .Q (___9_____39355));
  nor2s1 _____________496045(.DIN1
       (______________________________________________21906), .DIN2
       (___9__9__39305), .Q (___9_____39354));
  nor2s1 ______9______496046(.DIN1 (___9_____39303), .DIN2
       (___9_____39333), .Q (___9_9___39431));
  nor2s1 _____90______496047(.DIN1 (___9__0__39228), .DIN2
       (___9__9__39324), .Q (___9_____39353));
  or2s1 _____________496048(.DIN1 (___9_____39667), .DIN2
       (___9_____39326), .Q (___9__0__39352));
  nnd2s1 __________9__496049(.DIN1 (___9_____39358), .DIN2
       (___9_____39140), .Q (___9_09__39351));
  nnd2s1 ___________0_496050(.DIN1 (___9_____39358), .DIN2
       (___9__0__39209), .Q (___9_0___39350));
  nnd2s1 _____9_______496051(.DIN1 (___9_____39358), .DIN2
       (___9_____39210), .Q (___9_____39368));
  nor2s1 _____9______496052(.DIN1 (___9_____39175), .DIN2
       (___9__9__39305), .Q (___9_____39385));
  nor2s1 _____9____0__496053(.DIN1 (___9_____39176), .DIN2
       (___9__9__39305), .Q (___9_____39382));
  dffacs1 ________________496054(.CLRB (reset), .CLK (clk), .DIN
       (___9__0__39325), .Q (outData[24]));
  nor2s1 ___________0_496055(.DIN1 (_________38646), .DIN2
       (___9_____39328), .Q (___9__0__39380));
  nor2s1 _____00____9_496056(.DIN1 (___9_0___39349), .DIN2
       (___9_____39358), .Q (___9_____39386));
  nor2s1 ____0_9______496057(.DIN1 (____9___22737), .DIN2
       (___9_____39321), .Q (___9_0___39348));
  nor2s1 ____09______496058(.DIN1 (___9_____39743), .DIN2
       (___9_____39322), .Q (___9_0___39347));
  xor2s1 __________0_496059(.DIN1 (___9_____39308), .DIN2
       (___9__9__39234), .Q (___9_0___39346));
  or2s1 ______0______496060(.DIN1 (___9_0___39344), .DIN2
       (___9_____39323), .Q (___9_0___39345));
  or2s1 _________990_496061(.DIN1 (___9_99__39341), .DIN2
       (___9_00__39342), .Q (___9_0___39343));
  and2s1 ____________496062(.DIN1 (___9_00__39342), .DIN2
       (___9_99__39341), .Q (___9_____39373));
  or2s1 _____09____9_496063(.DIN1 (___9_9___39339), .DIN2
       (___9_____39316), .Q (___9_9___39340));
  nnd2s1 _____0_______496064(.DIN1 (___9_____39313), .DIN2
       (___9_____39644), .Q (___9_9___39338));
  nnd2s1 _____9_______496065(.DIN1 (___9_9___39336), .DIN2
       (___9_9___39335), .Q (___9_9___39337));
  xor2s1 _____________496066(.DIN1 (_________38665), .DIN2
       (___9_____39327), .Q (___9_90__39334));
  nnd2s1 _________9___496067(.DIN1 (___9_____39714), .DIN2
       (___9_____39307), .Q (___9_____39399));
  dffacs1 ______________9_496068(.CLRB (reset), .CLK (clk), .DIN
       (___9__9__39314), .QN (outData[19]));
  xor2s1 ___________496069(.DIN1 (___9_____39294), .DIN2
       (___9_____39332), .Q (___9_____39333));
  nor2s1 _____________496070(.DIN1 (___9_____39310), .DIN2
       (___9_____39285), .Q (___9_____39331));
  xor2s1 __________496071(.DIN1 (___9__0__39289), .DIN2
       (___00____39910), .Q (___9_____39330));
  nor2s1 ___________9_496072(.DIN1 (___9_____39267), .DIN2
       (___9_____39309), .Q (___9__0__39361));
  xor2s1 _____________496073(.DIN1 (___9_____39287), .DIN2
       (___9_____39177), .Q (___9_____39364));
  xor2s1 _____0_______496074(.DIN1 (___9__9__39298), .DIN2
       (___9__0__39136), .Q (___0__0__40291));
  nnd2s1 _____________496075(.DIN1 (___9_9___39611), .DIN2
       (___9_____39300), .Q (___9_____39329));
  and2s1 _____________496076(.DIN1 (___9_____39327), .DIN2
       (______0__38648), .Q (___9_____39328));
  xor2s1 __________9__496077(.DIN1 (___9__0__39299), .DIN2
       (_________38858), .Q (___9_____39326));
  nnd2s1 ______0____0_496078(.DIN1 (_________38834), .DIN2
       (___9_____39304), .Q (___9__0__39325));
  hi1s1 _______496079(.DIN (___9__9__39324), .Q (___9_____39358));
  nnd2s1 _____________496080(.DIN1 (________24580), .DIN2
       (___9_____39293), .Q (___9_____39323));
  xor2s1 ______9_____496081(.DIN1 (___9_____39269), .DIN2
       (____00___40726), .Q (___9_____39322));
  nor2s1 ____099(.DIN1 (___90____38993), .DIN2 (___9_____39286), .Q
       (___9_____39321));
  nor2s1 _______496082(.DIN1 (___9_____39319), .DIN2 (___9_____39317),
       .Q (___9_____39320));
  nnd2s1 ______496083(.DIN1 (___9_____39317), .DIN2 (___9_____39319),
       .Q (___9_____39318));
  nnd2s1 _______496084(.DIN1 (___9_____39752), .DIN2 (___9_____39215),
       .Q (___9_____39714));
  nor2s1 _______496085(.DIN1 (_____0__27317), .DIN2 (___9_____39752),
       .Q (___9_____39316));
  nnd2s1 _______496086(.DIN1 (___9_____39752), .DIN2 (___9_9___39696),
       .Q (___9__0__39315));
  nnd2s1 ______496087(.DIN1 (_____0___38231), .DIN2 (___9_____39296),
       .Q (___9__9__39314));
  nor2s1 _______496088(.DIN1 (________26192), .DIN2 (___9_____39297),
       .Q (___9_____39313));
  xor2s1 _______496089(.DIN1 (___9__9__39279), .DIN2 (___9_____39312),
       .Q (___9_9___39336));
  hi1s1 ______496090(.DIN (___9__9__39305), .Q (___9__9__39324));
  xor2s1 _____99(.DIN1 (___9_____39277), .DIN2 (___9_____39263), .Q
       (___9_00__39342));
  nor2s1 ______496091(.DIN1 (___0____24203), .DIN2 (___9_____39266), .Q
       (___9_____39311));
  and2s1 ______496092(.DIN1 (___9_____39265), .DIN2
       (_____________________________________9_______21884), .Q
       (___9_____39310));
  nor2s1 _______496093(.DIN1 (____00___40726), .DIN2 (___9_____39268),
       .Q (___9_____39309));
  xor2s1 _____9_496094(.DIN1 (___9__9__39288), .DIN2 (____0____38091),
       .Q (___9_____39308));
  nnd2s1 ______496095(.DIN1 (___99_0__39827), .DIN2 (___9_____39217),
       .Q (___9_____39307));
  nnd2s1 ______496096(.DIN1 (___9__0__39270), .DIN2 (_____9___38797),
       .Q (___9_____39327));
  nor2s1 _____9_496097(.DIN1 (___9_00__39251), .DIN2 (___9_____39272),
       .Q (___9_____39359));
  nnd2s1 _______496098(.DIN1 (___99_0__39827), .DIN2
       (______________________________________________21906), .Q
       (___9__0__39306));
  xor2s1 _______496099(.DIN1 (___9_09__39260), .DIN2 (________27668),
       .Q (___9__9__39305));
  nnd2s1 _______496100(.DIN1 (___9_____39281), .DIN2 (inData[0]), .Q
       (___9_____39304));
  xor2s1 _______496101(.DIN1 (___9_____39264), .DIN2 (____9____38944),
       .Q (___9_____39303));
  xor2s1 ______496102(.DIN1
       (______________________________________________21915), .DIN2
       (______________________________________________21917), .Q
       (___9_____39300));
  xnr2s1 ______496103(.DIN1 (___9_0___39077), .DIN2 (____00___40728),
       .Q (___9__0__39299));
  xor2s1 _______496104(.DIN1 (___9_____39273), .DIN2 (___9_0___39533),
       .Q (___9__9__39298));
  nor2s1 ______496105(.DIN1
       (______________________________________________21917), .DIN2
       (___00_0__39902), .Q (___9_____39297));
  nnd2s1 _______496106(.DIN1 (___9_0___39257), .DIN2 (_________38833),
       .Q (___9_____39296));
  nor2s1 _______496107(.DIN1 (_______22219), .DIN2 (___9_0___39259), .Q
       (___9_____39295));
  nnd2s1 _______496108(.DIN1 (___9_____39262), .DIN2 (___9_____39275),
       .Q (___9_____39294));
  hi1s1 _______496109(.DIN (___99_0__39827), .Q (___9_____39752));
  nnd2s1 _____0_496110(.DIN1 (___9_____39183), .DIN2 (___9_____39284),
       .Q (___9_____39293));
  or2s1 ______496111(.DIN1 (___9_____39291), .DIN2 (___9_____39290), .Q
       (___9_____39292));
  nor2s1 ______496112(.DIN1 (___9_____39282), .DIN2 (___9__9__39288),
       .Q (___9__0__39289));
  xor2s1 _____9_496113(.DIN1 (___9_0___39252), .DIN2 (___9_____39271),
       .Q (___9_____39287));
  xor2s1 _______496114(.DIN1 (___9_9___39248), .DIN2 (____9_0__38941),
       .Q (___9_____39286));
  nor2s1 ______496115(.DIN1 (___9_____39284), .DIN2 (___9_____39283),
       .Q (___9_____39285));
  nnd2s1 _______496116(.DIN1 (___9__9__39288), .DIN2 (___9_____39282),
       .Q (___9_____39317));
  dffacs1 __________________________________________0_____496117(.CLRB
       (reset), .CLK (clk), .DIN (___9__0__39261), .Q
       (______________________________________0_______21893));
  nor2s1 _______496118(.DIN1 (___9_0___39254), .DIN2 (____009__38047),
       .Q (___9_____39281));
  xor2s1 _______496119(.DIN1 (___9_99__39341), .DIN2 (___9_____39274),
       .Q (___9__0__39280));
  nor2s1 _______496120(.DIN1 (_________38766), .DIN2 (___9_____39278),
       .Q (___9__9__39279));
  xor2s1 _______496121(.DIN1 (___9_____39276), .DIN2 (___9_____39275),
       .Q (___9_____39277));
  xor2s1 ______496122(.DIN1 (___9_____39241), .DIN2 (___9_____39274),
       .Q (___9_9___39335));
  nnd2s1 _______496123(.DIN1 (___9_____39273), .DIN2 (___9__9__39135),
       .Q (___9_____39302));
  nor2s1 _______496124(.DIN1 (___9_0___39253), .DIN2 (___9_____39271),
       .Q (___9_____39272));
  nnd2s1 ______496125(.DIN1 (_____9___38796), .DIN2 (____00___40728),
       .Q (___9__0__39270));
  or2s1 _______496126(.DIN1 (___9_____39268), .DIN2 (___9_____39267),
       .Q (___9_____39269));
  nor2s1 _____0_496127(.DIN1 (_________22036), .DIN2 (________25394),
       .Q (___9_____39266));
  nnd2s1 _____0_496128(.DIN1 (____9____34315), .DIN2 (_________22036),
       .Q (___9_____39265));
  xnr2s1 _______496129(.DIN1 (___9_0___39258), .DIN2 (________26351),
       .Q (___99_0__39827));
  or2s1 _______496130(.DIN1 (___9_____39263), .DIN2 (___9_____39276),
       .Q (___9_____39264));
  nnd2s1 _______496131(.DIN1 (___9_____39276), .DIN2 (___9_____39263),
       .Q (___9_____39262));
  nnd2s1 _______496132(.DIN1 (___9_9___39246), .DIN2 (________28493),
       .Q (___9__0__39261));
  xor2s1 _______496133(.DIN1 (___9_____39230), .DIN2 (______9__22017),
       .Q (___9_09__39260));
  nor2s1 _______496134(.DIN1 (____9__22214), .DIN2 (___9_0___39258), .Q
       (___9_0___39259));
  xor2s1 ______496135(.DIN1 (___9__0__39235), .DIN2 (____9____38904),
       .Q (___9__9__39288));
  nnd2s1 _______496136(.DIN1 (___9_____39242), .DIN2 (inData[20]), .Q
       (___9_0___39257));
  hi1s1 _____9_496137(.DIN (___9_____39278), .Q (___9_0___39256));
  hi1s1 _______496138(.DIN (_________22036), .Q (___9_____39284));
  and2s1 _______496139(.DIN1 (___9_0___39255), .DIN2
       (_______________________________________________________________),
       .Q (___9_____39290));
  nor2s1 _______496140(.DIN1
       (_______________________________________________________________),
       .DIN2 (___9_0___39255), .Q (___9_____39291));
  dffacs1 ________________________________________________496141(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39243), .Q
       (______________________________________________21917));
  dffacs1 ________________________________________________496142(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39239), .Q
       (______________________________________________21955));
  xnr2s1 _____9_496143(.DIN1 (outData[28]), .DIN2 (outData[19]), .Q
       (___9_0___39254));
  nor2s1 _______496144(.DIN1 (___9_99__39250), .DIN2 (___9_0___39252),
       .Q (___9_0___39253));
  and2s1 _______496145(.DIN1 (___9_0___39252), .DIN2 (___9_99__39250),
       .Q (___9_00__39251));
  nor2s1 _______496146(.DIN1 (___9_____39212), .DIN2 (___9_____39237),
       .Q (___9_____39271));
  hi1s1 _____9_496147(.DIN (___9_____39276), .Q (___990___39802));
  xor2s1 _____9_496148(.DIN1 (___9_____39224), .DIN2 (___9_____39149),
       .Q (___9_9___39248));
  nnd2s1 _____0_496149(.DIN1 (___9_____39233), .DIN2 (___9_____39111),
       .Q (___9_____39273));
  nor2s1 _______496150(.DIN1
       (_______________________________________________________________9__21995),
       .DIN2 (___9_9___39247), .Q (___9_____39267));
  and2s1 _______496151(.DIN1 (___9_9___39247), .DIN2
       (_______________________________________________________________9__21995),
       .Q (___9_____39268));
  dffacs1 _________________________________________9___0_(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39238), .QN
       (_________22036));
  xor2s1 _____0_496152(.DIN1 (___9_____39240), .DIN2 (_________38842),
       .Q (___9_____39278));
  nnd2s1 _______496153(.DIN1 (___9_____39225), .DIN2 (___9_90__39245),
       .Q (___9_9___39246));
  and2s1 _______496154(.DIN1 (outData[19]), .DIN2 (outData[28]), .Q
       (___9__9__39244));
  nnd2s1 _______496155(.DIN1 (___9_____39223), .DIN2 (________27377),
       .Q (___9_____39243));
  and2s1 _______496156(.DIN1 (________24912), .DIN2 (outData[28]), .Q
       (___9_____39242));
  nor2s1 _____0_496157(.DIN1 (____9____38903), .DIN2 (___9_____39226),
       .Q (___9_99__39341));
  xor2s1 _____0_496158(.DIN1 (___9__9__39153), .DIN2 (___9_____39232),
       .Q (___9_____39276));
  nnd2s1 _______496159(.DIN1 (___9_____39240), .DIN2 (_____0___38806),
       .Q (___9_____39241));
  nnd2s1 _____0_496160(.DIN1 (___0_0__28796), .DIN2 (___9_____39220),
       .Q (___9_____39239));
  or2s1 _______496161(.DIN1 (___9_____39216), .DIN2 (___9__9__39650),
       .Q (___9_____39557));
  dffacs1 __________________________________________0___0_(.CLRB
       (reset), .CLK (clk), .DIN (___9__9__39227), .QN
       (______________________________________0___0_));
  nor2s1 _______496162(.DIN1 (__9_____29953), .DIN2 (___9_____39222),
       .Q (___9_0___39258));
  xor2s1 ______496163(.DIN1 (___9_____39214), .DIN2 (___9_____39236),
       .Q (___9_0___39255));
  nnd2s1 _______496164(.DIN1 (___9_____39213), .DIN2 (____0_0__34423),
       .Q (___9_____39238));
  nor2s1 _______496165(.DIN1 (___9_____39199), .DIN2 (___9_____39236),
       .Q (___9_____39237));
  xor2s1 _____00(.DIN1 (___99____39834), .DIN2 (____9_9__38905), .Q
       (___9__0__39235));
  xor2s1 _______496166(.DIN1 (___9_____39197), .DIN2 (_________36856),
       .Q (___9_9___39247));
  hi1s1 ______496167(.DIN (___9__9__39234), .Q (___9_____39282));
  xor2s1 _____0_496168(.DIN1 (___9__9__39201), .DIN2 (_________38813),
       .Q (___9_0___39252));
  or2s1 _______496169(.DIN1 (___9_____39084), .DIN2 (___9_____39232),
       .Q (___9_____39233));
  xor2s1 ______496170(.DIN1 (___9_____39221), .DIN2 (___0_____40583),
       .Q (___9_____39230));
  nnd2s1 ______496171(.DIN1 (___9__0__39202), .DIN2 (___9__0__39228),
       .Q (___9_9___39249));
  nnd2s1 _______496172(.DIN1 (___9_____39190), .DIN2 (_________38713),
       .Q (___9__9__39227));
  nor2s1 _______496173(.DIN1 (____9_0__38906), .DIN2 (___99____39834),
       .Q (___9_____39226));
  xor2s1 _______496174(.DIN1 (___9__0__39172), .DIN2 (___9_____39231),
       .Q (___9_____39225));
  xor2s1 _______496175(.DIN1
       (______________________________________________21932), .DIN2
       (____0_0__40730), .Q (___9_____39224));
  or2s1 _______496176(.DIN1 (___9_____39667), .DIN2 (___9_____39189),
       .Q (___9_____39223));
  and2s1 _______496177(.DIN1 (___9_____39221), .DIN2 (__9_____29952),
       .Q (___9_____39222));
  nnd2s1 _______496178(.DIN1 (___9_____39196), .DIN2 (___9_____39200),
       .Q (___9__9__39234));
  nnd2s1 _______496179(.DIN1 (___9_____39219), .DIN2 (___0_____40429),
       .Q (___9_____39220));
  xor2s1 _______496180(.DIN1 (___9_09__39171), .DIN2 (___9__0__41371),
       .Q (___9_____39240));
  dffacs1 ________________________________________________496181(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39194), .Q
       (_______________________________________________________________));
  nor2s1 ______496182(.DIN1 (___9__9__39218), .DIN2 (___9_____39217),
       .Q (___9__9__39650));
  dffacs1 ________________496183(.CLRB (reset), .CLK (clk), .DIN
       (___9__9__39191), .Q (outData[28]));
  dffacs1 ________________________________________________496184(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39193), .QN
       (______________________________________________21916));
  dffacs1 ________________________________________________496185(.CLRB
       (reset), .CLK (clk), .DIN (___9__0__39192), .Q (___0_____40436));
  nor2s1 ______496186(.DIN1 (___90____38999), .DIN2 (___9_____39215),
       .Q (___9_____39216));
  xor2s1 _______496187(.DIN1 (___9_____39198), .DIN2 (___9_____39211),
       .Q (___9_____39214));
  and2s1 _______496188(.DIN1 (___9_____39186), .DIN2 (___9_____39283),
       .Q (___9_____39213));
  nor2s1 _____9_496189(.DIN1 (___9_____39211), .DIN2 (___9_____39187),
       .Q (___9_____39212));
  hi1s1 _______496190(.DIN (___9__0__39209), .Q (___9_____39210));
  nor2s1 ______496191(.DIN1 (___9_____39147), .DIN2 (____0_0__40730),
       .Q (___9_____39229));
  nor2s1 _____0_496192(.DIN1 (___90____39012), .DIN2 (___9_____39179),
       .Q (___9_____39236));
  and2s1 _______496193(.DIN1 (___9_____39203), .DIN2 (___9_____39207),
       .Q (___9_____39208));
  nor2s1 _______496194(.DIN1 (___9_____39207), .DIN2 (___9_____39203),
       .Q (___9_____39204));
  xor2s1 _______496195(.DIN1 (___9_9___39155), .DIN2 (____9____38948),
       .Q (___9__0__39202));
  nor2s1 ______496196(.DIN1 (___9_____39092), .DIN2 (___9_____39174),
       .Q (___9_____39232));
  dffacs1 _______________________________________________496197(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39185), .Q
       (_____________________________________________21875));
  and2s1 _______496198(.DIN1 (___9_____39200), .DIN2 (___9_____39195),
       .Q (___9__9__39201));
  nor2s1 _____9_496199(.DIN1 (____9_9__38959), .DIN2 (___9_____39198),
       .Q (___9_____39199));
  xor2s1 _____496200(.DIN1 (___90____39039), .DIN2 (___9_____39178), .Q
       (___9_____39197));
  nnd2s1 _______496201(.DIN1 (___9_____39195), .DIN2 (_________38812),
       .Q (___9_____39196));
  dffacs1 ________________________________________________496202(.CLRB
       (reset), .CLK (clk), .DIN (___9_0___39164), .QN
       (___0_____40429));
  nnd2s1 _______496203(.DIN1 (___9_9___39160), .DIN2 (______0__37731),
       .Q (___9_____39194));
  xor2s1 _______496204(.DIN1 (___9_____39143), .DIN2 (____0_0__38064),
       .Q (___9__0__39209));
  xor2s1 _______496205(.DIN1 (___9_____39093), .DIN2 (___9_____39173),
       .Q (___99____39834));
  nnd2s1 _______496206(.DIN1 (___9_9___39154), .DIN2 (___9____24092),
       .Q (___9_____39193));
  nnd2s1 _______496207(.DIN1 (_________38814), .DIN2 (___9_0___39165),
       .Q (___9__0__39192));
  nnd2s1 ______496208(.DIN1 (___9_____39152), .DIN2 (___0____24186), .Q
       (___9__9__39191));
  nnd2s1 _______496209(.DIN1 (___9_9___39157), .DIN2 (___90____39040),
       .Q (___9_____39190));
  xor2s1 ______496210(.DIN1 (_________38459), .DIN2 (___9_0___39168),
       .Q (___9_____39189));
  or2s1 _______496211(.DIN1 (___9_____39207), .DIN2 (___9_0___39167),
       .Q (___9_____39188));
  nor2s1 _______496212(.DIN1 (___9_____39134), .DIN2 (___9_9___39159),
       .Q (___9_____39221));
  hi1s1 _______496213(.DIN (___9_____39215), .Q (___9_____39217));
  hi1s1 _______496214(.DIN (___9_____39198), .Q (___9_____39187));
  nor2s1 _____0_496215(.DIN1 (____0___23974), .DIN2 (___9_____39148),
       .Q (___9_____39186));
  or2s1 _______496216(.DIN1 (_________38751), .DIN2 (___9_____39151),
       .Q (___9_____39185));
  nnd2s1 _______496217(.DIN1 (___9__9__39145), .DIN2 (___9_____39183),
       .Q (___9_____39184));
  nor2s1 _______496218(.DIN1 (___9__9__39181), .DIN2 (___9_____39180),
       .Q (___9__0__39182));
  nor2s1 _______496219(.DIN1 (___90_9__39061), .DIN2 (___9_____39178),
       .Q (___9_____39179));
  xor2s1 _______496220(.DIN1 (___9_99__39250), .DIN2 (_____99__36913),
       .Q (___9_____39177));
  hi1s1 _____0_496221(.DIN (___9_____39175), .Q (___9_____39176));
  nor2s1 _______496222(.DIN1 (___9_____39091), .DIN2 (___9_____39173),
       .Q (___9_____39174));
  xor2s1 _______496223(.DIN1 (___9_____39139), .DIN2 (___9__0__41371),
       .Q (___9__0__39172));
  xor2s1 _______496224(.DIN1 (___9_____39128), .DIN2 (___9_0___39170),
       .Q (___9_09__39171));
  xor2s1 _______496225(.DIN1 (___9_00__39162), .DIN2 (___9_9__27761),
       .Q (___9_0___39169));
  or2s1 _______496226(.DIN1 (_________38441), .DIN2 (___9_0___39168),
       .Q (___9_____39205));
  hi1s1 _______496227(.DIN (___9_0___39167), .Q (___9_____39203));
  xnr2s1 ______496228(.DIN1 (___9_0___39166), .DIN2 (___9_____39127),
       .Q (___9_____39215));
  nnd2s1 _____9_496229(.DIN1 (___90____39051), .DIN2 (___9_____39129),
       .Q (___9_0___39165));
  nnd2s1 _____496230(.DIN1 (___9_____39130), .DIN2 (___0_90__40168), .Q
       (___9_0___39164));
  nor2s1 _______496231(.DIN1
       (______________________________________________21958), .DIN2
       (___9_00__39162), .Q (___9_0___39163));
  nnd2s1 _______496232(.DIN1 (___9_00__39162), .DIN2
       (______________________________________________21958), .Q
       (___9_99__39161));
  nor2s1 _____9_496233(.DIN1 (___0_____30689), .DIN2 (___9_____39132),
       .Q (___9_9___39160));
  nor2s1 _____9_496234(.DIN1 (___9_____39397), .DIN2 (___9_____39131),
       .Q (___9_9___39159));
  nnd2s1 _______496235(.DIN1 (___9_00__39162), .DIN2 (___9_9___39158),
       .Q (___9_____39200));
  or2s1 _______496236(.DIN1 (___9_9___39158), .DIN2 (___9_00__39162),
       .Q (___9_____39195));
  xor2s1 _______496237(.DIN1 (___9_____39116), .DIN2 (_________38491),
       .Q (___9_____39198));
  xor2s1 _____09(.DIN1 (___9_____39110), .DIN2 (___9_9___39790), .Q
       (___9_9___39157));
  nor2s1 _______496238(.DIN1 (___9_____39141), .DIN2 (___9__0__41371),
       .Q (___9_9___39156));
  nnd2s1 _______496239(.DIN1 (___9_____39127), .DIN2 (___9_____39100),
       .Q (___9_9___39155));
  nnd2s1 _____0_496240(.DIN1 (___9_____39124), .DIN2 (________23899),
       .Q (___9_9___39154));
  xor2s1 _______496241(.DIN1 (___9_____39112), .DIN2 (_________38385),
       .Q (___9__9__39153));
  nnd2s1 _____496242(.DIN1 (___9_____39127), .DIN2 (____9____38949), .Q
       (___9_____39152));
  nor2s1 _______496243(.DIN1 (_________41264), .DIN2 (___9_____39464),
       .Q (___9_0___39167));
  nnd2s1 ______496244(.DIN1 (___9_____39127), .DIN2 (___9__0__39126),
       .Q (___9_____39175));
  dffacs1 _________________________________________9___9_(.CLRB
       (reset), .CLK (clk), .DIN (___9_____39133), .QN
       (___0_____40624));
  nor2s1 _______496245(.DIN1 (____9____38898), .DIN2 (___9_____39121),
       .Q (___9_____39151));
  or2s1 ______496246(.DIN1 (___9__0__39146), .DIN2 (___9_____39149), .Q
       (___9_____39150));
  nnd2s1 _______496247(.DIN1 (___9_____39120), .DIN2 (___9_0__25087),
       .Q (___9_____39148));
  and2s1 _____0_496248(.DIN1 (___9_____39149), .DIN2 (___9__0__39146),
       .Q (___9_____39147));
  xor2s1 ______496249(.DIN1 (____0___28556), .DIN2 (___9_____39109), .Q
       (___9__9__39145));
  xor2s1 _______496250(.DIN1 (____0____40732), .DIN2 (___9_____39738),
       .Q (___9_____39178));
  nor2s1 _______496251(.DIN1
       (______________________________________________21957), .DIN2
       (___9_____39119), .Q (___9_____39180));
  nor2s1 _____9_496252(.DIN1 (___9_9___39696), .DIN2 (___9_____39142),
       .Q (___9_____39144));
  nnd2s1 _____0_496253(.DIN1 (___9_____39142), .DIN2 (___9_____39141),
       .Q (___9_____39143));
  nnd2s1 _____0_496254(.DIN1 (___9_____39142), .DIN2 (___9_____39139),
       .Q (___9_____39140));
  nnd2s1 _____9_496255(.DIN1 (___9_____39142), .DIN2 (___9_9___39696),
       .Q (___9_____39138));
  nor2s1 ______496256(.DIN1 (___9__0__39136), .DIN2 (___9_0___39533),
       .Q (___9_____39137));
  nnd2s1 _______496257(.DIN1 (___9_0___39533), .DIN2 (___0_9___40653),
       .Q (___9__9__39135));
  nor2s1 _______496258(.DIN1 (____9____38908), .DIN2 (___9_____39114),
       .Q (___9_____39173));
  nor2s1 _______496259(.DIN1 (_________38396), .DIN2 (___9__0__39118),
       .Q (___9_0___39168));
  nor2s1 _______496260(.DIN1 (_________________0_), .DIN2
       (___9__0__39099), .Q (___9_____39134));
  nnd2s1 _______496261(.DIN1 (___9_____39106), .DIN2 (_________38856),
       .Q (___9_____39133));
  nor2s1 _______496262(.DIN1
       (______________________________________________21914), .DIN2
       (_________38377), .Q (___9_____39132));
  nor2s1 _______496263(.DIN1 (___0____22311), .DIN2 (___9_____39104),
       .Q (___9_____39131));
  xor2s1 _______496264(.DIN1 (___9_____39096), .DIN2 (___9__9__39088),
       .Q (___9_____39130));
  nnd2s1 _______496265(.DIN1 (_________41337), .DIN2
       (______________________________________________21914), .Q
       (___9_____39129));
  nor2s1 _____496266(.DIN1 (_________38762), .DIN2 (___9_____39105), .Q
       (___9_99__39250));
  xor2s1 _______496267(.DIN1 (____99___38973), .DIN2 (___9_____39113),
       .Q (___9_00__39162));
  nnd2s1 _______496268(.DIN1 (___9_____39102), .DIN2 (___9_____39101),
       .Q (___9_____39128));
  xor2s1 _______496269(.DIN1 (___9_____39087), .DIN2 (___9__9__39125),
       .Q (___9__0__39126));
  xor2s1 _______496270(.DIN1 (___9__9__39117), .DIN2 (_________38397),
       .Q (___9_____39124));
  or2s1 _______496271(.DIN1 (___9_____39086), .DIN2 (___9_09__39535),
       .Q (___9_____39464));
  dffacs1 _____________________________________________0_(.CLRB
       (reset), .CLK (clk), .DIN (___9__9__39107), .QN
       (___0_00__40461));
  hi1s1 _______496272(.DIN (___9_____39142), .Q (___9_____39127));
  hi1s1 _______496273(.DIN (___9_____39142), .Q (___9__0__41371));
  dffacs1 _____________________0_496274(.CLRB (reset), .CLK (clk), .DIN
       (___9__0__39108), .QN (_________________0___21728));
  xor2s1 _______496275(.DIN1 (________28882), .DIN2 (___9_0___39073),
       .Q (___9_____39121));
  nnd2s1 _______496276(.DIN1 (___9_____39094), .DIN2 (___9_____39183),
       .Q (___9_____39120));
  xor2s1 _______496277(.DIN1 (___9_____39115), .DIN2 (_________36973),
       .Q (___9_____39119));
  xor2s1 _______496278(.DIN1 (___9_09__39078), .DIN2 (____9____38939),
       .Q (___9_____39149));
  and2s1 _______496279(.DIN1 (___9__9__39117), .DIN2 (______0__38362),
       .Q (___9__0__39118));
  xor2s1 _______496280(.DIN1 (_________38783), .DIN2 (___9_____39115),
       .Q (___9_____39116));
  nor2s1 _______496281(.DIN1 (____90___38893), .DIN2 (___9_____39113),
       .Q (___9_____39114));
  nnd2s1 _______496282(.DIN1 (___9_____39111), .DIN2 (___9_____39085),
       .Q (___9_____39112));
  or2s1 _______496283(.DIN1 (___9_____39083), .DIN2 (___9_____39139),
       .Q (___9_____39110));
  xor2s1 _______496284(.DIN1 (____0____40734), .DIN2 (___9_0___39349),
       .Q (___9_0___39533));
  xnr2s1 ______496285(.DIN1 (___9__9__39098), .DIN2 (___9_____39103),
       .Q (___9_____39142));
  nor2s1 _____0_496286(.DIN1 (_____9__28341), .DIN2 (___9_____39081),
       .Q (___9_____39109));
  nnd2s1 _____9_496287(.DIN1 (_________33967), .DIN2 (___9_0___39075),
       .Q (___9__0__39108));
  nnd2s1 _____9_496288(.DIN1 (___9_0___39076), .DIN2 (_____9___38319),
       .Q (___9__9__39107));
  nor2s1 _______496289(.DIN1 (__9_0___29811), .DIN2 (___9__0__39079),
       .Q (___9_____39106));
  and2s1 ______496290(.DIN1 (___9_____39115), .DIN2 (______0__38760),
       .Q (___9_____39105));
  and2s1 _______496291(.DIN1 (___9_____39103), .DIN2 (________22503),
       .Q (___9_____39104));
  and2s1 _______496292(.DIN1 (___9_____39115), .DIN2
       (______________________________________________21957), .Q
       (___9__9__39181));
  nnd2s1 _____9_496293(.DIN1 (___9_0___39349), .DIN2 (___90____39022),
       .Q (___9_____39102));
  or2s1 _____9_496294(.DIN1 (___9_____39100), .DIN2 (___9_0___39349),
       .Q (___9_____39101));
  or2s1 _______496295(.DIN1 (___9__9__39098), .DIN2 (___9_____39103),
       .Q (___9__0__39099));
  dffacs1 ________________496296(.CLRB (reset), .CLK (clk), .DIN
       (___9_0___39349), .Q (outData[27]));
  dffacs1 ________________________________________________496297(.CLRB
       (reset), .CLK (clk), .DIN (___9_0___39072), .Q
       (______________________________________________21914));
  nnd2s1 _____496298(.DIN1 (___9_0___39349), .DIN2 (___90____39021), .Q
       (___9_____39141));
  dffacs1 _______________________________________________496299(.CLRB
       (reset), .CLK (clk), .DIN (___9_0___39074), .Q (___0__9__40430));
  nor2s1 _____0_496300(.DIN1 (____9____38965), .DIN2 (___9_0___39349),
       .Q (___9_09__39535));
  nor2s1 _______496301(.DIN1
       (______________________________________________21905), .DIN2
       (___9__0__39228), .Q (___9_____39097));
  and2s1 _______496302(.DIN1 (___9_____39095), .DIN2 (___9__0__39089),
       .Q (___9_____39096));
  xor2s1 _______496303(.DIN1 (__9_99), .DIN2 (___9_____39080), .Q
       (___9_____39094));
  or2s1 _______496304(.DIN1 (___9_____39092), .DIN2 (___9_____39091),
       .Q (___9_____39093));
  nnd2s1 _______496305(.DIN1 (___9__0__39228), .DIN2
       (______________________________________________21905), .Q
       (___9_____39090));
  and2s1 ______496306(.DIN1 (___9__0__39089), .DIN2 (___9__9__39088),
       .Q (___9_____39122));
  nor2s1 ______496307(.DIN1 (____9____38962), .DIN2 (___9099__39070),
       .Q (___9_____39113));
  and2s1 _____0_496308(.DIN1 (___9__0__39228), .DIN2 (___9_____39100),
       .Q (___9_____39087));
  nor2s1 _____9_496309(.DIN1 (____9____38953), .DIN2 (___9__0__39228),
       .Q (___9_____39086));
  hi1s1 _____496310(.DIN (___9_____39084), .Q (___9_____39085));
  nor2s1 _______496311(.DIN1 (___9_____39082), .DIN2 (___9__0__39228),
       .Q (___9_____39083));
  nnd2s1 _____0_496312(.DIN1 (___909___39066), .DIN2 (_____9___38323),
       .Q (___9__9__39117));
  and2s1 ______496313(.DIN1 (___9__0__39228), .DIN2 (___9_____39082),
       .Q (___9_____39139));
  dffacs1 __________________________________________0___9_(.CLRB
       (reset), .CLK (clk), .DIN (___909___39068), .Q
       (______________________________________0___9_));
  nor2s1 ______496314(.DIN1 (_____0__28324), .DIN2 (___9_____39080), .Q
       (___9_____39081));
  nor2s1 _____496315(.DIN1 (_________38743), .DIN2 (___9090__39062), .Q
       (___9__0__39079));
  xor2s1 ______496316(.DIN1 (___90____39049), .DIN2 (___9_0___39077),
       .Q (___9_09__39078));
  nor2s1 _______496317(.DIN1 (________23773), .DIN2 (___90_0__39054),
       .Q (___9_0___39076));
  nor2s1 _______496318(.DIN1 (___90____39059), .DIN2 (____9____32399),
       .Q (___9_0___39075));
  nnd2s1 _____9_496319(.DIN1 (___909___39063), .DIN2 (___9_9), .Q
       (___9_0___39074));
  nor2s1 _______496320(.DIN1 (___90____39036), .DIN2 (___90____39060),
       .Q (___9_0___39073));
  nnd2s1 ______496321(.DIN1 (___90____39052), .DIN2 (________26365), .Q
       (___9_0___39072));
  nnd2s1 _____496322(.DIN1 (___9_____39579), .DIN2 (___9_00__39071), .Q
       (___9_____39111));
  nor2s1 _____9_496323(.DIN1 (___9_00__39071), .DIN2 (___9_____39579),
       .Q (___9_____39084));
  dffacs1 __________________________________________0_____496324(.CLRB
       (reset), .CLK (clk), .DIN (___90_9__39053), .Q
       (______________________________________0_______21892));
  xor2s1 _____0_496325(.DIN1 (___90____39045), .DIN2 (___9_____39738),
       .Q (___9_____39103));
  xor2s1 ______496326(.DIN1 (___90____39047), .DIN2 (___909___39069),
       .Q (___9_____39115));
  hi1s1 ______496327(.DIN (___9__0__39228), .Q (___9_0___39349));
  nor2s1 _____9_496328(.DIN1 (___90____39048), .DIN2 (___909___39069),
       .Q (___9099__39070));
  nnd2s1 _______496329(.DIN1 (___90_0__39044), .DIN2 (_____0__26655),
       .Q (___909___39068));
  xor2s1 _____0_496330(.DIN1 (___90____39029), .DIN2 (______0__35711),
       .Q (___9_____39091));
  nnd2s1 _____0_496331(.DIN1 (___909___39067), .DIN2
       (______________________________________________21931), .Q
       (___9_____39095));
  or2s1 _____0_496332(.DIN1
       (______________________________________________21931), .DIN2
       (___909___39067), .Q (___9__0__39089));
  xnr2s1 _______496333(.DIN1 (___909___39065), .DIN2 (___90_9__39024),
       .Q (___909___39066));
  or2s1 _______496334(.DIN1 (___9_____39667), .DIN2 (___90____39043),
       .Q (___909___39064));
  dffacs1 ______________________________________496335(.CLRB (reset),
       .CLK (clk), .DIN (___90____39050), .QN (_____________22085));
  xnr2s1 _______496336(.DIN1 (___0_____40448), .DIN2 (___90____39020),
       .Q (___9__0__39228));
  nor2s1 _______496337(.DIN1 (___90_9__39034), .DIN2 (______0__38594),
       .Q (___909___39063));
  xor2s1 _______496338(.DIN1 (___90____39017), .DIN2 (____0____36215),
       .Q (___9090__39062));
  xor2s1 _______496339(.DIN1 (___90____39016), .DIN2 (___9__9__39731),
       .Q (___90_9__39061));
  and2s1 _______496340(.DIN1 (___90____39038), .DIN2 (___9_____39312),
       .Q (___90____39060));
  nor2s1 _______496341(.DIN1 (___90____39037), .DIN2 (____9____33386),
       .Q (___90____39059));
  and2s1 _______496342(.DIN1 (___90____39057), .DIN2 (___90____39027),
       .Q (___90____39058));
  nor2s1 _______496343(.DIN1 (_________________9___21749), .DIN2
       (___90____39033), .Q (___90_0__39054));
  nnd2s1 _______496344(.DIN1 (___90____39041), .DIN2 (________23838),
       .Q (___90_9__39053));
  or2s1 _______496345(.DIN1 (___90____39051), .DIN2 (___90____39030),
       .Q (___90____39052));
  nor2s1 ______496346(.DIN1 (___90____38989), .DIN2 (___90_0__39035),
       .Q (___9_____39080));
  xor2s1 _______496347(.DIN1 (____0____40736), .DIN2 (___9__9__39218),
       .Q (___9_____39579));
  nnd2s1 _______496348(.DIN1 (___90____39013), .DIN2 (_________38628),
       .Q (___90____39050));
  xor2s1 ______496349(.DIN1 (____9____38957), .DIN2 (___90____39031),
       .Q (___90____39049));
  and2s1 _______496350(.DIN1 (___90____39046), .DIN2 (___90____39009),
       .Q (___90____39048));
  nnd2s1 _______496351(.DIN1 (___90____39046), .DIN2 (___90____39018),
       .Q (___90____39047));
  xor2s1 _______496352(.DIN1 (___90_9__38997), .DIN2 (_________38825),
       .Q (___909___39067));
  nnd2s1 ______496353(.DIN1 (___90____39007), .DIN2 (___900___38983),
       .Q (___90____39045));
  nnd2s1 _______496354(.DIN1 (___90____39003), .DIN2 (___9__9__39459),
       .Q (___90_0__39044));
  xor2s1 ______496355(.DIN1 (_____99__38324), .DIN2 (___90____39023),
       .Q (___90____39043));
  or2s1 _______496356(.DIN1 (___90____39000), .DIN2 (___90____39057),
       .Q (___90____39042));
  nnd2s1 _______496357(.DIN1 (___900___38986), .DIN2 (___90____39040),
       .Q (___90____39041));
  xor2s1 _______496358(.DIN1 (___90_9__39014), .DIN2 (___90_0__39015),
       .Q (___90____39039));
  nnd2s1 _______496359(.DIN1 (___90____38995), .DIN2 (_____0__28872),
       .Q (___90____39038));
  nnd2s1 _______496360(.DIN1 (_________31846), .DIN2 (___90____38996),
       .Q (___90____39037));
  nor2s1 _______496361(.DIN1 (___9_____39312), .DIN2 (___90____39032),
       .Q (___90____39036));
  nor2s1 _______496362(.DIN1 (___90____38990), .DIN2 (______0__38780),
       .Q (___90_0__39035));
  nnd2s1 _______496363(.DIN1 (____9____38946), .DIN2 (___90____38994),
       .Q (___90_9__39034));
  and2s1 _____9_496364(.DIN1 (___90____39032), .DIN2 (___90____38992),
       .Q (___90____39033));
  nnd2s1 _______496365(.DIN1 (___90_0__38998), .DIN2 (___90____39031),
       .Q (___90____39056));
  dffacs1 ________________496366(.CLRB (reset), .CLK (clk), .DIN
       (___90_0__38988), .QN (outData[26]));
  xor2s1 ______496367(.DIN1 (____0____38079), .DIN2 (____99___38971),
       .Q (___90____39030));
  nnd2s1 _______496368(.DIN1 (___90____39028), .DIN2 (___90____39019),
       .Q (___90____39029));
  nnd2s1 _______496369(.DIN1 (___90____39026), .DIN2 (___90_0__39025),
       .Q (___90____39027));
  nnd2s1 ______496370(.DIN1 (___90____39023), .DIN2 (_____9___38322),
       .Q (___90_9__39024));
  hi1s1 _______496371(.DIN (___90____39021), .Q (___90____39022));
  nor2s1 _______496372(.DIN1 (___90____39006), .DIN2 (___900___38984),
       .Q (___90____39020));
  nor2s1 _______496373(.DIN1 (___90____39019), .DIN2 (___90____39028),
       .Q (___9_____39092));
  dffacs1 __________________________________________0_____496374(.CLRB
       (reset), .CLK (clk), .DIN (___9009__38987), .QN
       (______________________________________0_______21891));
  nnd2s1 _______496375(.DIN1 (____99___38975), .DIN2 (___90____39008),
       .Q (___90____39018));
  xor2s1 _____0_496376(.DIN1 (_________38781), .DIN2
       (_________________________________________9___21874), .Q
       (___90____39017));
  or2s1 _____0_496377(.DIN1 (___90_0__39015), .DIN2 (___90_9__39014),
       .Q (___90____39016));
  nnd2s1 ______496378(.DIN1 (____999__38977), .DIN2 (inData[18]), .Q
       (___90____39013));
  and2s1 _____9_496379(.DIN1 (___90_9__39014), .DIN2 (___90_0__39015),
       .Q (___90____39012));
  nnd2s1 _______496380(.DIN1 (___90____39010), .DIN2 (____9____38937),
       .Q (___90____39011));
  nnd2s1 _______496381(.DIN1 (___900___38980), .DIN2 (___90____39008),
       .Q (___90____39009));
  or2s1 _______496382(.DIN1 (___0_____40448), .DIN2 (___90____39006),
       .Q (___90____39007));
  nor2s1 _______496383(.DIN1 (___90_9__39004), .DIN2 (____990__38969),
       .Q (___90_0__39005));
  nor2s1 ______496384(.DIN1 (____9____38967), .DIN2 (___9_____39082),
       .Q (___90____39003));
  nor2s1 ______496385(.DIN1 (____9____38954), .DIN2 (___90____39000),
       .Q (___9_____39275));
  nnd2s1 _______496386(.DIN1 (_________41372), .DIN2 (___90____38999),
       .Q (___90____39021));
  and2s1 _____9_496387(.DIN1 (___9_____39207), .DIN2 (____99___38972),
       .Q (___90____39057));
  xor2s1 _______496388(.DIN1 (____9_9__38940), .DIN2 (_________35806),
       .Q (___90_0__38998));
  xor2s1 _____9_496389(.DIN1 (____9____38945), .DIN2 (______9__38826),
       .Q (___90_9__38997));
  nnd2s1 _____0_496390(.DIN1
       (_________________________________________9___21874), .DIN2
       (inData[17]), .Q (___90____38996));
  nnd2s1 _____496391(.DIN1 (___90____38991), .DIN2 (________28873), .Q
       (___90____38995));
  nnd2s1 _______496392(.DIN1 (___90____38993), .DIN2 (____9____38964),
       .Q (___90____38994));
  nnd2s1 _______496393(.DIN1 (___90____38991), .DIN2 (___900___38982),
       .Q (___90____38992));
  nor2s1 _______496394(.DIN1
       (_________________________________________9___21874), .DIN2
       (_________41367), .Q (___90____38990));
  and2s1 _______496395(.DIN1 (________27612), .DIN2
       (_________________________________________9___21874), .Q
       (___90____38989));
  nnd2s1 _______496396(.DIN1 (____9_0__38960), .DIN2 (_________38868),
       .Q (___90____39031));
  nnd2s1 _______496397(.DIN1 (____9_9__38950), .DIN2 (________27318),
       .Q (___90_0__38988));
  nnd2s1 ______496398(.DIN1 (____9____38955), .DIN2 (____9____38021),
       .Q (___9009__38987));
  xor2s1 _______496399(.DIN1 (____9____38935), .DIN2 (___900___38985),
       .Q (___900___38986));
  hi1s1 _______496400(.DIN (___900___38983), .Q (___900___38984));
  nnd2s1 _______496401(.DIN1 (___900___38979), .DIN2 (______0__41289),
       .Q (___90____39046));
  hi1s1 _______496402(.DIN (___90____39000), .Q (___90____39026));
  or2s1 ______496403(.DIN1 (___900___38982), .DIN2 (___90____38991), .Q
       (___90____39032));
  nnd2s1 _____0_496404(.DIN1 (____9____38956), .DIN2 (____99___38035),
       .Q (___90____39023));
  nnd2s1 _____496405(.DIN1 (____9____38952), .DIN2 (___9__9__39218), .Q
       (___9_____39100));
  hi1s1 _______496406(.DIN (___900___38981), .Q (___90____39028));
  hi1s1 _______496407(.DIN (___900___38979), .Q (___900___38980));
  nnd2s1 _____9_496408(.DIN1 (___9__9__39218), .DIN2
       (_______________________________________________________________9),
       .Q (___9000__38978));
  nor2s1 _______496409(.DIN1 (_____0___38616), .DIN2 (____9____38943),
       .Q (____999__38977));
  nor2s1 _____9_496410(.DIN1
       (_______________________________________________________________9),
       .DIN2 (___9__9__39218), .Q (____99___38976));
  xor2s1 _______496411(.DIN1 (____9____38961), .DIN2 (___9_____39401),
       .Q (____99___38975));
  nor2s1 _______496412(.DIN1 (___90____38993), .DIN2 (____9____38938),
       .Q (____99___38974));
  xor2s1 _______496413(.DIN1 (____9____38918), .DIN2 (____90___38892),
       .Q (____99___38973));
  xor2s1 _____9_496414(.DIN1 (____0____40738), .DIN2 (____9____38934),
       .Q (___900___38981));
  nnd2s1 _______496415(.DIN1 (____9____38942), .DIN2
       (__________________________________________________________________22002),
       .Q (___90____39010));
  xor2s1 ______496416(.DIN1 (____9____38929), .DIN2 (_____00__38517),
       .Q (___90_9__39014));
  nnd2s1 _______496417(.DIN1 (___9__9__39218), .DIN2 (___9_____39414),
       .Q (____99___38972));
  xnr2s1 _______496418(.DIN1 (___090__23301), .DIN2 (____0_0__40740),
       .Q (____99___38971));
  nor2s1 _______496419(.DIN1 (____9____38919), .DIN2 (___9__9__39218),
       .Q (____99___38970));
  hi1s1 _______496420(.DIN (____9_9__38968), .Q (____990__38969));
  nor2s1 _____0_496421(.DIN1 (___90____38999), .DIN2 (____9____38933),
       .Q (____9____38967));
  nnd2s1 ______496422(.DIN1 (___9__9__39218), .DIN2 (____9_0__38951),
       .Q (___90____39002));
  nnd2s1 ______496423(.DIN1 (____9____38966), .DIN2
       (_____________22087), .Q (___900___38983));
  nor2s1 _____0_496424(.DIN1 (_____________22087), .DIN2
       (____9____38966), .Q (___90____39006));
  nor2s1 _______496425(.DIN1 (_________38745), .DIN2 (____9____38965),
       .Q (___90____39000));
  nor2s1 _____496426(.DIN1 (____9____38932), .DIN2 (___9__9__39218), .Q
       (___9_____39082));
  or2s1 _______496427(.DIN1 (____9____38963), .DIN2 (____9_0__38924),
       .Q (____9____38964));
  and2s1 _______496428(.DIN1 (___9_____39401), .DIN2 (____9____38961),
       .Q (____9____38962));
  nor2s1 _______496429(.DIN1 (_________38870), .DIN2 (____9____38928),
       .Q (____9_0__38960));
  hi1s1 _______496430(.DIN (___9_____39211), .Q (____9_9__38959));
  nnd2s1 ______496431(.DIN1 (____9____38957), .DIN2 (_________38765),
       .Q (____9____38958));
  dffacs1 ______________________________________________0_496432(.CLRB
       (reset), .CLK (clk), .DIN (____9____38925), .QN
       (__________________________________________________________________22009));
  xor2s1 _______496433(.DIN1 (____9____38910), .DIN2 (_________38271),
       .Q (___90____38991));
  dffacs1 _____________________________________________9_496434(.CLRB
       (reset), .CLK (clk), .DIN (____9____38926), .QN
       (_________________________________________9___21874));
  nnd2s1 ______496435(.DIN1 (____0_0__40740), .DIN2 (____99___38034),
       .Q (____9____38956));
  nnd2s1 _____496436(.DIN1 (____9____38921), .DIN2 (___9__9__39459), .Q
       (____9____38955));
  nor2s1 ______496437(.DIN1 (_________38725), .DIN2 (____9____38953),
       .Q (____9____38954));
  xor2s1 _______496438(.DIN1 (____9_0__38951), .DIN2 (_____0___36285),
       .Q (____9____38952));
  nnd2s1 _____9_496439(.DIN1 (___90____38999), .DIN2 (____9____38949),
       .Q (____9_9__38950));
  nor2s1 _______496440(.DIN1 (____9____38961), .DIN2 (___9_____39401),
       .Q (___900___38979));
  xor2s1 _______496441(.DIN1 (____9____38902), .DIN2 (____9____38948),
       .Q (____9_9__38968));
  dffacs1 _______________________________________________496442(.CLRB
       (reset), .CLK (clk), .DIN (____9____38927), .QN
       (___0__9__40480));
  nnd2s1 _______496443(.DIN1 (___90____38999), .DIN2 (_________38832),
       .Q (___9_____39207));
  hi1s1 _______496444(.DIN (___9_____39401), .Q (____9____38947));
  or2s1 _______496445(.DIN1 (____9____38913), .DIN2 (_________38471),
       .Q (____9____38946));
  xor2s1 _______496446(.DIN1 (____0____40742), .DIN2 (____9____38944),
       .Q (____9____38945));
  nnd2s1 ______496447(.DIN1 (________25800), .DIN2 (____9____38914), .Q
       (____9____38943));
  xor2s1 _______496448(.DIN1 (____9____38922), .DIN2 (____9_0__38941),
       .Q (____9____38942));
  nnd2s1 _______496449(.DIN1 (____9_9__38923), .DIN2 (____9____38939),
       .Q (____9_9__38940));
  xor2s1 _______496450(.DIN1 (____9____38897), .DIN2 (______9__38864),
       .Q (____9____38938));
  hi1s1 _____9_496451(.DIN (____9____38936), .Q (____9____38937));
  nnd2s1 _____9_496452(.DIN1 (____9_0__38916), .DIN2 (_____0___38518),
       .Q (___9_____39211));
  xor2s1 _______496453(.DIN1 (____9____38920), .DIN2 (____9____38934),
       .Q (____9____38935));
  hi1s1 _______496454(.DIN (____9____38932), .Q (____9____38933));
  dffacs1 ________________________________________________496455(.CLRB
       (reset), .CLK (clk), .DIN (____9____38917), .Q
       (______________________________________________21913));
  xor2s1 _______496456(.DIN1 (____90___38894), .DIN2 (___9_____39312),
       .Q (____9____38966));
  dffacs1 ________________________________________________496457(.CLRB
       (reset), .CLK (clk), .DIN (____9____38911), .QN
       (______________________________________________21903));
  dffacs1 ______________________________________496458(.CLRB (reset),
       .CLK (clk), .DIN (____9____38912), .QN (___0_____40584));
  hi1s1 ______496459(.DIN (___90____38999), .Q (___9__9__39218));
  xor2s1 _______496460(.DIN1 (______0__38477), .DIN2 (____9_9__38915),
       .Q (____9____38929));
  and2s1 _______496461(.DIN1 (____0____40742), .DIN2 (______0__38827),
       .Q (____9____38928));
  nnd2s1 _______496462(.DIN1 (____9____38899), .DIN2 (________25912),
       .Q (____9____38927));
  nor2s1 _______496463(.DIN1 (_________38583), .DIN2 (____9____38901),
       .Q (____9____38926));
  nnd2s1 _______496464(.DIN1 (________23899), .DIN2
       (__________________________________________0___21944), .Q
       (____9____38925));
  nor2s1 ______496465(.DIN1
       (__________________________________________0___21944), .DIN2
       (_________38348), .Q (____9_0__38924));
  hi1s1 _______496466(.DIN (____9_9__38923), .Q (____9____38957));
  nor2s1 _____0_496467(.DIN1
       (__________________________________________________________________22002),
       .DIN2 (____9____38922), .Q (____9____38936));
  xor2s1 _______496468(.DIN1 (____0____40744), .DIN2 (_________38729),
       .Q (___9_____39401));
  nor2s1 _______496469(.DIN1 (____909__38895), .DIN2 (____9____38920),
       .Q (____9____38921));
  xor2s1 ______496470(.DIN1 (___9__9__39487), .DIN2 (____9____38944),
       .Q (____9____38918));
  dffacs1 _____________________________________________9_496471(.CLRB
       (reset), .CLK (clk), .DIN (____90___38891), .QN
       (_________________________________________9___21901));
  nnd2s1 _______496472(.DIN1 (____9____38920), .DIN2 (____90___38890),
       .Q (____9____38932));
  xor2s1 ______496473(.DIN1 (_________38456), .DIN2 (____9____38934),
       .Q (____9____38953));
  dffacs1 _________________________________________9_____496474(.CLRB
       (reset), .CLK (clk), .DIN (____9____38900), .Q
       (_____________________________________9_______21883));
  xor2s1 _______496475(.DIN1 (_____9___38884), .DIN2 (_________38301),
       .Q (___90____38999));
  nnd2s1 _______496476(.DIN1 (_____9___38886), .DIN2 (________24493),
       .Q (____9____38917));
  nnd2s1 _______496477(.DIN1 (____9_9__38915), .DIN2 (_____99__38516),
       .Q (____9_0__38916));
  xor2s1 _______496478(.DIN1 (______9__38879), .DIN2 (___0____22347),
       .Q (____9____38914));
  hi1s1 _______496479(.DIN
       (__________________________________________0___21944), .Q
       (____9____38913));
  or2s1 _______496480(.DIN1 (_____9___38885), .DIN2 (_________38787),
       .Q (____9____38912));
  nnd2s1 ______496481(.DIN1 (_____9___38887), .DIN2 (________27100), .Q
       (____9____38911));
  nor2s1 _____0_496482(.DIN1 (_____9__28998), .DIN2 (____90___38889),
       .Q (____9____38910));
  xor2s1 _______496483(.DIN1 (_________38878), .DIN2 (____9____38909),
       .Q (____9_9__38923));
  dffacs1 ________________496484(.CLRB (reset), .CLK (clk), .DIN
       (____9____38934), .Q (outData[25]));
  nor2s1 _______496485(.DIN1 (____0____38099), .DIN2 (___9__9__39487),
       .Q (____9____38908));
  nnd2s1 _______496486(.DIN1 (____9____38934), .DIN2 (______9__38854),
       .Q (____9____38907));
  nor2s1 _______496487(.DIN1 (____9_9__38905), .DIN2 (____9____38904),
       .Q (____9_0__38906));
  and2s1 _______496488(.DIN1 (____9____38904), .DIN2 (____9_9__38905),
       .Q (____9____38903));
  nor2s1 _______496489(.DIN1 (_________33049), .DIN2 (____9____38934),
       .Q (____9____38902));
  nnd2s1 _____9_496490(.DIN1 (____9____38934), .DIN2 (_________38853),
       .Q (____9____38919));
  nor2s1 _____9_496491(.DIN1 (_________38851), .DIN2 (____9____38934),
       .Q (____9_0__38951));
  nor2s1 _____9_496492(.DIN1 (_________38852), .DIN2 (____9____38934),
       .Q (____9____38930));
  xor2s1 _______496493(.DIN1 (____9___29000), .DIN2 (____900__38888),
       .Q (____9____38901));
  nnd2s1 _______496494(.DIN1 (_____9___38608), .DIN2 (_________38875),
       .Q (____9____38900));
  or2s1 _______496495(.DIN1 (____9____38898), .DIN2 (_____9___38881),
       .Q (____9____38899));
  nnd2s1 _______496496(.DIN1 (____9_0__38896), .DIN2 (______9__38844),
       .Q (____9____38897));
  nnd2s1 _______496497(.DIN1 (______0__38865), .DIN2 (____9_0__38896),
       .Q (___9__9__39088));
  hi1s1 ______496498(.DIN (____9_9__38915), .Q (____9____38922));
  dffacs1 ______________________________________________0_496499(.CLRB
       (reset), .CLK (clk), .DIN (_____90__38880), .Q
       (__________________________________________0___21944));
  xor2s1 _______496500(.DIN1 (_________38848), .DIN2 (___9_____39384),
       .Q (____909__38895));
  nor2s1 _____0_496501(.DIN1 (________23004), .DIN2 (_________38874),
       .Q (____90___38894));
  nor2s1 _______496502(.DIN1 (____90___38892), .DIN2 (_____9___38883),
       .Q (____90___38893));
  nnd2s1 _______496503(.DIN1 (_____9___38882), .DIN2 (_________37539),
       .Q (____90___38891));
  nor2s1 _______496504(.DIN1
       (__________________________________________________________________21989),
       .DIN2 (____90___38890), .Q (___90_9__39004));
  xor2s1 _____9_496505(.DIN1 (_________38849), .DIN2 (___9_____39511),
       .Q (____9____38920));
  nor2s1 _______496506(.DIN1 (____90__28999), .DIN2 (____900__38888),
       .Q (____90___38889));
  nnd2s1 _______496507(.DIN1 (_________38861), .DIN2 (inData[22]), .Q
       (_____9___38887));
  nnd2s1 _______496508(.DIN1 (_________38859), .DIN2 (________23899),
       .Q (_____9___38886));
  nnd2s1 ______496509(.DIN1 (______0__38631), .DIN2 (_________38862),
       .Q (_____9___38885));
  xor2s1 _______496510(.DIN1 (_________38840), .DIN2 (_____9___38793),
       .Q (____9_9__38915));
  xor2s1 ______496511(.DIN1 (________23005), .DIN2 (______0__38873), .Q
       (_____9___38884));
  dffacs1 _______________________________________________496512(.CLRB
       (reset), .CLK (clk), .DIN (_________38863), .Q (___0_0___40462));
  nnd2s1 _______496513(.DIN1 (___9_____39263), .DIN2 (_________38850),
       .Q (____9____38904));
  dffacs1 __________________________________________0_____496514(.CLRB
       (reset), .CLK (clk), .DIN (______0__38855), .Q (___0__0__40619));
  dffacs1 _________________________________________9_____496515(.CLRB
       (reset), .CLK (clk), .DIN (_________38857), .Q (___0_9___40455));
  hi1s1 _______496516(.DIN (_____9___38883), .Q (___9__9__39487));
  hi1s1 _______496517(.DIN (____90___38890), .Q (____9____38934));
  nnd2s1 _____9_496518(.DIN1 (______0__38770), .DIN2 (_________38846),
       .Q (_____9___38882));
  xor2s1 _______496519(.DIN1 (_________38823), .DIN2 (________27618),
       .Q (_____9___38881));
  nnd2s1 _____496520(.DIN1 (_________38839), .DIN2 (_________38567), .Q
       (_____90__38880));
  xor2s1 _____9_496521(.DIN1 (______9__22034), .DIN2 (___0_9___40456),
       .Q (______9__38879));
  xor2s1 _____9_496522(.DIN1 (______0__38820), .DIN2 (_________38830),
       .Q (_________38878));
  nnd2s1 _____0_496523(.DIN1 (______0__38845), .DIN2
       (______________________________________________21930), .Q
       (____9_0__38896));
  dffacs1 ________________________________________________496524(.CLRB
       (reset), .CLK (clk), .DIN (_________38835), .QN
       (____________________________________________));
  nnd2s1 _____0_496525(.DIN1 (______0__38837), .DIN2 (inData[22]), .Q
       (_________38875));
  nor2s1 _______496526(.DIN1 (________23003), .DIN2 (______0__38873),
       .Q (_________38874));
  xor2s1 _______496527(.DIN1 (_________38736), .DIN2 (___9_____39414),
       .Q (_____9___38883));
  xor2s1 _______496528(.DIN1 (_________38815), .DIN2
       (______________22111), .Q (____90___38890));
  nor2s1 _______496529(.DIN1 (______9__38819), .DIN2 (_________38831),
       .Q (___90_0__39015));
  nor2s1 _______496530(.DIN1 (_________38869), .DIN2 (_________38867),
       .Q (_________38870));
  nnd2s1 _______496531(.DIN1 (_________38867), .DIN2 (_________38869),
       .Q (_________38868));
  xor2s1 _____496532(.DIN1 (_____0___38807), .DIN2
       (______________________________________________21956), .Q
       (_________38866));
  or2s1 _______496533(.DIN1 (_________38843), .DIN2 (______9__38864),
       .Q (______0__38865));
  or2s1 _____496534(.DIN1 (_________38633), .DIN2 (_________38821), .Q
       (_________38863));
  or2s1 _____0_496535(.DIN1 (______9__22034), .DIN2 (______0__38711),
       .Q (_________38862));
  nor2s1 _____0_496536(.DIN1 (_________38816), .DIN2 (_________36753),
       .Q (_________38861));
  xor2s1 _____9_496537(.DIN1 (______0__38810), .DIN2 (_________38860),
       .Q (____900__38888));
  xor2s1 _______496538(.DIN1 (_________38778), .DIN2 (_________38828),
       .Q (_________38859));
  xor2s1 _______496539(.DIN1 (_____9___38798), .DIN2 (___9_____39738),
       .Q (_________38858));
  nnd2s1 ______496540(.DIN1 (_________38818), .DIN2 (_________38856),
       .Q (_________38857));
  nnd2s1 _______496541(.DIN1 (_________38817), .DIN2 (________25276),
       .Q (______0__38855));
  hi1s1 _______496542(.DIN (_________38853), .Q (______9__38854));
  hi1s1 _______496543(.DIN (_________38851), .Q (_________38852));
  nnd2s1 _______496544(.DIN1 (___9_____39414), .DIN2 (_____9___41370),
       .Q (_________38850));
  nor2s1 _______496545(.DIN1 (_________38847), .DIN2 (___9_____39414),
       .Q (_________38849));
  nnd2s1 _______496546(.DIN1 (___9_____39414), .DIN2 (_________38847),
       .Q (_________38848));
  dffacs1 _______________________________________________496547(.CLRB
       (reset), .CLK (clk), .DIN (_________38824), .QN
       (_____________________________________________21845));
  nnd2s1 _______496548(.DIN1 (_____0___38802), .DIN2 (_________38811),
       .Q (_________38846));
  xor2s1 _______496549(.DIN1 (___09____40665), .DIN2 (_________41264),
       .Q (______0__38845));
  hi1s1 _______496550(.DIN (_________38843), .Q (______9__38844));
  nor2s1 _______496551(.DIN1 (_____9___38794), .DIN2 (______9__38836),
       .Q (_________38840));
  nnd2s1 _______496552(.DIN1 (_____0___38808), .DIN2 (_________38838),
       .Q (_________38839));
  nor2s1 _______496553(.DIN1 (_____0___38803), .DIN2 (_________38638),
       .Q (______0__38837));
  nor2s1 _______496554(.DIN1 (______9__38836), .DIN2 (_____9___38795),
       .Q (___909___39069));
  nnd2s1 _______496555(.DIN1 (_____09__38809), .DIN2 (_____0__26794),
       .Q (_________38835));
  or2s1 _______496556(.DIN1 (_________38833), .DIN2 (_________38832),
       .Q (_________38834));
  and2s1 _______496557(.DIN1 (_____0___38805), .DIN2 (_________38830),
       .Q (_________38831));
  nnd2s1 _______496558(.DIN1 (_________38832), .DIN2 (_________38748),
       .Q (_________38829));
  nor2s1 _______496559(.DIN1 (_________38737), .DIN2 (_________38832),
       .Q (_________38877));
  nor2s1 _______496560(.DIN1 (_________38738), .DIN2 (_________38832),
       .Q (_________38851));
  nnd2s1 _______496561(.DIN1 (_________38832), .DIN2 (_________38747),
       .Q (_________38853));
  nnd2s1 _______496562(.DIN1 (_________38764), .DIN2 (_________38828),
       .Q (_________38872));
  nor2s1 _______496563(.DIN1 (_____0__22519), .DIN2 (_____00__38800),
       .Q (______0__38873));
  nnd2s1 _______496564(.DIN1 (_________38832), .DIN2 (_____0___38708),
       .Q (___9_____39263));
  nnd2s1 _______496565(.DIN1 (______9__38826), .DIN2 (_________38825),
       .Q (______0__38827));
  or2s1 _____0_496566(.DIN1 (____0___24937), .DIN2 (_________38785), .Q
       (_________38824));
  xor2s1 _______496567(.DIN1
       (_____________________________________________21845), .DIN2
       (_________38775), .Q (_________38823));
  nor2s1 _______496568(.DIN1 (___9_0__25988), .DIN2 (_________38786),
       .Q (_________38821));
  or2s1 ______496569(.DIN1 (_________38825), .DIN2 (______9__38826), .Q
       (_________38867));
  dffacs1 _________________________________________9_____496570(.CLRB
       (reset), .CLK (clk), .DIN (_________38788), .QN
       (______9__22034));
  nor2s1 _______496571(.DIN1
       (______________________________________________21930), .DIN2
       (___09____40665), .Q (_________38843));
  nor2s1 _______496572(.DIN1 (_____0___38804), .DIN2 (______9__38819),
       .Q (______0__38820));
  and2s1 _______496573(.DIN1 (______9__38779), .DIN2 (____9___25857),
       .Q (_________38818));
  nnd2s1 ______496574(.DIN1 (_________38777), .DIN2 (___9__9__39459),
       .Q (_________38817));
  xor2s1 _______496575(.DIN1
       (_________________________________________9___21901), .DIN2
       (_____0___38801), .Q (_________38816));
  xor2s1 _______496576(.DIN1 (_____________22085), .DIN2
       (_____99__38799), .Q (_________38815));
  or2s1 _____0_496577(.DIN1 (___90____39051), .DIN2 (_________38782),
       .Q (_________38814));
  dffacs1 ________________________________________________496578(.CLRB
       (reset), .CLK (clk), .DIN (_________38784), .Q
       (______________________________________________21912));
  dffacs1 __________________________________________0_____496579(.CLRB
       (reset), .CLK (clk), .DIN (______9__38789), .QN
       (______________________________________0_______21890));
  hi1s1 _______496580(.DIN (_________38832), .Q (___9_____39414));
  xor2s1 ______496581(.DIN1 (_________38812), .DIN2 (___9_0___39624),
       .Q (_________38813));
  nnd2s1 _______496582(.DIN1 (_________38768), .DIN2 (____9____37062),
       .Q (_________38811));
  nnd2s1 ______496583(.DIN1 (_________38755), .DIN2 (_________38773),
       .Q (______0__38810));
  nnd2s1 _______496584(.DIN1 (_________38771), .DIN2 (inData[26]), .Q
       (_____09__38809));
  xor2s1 _______496585(.DIN1 (______0__38750), .DIN2 (______0__38721),
       .Q (_____0___38808));
  xor2s1 ______496586(.DIN1 (_____9___38791), .DIN2 (____0_0__38084),
       .Q (_____0___38807));
  and2s1 _______496587(.DIN1 (_____0___38806), .DIN2 (______0__37450),
       .Q (______9__38836));
  nnd2s1 _______496588(.DIN1 (______9__38769), .DIN2 (_________38642),
       .Q (_________38841));
  hi1s1 ______496589(.DIN (_____0___38804), .Q (_____0___38805));
  xnr2s1 _______496590(.DIN1 (_____________22087), .DIN2
       (_________38649), .Q (_____0___38803));
  nnd2s1 _______496591(.DIN1 (_____0___38801), .DIN2 (_________38767),
       .Q (_____0___38802));
  nor2s1 _____0_496592(.DIN1 (____0__22281), .DIN2 (_____99__38799), .Q
       (_____00__38800));
  nnd2s1 _______496593(.DIN1 (_____9___38797), .DIN2 (_____9___38796),
       .Q (_____9___38798));
  nnd2s1 _______496594(.DIN1 (_________38758), .DIN2 (______9__37240),
       .Q (_________38828));
  dffacs1 _____________________________________________0_496595(.CLRB
       (reset), .CLK (clk), .DIN (_________38774), .Q
       (_________________________________________0___21862));
  xnr2s1 _____9_496596(.DIN1 (______________22110), .DIN2
       (______9__38739), .Q (_________38832));
  nor2s1 _______496597(.DIN1 (_____9___38794), .DIN2 (_____9___38793),
       .Q (_____9___38795));
  nor2s1 _______496598(.DIN1
       (______________________________________________21956), .DIN2
       (_____9___38791), .Q (_____9___38792));
  and2s1 _______496599(.DIN1 (_____9___38791), .DIN2
       (______________________________________________21956), .Q
       (_____90__38790));
  nnd2s1 ______496600(.DIN1 (______9__38749), .DIN2 (___00___24172), .Q
       (______9__38789));
  or2s1 _______496601(.DIN1 (_________38787), .DIN2 (_________38756),
       .Q (_________38788));
  nor2s1 _______496602(.DIN1 (_________38752), .DIN2 (_________38772),
       .Q (_________38786));
  nor2s1 ______496603(.DIN1 (____9____38898), .DIN2 (_________38753),
       .Q (_________38785));
  and2s1 ______496604(.DIN1 (_____9___38791), .DIN2 (_________38776),
       .Q (______9__38819));
  xor2s1 _______496605(.DIN1 (_________38734), .DIN2 (_________38358),
       .Q (______9__38826));
  or2s1 _____0_496606(.DIN1 (_____9__26194), .DIN2 (_________38742), .Q
       (_________38784));
  xor2s1 _____9_496607(.DIN1 (_________38761), .DIN2 (______0__37673),
       .Q (_________38783));
  xor2s1 _______496608(.DIN1 (_________37263), .DIN2 (_________38757),
       .Q (_________38782));
  xor2s1 _______496609(.DIN1 (________27618), .DIN2 (______0__38780),
       .Q (_________38781));
  nor2s1 _____0_496610(.DIN1 (________26535), .DIN2 (_________38744),
       .Q (______9__38779));
  xor2s1 _____496611(.DIN1 (_________37531), .DIN2
       (__________________________________________________________________21984),
       .Q (_________38778));
  nnd2s1 _______496612(.DIN1 (_________38847), .DIN2 (_________38741),
       .Q (_________38777));
  nnd2s1 _______496613(.DIN1 (____9_9__38905), .DIN2 (_________38746),
       .Q (___9_9___39158));
  nor2s1 _____9_496614(.DIN1 (_________38776), .DIN2 (_____9___38791),
       .Q (_____0___38804));
  nnd2s1 _____9_496615(.DIN1 (_________38754), .DIN2 (_________38724),
       .Q (_________38822));
  dffacs1 _____________________________________________9_496616(.CLRB
       (reset), .CLK (clk), .DIN (______0__38740), .QN
       (___0_____40504));
  xor2s1 _______496617(.DIN1 (_____00__38702), .DIN2 (___9__9__39125),
       .Q (_________38775));
  nnd2s1 _______496618(.DIN1 (_________38732), .DIN2 (________26642),
       .Q (_________38774));
  nnd2s1 _______496619(.DIN1 (_________38772), .DIN2 (_________38591),
       .Q (_________38773));
  and2s1 _____0_496620(.DIN1 (______0__38770), .DIN2
       (__________________________________________________________________21984),
       .Q (_________38771));
  xor2s1 ______496621(.DIN1 (_________38717), .DIN2 (___9_____39582),
       .Q (______9__38769));
  nnd2s1 _____0_496622(.DIN1
       (__________________________________________________________________21984),
       .DIN2 (_________38767), .Q (_________38768));
  xor2s1 _____9_496623(.DIN1 (_________38766), .DIN2 (_____9___41303),
       .Q (_____0___38806));
  hi1s1 ______496624(.DIN (_________38765), .Q (____9____38939));
  dffacs1 _______________________________________496625(.CLRB (reset),
       .CLK (clk), .DIN (______0__38731), .QN (______________22112));
  or2s1 _______496626(.DIN1
       (__________________________________________________________________21984),
       .DIN2 (_________37617), .Q (_________38764));
  and2s1 _______496627(.DIN1 (_________37531), .DIN2
       (__________________________________________________________________21984),
       .Q (_________38763));
  and2s1 _______496628(.DIN1 (_________38761), .DIN2 (______9__38759),
       .Q (_________38762));
  or2s1 _______496629(.DIN1 (______9__38759), .DIN2 (_________38761),
       .Q (______0__38760));
  or2s1 _____496630(.DIN1 (_________37239), .DIN2 (_________38757), .Q
       (_________38758));
  nor2s1 _______496631(.DIN1 (____0), .DIN2 (_________38728), .Q
       (_____99__38799));
  and2s1 _______496632(.DIN1
       (__________________________________________________________________21984),
       .DIN2 (____________________________________________), .Q
       (_____0___38801));
  xor2s1 ______496633(.DIN1 (_____0___38703), .DIN2 (_________37864),
       .Q (_____9___38797));
  nnd2s1 _____0_496634(.DIN1 (_________38268), .DIN2 (_________38712),
       .Q (_________38756));
  nnd2s1 _______496635(.DIN1 (_________38723), .DIN2 (_________36291),
       .Q (_________38755));
  xor2s1 ______496636(.DIN1 (______9__38682), .DIN2 (____9_0__38941),
       .Q (_________38754));
  xor2s1 _______496637(.DIN1 (_____9___38694), .DIN2 (________22381),
       .Q (_________38753));
  nor2s1 _______496638(.DIN1 (_________38715), .DIN2 (_________38627),
       .Q (_________38752));
  nor2s1 _____496639(.DIN1 (___09____40664), .DIN2 (___9____25081), .Q
       (_________38751));
  xor2s1 _______496640(.DIN1 (_____9___38697), .DIN2 (___0_____40433),
       .Q (______0__38750));
  nnd2s1 _____0_496641(.DIN1 (_____09__38710), .DIN2 (___90____39040),
       .Q (______9__38749));
  nor2s1 ______496642(.DIN1 (_________37541), .DIN2 (_________38766),
       .Q (_____9___38794));
  xor2s1 _______496643(.DIN1 (_____90__38693), .DIN2 (____9____38007),
       .Q (_____9___38796));
  nor2s1 _____9_496644(.DIN1 (_________38357), .DIN2 (_________38718),
       .Q (_________38765));
  nor2s1 _______496645(.DIN1 (_________38670), .DIN2 (_________38722),
       .Q (______9__38864));
  hi1s1 _______496646(.DIN (_________38747), .Q (_________38748));
  nnd2s1 _____9_496647(.DIN1 (_________38745), .DIN2 (___09_9__40689),
       .Q (_________38746));
  nor2s1 _______496648(.DIN1 (_________38743), .DIN2 (_____9___38700),
       .Q (_________38744));
  nor2s1 ______496649(.DIN1 (___90____39051), .DIN2 (_____99__38701),
       .Q (_________38742));
  nnd2s1 _______496650(.DIN1 (_____0___38706), .DIN2 (_________38636),
       .Q (_________38741));
  nnd2s1 _______496651(.DIN1 (_____0___38707), .DIN2 (_________38550),
       .Q (______0__38740));
  xor2s1 _______496652(.DIN1 (___0_____40584), .DIN2 (_________38727),
       .Q (______9__38739));
  hi1s1 _______496653(.DIN (_________38737), .Q (_________38738));
  nor2s1 _______496654(.DIN1 (_________38686), .DIN2 (_____0___38709),
       .Q (_________38736));
  xor2s1 _______496655(.DIN1 (_________38726), .DIN2 (_________37884),
       .Q (_________38812));
  dffacs1 ______________________________________496656(.CLRB (reset),
       .CLK (clk), .DIN (_____0___38704), .QN (_____________22087));
  xor2s1 _______496657(.DIN1 (_________38592), .DIN2 (_________38681),
       .Q (_____9___38791));
  xor2s1 _____9_496658(.DIN1 (_________38719), .DIN2 (_________38643),
       .Q (_________38735));
  xor2s1 _____9_496659(.DIN1 (_________38733), .DIN2 (_________38359),
       .Q (_________38734));
  nnd2s1 _____496660(.DIN1 (_____9___38695), .DIN2 (_____9___37943), .Q
       (_________38732));
  nnd2s1 _______496661(.DIN1 (________26558), .DIN2 (_____9___38699),
       .Q (______0__38731));
  and2s1 _______496662(.DIN1 (___0_____40380), .DIN2 (_________38691),
       .Q (______9__38730));
  nor2s1 _______496663(.DIN1 (_________38714), .DIN2 (______9__38672),
       .Q (_________38772));
  nnd2s1 _______496664(.DIN1 (_____0___38705), .DIN2 (_________38729),
       .Q (_________38847));
  nor2s1 _______496665(.DIN1 (_______22236), .DIN2 (_________38727), .Q
       (_________38728));
  nnd2s1 ______496666(.DIN1 (_________38685), .DIN2 (_________38636),
       .Q (_________38747));
  nnd2s1 _______496667(.DIN1 (______0__38683), .DIN2 (_________38729),
       .Q (_________38737));
  nor2s1 ____9__496668(.DIN1 (_________38600), .DIN2 (_________38677),
       .Q (_________38757));
  nor2s1 _______496669(.DIN1 (________29221), .DIN2 (_________38679),
       .Q (______0__38780));
  or2s1 _______496670(.DIN1 (_________38687), .DIN2 (_________38726),
       .Q (_________38761));
  nnd2s1 ____90_496671(.DIN1 (_________38725), .DIN2 (_________38724),
       .Q (____9_9__38905));
  dffacs1 ________________________________________________496672(.CLRB
       (reset), .CLK (clk), .DIN (______9__38692), .QN
       (__________________________________________________________________21984));
  nnd2s1 _____496673(.DIN1 (______0__38673), .DIN2 (_________38688), .Q
       (_________38723));
  and2s1 _______496674(.DIN1 (______0__38721), .DIN2 (_________38668),
       .Q (_________38722));
  nor2s1 ______496675(.DIN1 (_________38716), .DIN2 (_________38719),
       .Q (______9__38720));
  and2s1 _______496676(.DIN1 (_________38733), .DIN2 (_________38360),
       .Q (_________38718));
  nnd2s1 _______496677(.DIN1 (_________38719), .DIN2 (_________38716),
       .Q (_________38717));
  hi1s1 _______496678(.DIN (_________38714), .Q (_________38715));
  nnd2s1 _______496679(.DIN1 (_____9___38509), .DIN2 (_________38674),
       .Q (_________38713));
  nnd2s1 _______496680(.DIN1 (______0__38711), .DIN2 (_________38667),
       .Q (_________38712));
  xor2s1 _______496681(.DIN1 (_________38689), .DIN2 (_________38690),
       .Q (_____09__38710));
  nor2s1 ______496682(.DIN1 (_________38659), .DIN2 (_____0___38708),
       .Q (_____0___38709));
  and2s1 ____9__496683(.DIN1 (______9__38647), .DIN2 (____0____40746),
       .Q (_____0___38707));
  hi1s1 ______496684(.DIN (_____0___38705), .Q (_____0___38706));
  or2s1 _______496685(.DIN1 (____0____40748), .DIN2 (______0__38664),
       .Q (_____0___38704));
  nnd2s1 _______496686(.DIN1 (_________38652), .DIN2
       (__________________________________________9_), .Q
       (_____0___38703));
  nor2s1 ______496687(.DIN1 (_____0___38619), .DIN2 (_________38661),
       .Q (_____00__38702));
  xor2s1 _____9_496688(.DIN1 (_____0___38614), .DIN2 (_________38676),
       .Q (_____99__38701));
  xor2s1 _____9_496689(.DIN1 (________29222), .DIN2 (_________38678),
       .Q (_____9___38700));
  nor2s1 ____90_496690(.DIN1 (_________38492), .DIN2 (_________38663),
       .Q (_____9___38793));
  hi1s1 ____9__496691(.DIN (_________38725), .Q (_________38745));
  xor2s1 _______496692(.DIN1 (______9__38506), .DIN2 (_____9___41370),
       .Q (_________38766));
  nnd2s1 _______496693(.DIN1 (_________38657), .DIN2 (inData[26]), .Q
       (_____9___38699));
  nnd2s1 ______496694(.DIN1 (______9__38655), .DIN2 (___9__9__39659),
       .Q (_____9___38698));
  xor2s1 _______496695(.DIN1 (_________38669), .DIN2 (_____9___38610),
       .Q (_____9___38697));
  nor2s1 _____9_496696(.DIN1 (_________38684), .DIN2 (_____9___41370),
       .Q (_____9___38696));
  xor2s1 _______496697(.DIN1 (______0__38640), .DIN2 (_________38660),
       .Q (_____9___38695));
  xor2s1 _______496698(.DIN1
       (_____________________________________________21828), .DIN2
       (______9__38602), .Q (_____9___38694));
  nor2s1 _______496699(.DIN1
       (__________________________________________9_), .DIN2
       (_____0___38708), .Q (_____90__38693));
  nnd2s1 _______496700(.DIN1 (_________38653), .DIN2 (___009__26959),
       .Q (______9__38692));
  nnd2s1 ______496701(.DIN1 (_________38654), .DIN2 (inData[2]), .Q
       (_________38691));
  nor2s1 _______496702(.DIN1 (_________38690), .DIN2 (_________38689),
       .Q (_____0___38705));
  dffacs1 _______________________________________________496703(.CLRB
       (reset), .CLK (clk), .DIN (______0__38656), .Q (___0_0___40463));
  nnd2s1 _______496704(.DIN1 (_________38671), .DIN2 (_________38688),
       .Q (_________38714));
  nor2s1 _____9_496705(.DIN1 (_________38386), .DIN2 (_____0___38708),
       .Q (_________38687));
  nor2s1 _____9_496706(.DIN1 (_________38645), .DIN2 (_________38689),
       .Q (_________38686));
  nnd2s1 _____496707(.DIN1 (_____0___38708), .DIN2 (_________38684), .Q
       (_________38685));
  nnd2s1 ____900(.DIN1 (_____9___41370), .DIN2 (_________38658), .Q
       (______0__38683));
  nor2s1 ____90_496708(.DIN1 (_________38439), .DIN2 (_____0___38708),
       .Q (______9__38682));
  xor2s1 ____90_496709(.DIN1 (_________38662), .DIN2 (_________38680),
       .Q (_________38681));
  dffacs1 ________________496710(.CLRB (reset), .CLK (clk), .DIN
       (_________38689), .Q (outData[22]));
  nor2s1 ____9__496711(.DIN1 (________29220), .DIN2 (_________38678),
       .Q (_________38679));
  nor2s1 ____9_0(.DIN1 (_____9___38605), .DIN2 (_________38676), .Q
       (_________38677));
  dffacs1 ________________________________________________496712(.CLRB
       (reset), .CLK (clk), .DIN (_________38644), .Q
       (______________________________________________21911));
  nor2s1 ____9__496713(.DIN1 (_________38625), .DIN2 (_________38651),
       .Q (_________38727));
  nor2s1 ____90_496714(.DIN1 (_____0___38330), .DIN2 (_____9___41370),
       .Q (_________38726));
  xor2s1 ____9_496715(.DIN1 (_________38729), .DIN2 (_________38675),
       .Q (_________38725));
  xor2s1 _____9_496716(.DIN1
       (______________________________________0_______21890), .DIN2
       (___0__9__40618), .Q (_________38674));
  nnd2s1 _______496717(.DIN1 (______9__38672), .DIN2 (_________38671),
       .Q (______0__38673));
  nor2s1 _______496718(.DIN1 (___0_____40433), .DIN2 (_________38669),
       .Q (_________38670));
  nnd2s1 _______496719(.DIN1 (_________38669), .DIN2 (___0_____40433),
       .Q (_________38668));
  nnd2s1 _______496720(.DIN1 (_________38641), .DIN2 (inData[24]), .Q
       (_________38667));
  xor2s1 _______496721(.DIN1 (______9__38630), .DIN2 (_________38666),
       .Q (_________38719));
  xor2s1 ______496722(.DIN1 (_________38629), .DIN2 (____0____38106),
       .Q (_________38733));
  xor2s1 ____9__496723(.DIN1
       (__________________________________________________________________21983),
       .DIN2 (_________38636), .Q (_________38665));
  nnd2s1 ____9__496724(.DIN1 (______9__38639), .DIN2 (___0_9__26131),
       .Q (______0__38664));
  nor2s1 ____9_496725(.DIN1 (_________38500), .DIN2 (_________38662),
       .Q (_________38663));
  and2s1 _____9_496726(.DIN1 (_________38660), .DIN2 (_____0___38620),
       .Q (_________38661));
  nnd2s1 ____9__496727(.DIN1 (_________38729), .DIN2 (_________38658),
       .Q (_________38659));
  dffacs1 ______________________________________496728(.CLRB (reset),
       .CLK (clk), .DIN (_________38637), .Q (_____________22086));
  and2s1 ____9__496729(.DIN1 (________24614), .DIN2 (______0__38622),
       .Q (_________38657));
  or2s1 ______496730(.DIN1 (____0____38052), .DIN2 (_________38635), .Q
       (______0__38656));
  xor2s1 _______496731(.DIN1 (_____0___38615), .DIN2 (___9_____39511),
       .Q (______9__38655));
  xor2s1 ____9__496732(.DIN1 (____90__22634), .DIN2 (_____9___38607),
       .Q (_________38654));
  nnd2s1 ____9__496733(.DIN1 (_________37538), .DIN2 (___0__9__40618),
       .Q (_________38653));
  nnd2s1 _______496734(.DIN1 (_________41367), .DIN2 (_________38634),
       .Q (_________38688));
  hi1s1 ____9__496735(.DIN (_________38652), .Q (_________38689));
  dffacs1 _____________________________________________9_496736(.CLRB
       (reset), .CLK (clk), .DIN (_________38632), .Q
       (_________________________________________9___21861));
  hi1s1 ____9__496737(.DIN (_________38652), .Q (_____9___41370));
  nb1s1 ____9__496738(.DIN (_________38652), .Q (_____0___38708));
  and2s1 ____9__496739(.DIN1 (_________38623), .DIN2 (_________38650),
       .Q (_________38651));
  nnd2s1 ____9_496740(.DIN1 (_________38636), .DIN2
       (__________________________________________________________________21983),
       .Q (______0__38648));
  nor2s1 ____9__496741(.DIN1 (_________38626), .DIN2 (_____09__38236),
       .Q (______9__38647));
  dffacs1 ________________496742(.CLRB (reset), .CLK (clk), .DIN
       (_________38636), .Q (outData[23]));
  nor2s1 ____9__496743(.DIN1
       (__________________________________________________________________21983),
       .DIN2 (_________38636), .Q (_________38646));
  nnd2s1 ____9__496744(.DIN1 (_________38636), .DIN2 (_________38684),
       .Q (_________38645));
  nnd2s1 ____0__496745(.DIN1 (_____09__38621), .DIN2 (________24407),
       .Q (_________38644));
  xor2s1 ____0__496746(.DIN1 (_____9___38609), .DIN2 (_________38860),
       .Q (_________38676));
  nor2s1 ____9__496747(.DIN1 (______9__38574), .DIN2 (_________38624),
       .Q (_________38678));
  xor2s1 ____9__496748(.DIN1 (_________38642), .DIN2 (___9_____39554),
       .Q (_________38643));
  xnr2s1 ____9_496749(.DIN1 (___0_9___40456), .DIN2 (___0_____40584),
       .Q (_________38641));
  dffacs1 _______________________________________________496750(.CLRB
       (reset), .CLK (clk), .DIN (_____0___38618), .QN
       (_____________________________________________21828));
  nor2s1 ____9_496751(.DIN1 (_________38581), .DIN2 (_____99__38612),
       .Q (_________38660));
  nnd2s1 _______496752(.DIN1 (_________38280), .DIN2 (___0__0__40481),
       .Q (_________38671));
  dffacs1 _________________________________________0_____(.CLRB
       (reset), .CLK (clk), .DIN (_____00__38613), .QN
       (___0_09__40570));
  xor2s1 ____90_496753(.DIN1 (_________38595), .DIN2 (_____09__38526),
       .Q (_________38669));
  xor2s1 ____9__496754(.DIN1 (_____9__28896), .DIN2 (__________22060),
       .Q (______0__38640));
  or2s1 ____9__496755(.DIN1 (_________38601), .DIN2 (_________38638),
       .Q (______9__38639));
  nnd2s1 ____9__496756(.DIN1 (____0___27121), .DIN2 (_____0___38617),
       .Q (_________38637));
  nor2s1 ____9_496757(.DIN1 (_________38468), .DIN2 (_____9___38604),
       .Q (_________38662));
  xor2s1 ____9__496758(.DIN1 (_________38590), .DIN2 (_________38869),
       .Q (_________38652));
  nnd2s1 ______496759(.DIN1 (_________38598), .DIN2 (___0_____30911),
       .Q (_________38635));
  hi1s1 ____90_496760(.DIN (___0__0__40481), .Q (_________38634));
  nor2s1 ____9_496761(.DIN1 (_________38597), .DIN2 (_________38576),
       .Q (_________38633));
  nnd2s1 ____9__496762(.DIN1 (_________38596), .DIN2 (_________38190),
       .Q (_________38632));
  nnd2s1 ____9__496763(.DIN1 (______0__38711), .DIN2 (___0_9___40456),
       .Q (______0__38631));
  xor2s1 ____9__496764(.DIN1 (_________38579), .DIN2 (_________37733),
       .Q (______9__38630));
  xor2s1 ____9__496765(.DIN1 (_____90__38603), .DIN2 (_________38566),
       .Q (_________38629));
  or2s1 ____9__496766(.DIN1 (___0_9___40456), .DIN2 (______0__38711),
       .Q (_________38628));
  dffacs1 __________________________________________0_____496767(.CLRB
       (reset), .CLK (clk), .DIN (______9__38593), .Q (___0__9__40618));
  hi1s1 ____9__496768(.DIN (_________38627), .Q (______9__38672));
  nor2s1 ____9__496769(.DIN1 (__________22060), .DIN2 (____09___37180),
       .Q (_________38626));
  nor2s1 ____9__496770(.DIN1 (_________38650), .DIN2 (_________38588),
       .Q (_________38625));
  nor2s1 ____9__496771(.DIN1 (_________38573), .DIN2 (_________38586),
       .Q (_________38624));
  nnd2s1 ____9__496772(.DIN1 (______0__38585), .DIN2 (________29157),
       .Q (_________38623));
  xor2s1 ____9__496773(.DIN1 (___0_____40448), .DIN2 (_____9___38606),
       .Q (______0__38622));
  nnd2s1 ____0__496774(.DIN1 (_________38589), .DIN2 (________23899),
       .Q (_____09__38621));
  nnd2s1 ____00_(.DIN1 (________27612), .DIN2 (__________22060), .Q
       (_____0___38620));
  nor2s1 ____00_496775(.DIN1 (__________22060), .DIN2 (________27618),
       .Q (_____0___38619));
  hi1s1 ____99_496776(.DIN (_________38729), .Q (_________38636));
  or2s1 ____9__496777(.DIN1 (___9____25082), .DIN2 (_________38580), .Q
       (_____0___38618));
  nnd2s1 ____9__496778(.DIN1 (_____0___38616), .DIN2 (______0__22035),
       .Q (_____0___38617));
  xor2s1 ____9__496779(.DIN1 (_________38570), .DIN2 (_________38563),
       .Q (_____0___38615));
  xor2s1 ____9__496780(.DIN1
       (__________________________________________________________________21987),
       .DIN2 (_________38599), .Q (_____0___38614));
  or2s1 ____909(.DIN1 (_________38577), .DIN2 (___9____25989), .Q
       (_____00__38613));
  and2s1 ____9__496781(.DIN1 (_________38582), .DIN2 (_____9___38611),
       .Q (_____99__38612));
  xor2s1 ____9_496782(.DIN1 (_________38560), .DIN2 (_____9___38610),
       .Q (_________38627));
  dffacs1 _______________________________________________496783(.CLRB
       (reset), .CLK (clk), .DIN (______9__38584), .QN
       (___0__0__40481));
  nor2s1 ____09_(.DIN1 (____9____37027), .DIN2 (_________38572), .Q
       (_____9___38609));
  or2s1 ____9__496784(.DIN1 (_________38743), .DIN2 (______0__38575),
       .Q (_____9___38608));
  and2s1 ____9__496785(.DIN1 (_____9___38606), .DIN2 (___0_____40447),
       .Q (_____9___38607));
  nor2s1 ____99_496786(.DIN1 (_____9___38606), .DIN2 (___09____40688),
       .Q (_____9___38605));
  and2s1 ____00_496787(.DIN1 (_____90__38603), .DIN2 (_________38541),
       .Q (_____9___38604));
  xor2s1 ____0__496788(.DIN1 (________27618), .DIN2 (_________38556),
       .Q (______9__38602));
  nnd2s1 ____9__496789(.DIN1 (_________38649), .DIN2 (______0__22035),
       .Q (_________38601));
  nor2s1 ____99_496790(.DIN1
       (__________________________________________________________________21987),
       .DIN2 (_________38599), .Q (_________38600));
  nnd2s1 ____9__496791(.DIN1 (_________38568), .DIN2 (____9____38001),
       .Q (_________38598));
  nor2s1 ____9__496792(.DIN1 (_________38562), .DIN2 (_________38543),
       .Q (_________38597));
  nnd2s1 ____9_496793(.DIN1 (_________38561), .DIN2 (_________38249),
       .Q (_________38596));
  xor2s1 ____9__496794(.DIN1 (___09____40666), .DIN2 (_________38306),
       .Q (_________38595));
  nor2s1 _______496795(.DIN1 (___90____38993), .DIN2 (_________38559),
       .Q (______0__38594));
  nnd2s1 ____9__496796(.DIN1 (_________38557), .DIN2 (________25876),
       .Q (______9__38593));
  nnd2s1 ____9_496797(.DIN1 (______0__38565), .DIN2 (_________38569),
       .Q (______0__38721));
  dffacs1 _________________________________________9_____496798(.CLRB
       (reset), .CLK (clk), .DIN (_________38558), .Q (___0_9___40456));
  xor2s1 ____00_496799(.DIN1 (_________38538), .DIN2 (_________38591),
       .Q (_________38592));
  xor2s1 ____00_496800(.DIN1 (______0__38537), .DIN2
       (______________22108), .Q (_________38590));
  xor2s1 _____0_496801(.DIN1 (____9____37063), .DIN2 (_________38571),
       .Q (_________38589));
  nnd2s1 ____0__496802(.DIN1 (_________38587), .DIN2 (__90____29684),
       .Q (_________38588));
  nor2s1 ____0__496803(.DIN1 (__9__9__30225), .DIN2 (_________38553),
       .Q (_________38586));
  or2s1 ____0__496804(.DIN1 (________29156), .DIN2 (_________38587), .Q
       (______0__38585));
  nnd2s1 ____0__496805(.DIN1 (______0__38555), .DIN2 (_____0___38522),
       .Q (_________38642));
  nnd2s1 ____0__496806(.DIN1 (______9__38554), .DIN2 (______9__38150),
       .Q (_________38825));
  dffacs1 _____________________________________________0_496807(.CLRB
       (reset), .CLK (clk), .DIN (_________38551), .Q
       (__________22060));
  or2s1 ____9__496808(.DIN1 (_________38583), .DIN2 (_________38548),
       .Q (______9__38584));
  nnd2s1 ____9__496809(.DIN1 (_________38547), .DIN2 (_____9___35561),
       .Q (_________38582));
  nor2s1 ____9_496810(.DIN1 (_____9___38611), .DIN2 (_________38542),
       .Q (_________38581));
  nor2s1 ____00_496811(.DIN1 (____9____38898), .DIN2 (_________38549),
       .Q (_________38580));
  xor2s1 ____0__496812(.DIN1 (_________38578), .DIN2 (______0__38161),
       .Q (_________38579));
  nor2s1 ____9__496813(.DIN1 (_________38544), .DIN2 (_________38576),
       .Q (_________38577));
  hi1s1 ____0__496814(.DIN
       (__________________________________________________________________21987),
       .Q (_____9___38606));
  xor2s1 ____0__496815(.DIN1 (_________38552), .DIN2 (_________38534),
       .Q (______0__38575));
  and2s1 ____0__496816(.DIN1 (_________38535), .DIN2 (_________38573),
       .Q (______9__38574));
  and2s1 _______496817(.DIN1 (_________38571), .DIN2 (____9____37025),
       .Q (_________38572));
  xor2s1 ____0__496818(.DIN1 (_____9___38514), .DIN2 (_________38533),
       .Q (_____90__38603));
  dffacs1 _________________________________________9_____496819(.CLRB
       (reset), .CLK (clk), .DIN (______9__38536), .QN
       (______0__22035));
  dffacs1 __________________________________________0_____496820(.CLRB
       (reset), .CLK (clk), .DIN (______9__38545), .Q
       (______________________________________0_____));
  dffacs1 ______________________________________________0_496821(.CLRB
       (reset), .CLK (clk), .DIN (_________38539), .QN
       (__________________________________________0_));
  and2s1 ____009(.DIN1 (______9__38564), .DIN2 (_________38569), .Q
       (_________38570));
  xor2s1 ____9__496822(.DIN1 (_________38505), .DIN2 (_________38529),
       .Q (_________38568));
  nnd2s1 ____9__496823(.DIN1 (_________38531), .DIN2 (inData[0]), .Q
       (_________38567));
  nnd2s1 ____9__496824(.DIN1 (_________38540), .DIN2 (_____0___38525),
       .Q (_________38566));
  nnd2s1 ____99_496825(.DIN1 (______9__38564), .DIN2 (_________38563),
       .Q (______0__38565));
  xnr2s1 ____999(.DIN1 (___0_09__40570), .DIN2 (_________38502), .Q
       (_________38562));
  xor2s1 ____000(.DIN1 (_________35611), .DIN2 (______0__38546), .Q
       (_________38561));
  nnd2s1 ____00_496826(.DIN1 (_________38530), .DIN2 (______9__38486),
       .Q (_________38560));
  xor2s1 ____9__496827(.DIN1 (_________38504), .DIN2 (_________41248),
       .Q (_________38559));
  or2s1 ____0__496828(.DIN1 (_________38787), .DIN2 (_________38532),
       .Q (_________38558));
  nnd2s1 ____0_9(.DIN1 (_____9___38513), .DIN2 (___90____39040), .Q
       (_________38557));
  xor2s1 ____0__496829(.DIN1 (_________38490), .DIN2 (_________38876),
       .Q (_________38556));
  nnd2s1 ____0__496830(.DIN1 (_____0___38333), .DIN2 (_________38528),
       .Q (______0__38555));
  nnd2s1 ____0__496831(.DIN1 (_________38578), .DIN2 (_________38148),
       .Q (______9__38554));
  nor2s1 ____0__496832(.DIN1 (____9___29273), .DIN2 (_________38552),
       .Q (_________38553));
  nnd2s1 ____0__496833(.DIN1 (_____0___38519), .DIN2 (_________38550),
       .Q (_________38551));
  nor2s1 ____0__496834(.DIN1 (_______22240), .DIN2 (_____0___38521), .Q
       (_________38587));
  dffacs1 ________________________________________________496835(.CLRB
       (reset), .CLK (clk), .DIN (_____0___38524), .Q
       (__________________________________________________________________21987));
  xor2s1 ____0__496836(.DIN1 (_________38478), .DIN2 (_____9___37002),
       .Q (_________38549));
  xor2s1 ____00_496837(.DIN1 (_________38481), .DIN2 (_________41264),
       .Q (_________38548));
  nnd2s1 ____0__496838(.DIN1 (______0__38546), .DIN2 (_____9___35562),
       .Q (_________38547));
  nnd2s1 ____0__496839(.DIN1 (____0____38119), .DIN2 (_____9___38510),
       .Q (______9__38545));
  nor2s1 ____9__496840(.DIN1 (_____90__38507), .DIN2 (_________38543),
       .Q (_________38544));
  or2s1 ____0_496841(.DIN1 (_________35610), .DIN2 (______0__38546), .Q
       (_________38542));
  nnd2s1 ____0_0(.DIN1 (_________38540), .DIN2 (_________38503), .Q
       (_________38541));
  nnd2s1 _______496842(.DIN1 (_________38493), .DIN2 (___09___27029),
       .Q (_________38539));
  nor2s1 ____0__496843(.DIN1 (_________38494), .DIN2 (_________38495),
       .Q (_________38538));
  xor2s1 ____0__496844(.DIN1 (_____0___38520), .DIN2
       (_____________22084), .Q (______0__38537));
  or2s1 ____0_496845(.DIN1 (_________38787), .DIN2 (_________38499), .Q
       (______9__38536));
  nor2s1 ____0__496846(.DIN1 (_________38534), .DIN2 (_____9___38511),
       .Q (_________38535));
  xor2s1 _______496847(.DIN1 (_________38479), .DIN2 (_________38533),
       .Q (_________38571));
  dffacs1 _______________________________________________496848(.CLRB
       (reset), .CLK (clk), .DIN (_____9___38508), .Q (_________22024));
  nnd2s1 ____0_496849(.DIN1 (_________38498), .DIN2 (_________37770),
       .Q (_________38716));
  dffacs1 _____________________________________________9_496850(.CLRB
       (reset), .CLK (clk), .DIN (______0__38497), .Q (___0_____40437));
  nnd2s1 ____0_496851(.DIN1 (_________38489), .DIN2 (________25512), .Q
       (_________38532));
  nor2s1 ____0__496852(.DIN1 (_________38838), .DIN2 (_________38485),
       .Q (_________38531));
  or2s1 ____0__496853(.DIN1 (_________38483), .DIN2 (_________38529),
       .Q (_________38530));
  nnd2s1 ____0__496854(.DIN1 (______0__38527), .DIN2 (_____09__38526),
       .Q (_________38528));
  nnd2s1 ____0_496855(.DIN1 (_________38484), .DIN2 (___909___39065),
       .Q (_____0___38525));
  nnd2s1 ____0__496856(.DIN1 (_________38480), .DIN2 (___0__9__40392),
       .Q (_____0___38524));
  nnd2s1 ____0__496857(.DIN1 (_________38488), .DIN2 (__900___29641),
       .Q (______9__38564));
  hi1s1 ____0__496858(.DIN (_____0___38523), .Q (_________38578));
  or2s1 ____0__496859(.DIN1 (_____09__38526), .DIN2 (______0__38527),
       .Q (_____0___38522));
  and2s1 ____0__496860(.DIN1 (_____0___38520), .DIN2 (____0__22205), .Q
       (_____0___38521));
  and2s1 ____0_496861(.DIN1 (______9__38476), .DIN2 (___9____25990), .Q
       (_____0___38519));
  nnd2s1 _____0_496862(.DIN1 (_____00__38517), .DIN2 (_____9___38515),
       .Q (_____0___38518));
  or2s1 _____0_496863(.DIN1 (_____9___38515), .DIN2 (_____00__38517),
       .Q (_____99__38516));
  nnd2s1 _______496864(.DIN1 (_________38474), .DIN2 (_________38393),
       .Q (_____9___38514));
  xor2s1 ____0_496865(.DIN1 (_________38460), .DIN2 (_____9___38512),
       .Q (_____9___38513));
  dffacs1 _______________________________________________496866(.CLRB
       (reset), .CLK (clk), .DIN (_________38475), .QN
       (_____________________________________________21910));
  hi1s1 ____0__496867(.DIN (_____9___38511), .Q (_________38552));
  nnd2s1 ____0__496868(.DIN1 (_____9___38509), .DIN2 (______9__38466),
       .Q (_____9___38510));
  nnd2s1 ____0_496869(.DIN1 (_________38472), .DIN2 (___9_9), .Q
       (_____9___38508));
  xor2s1 ____0__496870(.DIN1 (___0_____40496), .DIN2
       (_____________________________________________21860), .Q
       (_____90__38507));
  nor2s1 ____0__496871(.DIN1 (_________38440), .DIN2 (_________38469),
       .Q (______9__38506));
  xor2s1 ____0__496872(.DIN1 (______9__36859), .DIN2
       (_____________________________________________21860), .Q
       (_________38505));
  xor2s1 ____0_496873(.DIN1 (______0__38448), .DIN2 (________22439), .Q
       (_________38504));
  nnd2s1 ____0__496874(.DIN1 (_________38501), .DIN2 (___909___39065),
       .Q (_________38503));
  nor2s1 ____0_496875(.DIN1 (___0_0___40462), .DIN2 (_________38470),
       .Q (_________38502));
  or2s1 ____0__496876(.DIN1 (___909___39065), .DIN2 (_________38501),
       .Q (_________38540));
  nnd2s1 ____0__496877(.DIN1 (______0__38487), .DIN2
       (_________________________________________9___21929), .Q
       (_________38569));
  xor2s1 ____0__496878(.DIN1 (_________38454), .DIN2 (_________36527),
       .Q (______0__38546));
  nor2s1 ____496879(.DIN1 (_____90__37459), .DIN2 (___0_9___40653), .Q
       (_________38500));
  nnd2s1 ____09_496880(.DIN1 (_________38473), .DIN2 (_____0__25231),
       .Q (_________38499));
  nor2s1 ____09_496881(.DIN1 (_____00__38419), .DIN2 (_________38462),
       .Q (_________38498));
  nnd2s1 _____9_496882(.DIN1 (_________38455), .DIN2 (______9__38496),
       .Q (______0__38497));
  nor2s1 ____09_496883(.DIN1 (______0__37401), .DIN2 (___0_9___40653),
       .Q (_________38495));
  and2s1 ____09_496884(.DIN1 (___9__0__39136), .DIN2 (_________37333),
       .Q (_________38494));
  or2s1 _______496885(.DIN1 (___90____39051), .DIN2 (______0__38458),
       .Q (_________38493));
  and2s1 _____496886(.DIN1 (___9__0__39136), .DIN2 (_____0___37376), .Q
       (_________38492));
  xnr2s1 _____0_496887(.DIN1 (___0_____40308), .DIN2 (______9__38759),
       .Q (_________38491));
  nnd2s1 _______496888(.DIN1 (______9__38457), .DIN2 (_____9___38417),
       .Q (_________38490));
  xor2s1 ____0_496889(.DIN1 (_________38433), .DIN2 (______9__38447),
       .Q (_____0___38523));
  nnd2s1 ____09_496890(.DIN1 (_________38452), .DIN2 (_________38464),
       .Q (_____9___38511));
  nnd2s1 ____09_496891(.DIN1 (_________38446), .DIN2 (_____0___38616),
       .Q (_________38489));
  hi1s1 ____0__496892(.DIN (______0__38487), .Q (_________38488));
  nnd2s1 ____0__496893(.DIN1 (_________38482), .DIN2
       (_____________________________________________21860), .Q
       (______9__38486));
  nnd2s1 ____0__496894(.DIN1 (_________38453), .DIN2
       (____0_____________0___21723), .Q (_________38485));
  xor2s1 ____0__496895(.DIN1 (___9_00__39071), .DIN2 (______0__38467),
       .Q (_________38484));
  nor2s1 ____0_496896(.DIN1
       (_____________________________________________21860), .DIN2
       (_________38482), .Q (_________38483));
  xor2s1 ____0__496897(.DIN1 (_____0___38425), .DIN2 (_________37621),
       .Q (_________38481));
  nor2s1 ____0__496898(.DIN1 (________26397), .DIN2 (_________38449),
       .Q (_________38480));
  dffacs1 _____________________________________________9_496899(.CLRB
       (reset), .CLK (clk), .DIN (_________38445), .Q (___0_____40494));
  nor2s1 _______496900(.DIN1 (_________36843), .DIN2 (______0__38438),
       .Q (_________38479));
  xor2s1 _____0_496901(.DIN1 (_____9___38414), .DIN2
       (__________________________________9__________), .Q
       (_________38478));
  xor2s1 _____0_496902(.DIN1 (_________38444), .DIN2 (______0__36697),
       .Q (______0__38477));
  nor2s1 _______496903(.DIN1 (____9___26860), .DIN2 (_________38436),
       .Q (______9__38476));
  nnd2s1 _______496904(.DIN1 (_________38176), .DIN2 (_________38432),
       .Q (_________38475));
  nor2s1 _______496905(.DIN1 (______9__38390), .DIN2 (_________38434),
       .Q (_________38474));
  nnd2s1 _______496906(.DIN1 (_________38443), .DIN2 (______9__38400),
       .Q (_____0___38520));
  nnd2s1 _______496907(.DIN1 (______9__38759), .DIN2 (_____0___38426),
       .Q (_____00__38517));
  xor2s1 _______496908(.DIN1 (_________38461), .DIN2 (_________37773),
       .Q (______0__38527));
  nnd2s1 _______496909(.DIN1 (_____0___38424), .DIN2 (_____0___38616),
       .Q (_________38473));
  and2s1 ____0__496910(.DIN1 (_________38430), .DIN2 (_________38471),
       .Q (_________38472));
  hi1s1 ____0__496911(.DIN
       (_____________________________________________21860), .Q
       (_________38470));
  nor2s1 ____0__496912(.DIN1 (_________38724), .DIN2 (_________38465),
       .Q (_________38469));
  nor2s1 ____0__496913(.DIN1 (______0__38467), .DIN2 (___9_00__39071),
       .Q (_________38468));
  xor2s1 _____0_496914(.DIN1
       (______________________________________0_______21888), .DIN2
       (_________37822), .Q (______9__38466));
  nnd2s1 _____496915(.DIN1 (___9_00__39071), .DIN2 (______0__38467), .Q
       (_________38501));
  nnd2s1 ____0_496916(.DIN1 (_________38429), .DIN2 (______0__38286),
       .Q (______0__38487));
  nnd2s1 ______496917(.DIN1 (_________38465), .DIN2 (___09_9__40689),
       .Q (_________38684));
  or2s1 _______496918(.DIN1 (_________38463), .DIN2 (_____0___38423),
       .Q (_________38464));
  nor2s1 ______496919(.DIN1 (_________38214), .DIN2 (_________38461),
       .Q (_________38462));
  xor2s1 _______496920(.DIN1 (_________38431), .DIN2 (_________38724),
       .Q (_________38460));
  xor2s1 _______496921(.DIN1
       (______________________________________________21904), .DIN2
       (_________38724), .Q (_________38459));
  xor2s1 _______496922(.DIN1 (_________36865), .DIN2 (______9__38437),
       .Q (______0__38458));
  nnd2s1 _______496923(.DIN1 (_____0___38420), .DIN2 (_________38456),
       .Q (______9__38457));
  nor2s1 _______496924(.DIN1 (________24800), .DIN2 (_____0___38421),
       .Q (_________38455));
  dffacs1 _______________________________________________496925(.CLRB
       (reset), .CLK (clk), .DIN (_____9___38416), .Q (___0_____40438));
  dffacs1 _______________________________________________496926(.CLRB
       (reset), .CLK (clk), .DIN (_____9___38415), .QN
       (_____________________________________________21927));
  xor2s1 ______496927(.DIN1 (____0_0__40750), .DIN2 (_________38724),
       .Q (___9__0__39136));
  nor2s1 ______496928(.DIN1 (_________35453), .DIN2 (_________38407),
       .Q (_________38454));
  nnd2s1 ____0__496929(.DIN1 (_____90__38409), .DIN2 (_________38349),
       .Q (_________38453));
  nnd2s1 ______496930(.DIN1 (_________38403), .DIN2 (_________38463),
       .Q (_________38452));
  nnd2s1 _____0_496931(.DIN1 (_____0___38427), .DIN2 (_________38450),
       .Q (_________38451));
  and2s1 _______496932(.DIN1 (________26557), .DIN2
       (______________________________________0_______21888), .Q
       (_________38449));
  xor2s1 ____0__496933(.DIN1 (______0__38428), .DIN2 (____0____40752),
       .Q (______0__38448));
  nnd2s1 _______496934(.DIN1 (_________38392), .DIN2 (______9__38408),
       .Q (______9__38447));
  xor2s1 _______496935(.DIN1 (_________38384), .DIN2 (________27441),
       .Q (_________38446));
  nnd2s1 _______496936(.DIN1 (_____9___38411), .DIN2 (_________38262),
       .Q (_________38445));
  hi1s1 _______496937(.DIN (_________38444), .Q (_____9___38515));
  dffacs1 _______________________________________________496938(.CLRB
       (reset), .CLK (clk), .DIN (_____9___38410), .Q
       (_____________________________________________21860));
  nnd2s1 _______496939(.DIN1 (_________38398), .DIN2 (_____9___38412),
       .Q (_________38443));
  and2s1 _______496940(.DIN1 (_________38724), .DIN2
       (______________________________________________21904), .Q
       (_________38442));
  nor2s1 _______496941(.DIN1
       (______________________________________________21904), .DIN2
       (_________38724), .Q (_________38441));
  and2s1 _______496942(.DIN1 (_________38724), .DIN2 (_________38439),
       .Q (_________38440));
  and2s1 ______496943(.DIN1 (______9__38437), .DIN2 (_____0___36828),
       .Q (______0__38438));
  nor2s1 ______496944(.DIN1 (_________38435), .DIN2 (_________38399),
       .Q (_________38436));
  and2s1 _____0_496945(.DIN1 (_________38433), .DIN2 (______9__38351),
       .Q (_________38434));
  nnd2s1 _______496946(.DIN1 (________26394), .DIN2 (______0__38401),
       .Q (_________38432));
  nnd2s1 _______496947(.DIN1 (_________38724), .DIN2 (_________38431),
       .Q (_________38690));
  dffacs1 _____________________________________________0_496948(.CLRB
       (reset), .CLK (clk), .DIN (_________38405), .Q
       (__________22063));
  nnd2s1 _______496949(.DIN1 (_________38724), .DIN2 (_________38290),
       .Q (______9__38759));
  dffacs1 __________________________________________0_____496950(.CLRB
       (reset), .CLK (clk), .DIN (_________38404), .QN
       (______________________________________0_______21889));
  dffacs1 ________________496951(.CLRB (reset), .CLK (clk), .DIN
       (___09_9__40689), .Q (outData[21]));
  and2s1 ____0__496952(.DIN1 (____9____37976), .DIN2 (_________38387),
       .Q (_________38430));
  nnd2s1 ____090(.DIN1 (______0__38428), .DIN2 (_________38287), .Q
       (_________38429));
  nnd2s1 _______496953(.DIN1 (___09_9__40689), .DIN2 (_________38298),
       .Q (_____0___38426));
  xor2s1 _______496954(.DIN1 (___0_____40495), .DIN2 (_________38406),
       .Q (_____0___38425));
  nnd2s1 _______496955(.DIN1 (_________38402), .DIN2 (_________38389),
       .Q (_____0___38424));
  nor2s1 ______496956(.DIN1 (________28865), .DIN2 (_________38394), .Q
       (_____0___38423));
  xor2s1 _______496957(.DIN1 (_________38368), .DIN2 (___9_____39582),
       .Q (_________38465));
  xor2s1 _______496958(.DIN1 (_________38367), .DIN2 (_____0___38422),
       .Q (___9_00__39071));
  nor2s1 _______496959(.DIN1 (___0__0__39993), .DIN2 (_________38383),
       .Q (_____0___38421));
  nnd2s1 ______496960(.DIN1 (_________38382), .DIN2 (______9__35527),
       .Q (_____0___38420));
  nor2s1 _______496961(.DIN1 (_________37774), .DIN2 (_____99__38418),
       .Q (_____00__38419));
  or2s1 _____9_496962(.DIN1 (_________38456), .DIN2 (______9__38380),
       .Q (_____9___38417));
  or2s1 ______496963(.DIN1 (___9_____39575), .DIN2 (_________38379), .Q
       (_____9___38416));
  nnd2s1 _______496964(.DIN1 (__9__9__30149), .DIN2 (_________38378),
       .Q (_____9___38415));
  xor2s1 ______496965(.DIN1 (_________38355), .DIN2
       (_____________________________________________21815), .Q
       (_____9___38414));
  or2s1 ______496966(.DIN1 (_________38439), .DIN2 (___09_9__40689), .Q
       (_________38658));
  xor2s1 _______496967(.DIN1 (_____9___38413), .DIN2 (_________37769),
       .Q (_________38461));
  xor2s1 _______496968(.DIN1 (_________38354), .DIN2 (_____9___38412),
       .Q (_________38444));
  nor2s1 _______496969(.DIN1 (_____9___37944), .DIN2 (_________38356),
       .Q (_____9___38411));
  nor2s1 _______496970(.DIN1 (____0____38117), .DIN2 (_________38373),
       .Q (_____9___38410));
  nnd2s1 _______496971(.DIN1 (_________38374), .DIN2 (_________22024),
       .Q (_____90__38409));
  nnd2s1 _______496972(.DIN1 (_________38375), .DIN2 (_____00__35736),
       .Q (______9__38408));
  and2s1 _______496973(.DIN1 (_________38406), .DIN2 (_________35459),
       .Q (_________38407));
  nnd2s1 ______496974(.DIN1 (______9__38370), .DIN2 (_________38253),
       .Q (_________38405));
  nnd2s1 _______496975(.DIN1 (_________38366), .DIN2 (________25437),
       .Q (_________38404));
  dffacs1 __________________________________________0_____496976(.CLRB
       (reset), .CLK (clk), .DIN (______0__38371), .QN
       (______________________________________0_______21888));
  nnd2s1 ______496977(.DIN1 (_________37416), .DIN2 (_________38369),
       .Q (_____0___38427));
  hi1s1 _____9_496978(.DIN (_________38402), .Q (_________38403));
  xor2s1 _______496979(.DIN1 (_________22021), .DIN2 (_____0___37668),
       .Q (______0__38401));
  or2s1 _____9_496980(.DIN1 (_____9___38412), .DIN2 (______9__38361),
       .Q (______9__38400));
  xor2s1 _____496981(.DIN1 (_________35638), .DIN2 (______0__38381), .Q
       (_________38399));
  nnd2s1 _____496982(.DIN1 (_________38365), .DIN2 (___09___22356), .Q
       (_________38398));
  nor2s1 _____496983(.DIN1 (_________38396), .DIN2 (_________38363), .Q
       (_________38397));
  xor2s1 _______496984(.DIN1 (_________38346), .DIN2 (_________38395),
       .Q (_________38433));
  nor2s1 _______496985(.DIN1 (_________36839), .DIN2 (_________38353),
       .Q (______9__38437));
  hi1s1 _____9_496986(.DIN (___09_9__40689), .Q (_________38724));
  nor2s1 _______496987(.DIN1 (________28864), .DIN2 (_________38388),
       .Q (_________38394));
  nnd2s1 _______496988(.DIN1 (______0__38391), .DIN2 (_____00__35736),
       .Q (_________38393));
  nnd2s1 _______496989(.DIN1 (______0__38391), .DIN2
       (___________________), .Q (_________38392));
  nor2s1 _______496990(.DIN1 (_____00__35736), .DIN2 (______0__38391),
       .Q (______9__38390));
  or2s1 _____9_496991(.DIN1 (_________38376), .DIN2 (_________38388),
       .Q (_________38389));
  nnd2s1 _______496992(.DIN1 (___90____38993), .DIN2 (_________38347),
       .Q (_________38387));
  xor2s1 _____0_496993(.DIN1 (_________38386), .DIN2 (____0____38089),
       .Q (_________38776));
  nnd2s1 ______496994(.DIN1 (_________37432), .DIN2
       (_______________________________________________________________0__22006),
       .Q (_________38450));
  xor2s1 _______496995(.DIN1 (_________38340), .DIN2 (_________38385),
       .Q (______0__38428));
  xor2s1 _____0_496996(.DIN1 (_________38335), .DIN2 (___0_0___40465),
       .Q (_________38384));
  xor2s1 _____0_496997(.DIN1 (_________36840), .DIN2 (______0__38352),
       .Q (_________38383));
  or2s1 _______496998(.DIN1 (_____09__35574), .DIN2 (______0__38381),
       .Q (_________38382));
  nnd2s1 ______496999(.DIN1 (______0__38381), .DIN2 (_________35637),
       .Q (______9__38380));
  nnd2s1 _______497000(.DIN1 (_________38344), .DIN2 (____9___24837),
       .Q (_________38379));
  or2s1 _______497001(.DIN1 (_________22021), .DIN2 (_________38377),
       .Q (_________38378));
  hi1s1 ______497002(.DIN (_____9___38413), .Q (_____99__38418));
  nnd2s1 _____0_497003(.DIN1 (_________38388), .DIN2 (_________38376),
       .Q (_________38402));
  dffacs1 _______________________________________________497004(.CLRB
       (reset), .CLK (clk), .DIN (_________38345), .Q (___0_____40534));
  xor2s1 _____0_497005(.DIN1 (___90____39019), .DIN2 (_________38350),
       .Q (_________38375));
  hi1s1 _______497006(.DIN (_________38471), .Q (_________38374));
  xor2s1 _______497007(.DIN1 (_____0___38326), .DIN2 (_________38372),
       .Q (_________38373));
  nnd2s1 _______497008(.DIN1 (______0__38343), .DIN2 (_________37875),
       .Q (______0__38371));
  nor2s1 _______497009(.DIN1 (____00__25310), .DIN2 (_________38338),
       .Q (______9__38370));
  hi1s1 ______497010(.DIN
       (_______________________________________________________________0__22006),
       .Q (_________38369));
  nnd2s1 _____0_497011(.DIN1 (_________38341), .DIN2 (_____0___38331),
       .Q (_________38368));
  xor2s1 _____0_497012(.DIN1 (_____0___38328), .DIN2 (_________38311),
       .Q (_________38367));
  nnd2s1 _______497013(.DIN1 (_____0___38332), .DIN2 (_________37744),
       .Q (_________38366));
  nor2s1 _____497014(.DIN1 (_________38292), .DIN2 (______9__38342), .Q
       (_________38406));
  or2s1 _______497015(.DIN1 (____0___22367), .DIN2 (_________38364), .Q
       (_________38365));
  hi1s1 _______497016(.DIN (______0__38362), .Q (_________38363));
  nnd2s1 _______497017(.DIN1 (_________38364), .DIN2 (________22601),
       .Q (______9__38361));
  nnd2s1 _______497018(.DIN1 (_________38359), .DIN2 (_________38358),
       .Q (_________38360));
  nor2s1 _______497019(.DIN1 (_________38358), .DIN2 (_________38359),
       .Q (_________38357));
  nor2s1 _______497020(.DIN1 (_________38164), .DIN2 (_________38336),
       .Q (_________38356));
  xor2s1 _______497021(.DIN1 (_____9___38316), .DIN2 (_________38533),
       .Q (_________38355));
  nnd2s1 _______497022(.DIN1 (_________38386), .DIN2 (____0____38088),
       .Q (_________38354));
  dffacs1 ______________0_497023(.CLRB (reset), .CLK (clk), .DIN
       (_________38339), .Q (outData[20]));
  nor2s1 _______497024(.DIN1 (_________36838), .DIN2 (______0__38352),
       .Q (_________38353));
  xor2s1 _______497025(.DIN1 (_________38272), .DIN2 (_____9___38321),
       .Q (_____9___38413));
  or2s1 _______497026(.DIN1 (_________38350), .DIN2 (___90____39019),
       .Q (______9__38351));
  or2s1 _______497027(.DIN1 (_________22024), .DIN2 (_________38348),
       .Q (_________38349));
  nnd2s1 ______497028(.DIN1 (_____0___38329), .DIN2 (inData[4]), .Q
       (_________38347));
  xor2s1 ______497029(.DIN1 (______0__38295), .DIN2 (_________38242),
       .Q (______0__38362));
  dffacs1 _______________________________________________497030(.CLRB
       (reset), .CLK (clk), .DIN (_____0___38327), .QN
       (_______________________________________________________________0__22006));
  nnd2s1 _______497031(.DIN1 (___90____38993), .DIN2 (_________38348),
       .Q (_________38471));
  nor2s1 _______497032(.DIN1 (______0__38334), .DIN2 (_____00__38325),
       .Q (_________38388));
  nor2s1 _____9_497033(.DIN1 (_________38184), .DIN2 (_________38313),
       .Q (_________38346));
  or2s1 _______497034(.DIN1 (______9__38245), .DIN2 (______9__38314),
       .Q (_________38345));
  nnd2s1 _______497035(.DIN1 (_____90__38315), .DIN2 (________23899),
       .Q (_________38344));
  dffacs1 _______________________________________________497036(.CLRB
       (reset), .CLK (clk), .DIN (_________38312), .Q (_________22021));
  nor2s1 ______497037(.DIN1 (_________35529), .DIN2 (_____9___38318),
       .Q (______0__38381));
  and2s1 _______497038(.DIN1 (___90____39019), .DIN2 (_________38350),
       .Q (______0__38391));
  dffacs1 _______________________________________________497039(.CLRB
       (reset), .CLK (clk), .DIN (_____9___38320), .Q (___0_____40495));
  nnd2s1 ______497040(.DIN1 (_________38307), .DIN2 (___90____39040),
       .Q (______0__38343));
  nnd2s1 ______497041(.DIN1 (______9__38285), .DIN2 (_________38309),
       .Q (______9__38342));
  xor2s1 _______497042(.DIN1 (_________38291), .DIN2 (____9____38948),
       .Q (_________38341));
  xor2s1 _____0_497043(.DIN1 (_________38288), .DIN2 (____9____37970),
       .Q (_________38340));
  nnd2s1 _______497044(.DIN1 (_________38310), .DIN2 (________23353),
       .Q (_________38339));
  nor2s1 _______497045(.DIN1 (_____9__26765), .DIN2 (_________38303),
       .Q (_________38338));
  xor2s1 _______497046(.DIN1 (_________35531), .DIN2 (_____9___38317),
       .Q (_________38336));
  nor2s1 ______497047(.DIN1 (______0__38334), .DIN2 (______0__38305),
       .Q (_________38335));
  nor2s1 ______497048(.DIN1 (_________38296), .DIN2 (_________38431),
       .Q (_____0___38332));
  nor2s1 ______497049(.DIN1 (_________36470), .DIN2 (______9__38294),
       .Q (______0__38352));
  nor2s1 _______497050(.DIN1 (_________38270), .DIN2 (_________38302),
       .Q (_________38364));
  and2s1 _______497051(.DIN1 (_________38830), .DIN2 (_________38297),
       .Q (_________38359));
  nor2s1 _______497052(.DIN1 (_____0___38331), .DIN2 (_________38299),
       .Q (_________38439));
  hi1s1 _______497053(.DIN (_____0___38330), .Q (_________38386));
  nnd2s1 _______497054(.DIN1
       (_____________________________________________21942), .DIN2
       (___0__9__40430), .Q (_____0___38329));
  xor2s1 _______497055(.DIN1 (_________38264), .DIN2 (______9__37429),
       .Q (_____0___38328));
  or2s1 _____9_497056(.DIN1
       (_____________________________________________21942), .DIN2
       (___0__0__39993), .Q (_____0___38327));
  xor2s1 ______497057(.DIN1 (_________38308), .DIN2 (_________38284),
       .Q (_____0___38326));
  and2s1 _______497058(.DIN1 (______9__38304), .DIN2 (___0_0___40465),
       .Q (_____00__38325));
  nnd2s1 _______497059(.DIN1 (_____9___38323), .DIN2 (_____9___38322),
       .Q (_____99__38324));
  nnd2s1 _______497060(.DIN1 (_________38283), .DIN2 (______0__38141),
       .Q (_____0___38333));
  nor2s1 _____9_497061(.DIN1 (___0__9__40430), .DIN2
       (_____________________________________________21942), .Q
       (_________38348));
  dffacs1 _________________________________________9_____497062(.CLRB
       (reset), .CLK (clk), .DIN (_________38289), .QN
       (___0_____40621));
  nnd2s1 _____9_497063(.DIN1 (_________38278), .DIN2 (_____9___38224),
       .Q (_____9___38321));
  nnd2s1 _______497064(.DIN1 (______9__38275), .DIN2 (_____9___38319),
       .Q (_____9___38320));
  nor2s1 _______497065(.DIN1 (_________35530), .DIN2 (_____9___38317),
       .Q (_____9___38318));
  nor2s1 _____9_497066(.DIN1 (_________36590), .DIN2 (_________38277),
       .Q (_____9___38316));
  xor2s1 _______497067(.DIN1 (______9__36472), .DIN2 (_________38293),
       .Q (_____90__38315));
  nnd2s1 _______497068(.DIN1 (_________38274), .DIN2 (_____0__25711),
       .Q (______9__38314));
  nnd2s1 _______497069(.DIN1 (_________38273), .DIN2 (_________38183),
       .Q (_________38313));
  nnd2s1 _______497070(.DIN1 (_________38279), .DIN2 (_____9___37757),
       .Q (_________38312));
  xor2s1 _______497071(.DIN1 (_________38311), .DIN2 (___9_0___39166),
       .Q (_____0___38330));
  xor2s1 _______497072(.DIN1 (______9__38265), .DIN2 (________23513),
       .Q (___90____39019));
  nnd2s1 ______497073(.DIN1 (_________38311), .DIN2 (____9____38949),
       .Q (_________38310));
  or2s1 _______497074(.DIN1 (______0__38256), .DIN2 (_________38308),
       .Q (_________38309));
  xor2s1 _______497075(.DIN1 (_________38259), .DIN2 (_________38306),
       .Q (_________38307));
  hi1s1 ______497076(.DIN (______9__38304), .Q (______0__38305));
  xor2s1 _____497077(.DIN1 (_________36600), .DIN2 (______0__38276), .Q
       (_________38303));
  nor2s1 _____9_497078(.DIN1 (_________38301), .DIN2 (_________38269),
       .Q (_________38302));
  nor2s1 _____497079(.DIN1 (_____9___38219), .DIN2 (_________38311), .Q
       (_________38300));
  xor2s1 _______497080(.DIN1 (_____0___38230), .DIN2 (_________38282),
       .Q (_________38563));
  nor2s1 _____0_497081(.DIN1 (_____99__38226), .DIN2 (_________38298),
       .Q (_________38299));
  nnd2s1 _____0_497082(.DIN1 (_________38298), .DIN2 (______0__37643),
       .Q (_________38297));
  nor2s1 _____0_497083(.DIN1 (_____0___38232), .DIN2 (_____0___38331),
       .Q (_________38296));
  nnd2s1 _______497084(.DIN1 (_________38311), .DIN2
       (__________________________________________________________________21990),
       .Q (______0__38295));
  nor2s1 _______497085(.DIN1 (_________36471), .DIN2 (_________38293),
       .Q (______9__38294));
  nnd2s1 _____0_497086(.DIN1 (_________38213), .DIN2 (_________38311),
       .Q (_________38337));
  nor2s1 ______497087(.DIN1
       (__________________________________________________________________21990),
       .DIN2 (_________38311), .Q (_________38396));
  nor2s1 _______497088(.DIN1 (_____0___38233), .DIN2 (_________38311),
       .Q (_________38431));
  nor2s1 ______497089(.DIN1 (_________38257), .DIN2 (_________38267),
       .Q (_________38292));
  nor2s1 _____497090(.DIN1 (_____90__38218), .DIN2 (_________38290), .Q
       (_________38291));
  nnd2s1 _______497091(.DIN1 (_________38258), .DIN2 (_________40998),
       .Q (_________38289));
  xor2s1 _______497092(.DIN1 (______0__38237), .DIN2 (____9_0__37985),
       .Q (_________38288));
  nnd2s1 _______497093(.DIN1 (____0____40752), .DIN2
       (_____________________________________________21928), .Q
       (_________38287));
  or2s1 _______497094(.DIN1
       (_____________________________________________21928), .DIN2
       (____0____40752), .Q (______0__38286));
  nnd2s1 _____0_497095(.DIN1 (_________38284), .DIN2 (______9__38255),
       .Q (______9__38285));
  or2s1 _____0_497096(.DIN1 (_____0___38136), .DIN2 (_________38282),
       .Q (_________38283));
  nor2s1 _____9_497097(.DIN1
       (__________________________________9__________), .DIN2
       (_________38281), .Q (______0__38334));
  nnd2s1 _____9_497098(.DIN1 (_________38281), .DIN2 (_________38280),
       .Q (______9__38304));
  nnd2s1 _____0_497099(.DIN1 (_________38290), .DIN2
       (________________________________________________________________),
       .Q (_____9___38323));
  dffacs1 _______________________________________________497100(.CLRB
       (reset), .CLK (clk), .DIN (_________38260), .QN
       (_____________________________________________21942));
  or2s1 _____0_497101(.DIN1 (___90____39051), .DIN2 (_________38252),
       .Q (_________38279));
  nnd2s1 ______497102(.DIN1 (_________38251), .DIN2 (____9_9__38931),
       .Q (_________38278));
  nor2s1 _______497103(.DIN1 (______9__36588), .DIN2 (______0__38276),
       .Q (_________38277));
  nor2s1 _______497104(.DIN1 (________23467), .DIN2 (_________38250),
       .Q (______9__38275));
  nnd2s1 ______497105(.DIN1 (_________38247), .DIN2 (_________38177),
       .Q (_________38274));
  or2s1 _______497106(.DIN1 (_________38244), .DIN2 (_________38272),
       .Q (_________38273));
  xor2s1 _______497107(.DIN1 (_____9___38225), .DIN2 (_________38271),
       .Q (_____9___38322));
  nor2s1 ______497108(.DIN1 (_________38202), .DIN2 (_________38261),
       .Q (_____9___38317));
  dffacs1 _____________________________________________0_497109(.CLRB
       (reset), .CLK (clk), .DIN (______0__38246), .Q (___0_____40535));
  nnd2s1 _______497110(.DIN1 (_________38290), .DIN2 (_________37681),
       .Q (_________38830));
  dffacs1 _______________________________________________497111(.CLRB
       (reset), .CLK (clk), .DIN (_________38263), .QN
       (___0_____40505));
  dffacs1 ______________________________________________(.CLRB (reset),
       .CLK (clk), .DIN (_________38248), .QN
       (____________________________________________21847));
  dffacs1 _______________________________________________497112(.CLRB
       (reset), .CLK (clk), .DIN (_________38254), .QN
       (___0_____40536));
  nor2s1 _______497113(.DIN1 (_________35677), .DIN2 (_________38241),
       .Q (_________38270));
  nor2s1 _______497114(.DIN1 (___0_0), .DIN2 (_____0___38235), .Q
       (_________38269));
  nnd2s1 _______497115(.DIN1 (_________38238), .DIN2 (_____0___38616),
       .Q (_________38268));
  xor2s1 _______497116(.DIN1
       (_____________________________________________21844), .DIN2
       (_________38267), .Q (_________38308));
  hi1s1 _______497117(.DIN (______0__38266), .Q (_____0___38331));
  hi1s1 _______497118(.DIN (_________38290), .Q (_________38298));
  nb1s1 _______497119(.DIN (______0__38266), .Q (_________38311));
  xor2s1 _______497120(.DIN1 (______9__38198), .DIN2 (_________38193),
       .Q (______9__38265));
  nnd2s1 _______497121(.DIN1 (_____00__38227), .DIN2 (_________38210),
       .Q (_________38264));
  nor2s1 _______497122(.DIN1 (______9__36308), .DIN2 (_____0___38229),
       .Q (_________38293));
  dffacs1 ______________________________________________497123(.CLRB
       (reset), .CLK (clk), .DIN (_____9___38220), .QN
       (___0_____40548));
  dffacs1 ______________________________________________497124(.CLRB
       (reset), .CLK (clk), .DIN (_____9___38222), .Q
       (____________________________________________21789));
  dffacs1 ______________________________________________497125(.CLRB
       (reset), .CLK (clk), .DIN (_____9___38221), .QN
       (____________________________________________21864));
  dffacs1 _______________________________________________497126(.CLRB
       (reset), .CLK (clk), .DIN (_____0___38234), .QN
       (___0_____40517));
  dffacs1 _______________________________________________497127(.CLRB
       (reset), .CLK (clk), .DIN (_____9___38223), .QN
       (___0_0___40464));
  nnd2s1 _______497128(.DIN1 (______9__38217), .DIN2 (_________38262),
       .Q (_________38263));
  nor2s1 _______497129(.DIN1 (_________38200), .DIN2 (______0__38199),
       .Q (_________38261));
  or2s1 _______497130(.DIN1 (________23836), .DIN2 (_________38216), .Q
       (_________38260));
  xor2s1 _______497131(.DIN1 (_________38193), .DIN2 (_________38206),
       .Q (_________38259));
  nnd2s1 _______497132(.DIN1 (_________38215), .DIN2 (_________41345),
       .Q (_________38258));
  nnd2s1 _______497133(.DIN1 (______0__38256), .DIN2
       (_____________________________________________21844), .Q
       (_________38257));
  or2s1 ______497134(.DIN1
       (_____________________________________________21844), .DIN2
       (_________35404), .Q (______9__38255));
  nor2s1 _______497135(.DIN1 (____9____37986), .DIN2 (______9__38208),
       .Q (_________38282));
  nor2s1 _______497136(.DIN1 (______9__37909), .DIN2 (_________38212),
       .Q (_________38281));
  dffacs1 _______________________________________________497137(.CLRB
       (reset), .CLK (clk), .DIN (_________38195), .QN
       (___0_____40497));
  nnd2s1 ______497138(.DIN1 (_________38196), .DIN2 (_________38253),
       .Q (_________38254));
  xor2s1 _______497139(.DIN1 (_____0___38228), .DIN2 (_____9___36364),
       .Q (_________38252));
  nnd2s1 _______497140(.DIN1 (_________38243), .DIN2 (_________38204),
       .Q (_________38251));
  and2s1 _______497141(.DIN1 (_________38205), .DIN2 (_________38249),
       .Q (_________38250));
  nnd2s1 _______497142(.DIN1 (____9____34342), .DIN2 (_________38197),
       .Q (_________38248));
  xor2s1 _______497143(.DIN1 (_________38192), .DIN2 (________28894),
       .Q (_________38247));
  or2s1 _____497144(.DIN1 (______9__38245), .DIN2 (_________38194), .Q
       (______0__38246));
  and2s1 _____497145(.DIN1 (_________38243), .DIN2 (_________38186), .Q
       (_________38244));
  xor2s1 _______497146(.DIN1 (_________38180), .DIN2 (___9__9__39569),
       .Q (______0__38276));
  xor2s1 ______497147(.DIN1 (_________38239), .DIN2 (_________38240),
       .Q (______0__38266));
  xor2s1 _______497148(.DIN1 (_________38193), .DIN2 (_________38242),
       .Q (_________38290));
  nnd2s1 ______497149(.DIN1 (_________38240), .DIN2 (_________38239),
       .Q (_________38241));
  xor2s1 _______497150(.DIN1 (______0__37910), .DIN2 (_________38211),
       .Q (_________38238));
  xor2s1 _______497151(.DIN1 (_________38207), .DIN2 (____9_0__38941),
       .Q (______0__38237));
  nor2s1 _______497152(.DIN1 (_________38435), .DIN2 (______9__38188),
       .Q (_____09__38236));
  nor2s1 _______497153(.DIN1 (___0_0__22344), .DIN2 (_________38240),
       .Q (_____0___38235));
  nnd2s1 _______497154(.DIN1 (______0__38189), .DIN2 (_____9___38319),
       .Q (_____0___38234));
  hi1s1 _______497155(.DIN (_____0___38232), .Q (_____0___38233));
  nnd2s1 ______497156(.DIN1 (_____9___41369), .DIN2 (____9____34341),
       .Q (_____0___38231));
  xor2s1 _______497157(.DIN1 (_________38166), .DIN2 (___9__9__39125),
       .Q (_____0___38230));
  and2s1 _______497158(.DIN1 (_____0___38228), .DIN2 (_________36310),
       .Q (_____0___38229));
  nnd2s1 _______497159(.DIN1 (_____99__38226), .DIN2 (_____9___41369),
       .Q (_____00__38227));
  or2s1 _______497160(.DIN1
       (________________________________________________________________),
       .DIN2 (_____9___41369), .Q (_____9___38225));
  nnd2s1 _______497161(.DIN1 (_________38181), .DIN2 (_________38203),
       .Q (_____9___38224));
  nnd2s1 _______497162(.DIN1 (_________38185), .DIN2 (_________37722),
       .Q (_____9___38223));
  nnd2s1 ______497163(.DIN1 (_________33317), .DIN2 (______0__38179),
       .Q (_____9___38222));
  or2s1 _______497164(.DIN1 (_________38174), .DIN2 (_________38187),
       .Q (_____9___38221));
  nnd2s1 _______497165(.DIN1 (_________38191), .DIN2 (_________38172),
       .Q (_____9___38220));
  or2s1 _______497166(.DIN1 (_____90__38218), .DIN2 (_____9___41369),
       .Q (_____9___38219));
  nor2s1 _______497167(.DIN1 (____09__23701), .DIN2 (_________38165),
       .Q (______9__38217));
  nor2s1 _____497168(.DIN1 (___90____38993), .DIN2 (_________38167), .Q
       (_________38216));
  xor2s1 _______497169(.DIN1 (_____0___38133), .DIN2 (_________38214),
       .Q (_________38215));
  nor2s1 _______497170(.DIN1 (______0__38209), .DIN2 (_____99__38226),
       .Q (_________38213));
  nor2s1 _______497171(.DIN1 (_________37908), .DIN2 (_________38211),
       .Q (_________38212));
  nnd2s1 _______497172(.DIN1 (______0__38209), .DIN2 (_____90__38218),
       .Q (_________38210));
  nor2s1 _______497173(.DIN1 (____00___38040), .DIN2 (_________38207),
       .Q (______9__38208));
  nor2s1 ______497174(.DIN1 (_________38206), .DIN2 (______0__38209),
       .Q (_____0___38232));
  dffacs1 _______________________________________________497175(.CLRB
       (reset), .CLK (clk), .DIN (_________38171), .QN
       (_____________________________________________21844));
  dffacs1 ______________________________________________497176(.CLRB
       (reset), .CLK (clk), .DIN (_________38173), .QN
       (___0_____40532));
  or2s1 ______497177(.DIN1 (_________38158), .DIN2 (_________38201), .Q
       (_________38205));
  nnd2s1 _______497178(.DIN1 (_________38156), .DIN2 (_________38203),
       .Q (_________38204));
  and2s1 _______497179(.DIN1 (_________38201), .DIN2 (_________38200),
       .Q (_________38202));
  nor2s1 _____9_497180(.DIN1 (____0____35358), .DIN2 (______9__38160),
       .Q (______0__38199));
  nnd2s1 _____9_497181(.DIN1 (____99___38029), .DIN2 (_________38159),
       .Q (______9__38198));
  nnd2s1 _______497182(.DIN1 (_________38175), .DIN2 (inData[6]), .Q
       (_________38197));
  nor2s1 _______497183(.DIN1 (_____0___38138), .DIN2 (_________38162),
       .Q (_________38196));
  nnd2s1 _______497184(.DIN1 (_________38163), .DIN2 (____0____38108),
       .Q (_________38195));
  nnd2s1 _______497185(.DIN1 (_________38178), .DIN2 (_____0__25614),
       .Q (_________38194));
  nnd2s1 _______497186(.DIN1 (______0__38170), .DIN2 (____0____36245),
       .Q (_________38243));
  xnr2s1 _______497187(.DIN1 (______0__41339), .DIN2 (_____0___38137),
       .Q (_____09__38526));
  xor2s1 _______497188(.DIN1 (_________________0_), .DIN2
       (____0_9__38121), .Q (_________38192));
  nor2s1 _______497189(.DIN1 (_________38143), .DIN2 (_________33657),
       .Q (_________38191));
  nnd2s1 _____9_497190(.DIN1 (_____0___38134), .DIN2 (inData[16]), .Q
       (_________38190));
  nor2s1 _______497191(.DIN1 (_____0___38132), .DIN2 (_________37438),
       .Q (______0__38189));
  nnd2s1 _______497192(.DIN1 (_________38146), .DIN2 (____0____38048),
       .Q (_____0___38228));
  hi1s1 _____497193(.DIN (______0__38209), .Q (_________38193));
  dffacs1 _______________________________________________497194(.CLRB
       (reset), .CLK (clk), .DIN (_____0___38139), .Q (___0__0__40599));
  hi1s1 _____497195(.DIN (______0__38209), .Q (_____9___41369));
  xor2s1 _____0_497196(.DIN1 (____099__38130), .DIN2 (______0__38151),
       .Q (______9__38188));
  nnd2s1 ______497197(.DIN1 (____09___38127), .DIN2 (_________38144),
       .Q (_________38187));
  nnd2s1 ______497198(.DIN1 (______9__38169), .DIN2 (_________38203),
       .Q (_________38186));
  nor2s1 _______497199(.DIN1 (________24057), .DIN2 (_________38153),
       .Q (_________38185));
  nor2s1 ______497200(.DIN1 (____9_9__38931), .DIN2 (_________38182),
       .Q (_________38184));
  nnd2s1 _______497201(.DIN1 (_________38182), .DIN2 (____9_9__38931),
       .Q (_________38183));
  and2s1 _______497202(.DIN1 (_________38182), .DIN2 (_________32987),
       .Q (_________38181));
  nnd2s1 ______497203(.DIN1 (_________38152), .DIN2 (____0____38100),
       .Q (_________38180));
  nnd2s1 _______497204(.DIN1 (_________38145), .DIN2 (inData[14]), .Q
       (______0__38179));
  xor2s1 _______497205(.DIN1 (____09___38129), .DIN2 (___9_____39554),
       .Q (_________38240));
  nnd2s1 _______497206(.DIN1 (____0____38120), .DIN2 (_________38177),
       .Q (_________38178));
  or2s1 _____9_497207(.DIN1 (___90____39051), .DIN2 (____090__38122),
       .Q (_________38176));
  or2s1 _____0_497208(.DIN1 (____09___38124), .DIN2 (_________38174),
       .Q (_________38175));
  nnd2s1 _____0_497209(.DIN1 (____09___38123), .DIN2 (_________38172),
       .Q (_________38173));
  nor2s1 _____0_497210(.DIN1 (_________38583), .DIN2 (____0____38116),
       .Q (_________38171));
  hi1s1 _______497211(.DIN (______9__38169), .Q (______0__38170));
  xor2s1 ______497212(.DIN1 (____0____38092), .DIN2 (____0____38114),
       .Q (_________38167));
  xor2s1 ______497213(.DIN1 (_____9___37846), .DIN2 (_____09__38140),
       .Q (_________38166));
  dffacs1 _______________________________________________497214(.CLRB
       (reset), .CLK (clk), .DIN (____0____38118), .Q (___0_____40496));
  dffacs1 ____________________________________9_(.CLRB (reset), .CLK
       (clk), .DIN (____09___38128), .QN (___0_____40586));
  nor2s1 _____0_497215(.DIN1 (_________38164), .DIN2 (____0____38115),
       .Q (_________38165));
  and2s1 _______497216(.DIN1 (____09___38126), .DIN2 (____0_9__38083),
       .Q (_________38163));
  nnd2s1 _______497217(.DIN1 (_________37260), .DIN2 (____09___38125),
       .Q (_________38162));
  xor2s1 _______497218(.DIN1 (_________38149), .DIN2 (___9_____39627),
       .Q (______0__38161));
  nor2s1 _______497219(.DIN1 (_____0___35380), .DIN2 (_________38157),
       .Q (______9__38160));
  nor2s1 ______497220(.DIN1 (____9____38027), .DIN2 (_____00__38131),
       .Q (_________38159));
  nor2s1 _______497221(.DIN1 (_________38154), .DIN2 (_________38157),
       .Q (_________38158));
  xor2s1 _______497222(.DIN1 (____90___38892), .DIN2 (_________38142),
       .Q (_________38156));
  xor2s1 _______497223(.DIN1 (____0____38097), .DIN2 (_________38155),
       .Q (_________38211));
  and2s1 _______497224(.DIN1 (_________38157), .DIN2 (_________38154),
       .Q (_________38201));
  xor2s1 ______497225(.DIN1 (____0____40756), .DIN2 (____9____38909),
       .Q (_________38529));
  xor2s1 _______497226(.DIN1 (____0____40754), .DIN2 (_____99__37662),
       .Q (_________38207));
  xnr2s1 _______497227(.DIN1 (__________9___22107), .DIN2
       (____0_9__38111), .Q (______0__38209));
  nor2s1 _______497228(.DIN1 (_____9___37656), .DIN2 (____0____38103),
       .Q (_________38153));
  nnd2s1 _______497229(.DIN1 (______0__38151), .DIN2 (____0_0__38102),
       .Q (_________38152));
  nnd2s1 ______497230(.DIN1 (_________38147), .DIN2 (_________38149),
       .Q (______9__38150));
  or2s1 ______497231(.DIN1 (_________38149), .DIN2 (_________38147), .Q
       (_________38148));
  xor2s1 _______497232(.DIN1 (____0____38070), .DIN2 (___0_____40308),
       .Q (_________38146));
  nor2s1 _______497233(.DIN1 (____0____38095), .DIN2 (____9____34370),
       .Q (_________38145));
  or2s1 _____9_497234(.DIN1
       (____________________________________________21864), .DIN2
       (____0____40758), .Q (_________38144));
  nor2s1 _______497235(.DIN1 (____0____38096), .DIN2 (____0_9__38073),
       .Q (_________38143));
  nnd2s1 _______497236(.DIN1 (____90___38892), .DIN2 (_________38142),
       .Q (______9__38169));
  nor2s1 ______497237(.DIN1 (_________38142), .DIN2 (____90___38892),
       .Q (_________38182));
  nnd2s1 _____0_497238(.DIN1 (_____09__38140), .DIN2 (_____0___38135),
       .Q (______0__38141));
  nnd2s1 _______497239(.DIN1 (____0____38098), .DIN2 (________25250),
       .Q (_____0___38139));
  nor2s1 _______497240(.DIN1 (____0____38110), .DIN2 (______0__37872),
       .Q (_____0___38138));
  nnd2s1 _______497241(.DIN1 (____0____38107), .DIN2 (____0_0__40760),
       .Q (_____0___38137));
  nor2s1 _____0_497242(.DIN1 (_____0___38135), .DIN2 (_____09__38140),
       .Q (_____0___38136));
  nor2s1 _______497243(.DIN1 (________23372), .DIN2 (____0_0__38112),
       .Q (_____0___38134));
  xor2s1 _______497244(.DIN1 (____0____38080), .DIN2
       (_____________________________________________21872), .Q
       (_____0___38133));
  nor2s1 _______497245(.DIN1 (____0____38094), .DIN2 (_________38249),
       .Q (_____0___38132));
  dffacs1 _______________________________________________497246(.CLRB
       (reset), .CLK (clk), .DIN (____0____38113), .Q
       (_____________________________________________21815));
  dffacs1 _________________________________________9_____497247(.CLRB
       (reset), .CLK (clk), .DIN (____0____38105), .Q (___0_9___40457));
  dffacs1 _______________________________________________497248(.CLRB
       (reset), .CLK (clk), .DIN (____0____38109), .QN
       (___0_____40519));
  nor2s1 _______497249(.DIN1 (_________37597), .DIN2 (____0____38085),
       .Q (_____00__38131));
  xor2s1 _______497250(.DIN1 (____0_9__38101), .DIN2 (__________22062),
       .Q (____099__38130));
  nor2s1 _______497251(.DIN1 (__9_), .DIN2 (____0____38087), .Q
       (____09___38129));
  nnd2s1 _____0_497252(.DIN1 (____0____38075), .DIN2 (____0____38104),
       .Q (____09___38128));
  nor2s1 _____0_497253(.DIN1 (____0____38078), .DIN2 (______9__33102),
       .Q (____09___38127));
  nor2s1 _____497254(.DIN1 (____0____38076), .DIN2 (_________37934), .Q
       (____09___38126));
  nnd2s1 _____9_497255(.DIN1 (____0____37139), .DIN2 (____0____38077),
       .Q (____09___38125));
  xor2s1 _____9_497256(.DIN1 (____0____38090), .DIN2 (_____9___38611),
       .Q (_________38358));
  xor2s1 _____497257(.DIN1 (____00___38043), .DIN2 (_________36871), .Q
       (_____99__38226));
  nnd2s1 _______497258(.DIN1 (____0____38082), .DIN2 (____9____38025),
       .Q (_________38157));
  hi1s1 _______497259(.DIN (____0____40758), .Q (____09___38124));
  nor2s1 _______497260(.DIN1 (____0_0__38074), .DIN2 (______9__33706),
       .Q (____09___38123));
  xor2s1 _______497261(.DIN1 (____0____38049), .DIN2 (____0____38069),
       .Q (____090__38122));
  nor2s1 _______497262(.DIN1 (____0____38051), .DIN2 (____0____38072),
       .Q (____0_9__38121));
  xor2s1 _______497263(.DIN1 (____00___38046), .DIN2 (____0____38071),
       .Q (____0____38120));
  nnd2s1 _______497264(.DIN1 (____0____38081), .DIN2 (___90____39040),
       .Q (____0____38119));
  or2s1 _____0_497265(.DIN1 (____0____38117), .DIN2 (____0____38065),
       .Q (____0____38118));
  xor2s1 ______497266(.DIN1 (___09____40667), .DIN2
       (_____________________________________________21827), .Q
       (____0____38116));
  xor2s1 _______497267(.DIN1 (____0____38057), .DIN2 (_________35084),
       .Q (____0____38115));
  nor2s1 ______497268(.DIN1 (____0____38066), .DIN2 (____0____38114),
       .Q (_________38168));
  dffacs1 ______________________________________497269(.CLRB (reset),
       .CLK (clk), .DIN (____0_9__38063), .QN (_____________22083));
  nnd2s1 _____0_497270(.DIN1 (____0____38061), .DIN2 (____9_0__38009),
       .Q (____0____38113));
  xnr2s1 _______497271(.DIN1 (____99___38030), .DIN2 (___0_____40517),
       .Q (____0_0__38112));
  xor2s1 _______497272(.DIN1 (___0_____40586), .DIN2 (____0____38086),
       .Q (____0_9__38111));
  nnd2s1 _____9_497273(.DIN1 (________25354), .DIN2 (__________22062),
       .Q (____0____38110));
  nnd2s1 _____9_497274(.DIN1 (____0____38054), .DIN2 (____0____38108),
       .Q (____0____38109));
  nnd2s1 _______497275(.DIN1 (____0_0__38056), .DIN2 (____0____38106),
       .Q (____0____38107));
  nnd2s1 _____0_497276(.DIN1 (____0_9__38055), .DIN2 (____0____38104),
       .Q (____0____38105));
  xor2s1 ______497277(.DIN1 (____9____38020), .DIN2 (____0____38053),
       .Q (____0____38103));
  nnd2s1 _______497278(.DIN1 (____0_9__38101), .DIN2 (__________22062),
       .Q (____0_0__38102));
  or2s1 _______497279(.DIN1 (__________22062), .DIN2 (____0_9__38101),
       .Q (____0____38100));
  hi1s1 _______497280(.DIN (____0____38099), .Q (____90___38892));
  nnd2s1 _______497281(.DIN1 (____0____38050), .DIN2 (___9__9__39659),
       .Q (____0____38098));
  nor2s1 _______497282(.DIN1 (_________37790), .DIN2 (____0____38060),
       .Q (____0____38097));
  xor2s1 _______497283(.DIN1 (___0_____40532), .DIN2 (____9____38024),
       .Q (____0____38096));
  xor2s1 ______497284(.DIN1 (____9_9__38018), .DIN2 (___0_____40548),
       .Q (____0____38095));
  nor2s1 _______497285(.DIN1 (____0_0__38093), .DIN2 (____0____38058),
       .Q (____0____38094));
  xor2s1 _______497286(.DIN1 (____0____38067), .DIN2
       (_____________________________________________21927), .Q
       (____0____38092));
  xor2s1 _______497287(.DIN1 (____00___38039), .DIN2 (____0____38091),
       .Q (_____09__38140));
  nnd2s1 _______497288(.DIN1 (____0____38090), .DIN2 (____9____38026),
       .Q (_________38149));
  dffacs1 _______________________________________________497289(.CLRB
       (reset), .CLK (clk), .DIN (____00___38044), .QN
       (_____________________________________________21897));
  xnr2s1 _______497290(.DIN1 (_________38463), .DIN2 (____0____38088),
       .Q (____0____38089));
  and2s1 _____497291(.DIN1 (____0____38086), .DIN2 (_______22173), .Q
       (____0____38087));
  nnd2s1 _____497292(.DIN1 (____9_9__38028), .DIN2 (____0_0__38084), .Q
       (____0____38085));
  nnd2s1 _______497293(.DIN1 (____9____37998), .DIN2 (____9____38022),
       .Q (____0_9__38083));
  nnd2s1 _______497294(.DIN1 (____9____37989), .DIN2 (____000__38038),
       .Q (____0____38082));
  xor2s1 ______497295(.DIN1 (____00___38042), .DIN2 (____0____38088),
       .Q (____0____38081));
  xor2s1 _______497296(.DIN1 (____0____38059), .DIN2 (_________37789),
       .Q (____0____38080));
  xor2s1 _______497297(.DIN1 (____9___23128), .DIN2 (____0____38088),
       .Q (____0____38079));
  nor2s1 ______497298(.DIN1 (_________33293), .DIN2 (____0____38062),
       .Q (____0____38078));
  hi1s1 _______497299(.DIN (__________22062), .Q (____0____38077));
  xor2s1 _______497300(.DIN1 (_________37645), .DIN2 (____0____38088),
       .Q (____0____38099));
  nor2s1 ______497301(.DIN1 (_________36388), .DIN2 (____99___38032),
       .Q (______0__38151));
  and2s1 ______497302(.DIN1 (____9____38017), .DIN2 (___0_____40497),
       .Q (____0____38076));
  nor2s1 _______497303(.DIN1 (____9____37961), .DIN2 (____9____38023),
       .Q (____0____38075));
  nor2s1 _______497304(.DIN1 (____9____38014), .DIN2 (____0_9__38073),
       .Q (____0_0__38074));
  nor2s1 _______497305(.DIN1 (____9____38015), .DIN2 (____0____38071),
       .Q (____0____38072));
  nor2s1 ______497306(.DIN1 (____9____38013), .DIN2 (____0____38069),
       .Q (____0____38070));
  or2s1 _______497307(.DIN1
       (_____________________________________________21927), .DIN2
       (____0____38067), .Q (____0____38068));
  and2s1 ______497308(.DIN1 (____0____38067), .DIN2
       (_____________________________________________21927), .Q
       (____0____38066));
  xor2s1 _______497309(.DIN1 (____9____38003), .DIN2 (____0_0__38064),
       .Q (____0____38065));
  nnd2s1 _______497310(.DIN1 (____00___38041), .DIN2 (_____0__24945),
       .Q (____0_9__38063));
  nor2s1 _______497311(.DIN1 (_________37791), .DIN2 (____9____38011),
       .Q (____0____38114));
  nor2s1 _______497312(.DIN1
       (____________________________________________21846), .DIN2
       (____0____38062), .Q (_________38174));
  dffacs1 _______________________________________________497313(.CLRB
       (reset), .CLK (clk), .DIN (____99___38036), .Q
       (_____________________________________________21859));
  nnd2s1 _______497314(.DIN1 (____9_9__37992), .DIN2 (_____9___37752),
       .Q (____0____38061));
  nor2s1 _____0_497315(.DIN1 (______0__37786), .DIN2 (____0____38059),
       .Q (____0____38060));
  xnr2s1 _______497316(.DIN1
       (_____________________________________________21827), .DIN2
       (________22525), .Q (____0____38058));
  xor2s1 _______497317(.DIN1 (______0__36375), .DIN2 (____99___38031),
       .Q (____0____38057));
  nnd2s1 _____9_497318(.DIN1 (____9____38006), .DIN2 (____9____38005),
       .Q (____0_0__38056));
  nor2s1 _______497319(.DIN1 (____9_0__37968), .DIN2 (____9_0__38000),
       .Q (____0_9__38055));
  and2s1 ______497320(.DIN1 (____9____37051), .DIN2 (____9____38016),
       .Q (____0____38054));
  nor2s1 _______497321(.DIN1 (____9____38002), .DIN2 (____0____38052),
       .Q (____0____38108));
  dffacs1 _____________________________________________9_497322(.CLRB
       (reset), .CLK (clk), .DIN (____9____37995), .Q
       (__________22062));
  nor2s1 _______497323(.DIN1 (____9____37991), .DIN2 (____00___38045),
       .Q (____0____38051));
  xor2s1 _______497324(.DIN1 (_________37818), .DIN2 (____9____38010),
       .Q (____0____38050));
  and2s1 _______497325(.DIN1 (____9____38012), .DIN2 (____0____38048),
       .Q (____0____38049));
  xor2s1 _______497326(.DIN1
       (_________________________________________0___21786), .DIN2
       (____00___38045), .Q (____00___38046));
  nnd2s1 _______497327(.DIN1 (____9____37994), .DIN2 (_____90__36995),
       .Q (____00___38044));
  nor2s1 ______497328(.DIN1 (____0____38088), .DIN2 (_____0___37665),
       .Q (____00___38043));
  nnd2s1 _______497329(.DIN1 (____0____38088), .DIN2 (_________37233),
       .Q (____0____38090));
  nnd2s1 ______497330(.DIN1 (____00___38042), .DIN2 (____0____38088),
       .Q (_________38206));
  dffacs1 _________________________________________9_____497331(.CLRB
       (reset), .CLK (clk), .DIN (____9_9__38008), .Q
       (_____________________________________9_______21882));
  dffacs1 _____________________________________________0_497332(.CLRB
       (reset), .CLK (clk), .DIN (____9____37996), .QN
       (_________________________________________0___21814));
  dffacs1 ______________________________________________0_497333(.CLRB
       (reset), .CLK (clk), .DIN (____9_0__37993), .QN
       (__________________________________________________________________21988));
  nnd2s1 _____9_497334(.DIN1 (____9____37990), .DIN2 (inData[26]), .Q
       (____00___38041));
  xor2s1 _______497335(.DIN1 (____9____37971), .DIN2 (_________38200),
       .Q (____00___38040));
  xor2s1 _______497336(.DIN1 (____9____38004), .DIN2 (____9____37972),
       .Q (____00___38039));
  or2s1 _______497337(.DIN1
       (_____________________________________________21827), .DIN2
       (____999__38037), .Q (____000__38038));
  nnd2s1 _______497338(.DIN1 (_____9___37464), .DIN2 (____9____37987),
       .Q (____99___38036));
  or2s1 _______497339(.DIN1
       (______________________________________________21903), .DIN2
       (____99___38033), .Q (____99___38035));
  nnd2s1 _______497340(.DIN1 (____99___38033), .DIN2
       (______________________________________________21903), .Q
       (____99___38034));
  nor2s1 _______497341(.DIN1 (_________36346), .DIN2 (____99___38031),
       .Q (____99___38032));
  nor2s1 _______497342(.DIN1 (___0_____40495), .DIN2
       (_____________________________________________21827), .Q
       (____99___38030));
  nnd2s1 _______497343(.DIN1 (_________37648), .DIN2 (____99___38033),
       .Q (____99___38029));
  nnd2s1 _______497344(.DIN1 (____99___38033), .DIN2 (_________37598),
       .Q (____9_9__38028));
  nor2s1 _______497345(.DIN1 (____99___38033), .DIN2 (_________37619),
       .Q (____9____38027));
  nnd2s1 _______497346(.DIN1 (____99___38033), .DIN2 (_________37262),
       .Q (____9____38026));
  nnd2s1 _______497347(.DIN1 (____999__38037), .DIN2
       (_____________________________________________21827), .Q
       (____9____38025));
  nor2s1 _______497348(.DIN1 (____99___38033), .DIN2 (_________37618),
       .Q (_____90__38218));
  xor2s1 _______497349(.DIN1 (___09____40668), .DIN2 (_________37924),
       .Q (____0____38067));
  nor2s1 _______497350(.DIN1 (_________32032), .DIN2
       (_________________________________________0___21786), .Q
       (____9____38024));
  nnd2s1 _____497351(.DIN1 (_________37868), .DIN2 (____9____37982), .Q
       (____9____38023));
  nnd2s1 _____9_497352(.DIN1 (____9____37981), .DIN2 (inData[10]), .Q
       (____9____38022));
  nnd2s1 _____9_497353(.DIN1 (____9____37979), .DIN2 (inData[4]), .Q
       (____9____38021));
  nor2s1 _______497354(.DIN1 (____9____37997), .DIN2 (____9_0__38019),
       .Q (____9____38020));
  or2s1 _______497355(.DIN1
       (_________________________________________0___21786), .DIN2
       (___0_____40532), .Q (____9_9__38018));
  hi1s1 _______497356(.DIN (____9____38016), .Q (____9____38017));
  nor2s1 _______497357(.DIN1
       (_________________________________________0___21786), .DIN2
       (_________37715), .Q (____9____38015));
  nor2s1 ______497358(.DIN1 (__99_9__30508), .DIN2
       (_________________________________________0___21786), .Q
       (____9____38014));
  hi1s1 _____0_497359(.DIN (____9____38012), .Q (____9____38013));
  nor2s1 ______497360(.DIN1 (_________37800), .DIN2 (____9____38010),
       .Q (____9____38011));
  dffacs1 ________________497361(.CLRB (reset), .CLK (clk), .DIN
       (____99___38033), .Q (outData[18]));
  xor2s1 _______497362(.DIN1 (____9____37963), .DIN2 (___9_____39627),
       .Q (____0____38086));
  or2s1 _____497363(.DIN1 (___0_0___40465), .DIN2 (____009__38047), .Q
       (____0____38062));
  dffacs1 _______________________________________________497364(.CLRB
       (reset), .CLK (clk), .DIN (____9____37980), .QN
       (_____________________________________________21787));
  dffacs1 _____________________________________________9_497365(.CLRB
       (reset), .CLK (clk), .DIN (____9____37988), .QN
       (___0_____40549));
  dffacs1 _____________________________________________0_497366(.CLRB
       (reset), .CLK (clk), .DIN (____9____37983), .QN
       (_________________________________________0___21824));
  nnd2s1 _______497367(.DIN1 (____9____37959), .DIN2 (________22977),
       .Q (____9_0__38009));
  nnd2s1 _______497368(.DIN1 (____9____37969), .DIN2 (________25712),
       .Q (____9_9__38008));
  nor2s1 _______497369(.DIN1 (____9____37977), .DIN2 (____9____37973),
       .Q (____9____38006));
  or2s1 _______497370(.DIN1 (_________37616), .DIN2 (____9____38004),
       .Q (____9____38005));
  xor2s1 _______497371(.DIN1 (____90___37955), .DIN2 (____9_0__37043),
       .Q (____9____38003));
  nor2s1 _____9_497372(.DIN1 (____9____37966), .DIN2 (____9____38001),
       .Q (____9____38002));
  nnd2s1 _____9_497373(.DIN1 (_____9___37466), .DIN2 (____9_9__37974),
       .Q (____9_0__38000));
  nnd2s1 _____497374(.DIN1 (____9____37998), .DIN2 (____9____37964), .Q
       (____9____38016));
  xor2s1 _______497375(.DIN1 (____90___37953), .DIN2
       (___________________), .Q (____0____38059));
  hi1s1 _____497376(.DIN (____99___38033), .Q (____0____38088));
  nnd2s1 ______497377(.DIN1 (____9____37962), .DIN2 (________26461), .Q
       (____9____37996));
  nnd2s1 _______497378(.DIN1 (____9_9__37967), .DIN2 (_________38253),
       .Q (____9____37995));
  nnd2s1 ______497379(.DIN1 (______0__38770), .DIN2 (____9_0__37958),
       .Q (____9____37994));
  nnd2s1 _______497380(.DIN1 (____909__37957), .DIN2 (__9_____29949),
       .Q (____9_0__37993));
  xor2s1 _______497381(.DIN1 (_____0__28897), .DIN2 (_____9___37946),
       .Q (____9_9__37992));
  hi1s1 _______497382(.DIN
       (_________________________________________0___21786), .Q
       (____9____37991));
  xor2s1 _______497383(.DIN1 (______9__37938), .DIN2 (_________41343),
       .Q (____9____38012));
  xor2s1 ______497384(.DIN1 (_____9___37945), .DIN2 (____9_9__37984),
       .Q (____0____38053));
  dffacs1 _______________________________________________497385(.CLRB
       (reset), .CLK (clk), .DIN (____9____37965), .QN
       (_____________________________________________21802));
  dffacs1 ____________________________________0_497386(.CLRB (reset),
       .CLK (clk), .DIN (____9_0__37975), .QN (_________0_));
  and2s1 _______497387(.DIN1 (_____9__25785), .DIN2 (____90___37956),
       .Q (____9____37990));
  or2s1 _______497388(.DIN1 (______9__38245), .DIN2 (____900__37949),
       .Q (____9____37988));
  nnd2s1 _____9_497389(.DIN1 (____90___37950), .DIN2 (inData[20]), .Q
       (____9____37987));
  nor2s1 _______497390(.DIN1 (_________37889), .DIN2 (____9_0__37985),
       .Q (____9____37986));
  xnr2s1 _______497391(.DIN1 (___9_____39627), .DIN2 (_________37907),
       .Q (_________38272));
  xor2s1 _______497392(.DIN1 (_________37936), .DIN2 (____9_9__37984),
       .Q (____9____38010));
  dffacs1 _______________________________________________497393(.CLRB
       (reset), .CLK (clk), .DIN (____90___37954), .Q
       (_____________________________________________21827));
  nnd2s1 _______497394(.DIN1 (______0__36038), .DIN2 (_____9___37941),
       .Q (____9____37983));
  nnd2s1 ______497395(.DIN1 (______0__37929), .DIN2 (_____9___37947),
       .Q (____9____37982));
  or2s1 _______497396(.DIN1 (____9____37978), .DIN2 (___0_____40497),
       .Q (____9____37981));
  nnd2s1 _______497397(.DIN1 (_____9___37942), .DIN2 (________27076),
       .Q (____9____37980));
  nor2s1 ______497398(.DIN1 (_____9___37940), .DIN2 (___0____24191), .Q
       (____9____37979));
  nor2s1 _______497399(.DIN1 (____9____37978), .DIN2 (_________36937),
       .Q (____9____37997));
  xor2s1 ______497400(.DIN1 (_________37906), .DIN2 (_________38271),
       .Q (____99___38031));
  dffacs1 _______________________________________________497401(.CLRB
       (reset), .CLK (clk), .DIN (____90___37951), .Q (___0_0___40465));
  dffacs1 _____________________________________________0_497402(.CLRB
       (reset), .CLK (clk), .DIN (_____90__37939), .QN
       (_________________________________________0___21786));
  xnr2s1 _______497403(.DIN1 (___0_90__40451), .DIN2 (_________37915),
       .Q (____99___38033));
  nor2s1 _______497404(.DIN1 (_________37893), .DIN2 (_________37927),
       .Q (____9____37977));
  nnd2s1 _______497405(.DIN1 (_________37935), .DIN2 (_________38838),
       .Q (____9____37976));
  nnd2s1 _____9_497406(.DIN1 (____09__25687), .DIN2 (_________37930),
       .Q (____9_0__37975));
  or2s1 _______497407(.DIN1 (___0_9___40457), .DIN2 (____9____37960),
       .Q (____9_9__37974));
  nor2s1 ______497408(.DIN1 (____9____37972), .DIN2 (____90___37952),
       .Q (____9____37973));
  nor2s1 _______497409(.DIN1 (____9____37970), .DIN2 (_____99__37948),
       .Q (____9____37971));
  nnd2s1 _______497410(.DIN1 (______9__37928), .DIN2 (_________41345),
       .Q (____9____37969));
  nnd2s1 _____0_497411(.DIN1 (_________37933), .DIN2 (_________35142),
       .Q (____9____37989));
  xor2s1 _______497412(.DIN1 (___0_____40191), .DIN2 (_________37926),
       .Q (____9____38004));
  nor2s1 _____9_497413(.DIN1 (_________37923), .DIN2 (____0____40764),
       .Q (____9____37999));
  dffacs1 _________________________________________9_____497414(.CLRB
       (reset), .CLK (clk), .DIN (_________37931), .Q
       (_____________________________________9_______21881));
  nor2s1 _______497415(.DIN1 (______9__37919), .DIN2 (_________37834),
       .Q (____9_0__37968));
  nor2s1 _______497416(.DIN1 (_____9___41305), .DIN2 (_________37921),
       .Q (____9_9__37967));
  nnd2s1 _______497417(.DIN1 (___0_____40506), .DIN2 (___0_____40482),
       .Q (____9____37966));
  nnd2s1 _______497418(.DIN1 (____9____37068), .DIN2 (_________37916),
       .Q (____9____37965));
  nor2s1 ______497419(.DIN1 (___0_____40482), .DIN2 (___0_____40506),
       .Q (____9____37964));
  nor2s1 _______497420(.DIN1 (_________37913), .DIN2 (_________37917),
       .Q (____9____37963));
  nnd2s1 _______497421(.DIN1 (_________37911), .DIN2 (_________37717),
       .Q (____9____37962));
  nor2s1 _______497422(.DIN1 (______9__37891), .DIN2 (____9____37960),
       .Q (____9____37961));
  xor2s1 _______497423(.DIN1 (________22523), .DIN2 (_________37896),
       .Q (____9____37959));
  xor2s1 _______497424(.DIN1
       (_____________________________________________21898), .DIN2
       (_________35859), .Q (____9_0__37958));
  nor2s1 _______497425(.DIN1 (_________37912), .DIN2 (__9_9___29889),
       .Q (____909__37957));
  nor2s1 _______497426(.DIN1 (___0_____40482), .DIN2 (_________36992),
       .Q (____9_0__38019));
  dffacs1 _______________________________________________497427(.CLRB
       (reset), .CLK (clk), .DIN (_________37918), .QN
       (_____________________________________________21858));
  xor2s1 _______497428(.DIN1
       (_____________________________________9___0___21880), .DIN2
       (_________0_), .Q (____90___37956));
  xor2s1 _______497429(.DIN1
       (_____________________________________________21826), .DIN2
       (_________37932), .Q (____90___37955));
  nnd2s1 ______497430(.DIN1 (_________37902), .DIN2 (________23322), .Q
       (____90___37954));
  nor2s1 ______497431(.DIN1 (_____9__22662), .DIN2 (______0__37901), .Q
       (____90___37953));
  or2s1 _______497432(.DIN1 (________25781), .DIN2 (_________37897), .Q
       (____90___37951));
  nor2s1 _______497433(.DIN1 (_________37899), .DIN2 (_____0__23852),
       .Q (____90___37950));
  nnd2s1 _______497434(.DIN1 (_________37905), .DIN2 (________25612),
       .Q (____900__37949));
  hi1s1 _______497435(.DIN (___0_____40482), .Q (____9____37978));
  hi1s1 ______497436(.DIN (_____99__37948), .Q (____9_0__37985));
  nnd2s1 _____497437(.DIN1 (______0__37892), .DIN2 (inData[30]), .Q
       (_____9___37947));
  nor2s1 _____9_497438(.DIN1 (_____0___36638), .DIN2 (_________37904),
       .Q (_____9___37946));
  nnd2s1 _____9_497439(.DIN1 (_____99__37852), .DIN2 (_________37898),
       .Q (_____9___37945));
  nor2s1 _____497440(.DIN1 (____0____40762), .DIN2 (_____9___37943), .Q
       (_____9___37944));
  nnd2s1 _______497441(.DIN1 (_________37894), .DIN2 (_________38177),
       .Q (_____9___37942));
  nnd2s1 _______497442(.DIN1 (_________37895), .DIN2 (inData[6]), .Q
       (_____9___37941));
  xor2s1 _______497443(.DIN1 (___0_____40615), .DIN2
       (______________________________________0_______21889), .Q
       (_____9___37940));
  nnd2s1 _______497444(.DIN1 (_________37890), .DIN2 (_________41347),
       .Q (_____90__37939));
  nnd2s1 _______497445(.DIN1 (_________37937), .DIN2
       (_____________________________________________21898), .Q
       (______9__37938));
  or2s1 _____0_497446(.DIN1
       (_____________________________________________21898), .DIN2
       (_________37937), .Q (____0____38048));
  nnd2s1 _______497447(.DIN1 (_________37885), .DIN2 (_____0___37857),
       .Q (_________37936));
  nnd2s1 _____9_497448(.DIN1 (_____0___37859), .DIN2 (_________37887),
       .Q (_________37935));
  nor2s1 _______497449(.DIN1 (____9____37998), .DIN2 (_________37886),
       .Q (_________37934));
  or2s1 _______497450(.DIN1 (_________35135), .DIN2 (_________37932),
       .Q (_________37933));
  nnd2s1 _______497451(.DIN1 (_________37883), .DIN2 (_____9__26362),
       .Q (_________37931));
  or2s1 _______497452(.DIN1
       (_____________________________________9___0___21880), .DIN2
       (______0__37929), .Q (_________37930));
  xor2s1 _______497453(.DIN1 (_____0__22663), .DIN2 (______9__37900),
       .Q (______9__37928));
  nnd2s1 _______497454(.DIN1 (______0__37920), .DIN2 (_________37926),
       .Q (_________37927));
  nnd2s1 _______497455(.DIN1 (_________37922), .DIN2 (_________37924),
       .Q (_________37925));
  nor2s1 _______497456(.DIN1 (_________37924), .DIN2 (_________37922),
       .Q (_________37923));
  nnd2s1 _______497457(.DIN1 (_________37873), .DIN2 (___09___26136),
       .Q (_________37921));
  xor2s1 _______497458(.DIN1 (_____0___37856), .DIN2 (_________41252),
       .Q (_____99__37948));
  nor2s1 ______497459(.DIN1 (_________37926), .DIN2 (______0__37920),
       .Q (____90___37952));
  nor2s1 _______497460(.DIN1 (___99____39814), .DIN2 (_________37879),
       .Q (______9__37919));
  nnd2s1 _____9_497461(.DIN1 (_____9___37845), .DIN2 (_________37888),
       .Q (_________37918));
  nor2s1 _____9_497462(.DIN1 (___0_90__40451), .DIN2 (_________37914),
       .Q (_________37917));
  nnd2s1 _____9_497463(.DIN1 (_________37880), .DIN2 (________24882),
       .Q (_________37916));
  or2s1 _____9_497464(.DIN1 (_________37914), .DIN2 (_________37913),
       .Q (_________37915));
  nor2s1 _______497465(.DIN1 (___0_____40615), .DIN2 (_____9__28617),
       .Q (_________37912));
  xor2s1 ______497466(.DIN1 (_____0___36640), .DIN2 (_________37903),
       .Q (_________37911));
  or2s1 ______497467(.DIN1 (______9__37909), .DIN2 (_________37908), .Q
       (______0__37910));
  nor2s1 _______497468(.DIN1 (______0__37833), .DIN2 (_________37874),
       .Q (_________37907));
  nor2s1 _______497469(.DIN1 (_________37870), .DIN2 (______9__37871),
       .Q (_________37906));
  nnd2s1 _______497470(.DIN1 (______0__37929), .DIN2 (_________37869),
       .Q (____9____37960));
  dffacs1 _______________________________________________497471(.CLRB
       (reset), .CLK (clk), .DIN (______0__37882), .Q (___0_____40482));
  dffacs1 _______________________________________________497472(.CLRB
       (reset), .CLK (clk), .DIN (______9__37881), .QN
       (___0_____40516));
  nnd2s1 _______497473(.DIN1 (_________37865), .DIN2 (_________38177),
       .Q (_________37905));
  nor2s1 _______497474(.DIN1 (_____0___36639), .DIN2 (_________37903),
       .Q (_________37904));
  nnd2s1 _____0_497475(.DIN1 (_____0___37860), .DIN2 (_________38249),
       .Q (_________37902));
  nor2s1 ______497476(.DIN1 (________22661), .DIN2 (______9__37900), .Q
       (______0__37901));
  xor2s1 _______497477(.DIN1
       (_____________________________________________21873), .DIN2
       (____99___36174), .Q (_________37899));
  nnd2s1 _______497478(.DIN1 (_____00__37853), .DIN2 (_____9___34189),
       .Q (_________37898));
  hi1s1 _____0_497479(.DIN (______0__37920), .Q (___0_____40191));
  nor2s1 _______497480(.DIN1 (_________38833), .DIN2 (_____9___37848),
       .Q (_________37897));
  nnd2s1 _______497481(.DIN1 (_____0___37854), .DIN2
       (_____________________________________________21815), .Q
       (_________37896));
  nnd2s1 _______497482(.DIN1 (______9__37804), .DIN2 (_____09__37862),
       .Q (_________37895));
  xor2s1 ______497483(.DIN1 (_________37821), .DIN2 (_________37893),
       .Q (_________37894));
  nnd2s1 ______497484(.DIN1 (______9__37891), .DIN2 (_____9___37850),
       .Q (______0__37892));
  nnd2s1 _____497485(.DIN1 (_____9___37849), .DIN2 (____0_9__38073), .Q
       (_________37890));
  hi1s1 ______497486(.DIN (_________37889), .Q (____9____37970));
  dffacs1 _______________________________________________497487(.CLRB
       (reset), .CLK (clk), .DIN (_____0___37855), .QN
       (_____________________________________________21898));
  nnd2s1 ______497488(.DIN1 (_____0___37861), .DIN2 (____0____36220),
       .Q (_________37888));
  nnd2s1 _______497489(.DIN1 (_____9___37844), .DIN2 (_________37810),
       .Q (_________37887));
  xor2s1 ______497490(.DIN1 (_________37817), .DIN2 (_________37841),
       .Q (_________37886));
  xor2s1 ______497491(.DIN1 (_____0___37858), .DIN2 (_________37884),
       .Q (_________37885));
  nnd2s1 _______497492(.DIN1 (_________37840), .DIN2 (_________41345),
       .Q (_________37883));
  or2s1 _______497493(.DIN1 (____0____38052), .DIN2 (_________37830),
       .Q (______0__37882));
  nnd2s1 _______497494(.DIN1 (_________37839), .DIN2 (_________38550),
       .Q (______9__37881));
  nnd2s1 _______497495(.DIN1 (______0__37863), .DIN2 (_________37749),
       .Q (_________37880));
  nor2s1 ______497496(.DIN1 (_____________22082), .DIN2
       (_____9___37755), .Q (_________37879));
  or2s1 _______497497(.DIN1 (_________37877), .DIN2 (_________37876),
       .Q (_________37878));
  nor2s1 _______497498(.DIN1 (_________37801), .DIN2 (______9__37842),
       .Q (_________37932));
  dffacs1 _________________________________________9___0_497499(.CLRB
       (reset), .CLK (clk), .DIN (_____90__37843), .QN
       (_____________________________________9___0___21880));
  xor2s1 _______497500(.DIN1 (_________37812), .DIN2 (____9____38961),
       .Q (______0__37920));
  xor2s1 _______497501(.DIN1 (_________37811), .DIN2 (_____9___37851),
       .Q (_________37922));
  nnd2s1 _______497502(.DIN1 (_____9___38509), .DIN2 (______9__37823),
       .Q (_________37875));
  nnd2s1 _______497503(.DIN1 (______9__37832), .DIN2 (_____0___37664),
       .Q (_________37874));
  nnd2s1 _______497504(.DIN1 (_________37829), .DIN2 (______0__37872),
       .Q (_________37873));
  nor2s1 _______497505(.DIN1 (_____0___38422), .DIN2 (______0__37824),
       .Q (______9__37871));
  and2s1 _______497506(.DIN1 (_________37827), .DIN2 (_____0___38422),
       .Q (_________37870));
  and2s1 _______497507(.DIN1 (_____0___37764), .DIN2
       (_____________22082), .Q (_________37869));
  nnd2s1 _______497508(.DIN1 (_________37835), .DIN2 (___0_____40625),
       .Q (_________37868));
  nor2s1 _______497509(.DIN1 (_________37867), .DIN2
       (_____________________________________________21873), .Q
       (_________37908));
  and2s1 _______497510(.DIN1 (_________37866), .DIN2
       (_____________22082), .Q (_________37914));
  nnd2s1 ______497511(.DIN1 (_________37828), .DIN2 (_________37780),
       .Q (_________37889));
  dffacs1 __________________________________________0___0_497512(.CLRB
       (reset), .CLK (clk), .DIN (_________37819), .QN
       (___0_____40615));
  and2s1 _______497513(.DIN1 (_________37867), .DIN2
       (_____________________________________________21873), .Q
       (______9__37909));
  nor2s1 _______497514(.DIN1 (_____________22082), .DIN2
       (_________37866), .Q (_________37913));
  dffacs1 _______________________________________________497515(.CLRB
       (reset), .CLK (clk), .DIN (_________37838), .Q (___0_____40612));
  xor2s1 _______497516(.DIN1 (_________37771), .DIN2 (_________37864),
       .Q (_________37865));
  hi1s1 _______497517(.DIN (_____0___37861), .Q (_____09__37862));
  xor2s1 _______497518(.DIN1 (_________37825), .DIN2 (_________37826),
       .Q (_____0___37860));
  nnd2s1 _______497519(.DIN1 (_____0___37858), .DIN2 (_____0___37857),
       .Q (_____0___37859));
  xor2s1 _______497520(.DIN1 (_________37783), .DIN2 (______0__37776),
       .Q (_____0___37856));
  nor2s1 _______497521(.DIN1 (_____9___37564), .DIN2 (_________37816),
       .Q (______9__37900));
  nnd2s1 _______497522(.DIN1 (_________36807), .DIN2 (_________37803),
       .Q (_____0___37855));
  hi1s1 _______497523(.DIN
       (_____________________________________________21873), .Q
       (_____0___37854));
  nnd2s1 ______497524(.DIN1 (_________37808), .DIN2 (_________36566),
       .Q (_____00__37853));
  nnd2s1 _______497525(.DIN1 (_____9___37847), .DIN2 (_____9___37851),
       .Q (_____99__37852));
  hi1s1 _______497526(.DIN (_____________22082), .Q (_____9___37850));
  nnd2s1 ______497527(.DIN1 (___09____40669), .DIN2 (_________37820),
       .Q (_____9___37849));
  nor2s1 _____0_497528(.DIN1 (_________37809), .DIN2 (_____9___37847),
       .Q (_____9___37848));
  hi1s1 _____9_497529(.DIN (_____9___37846), .Q (_____0___38135));
  nor2s1 _______497530(.DIN1 (_________36785), .DIN2 (_________37806),
       .Q (_________37903));
  nor2s1 _______497531(.DIN1 (_________37798), .DIN2 (______0__37315),
       .Q (_____9___37845));
  nnd2s1 _____9_497532(.DIN1 (_____0___37857), .DIN2 (_________37797),
       .Q (_____9___37844));
  nnd2s1 ______497533(.DIN1 (_________37794), .DIN2 (________25648), .Q
       (_____90__37843));
  and2s1 _______497534(.DIN1 (_________37841), .DIN2 (_________37793),
       .Q (______9__37842));
  xor2s1 _______497535(.DIN1 (_____99__37565), .DIN2 (_________37815),
       .Q (_________37840));
  nor2s1 _______497536(.DIN1 (____09__26238), .DIN2 (_________37772),
       .Q (_________37839));
  or2s1 _____9_497537(.DIN1 (_________37837), .DIN2 (______9__37795),
       .Q (_________37838));
  nor2s1 _______497538(.DIN1 (_________37784), .DIN2 (________23533),
       .Q (_____0___37861));
  nor2s1 _______497539(.DIN1 (______9__37750), .DIN2 (______9__37785),
       .Q (______0__37863));
  hi1s1 _____9_497540(.DIN (_________37836), .Q (_________37876));
  dffacs1 _______________________________________________497541(.CLRB
       (reset), .CLK (clk), .DIN (_________37788), .QN
       (_____________________________________________21873));
  dffacs1 ______________________________________497542(.CLRB (reset),
       .CLK (clk), .DIN (_________37787), .Q (_____________22082));
  or2s1 _____0_497543(.DIN1 (______9__37891), .DIN2 (_________37834),
       .Q (_________37835));
  nor2s1 _____9_497544(.DIN1 (___090__23301), .DIN2 (_________37831),
       .Q (______0__37833));
  nnd2s1 _____9_497545(.DIN1 (_________37831), .DIN2 (___090__23301),
       .Q (______9__37832));
  nnd2s1 _____9_497546(.DIN1 (_________37781), .DIN2 (____0___25315),
       .Q (_________37830));
  xor2s1 _____497547(.DIN1 (______0__37805), .DIN2 (_________36786), .Q
       (_________37829));
  nnd2s1 _____0_497548(.DIN1 (_________37779), .DIN2 (_________37700),
       .Q (_________37828));
  and2s1 _____9_497549(.DIN1 (_________37826), .DIN2 (_________37825),
       .Q (_________37827));
  nor2s1 _____0_497550(.DIN1 (______0__37766), .DIN2 (______9__37775),
       .Q (______0__37824));
  xor2s1 _______497551(.DIN1 (_________22020), .DIN2 (_________37822),
       .Q (______9__37823));
  nnd2s1 _______497552(.DIN1 (_________37820), .DIN2 (________28328),
       .Q (_________37821));
  nnd2s1 _______497553(.DIN1 (_________37768), .DIN2 (______9__38496),
       .Q (_________37819));
  nnd2s1 _______497554(.DIN1 (_________37778), .DIN2 (_________37782),
       .Q (_____9___37846));
  xor2s1 _______497555(.DIN1 (_________37799), .DIN2
       (_____________________________________________21926), .Q
       (_________37818));
  xor2s1 _______497556(.DIN1 (______0__35032), .DIN2 (______09), .Q
       (_________37817));
  nor2s1 _______497557(.DIN1 (_____9___37563), .DIN2 (_________37815),
       .Q (_________37816));
  nor2s1 _______497558(.DIN1 (_________37725), .DIN2 (______9__37813),
       .Q (______0__37814));
  xor2s1 _____497559(.DIN1 (_____09__37765), .DIN2 (_____00__37663), .Q
       (_________37812));
  xor2s1 ______497560(.DIN1 (_________37739), .DIN2 (_________37737),
       .Q (_________37811));
  nor2s1 _____497561(.DIN1 (_________37810), .DIN2 (______0__37796), .Q
       (_____0___37858));
  xnr2s1 _______497562(.DIN1 (___9_0___39166), .DIN2 (_________37747),
       .Q (_________37836));
  and2s1 _______497563(.DIN1 (_________37807), .DIN2 (_________37802),
       .Q (_________37809));
  nnd2s1 _______497564(.DIN1 (_________37807), .DIN2 (_________36565),
       .Q (_________37808));
  and2s1 _______497565(.DIN1 (______0__37805), .DIN2 (_________36773),
       .Q (_________37806));
  nnd2s1 _______497566(.DIN1 (___09___24265), .DIN2 (_____0___37760),
       .Q (______9__37804));
  or2s1 ____9__497567(.DIN1 (_________22020), .DIN2 (________27099), .Q
       (_________37803));
  nor2s1 _______497568(.DIN1 (_________37802), .DIN2 (_________37807),
       .Q (_____9___37847));
  dffacs1 ______________________________________497569(.CLRB (reset),
       .CLK (clk), .DIN (_____0___37763), .Q (_____________22081));
  dffacs1 _______________________________________________497570(.CLRB
       (reset), .CLK (clk), .DIN (_____9___37758), .QN
       (_____________________________________________21785));
  dffacs1 _________________________________________9_____497571(.CLRB
       (reset), .CLK (clk), .DIN (_____0___37761), .Q (___0_____40623));
  nor2s1 _____0_497572(.DIN1 (______09), .DIN2 (_________37792), .Q
       (_________37801));
  nor2s1 _______497573(.DIN1
       (_____________________________________________21926), .DIN2
       (_________37799), .Q (_________37800));
  nor2s1 _______497574(.DIN1
       (_____________________________________________21872), .DIN2
       (___099__24266), .Q (_________37798));
  hi1s1 _______497575(.DIN (______0__37796), .Q (_________37797));
  nnd2s1 ______497576(.DIN1 (_____9___37756), .DIN2 (_____0__25882), .Q
       (______9__37795));
  nnd2s1 _______497577(.DIN1 (_____9___37754), .DIN2 (_________37834),
       .Q (_________37794));
  nnd2s1 _____0_497578(.DIN1 (_________37792), .DIN2 (______09), .Q
       (_________37793));
  and2s1 _______497579(.DIN1 (_________37799), .DIN2
       (_____________________________________________21926), .Q
       (_________37791));
  and2s1 _______497580(.DIN1 (_________37789), .DIN2
       (_____________________________________________21872), .Q
       (_________37790));
  nnd2s1 _______497581(.DIN1 (_____9___37753), .DIN2 (____99__22740),
       .Q (_________37788));
  or2s1 ______497582(.DIN1 (________26853), .DIN2 (______9__37740), .Q
       (_________37787));
  nor2s1 ______497583(.DIN1 (_________37789), .DIN2
       (_____________________________________________21872), .Q
       (______0__37786));
  nor2s1 _______497584(.DIN1 (_________37748), .DIN2 (_____90__37751),
       .Q (______9__37785));
  nnd2s1 _______497585(.DIN1
       (_____________________________________________21872), .DIN2
       (_____________________________________________21841), .Q
       (_________37784));
  nnd2s1 _______497586(.DIN1 (___09_9__40670), .DIN2
       (_____________________________________________21925), .Q
       (_____0___37857));
  and2s1 _______497587(.DIN1 (_________37782), .DIN2 (_________37777),
       .Q (_________37783));
  nnd2s1 _______497588(.DIN1 (_________37742), .DIN2 (____9____38001),
       .Q (_________37781));
  or2s1 _______497589(.DIN1 (___9_0___39170), .DIN2 (_________37738),
       .Q (_________37780));
  nnd2s1 _______497590(.DIN1 (_________37743), .DIN2 (_________37697),
       .Q (_________37779));
  nnd2s1 _______497591(.DIN1 (_________37777), .DIN2 (______0__37776),
       .Q (_________37778));
  nor2s1 _______497592(.DIN1 (_________37767), .DIN2 (_________37826),
       .Q (______9__37775));
  and2s1 ____9__497593(.DIN1 (_________37773), .DIN2 (_____0___37280),
       .Q (_________37774));
  nor2s1 _______497594(.DIN1 (_________38435), .DIN2 (______0__37741),
       .Q (_________37772));
  xor2s1 ______497595(.DIN1 (_________37716), .DIN2
       (_________________________________________9_), .Q
       (_________37771));
  or2s1 ____9__497596(.DIN1 (_________37769), .DIN2 (_________37773),
       .Q (_________37770));
  nor2s1 ______497597(.DIN1 (________23324), .DIN2 (_________37745), .Q
       (_________37768));
  nor2s1 _______497598(.DIN1 (_________37767), .DIN2 (______0__37766),
       .Q (_________37825));
  nnd2s1 _______497599(.DIN1 (_____99__37759), .DIN2 (________28979),
       .Q (_________37820));
  nnd2s1 _______497600(.DIN1 (_____09__37765), .DIN2 (_________37680),
       .Q (_________37831));
  xor2s1 _______497601(.DIN1 (_____0___37764), .DIN2 (___0_9___40457),
       .Q (______9__37891));
  nnd2s1 _______497602(.DIN1 (_________37728), .DIN2 (_________37554),
       .Q (_____0___37763));
  nnd2s1 _______497603(.DIN1 (_________37727), .DIN2 (______9__37652),
       .Q (_____0___37761));
  hi1s1 _______497604(.DIN
       (_____________________________________________21872), .Q
       (_____0___37760));
  nor2s1 ______497605(.DIN1 (______0__37411), .DIN2 (______9__37730),
       .Q (_________37815));
  xor2s1 ______497606(.DIN1 (______9__37710), .DIN2 (_________41248),
       .Q (______9__37813));
  xor2s1 _______497607(.DIN1 (_________37706), .DIN2 (____0_0__38084),
       .Q (______0__37796));
  nnd2s1 _______497608(.DIN1 (_________37718), .DIN2 (________25393),
       .Q (_____9___37758));
  nnd2s1 _______497609(.DIN1 (______0__37721), .DIN2 (_____0___36372),
       .Q (______0__37805));
  nor2s1 _______497610(.DIN1 (____0____35356), .DIN2 (_________37714),
       .Q (_________38284));
  dffacs1 __________________________________________0____(.CLRB
       (reset), .CLK (clk), .DIN (_________37724), .Q (_________22020));
  dffacs1 _______________________________________________497611(.CLRB
       (reset), .CLK (clk), .DIN (_________37732), .QN
       (_______________________________________________________________0__21998));
  nnd2s1 _______497612(.DIN1 (_________37719), .DIN2 (_________36488),
       .Q (_________37807));
  dffacs1 _______________________________________________497613(.CLRB
       (reset), .CLK (clk), .DIN (_________37723), .QN
       (___0_____40483));
  nnd2s1 _______497614(.DIN1 (___90____39051), .DIN2 (_________37708),
       .Q (_____9___37757));
  nnd2s1 _______497615(.DIN1 (______0__37711), .DIN2 (_________37230),
       .Q (_____9___37756));
  nor2s1 _______497616(.DIN1 (___0_9___40457), .DIN2 (___0_____40625),
       .Q (_____9___37755));
  xor2s1 ______497617(.DIN1 (___09____40672), .DIN2 (_________37729),
       .Q (_____9___37754));
  nnd2s1 _______497618(.DIN1 (_________37699), .DIN2 (_____9___37752),
       .Q (_____9___37753));
  or2s1 _______497619(.DIN1
       (_____________________________________________21813), .DIN2
       (_____________________________________________21802), .Q
       (_____90__37751));
  and2s1 ______497620(.DIN1
       (_____________________________________________21802), .DIN2
       (_____________________________________________21813), .Q
       (______9__37750));
  nnd2s1 _______497621(.DIN1 (_________37748), .DIN2
       (_____________________________________________21813), .Q
       (_________37749));
  nor2s1 _______497622(.DIN1
       (_________________________________________________________________22000),
       .DIN2 (_________37746), .Q (_________37747));
  and2s1 _______497623(.DIN1 (_________37746), .DIN2
       (_________________________________________________________________22000),
       .Q (_________37877));
  dffacs1 _______________________________________________497624(.CLRB
       (reset), .CLK (clk), .DIN (_________37709), .Q (______09));
  xor2s1 ______497625(.DIN1 (_________37691), .DIN2 (_________37638),
       .Q (_________37799));
  dffacs1 _______________________________________________497626(.CLRB
       (reset), .CLK (clk), .DIN (_________37712), .QN
       (_____________________________________________21872));
  and2s1 ____9__497627(.DIN1 (_________37698), .DIN2 (_________37744),
       .Q (_________37745));
  nnd2s1 _______497628(.DIN1 (______0__37702), .DIN2 (___9_0___39170),
       .Q (_________37743));
  xor2s1 _______497629(.DIN1 (____0____35357), .DIN2 (_________37713),
       .Q (_________37742));
  xor2s1 _______497630(.DIN1 (_________36405), .DIN2 (______9__37720),
       .Q (______0__37741));
  nor2s1 _______497631(.DIN1 (___0_____40625), .DIN2 (_____0__26599),
       .Q (______9__37740));
  nor2s1 _____9_497632(.DIN1 (______9__37701), .DIN2 (_________37736),
       .Q (_________37739));
  or2s1 ______497633(.DIN1 (_________37737), .DIN2 (_________37736), .Q
       (_________37738));
  and2s1 _____497634(.DIN1 (_________37735), .DIN2
       (_____________________________________________21813), .Q
       (_________37767));
  nor2s1 _______497635(.DIN1
       (_____________________________________________21813), .DIN2
       (_________37735), .Q (______0__37766));
  nnd2s1 _____9_497636(.DIN1 (_________37746), .DIN2 (_________37734),
       .Q (_________37777));
  xnr2s1 _____9_497637(.DIN1 (___9_9___39790), .DIN2 (_________37684),
       .Q (_____09__37765));
  nnd2s1 ____90_497638(.DIN1 (_________37704), .DIN2 (_____0___35475),
       .Q (_____99__37759));
  or2s1 ______497639(.DIN1 (_________37734), .DIN2 (_________37746), .Q
       (_________37782));
  nor2s1 ____9__497640(.DIN1 (______9__37682), .DIN2 (_________37733),
       .Q (_________37773));
  dffacs1 _____________________________________________9_497641(.CLRB
       (reset), .CLK (clk), .DIN (_________37707), .QN
       (_________22043));
  nnd2s1 _____9_497642(.DIN1 (_________37696), .DIN2 (______0__37731),
       .Q (_________37732));
  and2s1 _______497643(.DIN1 (_________37729), .DIN2 (_________37413),
       .Q (______9__37730));
  nnd2s1 ______497644(.DIN1 (________27402), .DIN2 (______0__37693), .Q
       (_________37728));
  nor2s1 _______497645(.DIN1 (______9__37692), .DIN2 (____0____37172),
       .Q (_________37727));
  hi1s1 _____9_497646(.DIN (_________37725), .Q (_________37726));
  nor2s1 _______497647(.DIN1 (_________37694), .DIN2 (_________37690),
       .Q (_____0___37762));
  hi1s1 _____9_497648(.DIN (___0_____40625), .Q (_____0___37764));
  nnd2s1 ____9__497649(.DIN1 (______0__37683), .DIN2 (_________37454),
       .Q (_________37724));
  nnd2s1 ____90_497650(.DIN1 (_________37685), .DIN2 (_________37722),
       .Q (_________37723));
  nnd2s1 ____90_497651(.DIN1 (______9__37720), .DIN2 (_________36389),
       .Q (______0__37721));
  nor2s1 ____90_497652(.DIN1 (______0__36481), .DIN2 (_________37689),
       .Q (_________37719));
  nnd2s1 ____9__497653(.DIN1 (_________37686), .DIN2 (_________37717),
       .Q (_________37718));
  xor2s1 ____9__497654(.DIN1 (_________37703), .DIN2 (_________37715),
       .Q (_________37716));
  nor2s1 ____90_497655(.DIN1 (____0____35355), .DIN2 (_________37713),
       .Q (_________37714));
  nnd2s1 ____90_497656(.DIN1 (_____0___37670), .DIN2 (________25790),
       .Q (_________37712));
  xor2s1 _______497657(.DIN1 (_____9___37659), .DIN2 (_________37580),
       .Q (______0__37711));
  nnd2s1 ____497658(.DIN1 (_________37705), .DIN2
       (_____________________________________________21954), .Q
       (______9__37710));
  or2s1 _______497659(.DIN1 (____0____38117), .DIN2 (_____09__37672),
       .Q (_________37709));
  nnd2s1 _____497660(.DIN1 (_________41337), .DIN2 (_____0___37669), .Q
       (_________37708));
  nnd2s1 ____497661(.DIN1 (_____0___37671), .DIN2 (_________37405), .Q
       (_________37707));
  nor2s1 _______497662(.DIN1
       (_____________________________________________21925), .DIN2
       (_________37695), .Q (_________37706));
  nor2s1 ____90_497663(.DIN1
       (_____________________________________________21954), .DIN2
       (_________37705), .Q (_________37725));
  nor2s1 _______497664(.DIN1 (_________37640), .DIN2 (_________37674),
       .Q (_________37810));
  dffacs1 __________________________________________0____497665(.CLRB
       (reset), .CLK (clk), .DIN (_____0___37667), .Q (___0_____40443));
  dffacs1 _________________________________________9___9_497666(.CLRB
       (reset), .CLK (clk), .DIN (_________37677), .Q (___0_____40625));
  dffacs1 _______________________________________________497667(.CLRB
       (reset), .CLK (clk), .DIN (_________37678), .Q
       (_____________________________________________21813));
  or2s1 ____9__497668(.DIN1 (_____0___35476), .DIN2 (_________37703),
       .Q (_________37704));
  nor2s1 ____9__497669(.DIN1 (_________36935), .DIN2 (_________37705),
       .Q (______0__37702));
  and2s1 ____9__497670(.DIN1 (_________37705), .DIN2 (_________37700),
       .Q (______9__37701));
  xor2s1 ____9__497671(.DIN1 (_________36487), .DIN2 (_________37688),
       .Q (_________37699));
  xor2s1 ____9__497672(.DIN1 (_________37644), .DIN2 (_________41341),
       .Q (_________37698));
  nnd2s1 ____9__497673(.DIN1 (_________37705), .DIN2 (____9____33397),
       .Q (_________37697));
  nor2s1 ____9_497674(.DIN1 (_________37700), .DIN2 (_________37705),
       .Q (_________37736));
  hi1s1 ____497675(.DIN (_________38147), .Q (_________37733));
  dffacs1 _______________________________________________497676(.CLRB
       (reset), .CLK (clk), .DIN (_________37675), .Q
       (_____________________________________________21826));
  xor2s1 ____9__497677(.DIN1 (_________37649), .DIN2 (_________37589),
       .Q (_________37746));
  dffacs1 _____________________________________________9_497678(.CLRB
       (reset), .CLK (clk), .DIN (_____0___37666), .QN
       (_________________________________________9___21803));
  dffacs1 __________________(.CLRB (reset), .CLK (clk), .DIN
       (_________37676), .QN (_______________22074));
  nor2s1 ____9__497679(.DIN1 (___000__26051), .DIN2 (_________37651),
       .Q (_________37696));
  xor2s1 _______497680(.DIN1 (_________37635), .DIN2 (___9_____39301),
       .Q (_________37694));
  or2s1 ____90_497681(.DIN1 (_________37634), .DIN2 (_____9___37660),
       .Q (______0__37693));
  nor2s1 ____9_497682(.DIN1 (_____9___37658), .DIN2 (______9__37555),
       .Q (______9__37692));
  xor2s1 _______497683(.DIN1 (_________37637), .DIN2 (_________37690),
       .Q (_________37691));
  and2s1 ____9__497684(.DIN1 (_________37688), .DIN2 (______0__36438),
       .Q (_________37689));
  nnd2s1 ____9__497685(.DIN1 (_____9___37655), .DIN2 (______0__37604),
       .Q (______9__37720));
  xor2s1 ____9__497686(.DIN1 (_________37624), .DIN2 (_________37687),
       .Q (_________37729));
  xor2s1 ____9__497687(.DIN1 (______9__37622), .DIN2 (________25804),
       .Q (_________37686));
  nor2s1 ____9__497688(.DIN1 (______0__41349), .DIN2 (_____9___37657),
       .Q (_________37685));
  nnd2s1 ____9__497689(.DIN1 (_________37650), .DIN2 (_________37544),
       .Q (_________37684));
  nor2s1 ____0_497690(.DIN1 (_________37646), .DIN2 (_________36956),
       .Q (______0__37683));
  nor2s1 ____99_497691(.DIN1 (_________37679), .DIN2 (_________37681),
       .Q (______9__37682));
  nnd2s1 ____00_497692(.DIN1 (____9____38961), .DIN2 (_________36739),
       .Q (_________37680));
  xor2s1 ____9__497693(.DIN1 (_________37628), .DIN2 (_____09__35744),
       .Q (_________37713));
  nnd2s1 ____0_497694(.DIN1 (_________37681), .DIN2 (_________37679),
       .Q (_________38147));
  dffacs1 _______________________________________________497695(.CLRB
       (reset), .CLK (clk), .DIN (_____9___37661), .QN
       (___0_____40484));
  dffacs1 ______________________________________497696(.CLRB (reset),
       .CLK (clk), .DIN (_____90__37653), .QN (___0_____40587));
  nnd2s1 ____9__497697(.DIN1 (_________37629), .DIN2 (_____9__22958),
       .Q (_________37678));
  nnd2s1 ____9__497698(.DIN1 (_________37641), .DIN2 (____0____38104),
       .Q (_________37677));
  nnd2s1 ____9__497699(.DIN1 (_________37630), .DIN2 (__90__), .Q
       (_________37676));
  nor2s1 ____9_497700(.DIN1 (_________38583), .DIN2 (_________37636),
       .Q (_________37675));
  xor2s1 ____9__497701(.DIN1 (_________37607), .DIN2 (______0__37673),
       .Q (_________37674));
  xor2s1 ____9__497702(.DIN1 (_________37606), .DIN2 (____9_0__36107),
       .Q (_____09__37672));
  dffacs1 __________________________________________0____497703(.CLRB
       (reset), .CLK (clk), .DIN (______9__37632), .Q
       (______________________________________0____));
  xor2s1 _____9_497704(.DIN1 (______0__37613), .DIN2 (______0__37584),
       .Q (_________37695));
  dffacs1 _____________________________________________0_497705(.CLRB
       (reset), .CLK (clk), .DIN (_________37631), .QN
       (_________________________________________0___21856));
  nor2s1 ____9__497706(.DIN1 (_________37626), .DIN2 (_________36335),
       .Q (_____0___37671));
  nnd2s1 ____9__497707(.DIN1 (_________37627), .DIN2 (______9__37314),
       .Q (_____0___37670));
  xor2s1 ____9__497708(.DIN1
       (_____________________________________________21909), .DIN2
       (_____0___37668), .Q (_____0___37669));
  nnd2s1 ____9_497709(.DIN1 (_________37625), .DIN2 (______9__38496),
       .Q (_____0___37667));
  nnd2s1 ____0__497710(.DIN1 (_________37620), .DIN2 (____90__23872),
       .Q (_____0___37666));
  xor2s1 ____99_497711(.DIN1 (_________37647), .DIN2 (_________37614),
       .Q (_____0___37665));
  nnd2s1 ____99_497712(.DIN1 (______9__37642), .DIN2 (_____00__37663),
       .Q (_____0___37664));
  xor2s1 ____497713(.DIN1 (______0__37594), .DIN2 (_____99__37662), .Q
       (_________37703));
  dffacs1 _______________________________________________497714(.CLRB
       (reset), .CLK (clk), .DIN (______0__37623), .QN
       (___0_____40525));
  xor2s1 ____9_497715(.DIN1 (_________37496), .DIN2 (_________37596),
       .Q (_________37705));
  nnd2s1 ____9__497716(.DIN1 (_________37605), .DIN2 (_____0___37283),
       .Q (_____9___37661));
  nnd2s1 ____9_497717(.DIN1 (_________37611), .DIN2 (_________37610),
       .Q (_____9___37660));
  xor2s1 ____9_497718(.DIN1 (_________37586), .DIN2 (_________37528),
       .Q (_____9___37659));
  xor2s1 ____9__497719(.DIN1 (___0_____40587), .DIN2 (______0__37633),
       .Q (_____9___37658));
  nor2s1 ____9__497720(.DIN1 (_____9___37656), .DIN2 (_________37591),
       .Q (_____9___37657));
  nnd2s1 ____9_497721(.DIN1 (_________37601), .DIN2 (_____9___37654),
       .Q (_____9___37655));
  nnd2s1 ____9_497722(.DIN1 (______9__37652), .DIN2 (_________37612),
       .Q (_____90__37653));
  nor2s1 ____9__497723(.DIN1 (______0__36385), .DIN2 (______9__37603),
       .Q (_________37688));
  nor2s1 ____9__497724(.DIN1 (____0____36193), .DIN2 (_________37609),
       .Q (_________37826));
  and2s1 ____99_497725(.DIN1 (___0_____30688), .DIN2
       (_____________________________________________21909), .Q
       (_________37651));
  nor2s1 ____99_497726(.DIN1 (_________37532), .DIN2 (_________37590),
       .Q (_________37650));
  nor2s1 ____00_497727(.DIN1 (_________37615), .DIN2 (_________37537),
       .Q (_________37649));
  and2s1 ____0__497728(.DIN1 (_________37647), .DIN2 (_________37202),
       .Q (_________37648));
  nor2s1 ____0__497729(.DIN1 (_________37588), .DIN2 (_________36670),
       .Q (_________37646));
  nnd2s1 ____0__497730(.DIN1 (_________37592), .DIN2 (_________37599),
       .Q (_________37645));
  or2s1 ____0__497731(.DIN1 (______9__37593), .DIN2 (____00___38042),
       .Q (_________37644));
  hi1s1 ____0__497732(.DIN (______0__37643), .Q (_________37681));
  dffacs1 _______________________________________________497733(.CLRB
       (reset), .CLK (clk), .DIN (_________37600), .Q
       (_____________________________________________21941));
  hi1s1 ____0__497734(.DIN (______9__37642), .Q (____9____38961));
  nor2s1 ____9__497735(.DIN1 (____9___26497), .DIN2 (_____0___37572),
       .Q (_________37641));
  nnd2s1 ____9__497736(.DIN1 (_________37582), .DIN2 (_________37529),
       .Q (_________37640));
  nnd2s1 ____9__497737(.DIN1 (_________37638), .DIN2 (_________37637),
       .Q (_________37639));
  xor2s1 ____9__497738(.DIN1 (_________36324), .DIN2 (_________37608),
       .Q (_________37636));
  nor2s1 ____9__497739(.DIN1 (_________37637), .DIN2 (_________37638),
       .Q (_________37635));
  and2s1 ____9__497740(.DIN1 (______0__37633), .DIN2 (___0_____40587),
       .Q (_________37634));
  nnd2s1 ____9__497741(.DIN1 (____9____36146), .DIN2 (_________37575),
       .Q (______9__37632));
  nnd2s1 ____9__497742(.DIN1 (____9____37085), .DIN2 (_________37577),
       .Q (_________37631));
  nnd2s1 ____9__497743(.DIN1 (_________37576), .DIN2 (_____0___37570),
       .Q (_________37630));
  nnd2s1 ____9__497744(.DIN1 (_____0___37568), .DIN2 (____0____37167),
       .Q (_________37629));
  nor2s1 ____9__497745(.DIN1 (___09_0__40671), .DIN2 (_________37585),
       .Q (_________37690));
  nnd2s1 ____0__497746(.DIN1 (______0__37574), .DIN2 (_________35176),
       .Q (_________37628));
  xor2s1 ____99_497747(.DIN1 (_________37602), .DIN2 (_____0___36458),
       .Q (_________37627));
  nor2s1 ____497748(.DIN1 (_________37578), .DIN2 (_________37317), .Q
       (_________37626));
  nor2s1 ____497749(.DIN1 (_____0___37571), .DIN2 (____0_9__37143), .Q
       (_________37625));
  nnd2s1 ____00_497750(.DIN1 (_________37517), .DIN2 (_____0___37567),
       .Q (_________37624));
  nnd2s1 ____99_497751(.DIN1 (_________37581), .DIN2 (_________37322),
       .Q (______0__37623));
  xor2s1 ____0__497752(.DIN1 (______9__37535), .DIN2 (_________37621),
       .Q (______9__37622));
  nnd2s1 ____0__497753(.DIN1 (_____00__37566), .DIN2 (_________37717),
       .Q (_________37620));
  hi1s1 ____0__497754(.DIN (_________37618), .Q (_________37619));
  xor2s1 ____0_497755(.DIN1 (_________37436), .DIN2 (_________37617),
       .Q (______9__37642));
  xor2s1 ____0__497756(.DIN1 (_________37617), .DIN2 (_________37616),
       .Q (______0__37643));
  nor2s1 ____0__497757(.DIN1 (_________37614), .DIN2 (_________37542),
       .Q (_________37615));
  nor2s1 ____9__497758(.DIN1 (___09_0__40671), .DIN2 (______9__37583),
       .Q (______0__37613));
  nor2s1 ____9__497759(.DIN1 (_____90__37556), .DIN2 (____9___25670),
       .Q (_________37612));
  nnd2s1 ____9__497760(.DIN1 (______0__37345), .DIN2 (_____9___37561),
       .Q (_________37611));
  or2s1 ____9__497761(.DIN1 (___0_____40587), .DIN2 (_____9___37560),
       .Q (_________37610));
  nor2s1 ____9_497762(.DIN1 (____0____36226), .DIN2 (_________37608),
       .Q (_________37609));
  nnd2s1 ____9__497763(.DIN1 (_____9___37559), .DIN2 (_________37579),
       .Q (_________37607));
  xor2s1 ____00_497764(.DIN1 (_________37522), .DIN2 (______0__37507),
       .Q (_________37606));
  nor2s1 ____0__497765(.DIN1 (________27329), .DIN2 (_________37550),
       .Q (_________37605));
  nnd2s1 ____0__497766(.DIN1 (_________37553), .DIN2 (_________34907),
       .Q (______0__37604));
  and2s1 ____0__497767(.DIN1 (_________37602), .DIN2 (_________36345),
       .Q (______9__37603));
  nnd2s1 ____0_497768(.DIN1 (______0__37546), .DIN2 (_____0___36548),
       .Q (_________37601));
  nnd2s1 ____9__497769(.DIN1 (_____9___37562), .DIN2 (_____9__25251),
       .Q (_________37600));
  dffacs1 _______________________________________________497770(.CLRB
       (reset), .CLK (clk), .DIN (_________37549), .QN
       (_____________________________________________21909));
  or2s1 ____497771(.DIN1 (_________37598), .DIN2 (_________37597), .Q
       (_________37599));
  nor2s1 ____0__497772(.DIN1 (_________37456), .DIN2 (_________37548),
       .Q (_________37596));
  nnd2s1 ____0_497773(.DIN1 (_________37597), .DIN2 (____9____38949),
       .Q (_________37595));
  nor2s1 ____0__497774(.DIN1 (_________37533), .DIN2 (______9__37545),
       .Q (______0__37594));
  nor2s1 ____09_497775(.DIN1 (_________37309), .DIN2 (_________37617),
       .Q (______9__37593));
  nnd2s1 ____09_497776(.DIN1 (_________37597), .DIN2 (_________37587),
       .Q (_________37592));
  xor2s1 ____0_497777(.DIN1 (_________35178), .DIN2 (_____09__37573),
       .Q (_________37591));
  nor2s1 ____0__497778(.DIN1 (_________37495), .DIN2 (_________37589),
       .Q (_________37590));
  and2s1 _______497779(.DIN1 (_________37822), .DIN2 (_________37540),
       .Q (_________37588));
  and2s1 _____0_497780(.DIN1 (_________37617), .DIN2 (_________37598),
       .Q (_________37647));
  nor2s1 _____0_497781(.DIN1 (_________37587), .DIN2 (_________37617),
       .Q (_________37618));
  nor2s1 _____0_497782(.DIN1 (_________37258), .DIN2 (_________37597),
       .Q (____00___38042));
  dffacs1 _______________________________________________497783(.CLRB
       (reset), .CLK (clk), .DIN (_____9___37557), .Q (___0_0___40466));
  dffacs1 _______________________________________________497784(.CLRB
       (reset), .CLK (clk), .DIN (_________37543), .Q
       (_____________________________________________21900));
  xor2s1 ____00_497785(.DIN1 (_____9___37558), .DIN2 (____9_0__38941),
       .Q (_________37586));
  nor2s1 ____9_497786(.DIN1 (______0__37584), .DIN2 (______9__37583),
       .Q (_________37585));
  nnd2s1 ____9__497787(.DIN1 (_________37527), .DIN2 (_________37199),
       .Q (_________37582));
  nor2s1 ____0_497788(.DIN1 (_________37530), .DIN2 (______0__35755),
       .Q (_________37581));
  xor2s1 ____00_497789(.DIN1 (_________37579), .DIN2 (___9_____39542),
       .Q (_________37580));
  xor2s1 ____0__497790(.DIN1
       (_________________________________________0___21856), .DIN2
       (_____0___37569), .Q (_________37578));
  nnd2s1 ____0__497791(.DIN1 (_________37576), .DIN2 (_________37520),
       .Q (_________37577));
  nnd2s1 ____0__497792(.DIN1 (____09__23606), .DIN2 (______9__37515),
       .Q (_________37575));
  nor2s1 ____0__497793(.DIN1 (___0_____40623), .DIN2 (______9__37525),
       .Q (______0__37633));
  nor2s1 ____9__497794(.DIN1 (____0____40766), .DIN2 (_________37519),
       .Q (_________37638));
  dffacs1 _____________________________________________9_497795(.CLRB
       (reset), .CLK (clk), .DIN (_________37518), .Q
       (_________________________________________9___21855));
  nnd2s1 ____0__497796(.DIN1 (_____09__37573), .DIN2 (_________35177),
       .Q (______0__37574));
  nor2s1 ____0__497797(.DIN1 (______0__37929), .DIN2 (_________37514),
       .Q (_____0___37572));
  nor2s1 ____0__497798(.DIN1 (______0__37516), .DIN2 (_________37744),
       .Q (_____0___37571));
  xnr2s1 ____0__497799(.DIN1 (_____0___37569), .DIN2 (_________22043),
       .Q (_____0___37570));
  xor2s1 ____0__497800(.DIN1 (_________37552), .DIN2 (_________37551),
       .Q (_____0___37568));
  or2s1 ____0__497801(.DIN1 (___00____39929), .DIN2 (_________37523),
       .Q (_____0___37567));
  xor2s1 _______497802(.DIN1 (_________37501), .DIN2 (________23821),
       .Q (_____00__37566));
  dffacs1 _______________________________________________497803(.CLRB
       (reset), .CLK (clk), .DIN (_________37512), .Q (_________22019));
  dffacs1 _______________________________________________497804(.CLRB
       (reset), .CLK (clk), .DIN (_________37524), .QN
       (___0_____40522));
  nor2s1 ____0__497805(.DIN1 (_____9___37564), .DIN2 (_____9___37563),
       .Q (_____99__37565));
  nnd2s1 ____99_497806(.DIN1 (_________37509), .DIN2 (___9__9__39659),
       .Q (_____9___37562));
  nor2s1 ____0_497807(.DIN1 (___0_____40623), .DIN2
       (_____________________________________9_______21879), .Q
       (_____9___37561));
  nnd2s1 ____0__497808(.DIN1
       (_____________________________________9_______21879), .DIN2
       (___0_____40623), .Q (_____9___37560));
  nnd2s1 ____0__497809(.DIN1 (_____9___37558), .DIN2 (_________22019),
       .Q (_____9___37559));
  nnd2s1 ____0__497810(.DIN1 (_________37499), .DIN2 (_____9___36996),
       .Q (_____9___37557));
  nor2s1 ____0__497811(.DIN1
       (_____________________________________9_______21879), .DIN2
       (______9__37555), .Q (_____90__37556));
  nnd2s1 ____0__497812(.DIN1 (______9__37555), .DIN2
       (_____________________________________9_______21879), .Q
       (_________37554));
  nor2s1 ____0__497813(.DIN1 (_________37552), .DIN2 (_________37551),
       .Q (_________37553));
  nor2s1 ____0__497814(.DIN1 (____0_0__37159), .DIN2 (_________37500),
       .Q (_________37550));
  or2s1 ____0__497815(.DIN1 (______9__37506), .DIN2 (_____0___36916),
       .Q (_________37549));
  and2s1 ____0__497816(.DIN1 (______0__37498), .DIN2 (_________37547),
       .Q (_________37548));
  nnd2s1 ____0__497817(.DIN1 (_________37551), .DIN2 (_____0___36547),
       .Q (______0__37546));
  nor2s1 ____0__497818(.DIN1 (_________37521), .DIN2 (_________37508),
       .Q (_________37608));
  xor2s1 ____0__497819(.DIN1 (______0__37478), .DIN2 (_____0___37475),
       .Q (_________37637));
  nor2s1 _______497820(.DIN1 (_________37621), .DIN2 (_________37534),
       .Q (______9__37545));
  nnd2s1 ____09_497821(.DIN1 (______0__37536), .DIN2 (_________37614),
       .Q (_________37544));
  nnd2s1 ____09_497822(.DIN1 (_____9__27279), .DIN2 (_________37503),
       .Q (_________37543));
  xor2s1 ____09_497823(.DIN1 (_________37541), .DIN2 (_________37494),
       .Q (_________37542));
  or2s1 _______497824(.DIN1
       (______________________________________0_____), .DIN2
       (___0__0__40441), .Q (_________37540));
  nnd2s1 _______497825(.DIN1 (_________37538), .DIN2 (___0__0__40441),
       .Q (_________37539));
  nor2s1 ____09_497826(.DIN1 (_________33729), .DIN2 (______0__37536),
       .Q (_________37537));
  nor2s1 _______497827(.DIN1 (_________37534), .DIN2 (_________37533),
       .Q (______9__37535));
  nor2s1 ____497828(.DIN1 (_________37614), .DIN2 (______0__37536), .Q
       (_________37532));
  nor2s1 _____0_497829(.DIN1 (______9__37458), .DIN2 (______9__37497),
       .Q (_________37589));
  xor2s1 _____0_497830(.DIN1 (_________37481), .DIN2 (_________37893),
       .Q (_________37602));
  nnd2s1 _______497831(.DIN1 (___0__0__40441), .DIN2
       (______________________________________0_____), .Q
       (_________37822));
  dffacs1 _______________________________________________497832(.CLRB
       (reset), .CLK (clk), .DIN (_________37505), .QN
       (_________22041));
  dffacs1 _______________________________________________497833(.CLRB
       (reset), .CLK (clk), .DIN (_________37511), .Q
       (_____________________________________________21940));
  nb1s1 _______497834(.DIN (_________37531), .Q (_________37617));
  hi1s1 _______497835(.DIN (_________37531), .Q (_________37597));
  nor2s1 ____0__497836(.DIN1 (______0__37488), .DIN2 (_________37223),
       .Q (_________37530));
  nnd2s1 ____0__497837(.DIN1 (______0__37526), .DIN2 (_________37528),
       .Q (_________37529));
  nor2s1 ____0__497838(.DIN1 (_________22019), .DIN2 (______0__37526),
       .Q (_________37527));
  hi1s1 ____0_497839(.DIN
       (_____________________________________9_______21879), .Q
       (______9__37525));
  nnd2s1 ____0__497840(.DIN1 (_________37482), .DIN2 (_________37504),
       .Q (_________37524));
  nor2s1 ____0__497841(.DIN1 (_____9___37365), .DIN2 (_________37491),
       .Q (_________37523));
  nor2s1 ____0__497842(.DIN1 (______9__37487), .DIN2 (_________37521),
       .Q (_________37522));
  xor2s1 ____0__497843(.DIN1 (_______________22074), .DIN2
       (___0_0___40467), .Q (_________37520));
  nor2s1 ____0__497844(.DIN1 (___0__9__40158), .DIN2 (_________37489),
       .Q (_________37519));
  nor2s1 ____00_497845(.DIN1 (_________37510), .DIN2 (_________37502),
       .Q (______9__37583));
  nnd2s1 ____0__497846(.DIN1 (____9____37035), .DIN2 (_________37483),
       .Q (_________37518));
  nnd2s1 ____0_497847(.DIN1 (_________37513), .DIN2 (___00____39929),
       .Q (_________37517));
  xor2s1 ____09_497848(.DIN1 (___0_____40442), .DIN2 (___99__22271), .Q
       (______0__37516));
  xor2s1 ____09_497849(.DIN1 (___0_____40442), .DIN2
       (______________________________________0______21887), .Q
       (______9__37515));
  nor2s1 _____497850(.DIN1 (_________37485), .DIN2 (_________37513), .Q
       (_________37514));
  nnd2s1 _______497851(.DIN1 (_____0___37473), .DIN2 (______0__37731),
       .Q (_________37512));
  xor2s1 _______497852(.DIN1 (_________37453), .DIN2 (___9_____39206),
       .Q (_________37531));
  nor2s1 _______497853(.DIN1 (_____00__35103), .DIN2 (_________37480),
       .Q (_____09__37573));
  nor2s1 _____0_497854(.DIN1 (_____09__37477), .DIN2 (_____0___37476),
       .Q (_________37924));
  dffacs1 _______________________________________________497855(.CLRB
       (reset), .CLK (clk), .DIN (_________37490), .Q (___0_____40506));
  nnd2s1 ____9_497856(.DIN1 (_____9___37465), .DIN2 (________27134), .Q
       (_________37511));
  xor2s1 ____0_497857(.DIN1 (_________37447), .DIN2 (_____00__37468),
       .Q (_________37509));
  and2s1 ____0__497858(.DIN1 (_________37486), .DIN2 (______0__37507),
       .Q (_________37508));
  nor2s1 _______497859(.DIN1 (_____9___37461), .DIN2 (_____0___33165),
       .Q (______9__37506));
  nnd2s1 _______497860(.DIN1 (_____9___37462), .DIN2 (_________37504),
       .Q (_________37505));
  nnd2s1 ______497861(.DIN1 (__9_9___29888), .DIN2 (___0_____40442), .Q
       (_________37503));
  nor2s1 ______497862(.DIN1 (___0_0___40467), .DIN2
       (_______________22076), .Q (_____9___37563));
  nnd2s1 ____0_497863(.DIN1 (_____0___37469), .DIN2 (_________37427),
       .Q (_________37579));
  hi1s1 ____0__497864(.DIN (______0__37526), .Q (_____9___37558));
  and2s1 _______497865(.DIN1 (_______________22076), .DIN2
       (___0_0___40467), .Q (_____9___37564));
  dffacs1 _________________________________________9_____497866(.CLRB
       (reset), .CLK (clk), .DIN (_____0___37470), .Q
       (_____________________________________9_______21879));
  xor2s1 _______497867(.DIN1 (_________37441), .DIN2 (_________37621),
       .Q (_________37501));
  xor2s1 _______497868(.DIN1 (_____0___35104), .DIN2 (_________37479),
       .Q (_________37500));
  nor2s1 _______497869(.DIN1 (________27223), .DIN2 (_____99__37467),
       .Q (_________37499));
  nnd2s1 _______497870(.DIN1 (_____9___37460), .DIN2 (______9__37334),
       .Q (______0__37498));
  and2s1 _______497871(.DIN1 (_________37496), .DIN2 (_________37457),
       .Q (______9__37497));
  nor2s1 _______497872(.DIN1 (_________37494), .DIN2 (_________37492),
       .Q (_________37495));
  or2s1 _______497873(.DIN1 (___0_0___40467), .DIN2
       (_______________22074), .Q (_____0___37569));
  and2s1 _______497874(.DIN1 (_________37493), .DIN2
       (_____________________________________________21770), .Q
       (_________37534));
  nor2s1 _______497875(.DIN1
       (_____________________________________________21770), .DIN2
       (_________37493), .Q (_________37533));
  nnd2s1 _______497876(.DIN1 (_________37492), .DIN2 (_________37494),
       .Q (______0__37536));
  dffacs1 __________________________________________0__9_(.CLRB
       (reset), .CLK (clk), .DIN (_________37455), .QN
       (___0__0__40441));
  nnd2s1 _______497877(.DIN1 (_____0___37471), .DIN2 (_________37418),
       .Q (_________37551));
  dffacs1 _______________________________________________497878(.CLRB
       (reset), .CLK (clk), .DIN (_________37451), .Q
       (_____________________________________________21784));
  nor2s1 _______497879(.DIN1 (_____9___37364), .DIN2 (_________37484),
       .Q (_________37491));
  or2s1 ____0_497880(.DIN1 (____0____38052), .DIN2 (_________37445), .Q
       (_________37490));
  nor2s1 ____0__497881(.DIN1 (_________37396), .DIN2 (_________37448),
       .Q (_________37489));
  xor2s1 _______497882(.DIN1 (_________37409), .DIN2 (________22660),
       .Q (______0__37488));
  hi1s1 _____0_497883(.DIN (_________37486), .Q (______9__37487));
  nor2s1 ______497884(.DIN1 (_____0___37472), .DIN2 (_________37484),
       .Q (_________37485));
  nnd2s1 ______497885(.DIN1 (___9____25039), .DIN2 (_________37443), .Q
       (_________37483));
  nor2s1 _______497886(.DIN1 (_________37442), .DIN2 (____0____36240),
       .Q (_________37482));
  nnd2s1 _______497887(.DIN1 (_________37446), .DIN2 (______0__37198),
       .Q (_________37502));
  xor2s1 ____0__497888(.DIN1 (______0__37430), .DIN2 (_________37386),
       .Q (_________37510));
  xor2s1 _____0_497889(.DIN1 (_________37421), .DIN2 (____0____37153),
       .Q (______0__37526));
  nnd2s1 ______497890(.DIN1 (_________37433), .DIN2 (______0__37382),
       .Q (_________37481));
  nor2s1 _______497891(.DIN1 (_____99__35102), .DIN2 (_________37479),
       .Q (_________37480));
  nor2s1 _______497892(.DIN1 (_____0___37474), .DIN2 (_____09__37477),
       .Q (______0__37478));
  nor2s1 _______497893(.DIN1 (_____0___37475), .DIN2 (_____0___37474),
       .Q (_____0___37476));
  nor2s1 _______497894(.DIN1 (___99___26048), .DIN2 (_________37437),
       .Q (_____0___37473));
  and2s1 _______497895(.DIN1 (_________37484), .DIN2 (_____0___37472),
       .Q (_________37513));
  hi1s1 ______497896(.DIN (_________37492), .Q (_________37541));
  nor2s1 _______497897(.DIN1 (______0__37440), .DIN2 (_________37435),
       .Q (____0____38071));
  dffacs1 _______________________________________________497898(.CLRB
       (reset), .CLK (clk), .DIN (______9__37439), .Q
       (_____________________________________________21843));
  dffacs1 ______________________________________497899(.CLRB (reset),
       .CLK (clk), .DIN (_________37444), .QN (___0_____40588));
  dffacs1 __________________497900(.CLRB (reset), .CLK (clk), .DIN
       (______9__37449), .QN (_______________22073));
  nnd2s1 _______497901(.DIN1 (_________37417), .DIN2 (_________37547),
       .Q (_____0___37471));
  nnd2s1 _______497902(.DIN1 (_________37423), .DIN2 (___09___28827),
       .Q (_____0___37470));
  or2s1 _______497903(.DIN1 (_________37425), .DIN2 (_____00__37468),
       .Q (_____0___37469));
  nor2s1 _______497904(.DIN1 (____0____37165), .DIN2 (_________37403),
       .Q (_____99__37467));
  nnd2s1 _______497905(.DIN1 (_________37422), .DIN2 (_________37834),
       .Q (_____9___37466));
  nor2s1 ____0__497906(.DIN1 (___9____26888), .DIN2 (______0__37420),
       .Q (_____9___37465));
  nnd2s1 ______497907(.DIN1 (_________37407), .DIN2 (_____9___37752),
       .Q (_____9___37464));
  nor2s1 _______497908(.DIN1
       (_____________________________________________21812), .DIN2
       (_____9___37463), .Q (_________37521));
  nnd2s1 ______497909(.DIN1 (_____9___37463), .DIN2
       (_____________________________________________21812), .Q
       (_________37486));
  dffacs1 __________________________________________0____497910(.CLRB
       (reset), .CLK (clk), .DIN (_________37404), .QN
       (___0_____40442));
  dffacs1 _______________________________________________497911(.CLRB
       (reset), .CLK (clk), .DIN (_________37406), .Q (___0_0___40467));
  nor2s1 _______497912(.DIN1 (_________37415), .DIN2 (_____9___36624),
       .Q (_____9___37462));
  xor2s1 _____497913(.DIN1
       (_____________________________________________21910), .DIN2
       (___0_____40614), .Q (_____9___37461));
  nnd2s1 _____9_497914(.DIN1 (_____90__37459), .DIN2 (_________36398),
       .Q (_____9___37460));
  nor2s1 _____9_497915(.DIN1 (_________37352), .DIN2 (_____90__37459),
       .Q (______9__37458));
  or2s1 _____9_497916(.DIN1 (_________37456), .DIN2 (_________37431),
       .Q (_________37457));
  nnd2s1 ______497917(.DIN1 (______9__37410), .DIN2 (_________37454),
       .Q (_________37455));
  xor2s1 _______497918(.DIN1 (_____0___37377), .DIN2 (_________37452),
       .Q (_________37453));
  nnd2s1 ______497919(.DIN1 (_________37408), .DIN2 (________27136), .Q
       (_________37451));
  xor2s1 _______497920(.DIN1 (_____0___37378), .DIN2 (_________38456),
       .Q (_________37493));
  xor2s1 _____0_497921(.DIN1 (_____0___37379), .DIN2 (____0____38106),
       .Q (_________37496));
  dffacs1 _______________________________________________497922(.CLRB
       (reset), .CLK (clk), .DIN (_________37428), .QN
       (___0_____40486));
  xnr2s1 _____0_497923(.DIN1 (_________36858), .DIN2 (______0__37450),
       .Q (_________37492));
  nnd2s1 _______497924(.DIN1 (______0__37391), .DIN2 (__9_____29964),
       .Q (______9__37449));
  nnd2s1 _______497925(.DIN1 (_________37399), .DIN2 (_________37387),
       .Q (_________37448));
  xor2s1 ______497926(.DIN1
       (_______________________________________________________________0__21998),
       .DIN2 (_________37426), .Q (_________37447));
  nor2s1 _______497927(.DIN1 (_________37200), .DIN2 (______9__37390),
       .Q (_________37446));
  nnd2s1 _______497928(.DIN1 (______9__37400), .DIN2 (___9____25100),
       .Q (_________37445));
  nnd2s1 _______497929(.DIN1 (______9__37652), .DIN2 (_________37397),
       .Q (_________37444));
  xor2s1 ______497930(.DIN1 (___0_0___40468), .DIN2 (_________36762),
       .Q (_________37443));
  nor2s1 _______497931(.DIN1 (_________37388), .DIN2 (_________37414),
       .Q (_________37442));
  dffacs1 _______________________________________________497932(.CLRB
       (reset), .CLK (clk), .DIN (_________37394), .Q
       (_____________________________________________21812));
  nor2s1 ______497933(.DIN1 (_____9___37271), .DIN2 (_________37393),
       .Q (_________37484));
  nor2s1 _____0_497934(.DIN1 (______0__37440), .DIN2 (_________37434),
       .Q (_________37441));
  nnd2s1 _______497935(.DIN1 (_________37385), .DIN2 (_____9__22978),
       .Q (______9__37439));
  and2s1 _______497936(.DIN1 (___09____40676), .DIN2 (_________38249),
       .Q (_________37438));
  nor2s1 ______497937(.DIN1 (___0_____40614), .DIN2 (_________38377),
       .Q (_________37437));
  xor2s1 _______497938(.DIN1 (______0__37354), .DIN2 (___9_____39461),
       .Q (_________37436));
  nor2s1 _____497939(.DIN1 (_________37621), .DIN2 (_________37434), .Q
       (_________37435));
  or2s1 _____0_497940(.DIN1 (_____0___37380), .DIN2 (____0_0__36219),
       .Q (_________37433));
  nor2s1 _______497941(.DIN1 (_________34947), .DIN2 (_________37384),
       .Q (_________37479));
  nnd2s1 _______497942(.DIN1 (___0_____40614), .DIN2 (____9___25676),
       .Q (_____0___37668));
  nor2s1 _____497943(.DIN1 (____9____37066), .DIN2 (_________37432), .Q
       (_____0___37474));
  dffacs1 _______________________________________________497944(.CLRB
       (reset), .CLK (clk), .DIN (_________37395), .QN
       (___0_____40485));
  and2s1 _______497945(.DIN1 (_________37402), .DIN2 (_________37547),
       .Q (_________37431));
  xor2s1 _______497946(.DIN1 (_________37398), .DIN2 (______9__37429),
       .Q (______0__37430));
  nnd2s1 ______497947(.DIN1 (_____9___37370), .DIN2 (____0____37173),
       .Q (_________37428));
  or2s1 _______497948(.DIN1 (_________37424), .DIN2 (_________37426),
       .Q (_________37427));
  and2s1 _______497949(.DIN1 (_________37426), .DIN2 (_________37424),
       .Q (_________37425));
  nnd2s1 _______497950(.DIN1 (_____99__37372), .DIN2 (______9__37555),
       .Q (_________37423));
  xor2s1 _____9_497951(.DIN1 (_____9___37273), .DIN2 (_________37392),
       .Q (_________37422));
  xor2s1 _____9_497952(.DIN1 (____0____37154), .DIN2 (_________37389),
       .Q (_________37421));
  nor2s1 ____0__497953(.DIN1 (______9__37419), .DIN2 (_____0___37374),
       .Q (______0__37420));
  nnd2s1 ______497954(.DIN1 (_____9___37366), .DIN2 (______9__37353),
       .Q (_________37418));
  nnd2s1 _____497955(.DIN1 (_____9___37368), .DIN2 (____0____36265), .Q
       (_________37417));
  nor2s1 _____9_497956(.DIN1 (_________37326), .DIN2 (_____00__37373),
       .Q (_____9___37463));
  nor2s1 _____9_497957(.DIN1 (____9____37067), .DIN2 (_________37416),
       .Q (_____09__37477));
  nor2s1 ______497958(.DIN1 (______9__37362), .DIN2 (_________37414),
       .Q (_________37415));
  nnd2s1 _______497959(.DIN1 (_________37412), .DIN2 (___0_0___40468),
       .Q (_________37413));
  nor2s1 ______497960(.DIN1 (_________37412), .DIN2 (___0_0___40468),
       .Q (______0__37411));
  nor2s1 _____9_497961(.DIN1 (____9___25853), .DIN2 (_________37359),
       .Q (______9__37410));
  and2s1 _______497962(.DIN1 (___0_0___40468), .DIN2 (___0_____40525),
       .Q (_________37409));
  nnd2s1 _______497963(.DIN1 (_________37355), .DIN2 (______0__37872),
       .Q (_________37408));
  xor2s1 _______497964(.DIN1 (______9__34948), .DIN2 (_________37383),
       .Q (_________37407));
  nnd2s1 _______497965(.DIN1 (_____9___37369), .DIN2 (_________37405),
       .Q (_________37406));
  nnd2s1 _______497966(.DIN1 (_________37360), .DIN2 (______9__38496),
       .Q (_________37404));
  xor2s1 _______497967(.DIN1 (____0____36221), .DIN2 (_____09__37381),
       .Q (_________37403));
  nor2s1 ______497968(.DIN1 (_________37547), .DIN2 (_________37402),
       .Q (_________37456));
  hi1s1 _______497969(.DIN (______0__37401), .Q (_____90__37459));
  dffacs1 _______________________________________________497970(.CLRB
       (reset), .CLK (clk), .DIN (_____90__37363), .Q
       (_____________________________________________21770));
  dffacs1 _______________________________________________497971(.CLRB
       (reset), .CLK (clk), .DIN (_________37357), .QN
       (_____________________________________________21783));
  dffacs1 _____________________________________________9_497972(.CLRB
       (reset), .CLK (clk), .DIN (_________37358), .Q
       (_________________________________________9_));
  nnd2s1 _______497973(.DIN1 (_________37349), .DIN2 (____9____38001),
       .Q (______9__37400));
  or2s1 ______497974(.DIN1 (_____9___36725), .DIN2 (_________37398), .Q
       (_________37399));
  and2s1 _____0_497975(.DIN1 (_________37346), .DIN2 (________25668),
       .Q (_________37397));
  nor2s1 _____0_497976(.DIN1 (___90____39055), .DIN2 (_________37348),
       .Q (_________37396));
  nnd2s1 _____0_497977(.DIN1 (_________37342), .DIN2 (____0____37147),
       .Q (_________37395));
  nnd2s1 _______497978(.DIN1 (_________37343), .DIN2 (______9__36755),
       .Q (_________37394));
  nor2s1 _______497979(.DIN1 (_____9___37272), .DIN2 (_________37392),
       .Q (_________37393));
  nnd2s1 _______497980(.DIN1 (__9_9___30364), .DIN2 (______9__37344),
       .Q (______0__37391));
  nor2s1 _______497981(.DIN1 (____0____37155), .DIN2 (_________37389),
       .Q (______9__37390));
  xnr2s1 _______497982(.DIN1 (_________37361), .DIN2 (_________22041),
       .Q (_________37388));
  nnd2s1 _______497983(.DIN1 (_________37356), .DIN2 (_________37386),
       .Q (_________37387));
  hi1s1 _______497984(.DIN (_________37416), .Q (_________37432));
  or2s1 _______497985(.DIN1 (_____9___37656), .DIN2 (_________37332),
       .Q (_________37385));
  nor2s1 _______497986(.DIN1 (_________34946), .DIN2 (_________37383),
       .Q (_________37384));
  or2s1 _______497987(.DIN1
       (_____________________________________________21858), .DIN2
       (_____09__37381), .Q (______0__37382));
  and2s1 _______497988(.DIN1 (_____09__37381), .DIN2
       (_____________________________________________21858), .Q
       (_____0___37380));
  nor2s1 _______497989(.DIN1 (_____00__37189), .DIN2 (_________37340),
       .Q (_____0___37379));
  nnd2s1 _____0_497990(.DIN1 (_________37337), .DIN2 (_____0___35382),
       .Q (_____0___37378));
  xor2s1 _______497991(.DIN1 (_________37306), .DIN2
       (______________22106), .Q (_____0___37377));
  xor2s1 ______497992(.DIN1 (_________37308), .DIN2 (_________37233),
       .Q (______0__37450));
  xor2s1 ______497993(.DIN1 (_____0___37376), .DIN2 (___0_____40308),
       .Q (______0__37401));
  and2s1 _______497994(.DIN1 (_____0___37375), .DIN2 (___0_____40549),
       .Q (_________37434));
  nor2s1 _______497995(.DIN1 (___0_____40549), .DIN2 (_____0___37375),
       .Q (______0__37440));
  dffacs1 _______________________________________________497996(.CLRB
       (reset), .CLK (clk), .DIN (______0__37335), .QN
       (___0_____40614));
  xor2s1 ______497997(.DIN1 (_________37329), .DIN2 (_________37301),
       .Q (_____0___37374));
  nor2s1 _______497998(.DIN1 (_________37327), .DIN2 (_____9___36629),
       .Q (_____00__37373));
  xor2s1 _______497999(.DIN1 (_________37303), .DIN2 (_________37296),
       .Q (_____99__37372));
  xor2s1 _______498000(.DIN1
       (_________________________________________________________________22001),
       .DIN2 (_________37350), .Q (_____9___37371));
  nor2s1 _______498001(.DIN1 (_________37328), .DIN2 (_________36489),
       .Q (_____9___37370));
  nor2s1 _______498002(.DIN1 (____9___29546), .DIN2 (_________37318),
       .Q (_____9___37369));
  nnd2s1 _______498003(.DIN1 (_____9___37367), .DIN2 (____0____36266),
       .Q (_____9___37368));
  nor2s1 _______498004(.DIN1 (______9__36295), .DIN2 (_____9___37367),
       .Q (_____9___37366));
  nor2s1 _______498005(.DIN1 (_____9___37365), .DIN2 (_____9___37364),
       .Q (_____0___37472));
  nor2s1 _____498006(.DIN1 (_____0___37196), .DIN2 (_________37330), .Q
       (_____00__37468));
  xor2s1 _______498007(.DIN1 (_____9___37274), .DIN2 (_________37339),
       .Q (_________37416));
  xor2s1 ______498008(.DIN1 (______9__37294), .DIN2 (_________37299),
       .Q (_________37426));
  dffacs1 _______________________________________________498009(.CLRB
       (reset), .CLK (clk), .DIN (______9__37324), .QN
       (___0__0__40431));
  nnd2s1 ______498010(.DIN1 (_________37312), .DIN2 (________27436), .Q
       (_____90__37363));
  and2s1 _______498011(.DIN1 (_________37331), .DIN2 (_________37361),
       .Q (______9__37362));
  nor2s1 _______498012(.DIN1 (________23379), .DIN2 (_________37316),
       .Q (_________37360));
  nor2s1 ______498013(.DIN1 (_________36955), .DIN2 (_________37310),
       .Q (_________37359));
  nnd2s1 _____9_498014(.DIN1 (_________37313), .DIN2 (_____9__26340),
       .Q (_________37358));
  nnd2s1 _____9_498015(.DIN1 (_________37319), .DIN2 (_________37221),
       .Q (_________37357));
  xor2s1 _______498016(.DIN1 (_____0___35383), .DIN2 (_________37336),
       .Q (_________37355));
  xor2s1 _______498017(.DIN1 (_____0___37281), .DIN2 (______9__37353),
       .Q (______0__37354));
  nor2s1 _______498018(.DIN1 (______9__37304), .DIN2 (_________37307),
       .Q (_________37866));
  xor2s1 _______498019(.DIN1 (_________37288), .DIN2 (________22381),
       .Q (_________37841));
  nnd2s1 _______498020(.DIN1 (_____0___37376), .DIN2 (_________37352),
       .Q (_________37402));
  dffacs1 _____________________________________________0_498021(.CLRB
       (reset), .CLK (clk), .DIN (_________37323), .QN
       (___0_0___40468));
  or2s1 _______498022(.DIN1
       (_________________________________________________________________22001),
       .DIN2 (_________37350), .Q (_________37351));
  xor2s1 ______498023(.DIN1 (___0_____40518), .DIN2 (_____9___36630),
       .Q (_________37349));
  or2s1 ______498024(.DIN1 (_________37341), .DIN2 (_________37350), .Q
       (_________37348));
  nnd2s1 _______498025(.DIN1 (_________37350), .DIN2
       (_________________________________________________________________22001),
       .Q (_________37347));
  nnd2s1 _______498026(.DIN1 (______0__37345), .DIN2 (______0__37295),
       .Q (_________37346));
  xor2s1 ______498027(.DIN1 (___0_0___40469), .DIN2 (___0_____40522),
       .Q (______9__37344));
  nnd2s1 _______498028(.DIN1 (_________37291), .DIN2 (_________38576),
       .Q (_________37343));
  nor2s1 _______498029(.DIN1 (_________37290), .DIN2 (_____90__36535),
       .Q (_________37342));
  nor2s1 _______498030(.DIN1 (_________37302), .DIN2 (_________37298),
       .Q (_________37392));
  dffacs1 _______________________________________________498031(.CLRB
       (reset), .CLK (clk), .DIN (______0__37286), .Q (______));
  xor2s1 _______498032(.DIN1 (_________37289), .DIN2 (_________37341),
       .Q (_________37398));
  nor2s1 _______498033(.DIN1 (_____0___37190), .DIN2 (_________37339),
       .Q (_________37340));
  and2s1 _______498034(.DIN1 (____9____37972), .DIN2 (_________37616),
       .Q (_________37338));
  nnd2s1 _______498035(.DIN1 (_________37336), .DIN2 (_____0___35381),
       .Q (_________37337));
  or2s1 _____9_498036(.DIN1 (_________32956), .DIN2 (_________37287),
       .Q (______0__37335));
  nnd2s1 _______498037(.DIN1 (_________37333), .DIN2 (_________37352),
       .Q (______9__37334));
  xor2s1 ______498038(.DIN1 (_________37261), .DIN2 (___90____39001),
       .Q (_________37332));
  xor2s1 _______498039(.DIN1 (_________37265), .DIN2 (______9__35584),
       .Q (_________37383));
  nnd2s1 _______498040(.DIN1 (_________37350), .DIN2 (_________37341),
       .Q (_________37356));
  nor2s1 _____498041(.DIN1 (_________37292), .DIN2 (_________37300), .Q
       (_________37389));
  and2s1 _______498042(.DIN1 (_____09__37285), .DIN2 (____0_0__40770),
       .Q (_____0___37375));
  nor2s1 _____498043(.DIN1 (_________37246), .DIN2 (_____0___37282), .Q
       (_____09__37381));
  dffacs1 _______________________________________________498044(.CLRB
       (reset), .CLK (clk), .DIN (_____0___37284), .Q
       (______0___22056));
  or2s1 _____9_498045(.DIN1 (___0_0___40469), .DIN2 (_________37321),
       .Q (_________37331));
  and2s1 _______498046(.DIN1 (_____0___37278), .DIN2 (_________37329),
       .Q (_________37330));
  nor2s1 _______498047(.DIN1 (_____99__37275), .DIN2 (____9_0__37080),
       .Q (_________37328));
  and2s1 _______498048(.DIN1 (______0__37325), .DIN2 (___0_____40518),
       .Q (_________37327));
  nor2s1 _______498049(.DIN1 (___0_____40518), .DIN2 (______0__37325),
       .Q (_________37326));
  or2s1 _____0_498050(.DIN1 (_________37837), .DIN2 (_____9___37270),
       .Q (______9__37324));
  nnd2s1 _____498051(.DIN1 (_____9___37268), .DIN2 (_________37322), .Q
       (_________37323));
  nnd2s1 _____0_498052(.DIN1 (_________37321), .DIN2 (___0_0___40469),
       .Q (_________37361));
  nor2s1 _____0_498053(.DIN1 (___0_0___40469), .DIN2 (_________37320),
       .Q (_____9___37365));
  and2s1 _____0_498054(.DIN1 (_________37320), .DIN2 (___0_0___40469),
       .Q (_____9___37364));
  nnd2s1 _____0_498055(.DIN1 (_____9___37269), .DIN2 (______0__36394),
       .Q (_____9___37367));
  nnd2s1 _______498056(.DIN1 (_________37264), .DIN2 (____99___37096),
       .Q (_________37319));
  and2s1 _______498057(.DIN1 (_____90__37267), .DIN2 (_________37317),
       .Q (_________37318));
  and2s1 _______498058(.DIN1 (______9__37266), .DIN2 (_________37744),
       .Q (_________37316));
  and2s1 _______498059(.DIN1 (_____00__37276), .DIN2 (______9__37314),
       .Q (______0__37315));
  nnd2s1 _______498060(.DIN1 (_________37311), .DIN2 (_________38177),
       .Q (_________37313));
  nnd2s1 _______498061(.DIN1 (_________37311), .DIN2 (______0__37872),
       .Q (_________37312));
  nor2s1 _____498062(.DIN1 (_________37241), .DIN2 (_________37309), .Q
       (_________37310));
  xnr2s1 _______498063(.DIN1 (_________38306), .DIN2 (____0____40768),
       .Q (_________37308));
  nor2s1 _______498064(.DIN1 (______________22106), .DIN2
       (______0__37305), .Q (_________37307));
  nor2s1 _______498065(.DIN1 (______0__37305), .DIN2 (______9__37304),
       .Q (_________37306));
  hi1s1 _______498066(.DIN (_________37333), .Q (_____0___37376));
  dffacs1 ______________________________________498067(.CLRB (reset),
       .CLK (clk), .DIN (_____0___37279), .QN (_____________22080));
  nor2s1 _____0_498068(.DIN1 (_________37302), .DIN2 (_________37297),
       .Q (_________37303));
  nor2s1 _______498069(.DIN1 (_____0___37277), .DIN2 (_________37255),
       .Q (_________37301));
  nor2s1 _____9_498070(.DIN1 (_________37299), .DIN2 (_________37293),
       .Q (_________37300));
  nor2s1 _____9_498071(.DIN1 (_________37297), .DIN2 (_________37296),
       .Q (_________37298));
  nnd2s1 _____9_498072(.DIN1 (_________37252), .DIN2 (inData[2]), .Q
       (______0__37295));
  or2s1 ______498073(.DIN1 (_________37293), .DIN2 (_________37292), .Q
       (______9__37294));
  xor2s1 _______498074(.DIN1 (______0__36499), .DIN2 (____0____40772),
       .Q (_________37291));
  nor2s1 _______498075(.DIN1 (_________37251), .DIN2 (____9____37049),
       .Q (_________37290));
  xor2s1 _______498076(.DIN1 (______0__37222), .DIN2 (______0__41289),
       .Q (_________37333));
  dffacs1 _______________________________________________498077(.CLRB
       (reset), .CLK (clk), .DIN (_________37250), .QN
       (___0__9__40550));
  hi1s1 _______498078(.DIN (_________37289), .Q (_________37350));
  nor2s1 _______498079(.DIN1 (______0__34915), .DIN2 (_________37243),
       .Q (_________37288));
  nnd2s1 ______498080(.DIN1 (_________37253), .DIN2 (________24827), .Q
       (_________37287));
  nnd2s1 _______498081(.DIN1 (_________37249), .DIN2 (______9__38496),
       .Q (______0__37286));
  nnd2s1 _______498082(.DIN1 (_________37235), .DIN2 (_________37547),
       .Q (_____09__37285));
  nnd2s1 _______498083(.DIN1 (_________37237), .DIN2 (_____0___37283),
       .Q (_____0___37284));
  nor2s1 _______498084(.DIN1 (______0__37248), .DIN2 (_________36041),
       .Q (_____0___37282));
  nnd2s1 _______498085(.DIN1 (_________37236), .DIN2 (_________37238),
       .Q (_____0___37281));
  or2s1 _____0_498086(.DIN1 (________24683), .DIN2 (_________37769), .Q
       (_____0___37280));
  nor2s1 _____498087(.DIN1 (____0____35337), .DIN2 (______0__37257), .Q
       (_________37336));
  nor2s1 _______498088(.DIN1 (____00___37106), .DIN2 (_________37254),
       .Q (_________37339));
  nor2s1 _______498089(.DIN1 (_________37244), .DIN2 (_________37769),
       .Q (____9____37972));
  or2s1 _______498090(.DIN1 (____9___23688), .DIN2 (_________37228), .Q
       (_____0___37279));
  or2s1 _______498091(.DIN1 (_________37229), .DIN2 (_____0___37277),
       .Q (_____0___37278));
  xor2s1 _______498092(.DIN1 (_________37206), .DIN2 (_________34991),
       .Q (_____00__37276));
  xor2s1 _______498093(.DIN1 (___0__9__40500), .DIN2 (___0__0__40471),
       .Q (_____99__37275));
  xor2s1 ______498094(.DIN1 (_________37213), .DIN2 (___009___39979),
       .Q (_____9___37274));
  or2s1 ______498095(.DIN1 (_____9___37272), .DIN2 (_____9___37271), .Q
       (_____9___37273));
  nnd2s1 ______498096(.DIN1 (______9__37231), .DIN2 (________25880), .Q
       (_____9___37270));
  nnd2s1 _______498097(.DIN1 (____0____40772), .DIN2 (_____99__36366),
       .Q (_____9___37269));
  and2s1 _______498098(.DIN1 (_________37224), .DIN2 (__9_____29764),
       .Q (_____9___37268));
  xor2s1 _______498099(.DIN1 (______9__37214), .DIN2 (____0____40782),
       .Q (_________37289));
  dffacs1 _______________________________________________498100(.CLRB
       (reset), .CLK (clk), .DIN (_________37227), .QN
       (___0_____40518));
  dffacs1 _____________________________________________9_498101(.CLRB
       (reset), .CLK (clk), .DIN (_________37226), .QN
       (___0_0___40469));
  xor2s1 _______498102(.DIN1 (_________36042), .DIN2 (______9__37247),
       .Q (_____90__37267));
  xor2s1 _______498103(.DIN1 (_________37216), .DIN2 (____0_9__36267),
       .Q (______9__37266));
  nnd2s1 _______498104(.DIN1 (_________37220), .DIN2 (____09___37184),
       .Q (_________37265));
  xor2s1 _____0_498105(.DIN1 (______9__37256), .DIN2 (_________35428),
       .Q (_________37264));
  xor2s1 _____0_498106(.DIN1 (_________31820), .DIN2 (_________37262),
       .Q (_________37263));
  xor2s1 _____0_498107(.DIN1 (_________34955), .DIN2 (_________37242),
       .Q (_________37261));
  dffacs1 ________________498108(.CLRB (reset), .CLK (clk), .DIN
       (_________37201), .Q (outData[16]));
  nnd2s1 _______498109(.DIN1 (_________37218), .DIN2 (______0__37872),
       .Q (_________37260));
  nor2s1 _______498110(.DIN1 (_____________22081), .DIN2
       (_________37259), .Q (______9__37304));
  and2s1 _______498111(.DIN1 (_________37259), .DIN2
       (_____________22081), .Q (______0__37305));
  hi1s1 ______498112(.DIN (_________37258), .Q (_________37309));
  xor2s1 _______498113(.DIN1 (_________37203), .DIN2 (___0_____40308),
       .Q (_________37311));
  dffacs1 _______________________________________________498114(.CLRB
       (reset), .CLK (clk), .DIN (_________37219), .Q
       (__________22059));
  and2s1 _______498115(.DIN1 (______9__37256), .DIN2 (____0____35336),
       .Q (______0__37257));
  and2s1 _______498116(.DIN1 (_________37211), .DIN2 (___9_0___39619),
       .Q (_________37255));
  nor2s1 _____9_498117(.DIN1 (_________37210), .DIN2 (____0____40782),
       .Q (_________37254));
  nnd2s1 _____9_498118(.DIN1 (_________37207), .DIN2 (___99____39861),
       .Q (_________37253));
  xor2s1 _______498119(.DIN1 (_____________22080), .DIN2
       (___0_9___40458), .Q (_________37252));
  xor2s1 _______498120(.DIN1 (___0_09__40470), .DIN2 (___0_____40499),
       .Q (_________37251));
  nnd2s1 ______498121(.DIN1 (_________37212), .DIN2 (_____9___38319),
       .Q (_________37250));
  nor2s1 _______498122(.DIN1 (____90__24925), .DIN2 (_________37208),
       .Q (_________37249));
  nor2s1 _______498123(.DIN1 (_________37245), .DIN2 (______9__37247),
       .Q (______0__37248));
  and2s1 _______498124(.DIN1 (______9__37247), .DIN2 (_________37245),
       .Q (_________37246));
  dffacs1 _______________________________________________498125(.CLRB
       (reset), .CLK (clk), .DIN (_________37217), .QN
       (_____________________________________________21857));
  nor2s1 _______498126(.DIN1 (___0__0__40471), .DIN2
       (_______________22073), .Q (_________37297));
  nor2s1 ______498127(.DIN1 (____0____37176), .DIN2 (_________37215),
       .Q (_________37293));
  and2s1 _______498128(.DIN1 (_______________22073), .DIN2
       (___0__0__40471), .Q (_________37302));
  nor2s1 _______498129(.DIN1 (____9____37073), .DIN2 (_________37233),
       .Q (_________37244));
  nor2s1 _______498130(.DIN1 (_____9___34928), .DIN2 (_________37242),
       .Q (_________37243));
  nor2s1 _______498131(.DIN1 (_________37233), .DIN2 (_________37234),
       .Q (_________37241));
  nnd2s1 _______498132(.DIN1 (_________37233), .DIN2
       (______________________________________________21902), .Q
       (______9__37240));
  nor2s1 ______498133(.DIN1
       (______________________________________________21902), .DIN2
       (_________37233), .Q (_________37239));
  nnd2s1 _______498134(.DIN1 (_________37233), .DIN2 (______0__37232),
       .Q (_________37238));
  nor2s1 _______498135(.DIN1 (________28390), .DIN2 (______0__37205),
       .Q (_________37237));
  nnd2s1 _______498136(.DIN1 (_________37262), .DIN2 (____0____37161),
       .Q (_________37236));
  nnd2s1 _______498137(.DIN1 (_________37204), .DIN2 (____099__35378),
       .Q (_________37235));
  nnd2s1 _______498138(.DIN1 (_________37234), .DIN2 (_________37233),
       .Q (_________37258));
  nor2s1 _______498139(.DIN1 (______0__37232), .DIN2 (_________37262),
       .Q (_________37587));
  nnd2s1 ______498140(.DIN1 (____0____37162), .DIN2 (_________37262),
       .Q (_________37598));
  nor2s1 _______498141(.DIN1 (____9____37026), .DIN2 (_________37262),
       .Q (_________37769));
  nnd2s1 _______498142(.DIN1 (_____0___37194), .DIN2 (_________37230),
       .Q (______9__37231));
  and2s1 _______498143(.DIN1 (_________37225), .DIN2 (___9_0___39619),
       .Q (_________37229));
  nor2s1 _____9_498144(.DIN1 (___0_9___40458), .DIN2 (____9_9__37052),
       .Q (_________37228));
  or2s1 _______498145(.DIN1 (____0____38117), .DIN2 (_____0___37192),
       .Q (_________37227));
  nnd2s1 ______498146(.DIN1 (_____0___37191), .DIN2 (_________37504),
       .Q (_________37226));
  and2s1 _______498147(.DIN1
       (_______________________________________________________________________________________),
       .DIN2 (___0_09__40470), .Q (_____9___37272));
  nor2s1 _______498148(.DIN1 (___0_09__40470), .DIN2
       (_______________________________________________________________________________________),
       .Q (_____9___37271));
  nor2s1 ______498149(.DIN1 (____0____37177), .DIN2 (____0____40774),
       .Q (_________37292));
  nor2s1 _______498150(.DIN1 (___9_0___39619), .DIN2 (_________37225),
       .Q (_____0___37277));
  nnd2s1 _____0_498151(.DIN1 (_____0___37193), .DIN2 (_________37223),
       .Q (_________37224));
  xor2s1 ______498152(.DIN1 (____0_9__37158), .DIN2 (___09____40688),
       .Q (______0__37222));
  nnd2s1 _______498153(.DIN1 (____09__25318), .DIN2 (____09___37185),
       .Q (_________37221));
  or2s1 ______498154(.DIN1 (_________36680), .DIN2 (____09___37187), .Q
       (_________37220));
  nnd2s1 _______498155(.DIN1 (____09___37181), .DIN2 (_________38550),
       .Q (_________37219));
  xor2s1 _____9_498156(.DIN1 (_________35430), .DIN2 (____0____40776),
       .Q (_________37218));
  nor2s1 _____0_498157(.DIN1 (____0____37132), .DIN2 (____09___37182),
       .Q (_________37259));
  dffacs1 ______________________________________________498158(.CLRB
       (reset), .CLK (clk), .DIN (____09___37183), .QN (________));
  dffacs1 _______________________________________________498159(.CLRB
       (reset), .CLK (clk), .DIN (____090__37179), .QN
       (__________22061));
  nnd2s1 _______498160(.DIN1 (____0____37166), .DIN2 (__9_____30145),
       .Q (_________37217));
  nnd2s1 _______498161(.DIN1 (____0_9__37178), .DIN2 (____99___37094),
       .Q (_________37216));
  hi1s1 _____9_498162(.DIN (____0____40774), .Q (_________37215));
  nnd2s1 _____0_498163(.DIN1 (_________37209), .DIN2 (____0____37171),
       .Q (______9__37214));
  xor2s1 _____0_498164(.DIN1 (____909__36106), .DIN2 (______0__38467),
       .Q (_________37213));
  and2s1 _______498165(.DIN1 (____0_9__37168), .DIN2 (___0____24245),
       .Q (_________37212));
  xor2s1 _______498166(.DIN1
       (__________________________________________________________________21992),
       .DIN2 (_____0___37195), .Q (_________37211));
  and2s1 _______498167(.DIN1 (_________37209), .DIN2 (____0____37164),
       .Q (_________37210));
  nor2s1 _______498168(.DIN1 (___0__0__39993), .DIN2 (____0____37163),
       .Q (_________37208));
  xor2s1 _______498169(.DIN1 (____0____37141), .DIN2 (___9_____39372),
       .Q (_________37207));
  nnd2s1 _______498170(.DIN1 (____0____37170), .DIN2 (_________35800),
       .Q (______9__37247));
  dffacs1 _______________________________________________498171(.CLRB
       (reset), .CLK (clk), .DIN (____0____37174), .Q (___0__0__40471));
  xor2s1 ______498172(.DIN1 (____09___37186), .DIN2 (_________38395),
       .Q (_________37206));
  nnd2s1 _______498173(.DIN1 (____0____37160), .DIN2 (_____9__27362),
       .Q (______0__37205));
  nnd2s1 _______498174(.DIN1 (____0____40776), .DIN2 (_____00__35379),
       .Q (_________37204));
  xor2s1 _____0_498175(.DIN1 (________29292), .DIN2 (____0_0__37144),
       .Q (_________37203));
  hi1s1 _______498176(.DIN (_________37201), .Q (_________37233));
  xor2s1 _______498177(.DIN1 (____0_0__37134), .DIN2 (_________37202),
       .Q (______9__37256));
  xor2s1 _______498178(.DIN1 (____0_9__37133), .DIN2 (____9____38948),
       .Q (_________37242));
  dffacs1 _________________________________________9_____498179(.CLRB
       (reset), .CLK (clk), .DIN (____0____37175), .Q (___0_____40622));
  nb1s1 _____9_498180(.DIN (_________37201), .Q (_________37262));
  nor2s1 ______498181(.DIN1 (_________37199), .DIN2 (_____09__37197),
       .Q (_________37200));
  nnd2s1 ______498182(.DIN1 (_____09__37197), .DIN2 (_________37199),
       .Q (______0__37198));
  and2s1 _______498183(.DIN1 (_____0___37195), .DIN2
       (__________________________________________________________________21992),
       .Q (_____0___37196));
  xor2s1 _______498184(.DIN1 (____0____37130), .DIN2 (____0_0__40780),
       .Q (_____0___37194));
  xor2s1 _______498185(.DIN1 (_____90__35823), .DIN2 (____0_0__37169),
       .Q (_____0___37193));
  xor2s1 _____9_498186(.DIN1 (____0____37131), .DIN2 (___90_0__39025),
       .Q (_____0___37192));
  nor2s1 ______498187(.DIN1 (__9__9__29886), .DIN2 (____0____37152), .Q
       (_____0___37191));
  nnd2s1 ______498188(.DIN1 (____0____37150), .DIN2 (____0____37115),
       .Q (_________37329));
  dffacs1 _________________________________________9_____498189(.CLRB
       (reset), .CLK (clk), .DIN (____0_0__37151), .Q (___0_9___40458));
  or2s1 _______498190(.DIN1
       (__________________________________________________________________21992),
       .DIN2 (_____0___37195), .Q (_________37225));
  dffacs1 _______________________________________________498191(.CLRB
       (reset), .CLK (clk), .DIN (____0____37148), .QN
       (___0_09__40470));
  nor2s1 ______498192(.DIN1 (____099__37188), .DIN2 (______0__38467),
       .Q (_____0___37190));
  and2s1 _______498193(.DIN1 (______0__38467), .DIN2 (____099__37188),
       .Q (_____00__37189));
  nor2s1 _______498194(.DIN1
       (_____________________________________________21842), .DIN2
       (____09___37186), .Q (____09___37187));
  nor2s1 ______498195(.DIN1 (____0____37142), .DIN2 (________25930), .Q
       (____09___37185));
  nnd2s1 _______498196(.DIN1 (____09___37186), .DIN2
       (_____________________________________________21842), .Q
       (____09___37184));
  nnd2s1 _______498197(.DIN1 (____9____33373), .DIN2 (____0____37145),
       .Q (____09___37183));
  and2s1 _______498198(.DIN1 (____0____37146), .DIN2 (____9____38007),
       .Q (____09___37182));
  and2s1 ______498199(.DIN1 (____0____37136), .DIN2 (____09___37180),
       .Q (____09___37181));
  nnd2s1 _______498200(.DIN1 (____0____37140), .DIN2 (_________38253),
       .Q (____090__37179));
  hi1s1 _______498201(.DIN (____0_9__37178), .Q (_________37234));
  nor2s1 _______498202(.DIN1 (____9____36143), .DIN2 (____0____37138),
       .Q (____0____38069));
  xor2s1 _______498203(.DIN1 (___09____40686), .DIN2 (___0_____40650),
       .Q (_________37201));
  dffacs1 _______________________________________________498204(.CLRB
       (reset), .CLK (clk), .DIN (____0____37135), .QN
       (_____________________________________________21769));
  hi1s1 _____9_498205(.DIN (____0____37176), .Q (____0____37177));
  nnd2s1 _______498206(.DIN1 (____0____37128), .DIN2 (______9__37652),
       .Q (____0____37175));
  nnd2s1 ______498207(.DIN1 (____0____37127), .DIN2 (____0____37173),
       .Q (____0____37174));
  nor2s1 _______498208(.DIN1 (______0__37345), .DIN2 (____0____37126),
       .Q (____0____37172));
  or2s1 _______498209(.DIN1 (_____0___38422), .DIN2 (____0____37125),
       .Q (____0____37171));
  nnd2s1 _______498210(.DIN1 (_________35801), .DIN2 (____0_0__37169),
       .Q (____0____37170));
  nnd2s1 ______498211(.DIN1 (____0____37122), .DIN2 (____0____37167),
       .Q (____0_9__37168));
  or2s1 _____9_498212(.DIN1 (____0____37165), .DIN2 (____0_9__37123),
       .Q (____0____37166));
  or2s1 _____9_498213(.DIN1 (_____0___38422), .DIN2 (____0____37156),
       .Q (____0____37164));
  xor2s1 _____498214(.DIN1 (____9____36144), .DIN2 (____0____37137), .Q
       (____0____37163));
  xor2s1 _____0_498215(.DIN1 (____0____37161), .DIN2 (_________38203),
       .Q (____0____37162));
  or2s1 _______498216(.DIN1 (____0_0__37159), .DIN2 (____0____37119),
       .Q (____0____37160));
  nnd2s1 _____0_498217(.DIN1 (____00___37105), .DIN2 (____0____37121),
       .Q (____0_9__37158));
  dffacs1 _____________________________________________0_498218(.CLRB
       (reset), .CLK (clk), .DIN (____0_0__37124), .Q
       (_________________________________________0___21939));
  nnd2s1 _____0_498219(.DIN1 (____0____37156), .DIN2 (_____0___38422),
       .Q (_________37209));
  xor2s1 ______498220(.DIN1 (____000__37100), .DIN2 (______0__37673),
       .Q (____0_9__37178));
  dffacs1 _______________________________________________498221(.CLRB
       (reset), .CLK (clk), .DIN (____0____37120), .Q
       (_____________________________________________21842));
  and2s1 _____498222(.DIN1 (____0____37154), .DIN2 (____0____37153), .Q
       (____0____37155));
  nor2s1 _____9_498223(.DIN1 (_________41090), .DIN2 (____00___37107),
       .Q (____0____37152));
  nnd2s1 _______498224(.DIN1 (____0____37117), .DIN2 (______0__36932),
       .Q (____0_0__37151));
  nnd2s1 ______498225(.DIN1 (____0_0__37116), .DIN2 (____0____37129),
       .Q (____0____37150));
  nnd2s1 _______498226(.DIN1 (____0____37110), .DIN2 (____0____37147),
       .Q (____0____37148));
  or2s1 _______498227(.DIN1 (____0____37153), .DIN2 (____0____37154),
       .Q (_____09__37197));
  nor2s1 _______498228(.DIN1 (_________36887), .DIN2 (____0____37112),
       .Q (_________37296));
  xor2s1 _____498229(.DIN1 (____9____37084), .DIN2 (_________38650), .Q
       (____0____37176));
  xor2s1 _______498230(.DIN1 (____9____37083), .DIN2 (_________36952),
       .Q (_____0___37195));
  dffacs1 __________________________________________0____498231(.CLRB
       (reset), .CLK (clk), .DIN (____00___37103), .QN
       (______________________________________0______21886));
  xor2s1 _______498232(.DIN1 (____9____37074), .DIN2 (_____9___38512),
       .Q (______0__38467));
  nnd2s1 _______498233(.DIN1 (____9_9__37089), .DIN2 (___0____22301),
       .Q (____0____37146));
  nnd2s1 _______498234(.DIN1 (___9____25093), .DIN2 (____00___37104),
       .Q (____0____37145));
  xor2s1 _____9_498235(.DIN1 (____0____40778), .DIN2 (_________36087),
       .Q (____0_0__37144));
  and2s1 _______498236(.DIN1 (____999__37099), .DIN2 (_________37744),
       .Q (____0_9__37143));
  xor2s1 _______498237(.DIN1 (_______22212), .DIN2 (____9____37071), .Q
       (____0____37142));
  xor2s1 _______498238(.DIN1 (____9____37061), .DIN2 (____0_0__36201),
       .Q (____0____37141));
  nor2s1 _______498239(.DIN1 (____0____37139), .DIN2 (____99___37095),
       .Q (____0____37140));
  nor2s1 _______498240(.DIN1 (____9____36142), .DIN2 (____0____37137),
       .Q (____0____37138));
  and2s1 _______498241(.DIN1 (____99___37097), .DIN2 (____9___26225),
       .Q (____0____37136));
  nnd2s1 _______498242(.DIN1 (____990__37090), .DIN2 (_____0__27401),
       .Q (____0____37135));
  nor2s1 _______498243(.DIN1 (____9____37017), .DIN2 (____00___37101),
       .Q (____0_0__37134));
  nnd2s1 _______498244(.DIN1 (____99___37093), .DIN2 (_________35006),
       .Q (____0_9__37133));
  nor2s1 _______498245(.DIN1 (____9____38007), .DIN2 (____9____37087),
       .Q (____0____37132));
  nnd2s1 ______498246(.DIN1 (____0_0__37109), .DIN2 (_________34787),
       .Q (____09___37186));
  dffacs1 ______________________________________________498247(.CLRB
       (reset), .CLK (clk), .DIN (____99___37091), .QN
       (____________________________________________21790));
  xor2s1 _____498248(.DIN1 (_____0___36284), .DIN2 (____00___37102), .Q
       (____0____37131));
  xor2s1 _______498249(.DIN1 (________27669), .DIN2 (____0____37129),
       .Q (____0____37130));
  and2s1 _______498250(.DIN1 (____9____37082), .DIN2 (________26244),
       .Q (____0____37128));
  nor2s1 _______498251(.DIN1 (__9_____30166), .DIN2 (____9____37081),
       .Q (____0____37127));
  xor2s1 _____9_498252(.DIN1 (______9__36888), .DIN2 (____0____37111),
       .Q (____0____37126));
  xor2s1 _____0_498253(.DIN1 (____0____37118), .DIN2 (_________38350),
       .Q (____0____37125));
  nnd2s1 _______498254(.DIN1 (____9_9__37079), .DIN2 (________28136),
       .Q (____0_0__37124));
  nnd2s1 _______498255(.DIN1 (____9____37078), .DIN2 (______0__35701),
       .Q (____0_0__37169));
  dffacs1 _______________________________________________498256(.CLRB
       (reset), .CLK (clk), .DIN (____9_0__37070), .QN
       (___0_____40537));
  xor2s1 ______498257(.DIN1 (_________34822), .DIN2 (____009__37108),
       .Q (____0_9__37123));
  xor2s1 _______498258(.DIN1 (____9____37044), .DIN2 (____0_0__40790),
       .Q (____0____37122));
  xor2s1 _______498259(.DIN1 (____9____37038), .DIN2 (_________38372),
       .Q (____0____37121));
  nnd2s1 _______498260(.DIN1 (____9_9__37069), .DIN2 (________23839),
       .Q (____0____37120));
  xor2s1 _______498261(.DIN1 (______9__35007), .DIN2 (____99___37092),
       .Q (____0____37119));
  nor2s1 _____9_498262(.DIN1 (_________38599), .DIN2 (____9____37065),
       .Q (____0____37157));
  nor2s1 ______498263(.DIN1 (____0____37118), .DIN2 (____9____37076),
       .Q (____0____37156));
  xor2s1 _______498264(.DIN1 (____9____37086), .DIN2 (______0__38256),
       .Q (_________37926));
  nor2s1 _______498265(.DIN1 (_____9__25527), .DIN2 (____9_0__37053),
       .Q (____0____37117));
  nnd2s1 _______498266(.DIN1 (____0_0__40780), .DIN2
       (_____________________________________________21924), .Q
       (____0_0__37116));
  or2s1 _______498267(.DIN1
       (_____________________________________________21924), .DIN2
       (____0_0__40780), .Q (____0____37115));
  nor2s1 _______498268(.DIN1 (_________36886), .DIN2 (____0____37111),
       .Q (____0____37112));
  nor2s1 _______498269(.DIN1 (_________36501), .DIN2 (____9____37050),
       .Q (____0____37110));
  or2s1 ______498270(.DIN1 (_________34788), .DIN2 (____009__37108), .Q
       (____0_0__37109));
  xor2s1 ______498271(.DIN1 (_________35702), .DIN2 (____9____37077),
       .Q (____00___37107));
  nor2s1 _______498272(.DIN1 (_________36022), .DIN2 (_________38350),
       .Q (____00___37106));
  xor2s1 _______498273(.DIN1 (____9_9__37022), .DIN2 (___9_____39784),
       .Q (____00___37105));
  nnd2s1 _______498274(.DIN1 (____9____37055), .DIN2 (____90__26673),
       .Q (____00___37104));
  nnd2s1 ______498275(.DIN1 (_________36422), .DIN2 (____9____37054),
       .Q (____00___37103));
  nor2s1 ______498276(.DIN1 (____00___37102), .DIN2 (_________36339),
       .Q (____0____37149));
  xor2s1 _______498277(.DIN1 (____9____37034), .DIN2 (_________36531),
       .Q (____0____37154));
  nor2s1 ______498278(.DIN1 (____9____37046), .DIN2 (____0_0__40790),
       .Q (____00___37101));
  nor2s1 _____498279(.DIN1 (_________38599), .DIN2 (____99___37098), .Q
       (____000__37100));
  nnd2s1 _______498280(.DIN1 (____99___37098), .DIN2 (____9____37024),
       .Q (____999__37099));
  nnd2s1 _______498281(.DIN1 (____9____37040), .DIN2 (____99___37096),
       .Q (____99___37097));
  nnd2s1 _______498282(.DIN1 (____9____37041), .DIN2 (________25657),
       .Q (____99___37095));
  nnd2s1 _______498283(.DIN1 (____99___37098), .DIN2 (_________38599),
       .Q (____99___37094));
  or2s1 _______498284(.DIN1 (_________34985), .DIN2 (____99___37092),
       .Q (____99___37093));
  nnd2s1 _______498285(.DIN1 (_____99__33813), .DIN2 (____9_9__37042),
       .Q (____99___37091));
  nnd2s1 _______498286(.DIN1 (____9____37039), .DIN2 (_____9___37943),
       .Q (____990__37090));
  or2s1 ______498287(.DIN1 (________22527), .DIN2 (____9____37088), .Q
       (____9_9__37089));
  nnd2s1 _______498288(.DIN1 (____9____37088), .DIN2 (_____0__22654),
       .Q (____9____37087));
  nor2s1 _____9_498289(.DIN1 (____9____37058), .DIN2 (____9____37086),
       .Q (_________37734));
  nor2s1 _____498290(.DIN1 (____9_0__37060), .DIN2 (____9____37057), .Q
       (____0____37137));
  dffacs1 _______________________________________________498291(.CLRB
       (reset), .CLK (clk), .DIN (____9____37048), .QN
       (___0_____40487));
  nor2s1 _____0_498292(.DIN1 (_________38599), .DIN2 (____9____37064),
       .Q (____0____37161));
  nnd2s1 _____0_498293(.DIN1 (______0__37776), .DIN2 (____9_0__37023),
       .Q (_________37700));
  nnd2s1 _______498294(.DIN1 (____9____37031), .DIN2 (_________37317),
       .Q (____9____37085));
  xor2s1 _____0_498295(.DIN1 (____90___37010), .DIN2 (______0__36985),
       .Q (____9____37084));
  xor2s1 _____0_498296(.DIN1 (_________36953), .DIN2 (____9____37047),
       .Q (____9____37083));
  nnd2s1 _______498297(.DIN1 (____9____37029), .DIN2 (______9__37555),
       .Q (____9____37082));
  and2s1 _______498298(.DIN1 (____9____37030), .DIN2 (____9_0__37080),
       .Q (____9____37081));
  nnd2s1 _______498299(.DIN1 (____9____37028), .DIN2 (_________37230),
       .Q (____9_9__37079));
  or2s1 _______498300(.DIN1 (_____0___35655), .DIN2 (____9____37077),
       .Q (____9____37078));
  hi1s1 ______498301(.DIN (_________38350), .Q (____9____37076));
  nnd2s1 ______498302(.DIN1 (____9____37072), .DIN2 (_________38599),
       .Q (____9____37075));
  xor2s1 _____9_498303(.DIN1 (_________36894), .DIN2 (____9____37073),
       .Q (____9____37074));
  nor2s1 _____9_498304(.DIN1 (___09____40688), .DIN2 (____9____37072),
       .Q (______0__37232));
  xor2s1 ______498305(.DIN1 (________), .DIN2 (____9____37045), .Q
       (____9____37071));
  nnd2s1 _______498306(.DIN1 (____9____37020), .DIN2 (_____9___38319),
       .Q (____9_0__37070));
  nnd2s1 _______498307(.DIN1 (____9____37019), .DIN2 (_____9___37752),
       .Q (____9_9__37069));
  nnd2s1 _______498308(.DIN1 (____9____37018), .DIN2 (____0____37167),
       .Q (____9____37068));
  hi1s1 _______498309(.DIN (____9____37066), .Q (____9____37067));
  hi1s1 _______498310(.DIN (____9____37064), .Q (____9____37065));
  xor2s1 _____9_498311(.DIN1 (____9____37062), .DIN2 (____9____37073),
       .Q (____9____37063));
  nor2s1 ______498312(.DIN1 (____9____37056), .DIN2 (____9_0__37060),
       .Q (____9____37061));
  dffacs1 _______________________________________________498313(.CLRB
       (reset), .CLK (clk), .DIN (____9____37021), .Q
       (_____________________________________________21841));
  nor2s1 ______498314(.DIN1 (____9____37037), .DIN2 (_________37679),
       .Q (____9____37058));
  nor2s1 _______498315(.DIN1 (____0____36235), .DIN2 (____9____37056),
       .Q (____9____37057));
  xor2s1 _______498316(.DIN1
       (____________________________________________21790), .DIN2
       (___0_9___40555), .Q (____9____37055));
  nnd2s1 _______498317(.DIN1 (______9__36994), .DIN2 (inData[30]), .Q
       (____9____37054));
  nor2s1 _______498318(.DIN1 (____9_9__37052), .DIN2 (_____99__37003),
       .Q (____9_0__37053));
  nnd2s1 _______498319(.DIN1 (____900__37004), .DIN2 (____9____38001),
       .Q (____9____37051));
  and2s1 _______498320(.DIN1 (____90___37005), .DIN2 (____9____37049),
       .Q (____9____37050));
  nnd2s1 ______498321(.DIN1 (_________36965), .DIN2 (____90___37008),
       .Q (____9____37048));
  nnd2s1 _______498322(.DIN1 (____90___37011), .DIN2 (_________36524),
       .Q (______0__37584));
  nor2s1 _______498323(.DIN1 (______0__36951), .DIN2 (____9____37047),
       .Q (____0____37114));
  nor2s1 _______498324(.DIN1 (_________36645), .DIN2 (____9_0__37014),
       .Q (____0____37111));
  nor2s1 _______498325(.DIN1 (_________34824), .DIN2 (_____9___36999),
       .Q (____009__37108));
  nor2s1 _____0_498326(.DIN1 (_________36968), .DIN2 (_____9___37001),
       .Q (____00___37102));
  xor2s1 _______498327(.DIN1 (_________36983), .DIN2 (______0__36970),
       .Q (____0____37129));
  xor2s1 _____0_498328(.DIN1 (____0____40784), .DIN2 (_________36864),
       .Q (_________38350));
  nor2s1 _____0_498329(.DIN1 (____9____37045), .DIN2 (_________35157),
       .Q (____9____37046));
  xor2s1 _______498330(.DIN1 (____9_0__37043), .DIN2 (___0_9___40555),
       .Q (____9____37044));
  nnd2s1 _____0_498331(.DIN1 (_____0___36728), .DIN2 (____9____37045),
       .Q (____9_9__37042));
  nnd2s1 _____9_498332(.DIN1 (_________36993), .DIN2 (______0__37872),
       .Q (____9____37041));
  xor2s1 _____498333(.DIN1 (_________35411), .DIN2 (____9____37015), .Q
       (____9____37040));
  xor2s1 _____0_498334(.DIN1 (____9____37016), .DIN2 (_________36885),
       .Q (____9____37039));
  nor2s1 _______498335(.DIN1 (_________36834), .DIN2 (____9____37073),
       .Q (____9____37038));
  nor2s1 _______498336(.DIN1 (_________34785), .DIN2 (_________36990),
       .Q (____99___37092));
  nor2s1 _______498337(.DIN1 (______0__36833), .DIN2 (____9____37073),
       .Q (____9____37064));
  and2s1 _______498338(.DIN1 (_________37679), .DIN2 (____9____37037),
       .Q (____9____37086));
  dffacs1 _______________________________________________498339(.CLRB
       (reset), .CLK (clk), .DIN (_____9___37000), .QN
       (_____________________________________________21801));
  xor2s1 _______498340(.DIN1 (_________36980), .DIN2 (____9____37036),
       .Q (____9____37066));
  nnd2s1 _______498341(.DIN1 (____9____37073), .DIN2 (_________36805),
       .Q (______0__37776));
  dffacs1 _______________________________________________498342(.CLRB
       (reset), .CLK (clk), .DIN (____90___37007), .QN
       (___0__9__40510));
  nor2s1 _______498343(.DIN1 (_________36959), .DIN2 (_________36991),
       .Q (____9____37088));
  nnd2s1 _______498344(.DIN1 (____9____37073), .DIN2 (_____9___36909),
       .Q (____99___37098));
  dffacs1 __________________498345(.CLRB (reset), .CLK (clk), .DIN
       (_____9___36997), .QN
       (_______________________________________________________________________________________));
  nnd2s1 ______498346(.DIN1 (_________36988), .DIN2 (_________37223),
       .Q (____9____37035));
  xor2s1 _______498347(.DIN1 (_____9___36453), .DIN2 (____9_9__37032),
       .Q (____9____37034));
  xor2s1 _______498348(.DIN1 (_____9__26456), .DIN2 (____9_9__37032),
       .Q (____9_0__37033));
  xor2s1 _______498349(.DIN1 (_____9___36998), .DIN2 (_________34825),
       .Q (____9____37031));
  xor2s1 _______498350(.DIN1 (_________36958), .DIN2 (_____9___37851),
       .Q (____9____37030));
  xor2s1 _______498351(.DIN1 (_________36763), .DIN2 (____909__37013),
       .Q (____9____37029));
  xor2s1 _____498352(.DIN1 (_________36974), .DIN2 (_____0___36921), .Q
       (____9____37028));
  nor2s1 _______498353(.DIN1
       (____________________________________________), .DIN2
       (____9____37026), .Q (____9____37027));
  nnd2s1 _______498354(.DIN1 (____9____37026), .DIN2
       (____________________________________________), .Q
       (____9____37025));
  nnd2s1 ______498355(.DIN1 (____9____37026), .DIN2 (_________36855),
       .Q (____9____37024));
  nor2s1 ______498356(.DIN1 (______9__35405), .DIN2 (_________36982),
       .Q (____9____37077));
  nnd2s1 _______498357(.DIN1 (_________36987), .DIN2 (____90___37009),
       .Q (____0____37153));
  nnd2s1 ______498358(.DIN1 (____9____37026), .DIN2 (______0__36775),
       .Q (____9_0__37023));
  nor2s1 _______498359(.DIN1 (_________36861), .DIN2 (____9____37026),
       .Q (____9_9__37022));
  dffacs1 ________________498360(.CLRB (reset), .CLK (clk), .DIN
       (____9____37026), .Q (outData[14]));
  nnd2s1 ______498361(.DIN1 (______9__36977), .DIN2 (____9___23873), .Q
       (____9____37021));
  nor2s1 _____9_498362(.DIN1 (_____9__26167), .DIN2 (_________36981),
       .Q (____9____37020));
  xor2s1 _____498363(.DIN1 (_________34807), .DIN2 (_________36989), .Q
       (____9____37019));
  xor2s1 _____0_498364(.DIN1 (______0__36961), .DIN2 (_________35158),
       .Q (____9____37018));
  nor2s1 _____0_498365(.DIN1 (___0_9___40555), .DIN2 (____9_0__37043),
       .Q (____9____37017));
  nor2s1 _____0_498366(.DIN1 (___0_____40439), .DIN2 (_________36979),
       .Q (____9_0__37060));
  nor2s1 _______498367(.DIN1 (______0__36860), .DIN2 (____9____37026),
       .Q (____9____37072));
  nor2s1 _______498368(.DIN1 (_________35410), .DIN2 (____9____37015),
       .Q (____9____37059));
  dffacs1 __________________498369(.CLRB (reset), .CLK (clk), .DIN
       (______9__36984), .QN (___0__9__40412));
  nor2s1 _______498370(.DIN1 (______0__36660), .DIN2 (____909__37013),
       .Q (____9_0__37014));
  nnd2s1 _______498371(.DIN1 (____9_9__37032), .DIN2
       (__________________________________________________________________22005),
       .Q (____90___37012));
  or2s1 _______498372(.DIN1 (_________36532), .DIN2 (____9_9__37032),
       .Q (____90___37011));
  and2s1 _____9_498373(.DIN1 (_________36986), .DIN2 (____90___37009),
       .Q (____90___37010));
  nnd2s1 ______498374(.DIN1 (____9_9__36114), .DIN2 (_________36966),
       .Q (____90___37008));
  nnd2s1 _______498375(.DIN1 (_________36967), .DIN2 (______0__36924),
       .Q (____90___37007));
  or2s1 _______498376(.DIN1
       (__________________________________________________________________22005),
       .DIN2 (____9_9__37032), .Q (____90___37006));
  xor2s1 _______498377(.DIN1 (_________35407), .DIN2 (____0____40786),
       .Q (____90___37005));
  xor2s1 _______498378(.DIN1 (______9__36950), .DIN2 (_________36975),
       .Q (____900__37004));
  xor2s1 _______498379(.DIN1 (_________36947), .DIN2 (_____9___37002),
       .Q (_____99__37003));
  nor2s1 _______498380(.DIN1 (____9____36124), .DIN2 (_________36976),
       .Q (_____9___37001));
  nor2s1 _____0_498381(.DIN1 (___09____40673), .DIN2 (_________36971),
       .Q (____9____37047));
  dffacs1 ________________498382(.CLRB (reset), .CLK (clk), .DIN
       (_________38599), .Q (outData[15]));
  nnd2s1 ______498383(.DIN1 (______9__36960), .DIN2 (________24445), .Q
       (_____9___37000));
  and2s1 _______498384(.DIN1 (_____9___36998), .DIN2 (______9__34789),
       .Q (_____9___36999));
  nnd2s1 ______498385(.DIN1 (_____9___36996), .DIN2 (_________36957),
       .Q (_____9___36997));
  nnd2s1 _______498386(.DIN1 (_________37538), .DIN2 (___0_____40444),
       .Q (_____90__36995));
  and2s1 _____9_498387(.DIN1 (________24384), .DIN2 (___0_____40444),
       .Q (______9__36994));
  xor2s1 _______498388(.DIN1 (_________36992), .DIN2 (_________36944),
       .Q (_________36993));
  and2s1 ______498389(.DIN1 (_________36963), .DIN2 (___9_0___39077),
       .Q (_________36991));
  nor2s1 ______498390(.DIN1 (_________34793), .DIN2 (_________36989),
       .Q (_________36990));
  nor2s1 _____498391(.DIN1 (___9____27819), .DIN2 (______0__36978), .Q
       (____9____37056));
  hi1s1 _______498392(.DIN (___0_9___40555), .Q (____9____37045));
  xor2s1 _______498393(.DIN1 (___09____40688), .DIN2 (_________38573),
       .Q (_________37679));
  dffacs1 _______________________________________________498394(.CLRB
       (reset), .CLK (clk), .DIN (_________36962), .QN
       (_____________________________________________21823));
  hi1s1 _____9_498395(.DIN (____9____37026), .Q (____9____37073));
  xor2s1 _____9_498396(.DIN1 (_____9___36911), .DIN2 (____0____40792),
       .Q (_________36988));
  nnd2s1 _______498397(.DIN1 (_________36986), .DIN2 (______0__36985),
       .Q (_________36987));
  nnd2s1 _______498398(.DIN1 (_________36948), .DIN2 (__90____29645),
       .Q (______9__36984));
  nor2s1 _______498399(.DIN1 (______9__36969), .DIN2 (___09____40673),
       .Q (_________36983));
  nor2s1 ______498400(.DIN1 (_________35409), .DIN2 (____0____40786),
       .Q (_________36982));
  dffacs1 _______________________________________________498401(.CLRB
       (reset), .CLK (clk), .DIN (_________36949), .QN
       (_____________________________________________21811));
  and2s1 _______498402(.DIN1 (______9__36941), .DIN2 (_________38249),
       .Q (_________36981));
  nor2s1 _______498403(.DIN1 (_____0___36917), .DIN2 (_________37737),
       .Q (_________36980));
  hi1s1 ______498404(.DIN (______0__36978), .Q (_________36979));
  nnd2s1 _______498405(.DIN1 (______0__36942), .DIN2 (______9__37314),
       .Q (______9__36977));
  nor2s1 _______498406(.DIN1 (_________36943), .DIN2 (_________36938),
       .Q (____9____37016));
  nor2s1 _______498407(.DIN1 (______9__35121), .DIN2 (_________36940),
       .Q (____9____37015));
  dffacs1 _______________________________________________498408(.CLRB
       (reset), .CLK (clk), .DIN (_________36945), .Q (___0_9___40555));
  xnr2s1 _______498409(.DIN1 (___909___39065), .DIN2 (_____0___36920),
       .Q (____9____37026));
  and2s1 _____0_498410(.DIN1 (_________36975), .DIN2 (___0_____40538),
       .Q (_________36976));
  xor2s1 _____498411(.DIN1 (_____9__22567), .DIN2 (_________36898), .Q
       (_________36974));
  nor2s1 _______498412(.DIN1 (______0__36970), .DIN2 (______9__36969),
       .Q (_________36971));
  nor2s1 _____9_498413(.DIN1 (___0_____40538), .DIN2 (_________36975),
       .Q (_________36968));
  nor2s1 _______498414(.DIN1 (_____09__36923), .DIN2 (____0____35325),
       .Q (_________36967));
  nnd2s1 _______498415(.DIN1 (_________36926), .DIN2 (inData[8]), .Q
       (_________36966));
  nor2s1 _______498416(.DIN1 (_________36925), .DIN2 (____9_0__36115),
       .Q (_________36965));
  dffacs1 _________________________________________9_____498417(.CLRB
       (reset), .CLK (clk), .DIN (_________36933), .QN
       (___0_9___40459));
  nnd2s1 _______498418(.DIN1 (_________36964), .DIN2 (_________36595),
       .Q (____90___37009));
  nor2s1 _______498419(.DIN1 (______9__36931), .DIN2 (_________36927),
       .Q (____909__37013));
  xor2s1 _______498420(.DIN1 (______0__36897), .DIN2 (_________38142),
       .Q (____9_9__37032));
  nnd2s1 _______498421(.DIN1 (_____9___36908), .DIN2 (_______22178), .Q
       (_________36963));
  nnd2s1 _______498422(.DIN1 (______9__35896), .DIN2 (_____0___36919),
       .Q (_________36962));
  xor2s1 _____0_498423(.DIN1 (_________36939), .DIN2 (___0_____40308),
       .Q (______0__36961));
  nnd2s1 ______498424(.DIN1 (_____00__36914), .DIN2 (_________38576),
       .Q (______9__36960));
  nor2s1 _____9_498425(.DIN1 (___9_0___39077), .DIN2 (_____90__36904),
       .Q (_________36959));
  xor2s1 _____0_498426(.DIN1 (___0_____40485), .DIN2 (_________36892),
       .Q (_________36958));
  nor2s1 _______498427(.DIN1 (_____0___36918), .DIN2 (____09__27400),
       .Q (_________36957));
  nor2s1 ______498428(.DIN1 (_________36955), .DIN2 (_____9___36910),
       .Q (_________36956));
  xor2s1 _______498429(.DIN1 (______0__36889), .DIN2 (___009___39979),
       .Q (______0__36978));
  xnr2s1 _______498430(.DIN1 (_________35968), .DIN2 (_________36890),
       .Q (_____9___36998));
  nor2s1 _______498431(.DIN1 (_____0___34758), .DIN2 (_____9___36906),
       .Q (_________36989));
  dffacs1 __________________________________________0____498432(.CLRB
       (reset), .CLK (clk), .DIN (_____9___36912), .QN
       (___0_____40444));
  dffacs1 _______________________________________________498433(.CLRB
       (reset), .CLK (clk), .DIN (_________36934), .Q
       (_____________________________________________21908));
  hi1s1 _______498434(.DIN (___09____40688), .Q (_________38599));
  nnd2s1 _____0_498435(.DIN1 (_________36953), .DIN2 (_________36952),
       .Q (_________36954));
  nor2s1 _____0_498436(.DIN1 (_________36952), .DIN2 (_________36953),
       .Q (______0__36951));
  xor2s1 ______498437(.DIN1 (____9____36125), .DIN2 (___0_____40538),
       .Q (______9__36950));
  nnd2s1 _______498438(.DIN1 (_________36902), .DIN2 (_____0__24656),
       .Q (_________36949));
  nnd2s1 _______498439(.DIN1 (_________36901), .DIN2 (______0__36766),
       .Q (_________36948));
  nnd2s1 _______498440(.DIN1 (_________36930), .DIN2 (_________36893),
       .Q (_________36947));
  nnd2s1 _______498441(.DIN1 (_________36946), .DIN2 (_________36596),
       .Q (_________36986));
  nnd2s1 _______498442(.DIN1 (_________36891), .DIN2 (_________38550),
       .Q (_________36945));
  nor2s1 _______498443(.DIN1 (_________36943), .DIN2 (_________36936),
       .Q (_________36944));
  xor2s1 _____9_498444(.DIN1 (_________34792), .DIN2 (_____9___36905),
       .Q (______0__36942));
  xor2s1 _____498445(.DIN1 (_________36857), .DIN2 (______0__35087), .Q
       (______9__36941));
  nor2s1 _______498446(.DIN1 (_________35119), .DIN2 (_________36939),
       .Q (_________36940));
  nor2s1 ______498447(.DIN1 (_________36937), .DIN2 (_________36936),
       .Q (_________36938));
  dffacs1 _______________________________________________498448(.CLRB
       (reset), .CLK (clk), .DIN (______9__36896), .Q
       (_____________________________________________21808));
  hi1s1 _______498449(.DIN (_________36935), .Q (_________37737));
  dffacs1 _______________________________________________498450(.CLRB
       (reset), .CLK (clk), .DIN (_________36900), .QN
       (___0__9__40520));
  nnd2s1 _______498451(.DIN1 (_________36874), .DIN2 (________27369),
       .Q (_________36934));
  nnd2s1 _______498452(.DIN1 (_________36881), .DIN2 (______0__36932),
       .Q (_________36933));
  nor2s1 _______498453(.DIN1 (_________________0_), .DIN2
       (_________36930), .Q (______9__36931));
  nor2s1 ______498454(.DIN1 (___9_____39397), .DIN2 (_________36873),
       .Q (_________36927));
  and2s1 _______498455(.DIN1 (_____0___36922), .DIN2 (_________36853),
       .Q (_________36926));
  nor2s1 _______498456(.DIN1 (_________36852), .DIN2 (______0__36924),
       .Q (_________36925));
  nor2s1 _______498457(.DIN1 (_____0___36922), .DIN2 (_________36870),
       .Q (_____09__36923));
  nnd2s1 _______498458(.DIN1 (_________36877), .DIN2 (_________36849),
       .Q (_________37299));
  nor2s1 ______498459(.DIN1 (_________36771), .DIN2 (_________36899),
       .Q (______9__36969));
  hi1s1 _____9_498460(.DIN (_________36946), .Q (_________36964));
  nnd2s1 _______498461(.DIN1 (_____0___36921), .DIN2 (_________36875),
       .Q (_________36972));
  nor2s1 _______498462(.DIN1 (_____9___36818), .DIN2 (_________36872),
       .Q (_________36975));
  xor2s1 _____0_498463(.DIN1 (_____0___36829), .DIN2
       (______________22104), .Q (_____0___36920));
  nnd2s1 _______498464(.DIN1 (_________36867), .DIN2 (inData[20]), .Q
       (_____0___36919));
  and2s1 _______498465(.DIN1 (____0____37165), .DIN2 (_________36862),
       .Q (_____0___36918));
  nor2s1 ______498466(.DIN1 (______9__36903), .DIN2 (____9____37037),
       .Q (_____0___36917));
  nor2s1 _____498467(.DIN1 (______0__32803), .DIN2 (_________36866), .Q
       (_____0___36916));
  or2s1 _____9_498468(.DIN1 (___90____39055), .DIN2 (_________37386),
       .Q (_____0___36915));
  xor2s1 _____498469(.DIN1 (_____0___36827), .DIN2 (_____99__36913), .Q
       (_____00__36914));
  nnd2s1 _______498470(.DIN1 (______9__36868), .DIN2 (_________37454),
       .Q (_____9___36912));
  xor2s1 _____0_498471(.DIN1 (_____0___36826), .DIN2 (_________36778),
       .Q (_____9___36911));
  nor2s1 ______498472(.DIN1 (_________36836), .DIN2 (_____9___36909),
       .Q (_____9___36910));
  or2s1 _______498473(.DIN1 (_______22182), .DIN2 (_____9___36907), .Q
       (_____9___36908));
  nor2s1 _______498474(.DIN1 (_____0___34759), .DIN2 (_____9___36905),
       .Q (_____9___36906));
  nnd2s1 _______498475(.DIN1 (_____9___36907), .DIN2 (________22602),
       .Q (_____90__36904));
  nnd2s1 _______498476(.DIN1 (____9____37037), .DIN2 (______9__36903),
       .Q (_________36935));
  dffacs1 _______________________________________________498477(.CLRB
       (reset), .CLK (clk), .DIN (______9__36878), .QN
       (_____________________________________________21969));
  or2s1 _______498478(.DIN1 (_____9___37656), .DIN2 (_________36848),
       .Q (_________36902));
  nnd2s1 _______498479(.DIN1 (______0__36851), .DIN2 (inData[0]), .Q
       (_________36901));
  nnd2s1 _______498480(.DIN1 (______9__36850), .DIN2 (_________36621),
       .Q (_________36900));
  xor2s1 _______498481(.DIN1 (______0__36879), .DIN2 (___9__9__39125),
       .Q (_________36898));
  xor2s1 _______498482(.DIN1 (_________35900), .DIN2 (______0__36869),
       .Q (______0__36897));
  nnd2s1 ______498483(.DIN1 (____0____35335), .DIN2 (_________36845),
       .Q (______9__36896));
  xor2s1 _______498484(.DIN1 (_________36876), .DIN2 (______9__36328),
       .Q (_________36953));
  xor2s1 _______498485(.DIN1 (_____9___36819), .DIN2 (_________36764),
       .Q (_________36946));
  nor2s1 _______498486(.DIN1 (_________36804), .DIN2 (_____09__36832),
       .Q (_________36894));
  nnd2s1 _____9_498487(.DIN1 (_________36689), .DIN2 (_________36847),
       .Q (_________36893));
  nnd2s1 _____0_498488(.DIN1 (______0__36842), .DIN2 (___09____40674),
       .Q (_________36892));
  nor2s1 _______498489(.DIN1 (____9___26224), .DIN2 (______9__36841),
       .Q (_________36891));
  nnd2s1 _______498490(.DIN1 (_________36835), .DIN2 (_________36798),
       .Q (_________36890));
  nnd2s1 _______498491(.DIN1 (_____0___36831), .DIN2 (_________35860),
       .Q (______0__36889));
  nor2s1 ______498492(.DIN1 (_________36887), .DIN2 (_________36886),
       .Q (______9__36888));
  nor2s1 _______498493(.DIN1 (_________36884), .DIN2 (_________36863),
       .Q (_________36885));
  nor2s1 _______498494(.DIN1 (_________35072), .DIN2 (_____0___36825),
       .Q (_________36939));
  and2s1 _______498495(.DIN1 (_________36882), .DIN2 (_________36883),
       .Q (_________36943));
  nor2s1 _______498496(.DIN1 (_________36883), .DIN2 (_________36882),
       .Q (_________36936));
  dffacs1 _______________________________________________498497(.CLRB
       (reset), .CLK (clk), .DIN (_________36844), .QN
       (___0__9__40420));
  nor2s1 _______498498(.DIN1 (________25235), .DIN2 (_____9___36821),
       .Q (_________36881));
  nnd2s1 _______498499(.DIN1 (______0__36879), .DIN2
       (_______________________________________________________________0),
       .Q (_________36880));
  nnd2s1 _______498500(.DIN1 (_____9___36820), .DIN2 (________29316),
       .Q (______9__36878));
  or2s1 _______498501(.DIN1 (___9_____39123), .DIN2 (_________36876),
       .Q (_________36877));
  or2s1 _______498502(.DIN1
       (_______________________________________________________________0),
       .DIN2 (______0__36879), .Q (_________36875));
  nnd2s1 _______498503(.DIN1 (_________36808), .DIN2 (___9__9__39459),
       .Q (_________36874));
  nor2s1 ______498504(.DIN1 (_________36809), .DIN2 (_____9___36815),
       .Q (_________36873));
  nor2s1 _____9_498505(.DIN1 (_________36653), .DIN2 (_____9___36816),
       .Q (_________36872));
  xor2s1 ______498506(.DIN1 (______9__36792), .DIN2 (_________36871),
       .Q (_________36899));
  nor2s1 _______498507(.DIN1 (_____99__36822), .DIN2 (__99____30514),
       .Q (_____0___36922));
  or2s1 _______498508(.DIN1 (______9__36812), .DIN2 (_________36870),
       .Q (______0__36924));
  nor2s1 _______498509(.DIN1 (______0__36793), .DIN2 (_____90__36813),
       .Q (___0_____40130));
  nor2s1 _____0_498510(.DIN1 (_________36782), .DIN2 (______0__36869),
       .Q (_________36929));
  nnd2s1 _____0_498511(.DIN1 (_____9___36814), .DIN2 (_________36846),
       .Q (_________36930));
  dffacs1 __________________498512(.CLRB (reset), .CLK (clk), .DIN
       (_________36811), .QN
       (_________________________________________________________________________________________22091));
  nor2s1 _______498513(.DIN1 (_________36671), .DIN2 (______9__36802),
       .Q (______9__36868));
  and2s1 ______498514(.DIN1 (_________37576), .DIN2 (_________36801),
       .Q (_________36867));
  xor2s1 _______498515(.DIN1 (_________35887), .DIN2 (_____0___36830),
       .Q (_________36866));
  xor2s1 ______498516(.DIN1 (________24333), .DIN2 (_________36864), .Q
       (_________36865));
  nnd2s1 ______498517(.DIN1 (______0__36803), .DIN2 (inData[8]), .Q
       (_________36862));
  hi1s1 _____9_498518(.DIN (______0__36860), .Q (_________36861));
  xor2s1 ____9_498519(.DIN1 (_________38482), .DIN2 (_________36858),
       .Q (______9__36859));
  xor2s1 ____9_498520(.DIN1 (_____0___36824), .DIN2 (_________36856),
       .Q (_________36857));
  xor2s1 ____9__498521(.DIN1 (____0____40788), .DIN2 (_________41341),
       .Q (_____9___36905));
  hi1s1 _____9_498522(.DIN (_________36855), .Q (_____9___36909));
  nor2s1 ______498523(.DIN1 (___09___22358), .DIN2 (_________36800), .Q
       (_____9___36907));
  or2s1 _______498524(.DIN1 (_________36806), .DIN2 (_____0___37475),
       .Q (_________37386));
  dffacs1 _______________________________________________498525(.CLRB
       (reset), .CLK (clk), .DIN (_________36795), .Q (___0_____40538));
  xor2s1 _______498526(.DIN1 (_________36854), .DIN2 (_________36864),
       .Q (____9____37037));
  nnd2s1 _______498527(.DIN1 (_________36837), .DIN2 (_________36852),
       .Q (_________36853));
  nor2s1 _______498528(.DIN1 (_________36789), .DIN2 (_________36713),
       .Q (______0__36851));
  nor2s1 _______498529(.DIN1 (________27104), .DIN2 (_________36790),
       .Q (______9__36850));
  nor2s1 _______498530(.DIN1 (_________36325), .DIN2 (_________36791),
       .Q (_________36849));
  xor2s1 _____9_498531(.DIN1 (_________36654), .DIN2 (_____9___36817),
       .Q (_________36848));
  hi1s1 _______498532(.DIN (_________36846), .Q (_________36847));
  nnd2s1 _______498533(.DIN1 (_________36787), .DIN2 (inData[2]), .Q
       (_________36845));
  nnd2s1 ______498534(.DIN1 (_________36794), .DIN2 (___9909__39806),
       .Q (_________36844));
  nor2s1 ______498535(.DIN1
       (__________________________________________________________________21988),
       .DIN2 (_________36864), .Q (_________36843));
  nor2s1 _______498536(.DIN1 (_________38435), .DIN2 (_________36780),
       .Q (______9__36841));
  or2s1 _______498537(.DIN1 (_________36839), .DIN2 (_________36838),
       .Q (_________36840));
  nor2s1 _______498538(.DIN1 (______9__36903), .DIN2 (_________36788),
       .Q (_________36895));
  nor2s1 _______498539(.DIN1 (______9__34981), .DIN2 (_________36837),
       .Q (_________36886));
  nor2s1 _______498540(.DIN1 (_____00__36823), .DIN2 (_________36864),
       .Q (_________36836));
  nnd2s1 ______498541(.DIN1 (____0____40792), .DIN2 (_________36779),
       .Q (_________36835));
  hi1s1 _____9_498542(.DIN (______0__36833), .Q (_________36834));
  nor2s1 ____90_498543(.DIN1 (______0__36736), .DIN2 (_________36864),
       .Q (_____09__36832));
  or2s1 ____90_498544(.DIN1 (_________35763), .DIN2 (_____0___36830),
       .Q (_____0___36831));
  xor2s1 ____9__498545(.DIN1 (_____________22080), .DIN2
       (_________36799), .Q (_____0___36829));
  nnd2s1 ______498546(.DIN1 (_________36864), .DIN2
       (__________________________________________________________________21988),
       .Q (_____0___36828));
  xor2s1 ____9__498547(.DIN1 (_________36760), .DIN2 (_________34954),
       .Q (_____0___36827));
  xor2s1 ____9__498548(.DIN1 (_________36797), .DIN2 (___9_0___39077),
       .Q (_____0___36826));
  nor2s1 ____9__498549(.DIN1 (_________35071), .DIN2 (_____0___36824),
       .Q (_____0___36825));
  nnd2s1 ____9__498550(.DIN1 (_________36864), .DIN2 (_____00__36823),
       .Q (_________36855));
  nor2s1 ____9__498551(.DIN1 (_____09__36735), .DIN2 (_________36864),
       .Q (______0__36860));
  nor2s1 ____9__498552(.DIN1 (___0_0___40566), .DIN2 (_________38482),
       .Q (_________36863));
  nnd2s1 ____9__498553(.DIN1 (_________36777), .DIN2 (_________36703),
       .Q (_________36882));
  dffacs1 _______________________________________________498554(.CLRB
       (reset), .CLK (clk), .DIN (_________36776), .QN
       (_____________________________________________21767));
  nor2s1 _______498555(.DIN1
       (_____________________________________________21871), .DIN2
       (_____________________________________________21837), .Q
       (_____99__36822));
  nor2s1 _____9_498556(.DIN1 (____9_9__37052), .DIN2 (_________36769),
       .Q (_____9___36821));
  nnd2s1 _____9_498557(.DIN1 (_________36770), .DIN2 (___0_____40156),
       .Q (_____9___36820));
  xor2s1 _____0_498558(.DIN1 (_________36740), .DIN2 (_________38650),
       .Q (_____9___36819));
  nor2s1 _______498559(.DIN1
       (_____________________________________________21800), .DIN2
       (_____9___36817), .Q (_____9___36818));
  and2s1 ______498560(.DIN1 (_____9___36817), .DIN2
       (_____________________________________________21800), .Q
       (_____9___36816));
  nor2s1 _______498561(.DIN1 (_________36810), .DIN2 (_____9___36814),
       .Q (_____9___36815));
  nor2s1 _______498562(.DIN1 (_____________________21677), .DIN2
       (_________36768), .Q (_____90__36813));
  nnd2s1 _______498563(.DIN1
       (_____________________________________________21837), .DIN2
       (_____________________________________________21871), .Q
       (______9__36812));
  nnd2s1 _______498564(.DIN1 (_________36767), .DIN2 (__9_____29740),
       .Q (_________36811));
  nnd2s1 _______498565(.DIN1 (______0__36784), .DIN2 (____9____35235),
       .Q (______0__36842));
  nor2s1 _______498566(.DIN1 (_________36810), .DIN2 (_________36809),
       .Q (_________36846));
  nor2s1 _______498567(.DIN1
       (_____________________________________________21871), .DIN2
       (___0_____40411), .Q (_________36887));
  xor2s1 _____0_498568(.DIN1 (___0_____40125), .DIN2 (____9____36127),
       .Q (_________36876));
  xor2s1 ______498569(.DIN1 (_________36744), .DIN2 (_________36748),
       .Q (______0__36879));
  xor2s1 ____90_498570(.DIN1 (_____0___36732), .DIN2 (_____0___36733),
       .Q (_________36808));
  nnd2s1 _______498571(.DIN1 (_________36754), .DIN2 (inData[8]), .Q
       (_________36807));
  nor2s1 _____498572(.DIN1 (_________36446), .DIN2 (_________36805), .Q
       (_________36806));
  nor2s1 ____90_498573(.DIN1 (_____0___36731), .DIN2 (_________36796),
       .Q (_________36804));
  xor2s1 ____90_498574(.DIN1 (___0_____40523), .DIN2 (___0_____40498),
       .Q (______0__36803));
  nor2s1 _______498575(.DIN1 (_________36955), .DIN2 (_________36758),
       .Q (______9__36802));
  xor2s1 ____9_498576(.DIN1 (_______22242), .DIN2 (___0_____40498), .Q
       (_________36801));
  and2s1 ____9__498577(.DIN1 (_________36799), .DIN2 (_____0), .Q
       (_________36800));
  nnd2s1 ____9__498578(.DIN1 (_________35907), .DIN2 (_________36797),
       .Q (_________36798));
  dffacs1 ________________498579(.CLRB (reset), .CLK (clk), .DIN
       (_________36796), .Q (outData[13]));
  or2s1 _______498580(.DIN1 (____0____38117), .DIN2 (_________36759),
       .Q (_________36795));
  nor2s1 ____9__498581(.DIN1 (_____0___36730), .DIN2 (_________36796),
       .Q (______0__36833));
  nor2s1 ______498582(.DIN1 (_________36752), .DIN2 (______9__36765),
       .Q (______0__36869));
  nor2s1 ____9__498583(.DIN1 (_________36883), .DIN2 (______9__36774),
       .Q (_________36884));
  dffacs1 _____________________________________________0_498584(.CLRB
       (reset), .CLK (clk), .DIN (______0__36756), .QN
       (_________________________________________0___21840));
  dffacs1 __________________________________________0__0_(.CLRB
       (reset), .CLK (clk), .DIN (_________36757), .Q
       (______________________________________0__0_));
  and2s1 _______498585(.DIN1 (_________36751), .DIN2 (________28518),
       .Q (_________36794));
  nor2s1 _______498586(.DIN1 (___9_9___39790), .DIN2 (_________36747),
       .Q (______0__36793));
  nnd2s1 _______498587(.DIN1 (_________36749), .DIN2 (_________36742),
       .Q (______9__36792));
  and2s1 ______498588(.DIN1 (___0_____40125), .DIN2 (______0__36329),
       .Q (_________36791));
  nor2s1 _______498589(.DIN1 (_________36521), .DIN2 (_________36741),
       .Q (_________36790));
  xor2s1 _______498590(.DIN1
       (_____________________________________________21869), .DIN2
       (______0__36561), .Q (_________36789));
  xor2s1 ____90_498591(.DIN1 (_________36704), .DIN2 (_________38842),
       .Q (_________36788));
  nor2s1 _______498592(.DIN1 (_________36750), .DIN2 (_________36618),
       .Q (_________36787));
  nor2s1 _______498593(.DIN1 (_________36785), .DIN2 (_________36772),
       .Q (_________36786));
  nnd2s1 ____498594(.DIN1 (_________38142), .DIN2 (_________36781), .Q
       (______9__36783));
  nor2s1 ____90_498595(.DIN1 (_________36781), .DIN2 (_________38142),
       .Q (_________36782));
  hi1s1 _______498596(.DIN
       (_____________________________________________21871), .Q
       (_________36837));
  xor2s1 ____9__498597(.DIN1 (_________36705), .DIN2 (_________36648),
       .Q (_________36780));
  nnd2s1 ____9__498598(.DIN1 (_________36778), .DIN2 (___0_____40498),
       .Q (_________36779));
  or2s1 ____498599(.DIN1 (___99_0__39864), .DIN2 (_________36737), .Q
       (_________36777));
  nnd2s1 ____9__498600(.DIN1 (______9__36490), .DIN2 (_____0___36729),
       .Q (_________36776));
  xnr2s1 ____9__498601(.DIN1 (_____9___38512), .DIN2 (_________36709),
       .Q (_________36838));
  nor2s1 ____9__498602(.DIN1 (_________36683), .DIN2 (_____0___36734),
       .Q (_____0___36830));
  nor2s1 ____99_498603(.DIN1 (_____9___34926), .DIN2 (_____0___36727),
       .Q (_____0___36824));
  xor2s1 ____9__498604(.DIN1 (______9__36716), .DIN2 (_____00__35736),
       .Q (_________36839));
  nor2s1 ____9__498605(.DIN1 (_________36390), .DIN2 (______0__36775),
       .Q (_____0___37475));
  dffacs1 __________________________________________0____498606(.CLRB
       (reset), .CLK (clk), .DIN (_________36738), .Q
       (______________________________________0______21887));
  hi1s1 ____00_498607(.DIN (______9__36774), .Q (_________38482));
  hi1s1 ____9__498608(.DIN (_________36796), .Q (_________36864));
  hi1s1 ____9__498609(.DIN (_________36772), .Q (_________36773));
  xor2s1 _______498610(.DIN1 (______0__36746), .DIN2 (______9__36745),
       .Q (_________36770));
  xor2s1 _______498611(.DIN1 (_________36694), .DIN2 (_____9___37002),
       .Q (_________36769));
  nor2s1 ______498612(.DIN1 (_________36665), .DIN2 (_____9___36719),
       .Q (_________36768));
  nnd2s1 _______498613(.DIN1 (_________36714), .DIN2 (______0__36766),
       .Q (_________36767));
  nor2s1 ______498614(.DIN1 (_________36712), .DIN2 (_________36764),
       .Q (______9__36765));
  xor2s1 ____9__498615(.DIN1 (_________36698), .DIN2 (_________36762),
       .Q (_________36763));
  xor2s1 ____9__498616(.DIN1 (_________36691), .DIN2 (____9_0__38941),
       .Q (______0__36784));
  nor2s1 _______498617(.DIN1
       (_____________________________________________21869), .DIN2
       (_________36761), .Q (_________36810));
  and2s1 _______498618(.DIN1 (_________36761), .DIN2
       (_____________________________________________21869), .Q
       (_________36809));
  nor2s1 _______498619(.DIN1 (_________36695), .DIN2 (_____9___36722),
       .Q (_________36952));
  nor2s1 _____9_498620(.DIN1 (_________35821), .DIN2 (_____9___36718),
       .Q (_____9___36817));
  dffacs1 _______________________________________________498621(.CLRB
       (reset), .CLK (clk), .DIN (_________36715), .Q
       (_____________________________________________21871));
  xor2s1 ____0__498622(.DIN1
       (_____________________________________________21782), .DIN2
       (_____00__36726), .Q (_________36760));
  xor2s1 ____9__498623(.DIN1 (_____0___36550), .DIN2 (_________36681),
       .Q (_________36759));
  nor2s1 ____9__498624(.DIN1 (_____9___36723), .DIN2 (_____00__36823),
       .Q (_________36758));
  nnd2s1 ____9__498625(.DIN1 (_________35955), .DIN2 (_________36711),
       .Q (_________36757));
  nnd2s1 ____9__498626(.DIN1 (_________36701), .DIN2 (__9_____30135),
       .Q (______0__36756));
  nnd2s1 ____9__498627(.DIN1 (_________36700), .DIN2 (inData[10]), .Q
       (______9__36755));
  nor2s1 ____9__498628(.DIN1 (_________36708), .DIN2 (_________36753),
       .Q (_________36754));
  hi1s1 ____9__498629(.DIN (___0_____40498), .Q (_________36797));
  nnd2s1 ____99_498630(.DIN1 (_________36702), .DIN2 (_________36672),
       .Q (_________36799));
  hi1s1 ____00_498631(.DIN (_________36937), .Q (_________36992));
  hi1s1 ____9_498632(.DIN (______0__36775), .Q (_________36805));
  xnr2s1 ____0__498633(.DIN1 (____9_9__37984), .DIN2 (_________36675),
       .Q (______9__36774));
  xor2s1 ____9__498634(.DIN1 (_________22015), .DIN2 (_________36673),
       .Q (_________36796));
  dffacs1 _______________________________________________498635(.CLRB
       (reset), .CLK (clk), .DIN (_________36710), .QN
       (_____________________________________________21768));
  nor2s1 ____9_498636(.DIN1 (____90___32382), .DIN2 (_____00__37663),
       .Q (_________36752));
  nnd2s1 _______498637(.DIN1 (______9__36696), .DIN2 (___0_____40100),
       .Q (_________36751));
  xor2s1 ____9__498638(.DIN1
       (_________________________________________________________________________________________22091),
       .DIN2 (_________36658), .Q (_________36750));
  nnd2s1 _______498639(.DIN1 (_________36743), .DIN2 (_________36748),
       .Q (_________36749));
  nnd2s1 _______498640(.DIN1 (______0__36746), .DIN2 (______9__36745),
       .Q (_________36747));
  nnd2s1 _______498641(.DIN1 (_________36743), .DIN2 (_________36742),
       .Q (_________36744));
  xor2s1 ____498642(.DIN1 (_________35848), .DIN2 (_____90__36717), .Q
       (_________36741));
  xor2s1 ____9__498643(.DIN1 (____900__32381), .DIN2 (_________36739),
       .Q (_________36740));
  or2s1 ____9__498644(.DIN1 (________24499), .DIN2 (_________36690), .Q
       (_________36738));
  nor2s1 _____498645(.DIN1 (_________33014), .DIN2 (_________36693), .Q
       (_____0___36921));
  and2s1 ____9__498646(.DIN1 (____0_9__38101), .DIN2
       (_________________________________________9___21803), .Q
       (_________36785));
  nor2s1 ____9__498647(.DIN1
       (_________________________________________9___21803), .DIN2
       (____0_9__38101), .Q (_________36772));
  xor2s1 _______498648(.DIN1 (_____9___36720), .DIN2 (____99___36178),
       .Q (_________36771));
  xor2s1 ____9__498649(.DIN1 (_________36663), .DIN2 (____0____40796),
       .Q (___0_____40125));
  nor2s1 ____0_498650(.DIN1 (_________36567), .DIN2 (_________36678),
       .Q (_________36737));
  hi1s1 ____498651(.DIN (_____09__36735), .Q (______0__36736));
  nor2s1 ____00_498652(.DIN1 (_________36682), .DIN2 (_____0___36733),
       .Q (_____0___36734));
  nor2s1 ____0_498653(.DIN1 (_________36684), .DIN2 (_________36685),
       .Q (_____0___36732));
  hi1s1 ____498654(.DIN (_____0___36730), .Q (_____0___36731));
  nnd2s1 ____0__498655(.DIN1 (_____0___36728), .DIN2 (______9__36676),
       .Q (_____0___36729));
  nor2s1 ____0__498656(.DIN1 (_____9___34923), .DIN2 (_____00__36726),
       .Q (_____0___36727));
  xor2s1 ____9_498657(.DIN1 (_____9___36724), .DIN2 (_____9___36725),
       .Q (______0__36775));
  xor2s1 ____0__498658(.DIN1 (_________36656), .DIN2 (_________38242),
       .Q (_________36937));
  dffacs1 _____________________________________________9_498659(.CLRB
       (reset), .CLK (clk), .DIN (______9__36686), .Q (___0_____40498));
  dffacs1 _______________________________________________498660(.CLRB
       (reset), .CLK (clk), .DIN (_________36679), .Q
       (_____________________________________________21782));
  xor2s1 ____9__498661(.DIN1 (_________36475), .DIN2 (_____9___36724),
       .Q (_________38142));
  dffacs1 __________________498662(.CLRB (reset), .CLK (clk), .DIN
       (_________36692), .QN
       (_________________________________________________________________________________________22090));
  nor2s1 ____00_498663(.DIN1 (_________36441), .DIN2 (_____9___36724),
       .Q (_____9___36723));
  nor2s1 _______498664(.DIN1 (_____9___36721), .DIN2 (_____9___36720),
       .Q (_____9___36722));
  nor2s1 _______498665(.DIN1 (_________36667), .DIN2 (______9__36745),
       .Q (_____9___36719));
  and2s1 ____9_498666(.DIN1 (_____90__36717), .DIN2 (_____0___35837),
       .Q (_____9___36718));
  nnd2s1 ____99_498667(.DIN1 (_____9___36724), .DIN2 (_________38767),
       .Q (______9__36716));
  nnd2s1 ____9__498668(.DIN1 (______9__36668), .DIN2 (___0_____31340),
       .Q (_________36715));
  or2s1 ____9__498669(.DIN1 (_________36661), .DIN2 (_________36713),
       .Q (_________36714));
  nor2s1 ____9__498670(.DIN1 (____90___32384), .DIN2 (_________36739),
       .Q (_________36712));
  nnd2s1 ____9__498671(.DIN1 (______0__36669), .DIN2 (clk), .Q
       (_________36711));
  nnd2s1 ____9_498672(.DIN1 (_________36657), .DIN2 (________22827), .Q
       (_________36710));
  nor2s1 ____9_498673(.DIN1 (_________38767), .DIN2 (_____9___36724),
       .Q (_________36709));
  nor2s1 ____99_498674(.DIN1 (______9__36579), .DIN2 (_________36655),
       .Q (_________36764));
  dffacs1 _______________________________________________498675(.CLRB
       (reset), .CLK (clk), .DIN (_________36662), .QN
       (_____________________________________________21869));
  dffacs1 _____________________________________________0_498676(.CLRB
       (reset), .CLK (clk), .DIN (_________36664), .QN
       (___0__0__40521));
  dffacs1 ________________498677(.CLRB (reset), .CLK (clk), .DIN
       (______9__36706), .Q (outData[12]));
  xor2s1 ____0__498678(.DIN1 (______0__22018), .DIN2 (_____9__28972),
       .Q (_________36708));
  nnd2s1 ____0_498679(.DIN1 (______9__36706), .DIN2 (_________36699),
       .Q (______0__36707));
  xor2s1 ____0_498680(.DIN1 (______0__36677), .DIN2 (___0_____40308),
       .Q (_________36705));
  nnd2s1 ____0__498681(.DIN1 (_____9___36724), .DIN2 (______0__36428),
       .Q (_________36704));
  nnd2s1 ____0__498682(.DIN1 (_________36649), .DIN2 (___99_0__39864),
       .Q (_________36703));
  or2s1 ____0__498683(.DIN1 (_________22015), .DIN2 (_________36652),
       .Q (_________36702));
  or2s1 ____0__498684(.DIN1 (____0____37165), .DIN2 (_________36650),
       .Q (_________36701));
  nor2s1 ____0__498685(.DIN1 (_________36647), .DIN2 (________23452),
       .Q (_________36700));
  nor2s1 ____0__498686(.DIN1 (_________36699), .DIN2 (_____9___36724),
       .Q (_____0___36730));
  nor2s1 ____0__498687(.DIN1 (_________36429), .DIN2 (______9__36706),
       .Q (_____09__36735));
  nor2s1 ____0__498688(.DIN1 (_________36554), .DIN2 (______9__36706),
       .Q (_____00__36823));
  xor2s1 ____0_498689(.DIN1 (______9__36659), .DIN2 (______0__36697),
       .Q (_________36698));
  xor2s1 ____90_498690(.DIN1 (______9__36613), .DIN2 (_________36617),
       .Q (______9__36696));
  nnd2s1 ____9__498691(.DIN1 (______0__36642), .DIN2 (____99___36179),
       .Q (_________36695));
  xor2s1 ____9__498692(.DIN1 (_________36611), .DIN2 (___0_____40472),
       .Q (_________36694));
  nnd2s1 _______498693(.DIN1 (_____0___36635), .DIN2 (______9__32949),
       .Q (_________36693));
  nnd2s1 ____9__498694(.DIN1 (_________36643), .DIN2 (_____0___36637),
       .Q (_________36692));
  nnd2s1 ____99_498695(.DIN1 (_____0___36636), .DIN2 (_________36584),
       .Q (_________36691));
  and2s1 ____00_498696(.DIN1 (_____0___36634), .DIN2 (_________37744),
       .Q (_________36690));
  hi1s1 ____9__498697(.DIN (_________36689), .Q (_____9___36814));
  xor2s1 ____9__498698(.DIN1 (_________36666), .DIN2
       (_______________________________________________________________0__22010),
       .Q (______0__36746));
  or2s1 ____9_498699(.DIN1 (______0__36687), .DIN2 (_________36688), .Q
       (_________36743));
  nnd2s1 ____9_498700(.DIN1 (_________36688), .DIN2 (______0__36687),
       .Q (_________36742));
  hi1s1 ____00_498701(.DIN (_________36739), .Q (_____00__37663));
  dffacs1 _______________________________________________498702(.CLRB
       (reset), .CLK (clk), .DIN (_____9___36626), .Q (_________22044));
  xor2s1 ____0__498703(.DIN1 (_________36601), .DIN2 (_________36340),
       .Q (____0_9__38101));
  nnd2s1 ____0_498704(.DIN1 (_____99__36631), .DIN2 (_________37405),
       .Q (______9__36686));
  and2s1 ____0_498705(.DIN1 (______9__35888), .DIN2 (______0__22018),
       .Q (_________36685));
  nor2s1 ____0__498706(.DIN1 (______0__22018), .DIN2 (_________31938),
       .Q (_________36684));
  and2s1 ____0__498707(.DIN1 (_________31821), .DIN2 (______0__22018),
       .Q (_________36683));
  nor2s1 ____0__498708(.DIN1 (______0__22018), .DIN2 (_________32145),
       .Q (_________36682));
  xor2s1 ____0_498709(.DIN1 (_________36594), .DIN2 (_________36680),
       .Q (_________36681));
  nnd2s1 ____0__498710(.DIN1 (_____00__36632), .DIN2 (________23373),
       .Q (_________36679));
  nor2s1 ____0__498711(.DIN1 (_________36568), .DIN2 (______0__36677),
       .Q (_________36678));
  nnd2s1 ____0__498712(.DIN1 (_____9___36628), .DIN2 (____0____40794),
       .Q (______9__36676));
  nor2s1 ____09_498713(.DIN1 (________29497), .DIN2 (_____9___36625),
       .Q (_________36675));
  and2s1 ____0__498714(.DIN1 (______0__36651), .DIN2 (_________36672),
       .Q (_________36673));
  nor2s1 _______498715(.DIN1 (_________36576), .DIN2 (_____90__36623),
       .Q (_____00__36726));
  dffacs1 _______________________________________________498716(.CLRB
       (reset), .CLK (clk), .DIN (______9__36622), .QN
       (___0_____40507));
  dffacs2 __________________498717(.CLRB (reset), .CLK (clk), .DIN
       (_________36644), .QN
       (_________________________________________________________________________________________22094));
  nor2s1 ____0__498718(.DIN1 (_________36608), .DIN2 (_________36670),
       .Q (_________36671));
  nor2s1 ____0__498719(.DIN1 (______0__36604), .DIN2 (___0____24195),
       .Q (______0__36669));
  nnd2s1 ____9__498720(.DIN1 (_________36605), .DIN2 (_________36870),
       .Q (______9__36668));
  nor2s1 ____9__498721(.DIN1
       (_______________________________________________________________0__22010),
       .DIN2 (_________36666), .Q (_________36667));
  and2s1 ____9__498722(.DIN1 (_________36666), .DIN2
       (_______________________________________________________________0__22010),
       .Q (_________36665));
  nnd2s1 ____9__498723(.DIN1 (_________36606), .DIN2 (_____9___41307),
       .Q (_________36664));
  xor2s1 ____0__498724(.DIN1 (_________36577), .DIN2 (_________36578),
       .Q (_________36663));
  nnd2s1 ____0__498725(.DIN1 (_________36401), .DIN2 (_________36619),
       .Q (_________36662));
  xor2s1 ____0__498726(.DIN1 (________22491), .DIN2
       (_____________________________________________21870), .Q
       (_________36661));
  nnd2s1 ____99_498727(.DIN1 (_________36612), .DIN2 (_________36609),
       .Q (_________36689));
  xor2s1 ____9_498728(.DIN1 (_____09__36641), .DIN2 (_________35904),
       .Q (_____9___36720));
  xor2s1 ____0__498729(.DIN1 (_________36582), .DIN2 (___9_0___39624),
       .Q (_____90__36717));
  nnd2s1 ____9__498730(.DIN1 (_________36615), .DIN2 (_________36616),
       .Q (______9__36745));
  xor2s1 ____0__498731(.DIN1 (____0____40798), .DIN2 (______9__36903),
       .Q (_________36739));
  nor2s1 ____0__498732(.DIN1 (______9__36659), .DIN2
       (_______________22072), .Q (______0__36660));
  nnd2s1 ____0__498733(.DIN1 (_________36556), .DIN2 (______9__36659),
       .Q (_________36658));
  nnd2s1 ____0__498734(.DIN1 (_________36602), .DIN2 (____0____37167),
       .Q (_________36657));
  xor2s1 ______498735(.DIN1 (______0__36570), .DIN2 (_________38876),
       .Q (_________36656));
  nor2s1 ____0__498736(.DIN1 (______0__36580), .DIN2 (____0____40796),
       .Q (_________36655));
  xor2s1 ____0__498737(.DIN1
       (_____________________________________________21800), .DIN2
       (_________36653), .Q (_________36654));
  hi1s1 ____0__498738(.DIN (______0__36651), .Q (_________36652));
  xor2s1 _____0_498739(.DIN1 (_________34588), .DIN2 (____0_0__40800),
       .Q (_________36650));
  nor2s1 ______498740(.DIN1 (_________36648), .DIN2 (_________36620),
       .Q (_________36649));
  xnr2s1 _______498741(.DIN1 (_____9___36627), .DIN2
       (_____________________________________________21767), .Q
       (_________36647));
  hi1s1 ____0__498742(.DIN (_________36646), .Q (______9__36706));
  nb1s1 ____0__498743(.DIN (_________36646), .Q (_____9___36724));
  nor2s1 ____0__498744(.DIN1
       (_____________________________________________21870), .DIN2
       (_________36762), .Q (_________36645));
  nnd2s1 ____9__498745(.DIN1 (_________36643), .DIN2 (_________36591),
       .Q (_________36644));
  nnd2s1 ____00_498746(.DIN1 (_____09__36641), .DIN2 (____99___36173),
       .Q (______0__36642));
  nor2s1 ____0__498747(.DIN1 (_____0___36639), .DIN2 (_____0___36638),
       .Q (_____0___36640));
  nor2s1 ____0__498748(.DIN1 (_________36587), .DIN2 (__99____30477),
       .Q (_____0___36637));
  nnd2s1 ____0_498749(.DIN1 (_________36586), .DIN2 (____0____35309),
       .Q (_____0___36636));
  nor2s1 _____9_498750(.DIN1 (_________32806), .DIN2 (_________36593),
       .Q (_____0___36635));
  xor2s1 ____0__498751(.DIN1 (_________36555), .DIN2 (________22381),
       .Q (_____0___36634));
  or2s1 ____09_498752(.DIN1 (_____________22079), .DIN2
       (_____0___36633), .Q (_________36672));
  nnd2s1 ____498753(.DIN1 (_____0___36633), .DIN2 (_____________22079),
       .Q (______0__36651));
  xor2s1 ____0__498754(.DIN1 (_________36563), .DIN2
       (______________22103), .Q (_________36646));
  xor2s1 ____0__498755(.DIN1 (_________36559), .DIN2 (_____9___36540),
       .Q (______0__36687));
  nnd2s1 _______498756(.DIN1 (_________36571), .DIN2 (_________38249),
       .Q (_____00__36632));
  nor2s1 _____0_498757(.DIN1 (___90___29556), .DIN2 (_________36574),
       .Q (_____99__36631));
  xnr2s1 _______498758(.DIN1 (______0__37325), .DIN2 (_____9___36629),
       .Q (_____9___36630));
  or2s1 _______498759(.DIN1
       (_____________________________________________21767), .DIN2
       (_____9___36627), .Q (_____9___36628));
  nnd2s1 _______498760(.DIN1 (_________36572), .DIN2 (_________37722),
       .Q (_____9___36626));
  xor2s1 _______498761(.DIN1 (______0__36551), .DIN2 (____9____37036),
       .Q (_____9___36625));
  nor2s1 _____0_498762(.DIN1 (_________41090), .DIN2 (_________36575),
       .Q (_____9___36624));
  nor2s1 _______498763(.DIN1 (_________36573), .DIN2 (_____0___36549),
       .Q (_____90__36623));
  nnd2s1 _______498764(.DIN1 (______9__36569), .DIN2 (_________36621),
       .Q (______9__36622));
  and2s1 _______498765(.DIN1 (____0_0__40800), .DIN2 (_________34546),
       .Q (_________36674));
  dffacs1 _________________________________________9_____498766(.CLRB
       (reset), .CLK (clk), .DIN (_________36592), .Q
       (_____________________________________9_______21878));
  hi1s1 _______498767(.DIN (_________36620), .Q (______0__36677));
  dffacs1 _______________________________________________498768(.CLRB
       (reset), .CLK (clk), .DIN (_________36581), .QN
       (______0__22018));
  or2s1 ____0__498769(.DIN1 (_________36562), .DIN2 (_________36618),
       .Q (_________36619));
  nnd2s1 ____498770(.DIN1 (______0__36614), .DIN2 (_________36616), .Q
       (_________36617));
  nnd2s1 ____0__498771(.DIN1 (______0__36614), .DIN2 (______9__36613),
       .Q (_________36615));
  nnd2s1 ____0__498772(.DIN1 (_________36610), .DIN2 (___0_____40472),
       .Q (_________36612));
  and2s1 ____0__498773(.DIN1 (_________36610), .DIN2 (_________36609),
       .Q (_________36611));
  nor2s1 ____0__498774(.DIN1 (_____9__22432), .DIN2 (______9__36603),
       .Q (_________36608));
  nnd2s1 ____9_498775(.DIN1 (_________36564), .DIN2 (inData[6]), .Q
       (_________36607));
  nnd2s1 ____0__498776(.DIN1 (______9__36560), .DIN2 (______9__37314),
       .Q (_________36606));
  xor2s1 ____0__498777(.DIN1 (____990__35280), .DIN2 (_________36585),
       .Q (_________36605));
  nor2s1 ____0__498778(.DIN1 (_________36483), .DIN2 (______9__36603),
       .Q (______0__36604));
  hi1s1 ____0__498779(.DIN
       (_____________________________________________21870), .Q
       (______9__36659));
  hi1s1 ____0_498780(.DIN (_____09__36641), .Q (_________36666));
  xor2s1 _______498781(.DIN1 (_________36528), .DIN2 (_________36552),
       .Q (_________36602));
  xor2s1 _______498782(.DIN1 (______0__36526), .DIN2
       (__________________________________9__________), .Q
       (_________36601));
  xor2s1 ______498783(.DIN1
       (_________________________________________0___21814), .DIN2
       (______0__36589), .Q (_________36600));
  hi1s1 _______498784(.DIN (_________36595), .Q (_________36596));
  xor2s1 _______498785(.DIN1
       (_____________________________________________21781), .DIN2
       (_____9___36721), .Q (_________36594));
  nnd2s1 _______498786(.DIN1 (_________36553), .DIN2 (_________36412),
       .Q (_________36620));
  dffacs1 _______________________________________________498787(.CLRB
       (reset), .CLK (clk), .DIN (_________36557), .QN
       (___0_9___40556));
  nnd2s1 ____9_498788(.DIN1 (_____9___36542), .DIN2 (______9__32645),
       .Q (_________36593));
  nnd2s1 ____9__498789(.DIN1 (_____00__36544), .DIN2 (_____0__23797),
       .Q (_________36592));
  nor2s1 ____0_498790(.DIN1 (_____99__36543), .DIN2 (__99_0__30479), .Q
       (_________36591));
  and2s1 _______498791(.DIN1 (______0__36589), .DIN2
       (_________________________________________0___21814), .Q
       (_________36590));
  nor2s1 ______498792(.DIN1
       (_________________________________________0___21814), .DIN2
       (______0__36589), .Q (______9__36588));
  nor2s1 ____0__498793(.DIN1 (_____9___36536), .DIN2 (_________35966),
       .Q (_________36587));
  nnd2s1 ____0_498794(.DIN1 (_________36585), .DIN2 (_________36583),
       .Q (_________36586));
  or2s1 ____0__498795(.DIN1 (_________36583), .DIN2 (_________36585),
       .Q (_________36584));
  nor2s1 ____09_498796(.DIN1 (_________35686), .DIN2 (_____9___36539),
       .Q (_________36582));
  nnd2s1 ______498797(.DIN1 (_____0___36545), .DIN2 (________26826), .Q
       (_________36581));
  and2s1 _____0_498798(.DIN1 (_________37494), .DIN2 (_________32014),
       .Q (______0__36580));
  nor2s1 _____0_498799(.DIN1 (_________36578), .DIN2 (_________37494),
       .Q (______9__36579));
  and2s1 _______498800(.DIN1 (_________37494), .DIN2 (_____9___36725),
       .Q (_________36577));
  nnd2s1 ____0__498801(.DIN1 (_____9___36541), .DIN2 (_________36558),
       .Q (______0__36970));
  xor2s1 ____0__498802(.DIN1 (_________36514), .DIN2 (_____0___36462),
       .Q (_____09__36641));
  dffacs1 _______________________________________________498803(.CLRB
       (reset), .CLK (clk), .DIN (_____9___36537), .Q
       (_____________________________________________21870));
  nor2s1 _____498804(.DIN1
       (_____________________________________________21781), .DIN2
       (_________36680), .Q (_________36576));
  xor2s1 ______498805(.DIN1 (____09___34474), .DIN2 (_____0___36546),
       .Q (_________36575));
  and2s1 _______498806(.DIN1 (_________36529), .DIN2 (_________37317),
       .Q (_________36574));
  and2s1 _____9_498807(.DIN1 (_________36680), .DIN2
       (_____________________________________________21781), .Q
       (_________36573));
  nor2s1 ______498808(.DIN1 (________24521), .DIN2 (______9__36525), .Q
       (_________36572));
  xor2s1 _____0_498809(.DIN1 (_________35093), .DIN2 (____0____40804),
       .Q (_________36571));
  xor2s1 _____0_498810(.DIN1 (______0__35957), .DIN2 (____0____40802),
       .Q (______0__36570));
  nor2s1 _______498811(.DIN1 (___0_9__26991), .DIN2 (_________36522),
       .Q (______9__36569));
  nnd2s1 _______498812(.DIN1
       (_____________________________________________21781), .DIN2
       (____0_0__36258), .Q (_____9___36627));
  or2s1 _______498813(.DIN1 (_________36568), .DIN2 (_________36567),
       .Q (_________36648));
  nor2s1 _______498814(.DIN1 (___0_____40535), .DIN2 (______0__36589),
       .Q (_____0___36639));
  and2s1 _______498815(.DIN1 (______0__36589), .DIN2 (___0_____40535),
       .Q (_____0___36638));
  xor2s1 ______498816(.DIN1 (______9__36507), .DIN2 (___9_____39688),
       .Q (_________36595));
  nor2s1 _______498817(.DIN1 (________22417), .DIN2 (______9__36534),
       .Q (_____0___36633));
  nnd2s1 _______498818(.DIN1 (_________36566), .DIN2 (_________36565),
       .Q (_________37802));
  dffacs1 _______________________________________________498819(.CLRB
       (reset), .CLK (clk), .DIN (_________36530), .QN
       (_____________________________________________21800));
  nor2s1 ____9_498820(.DIN1 (_________36509), .DIN2 (___0_____40166),
       .Q (_________36564));
  xor2s1 _______498821(.DIN1 (___0_____40589), .DIN2 (_________36533),
       .Q (_________36563));
  xnr2s1 _____498822(.DIN1
       (_________________________________________________________________________________________22090),
       .DIN2 (______0__36561), .Q (_________36562));
  xor2s1 _______498823(.DIN1 (_________35687), .DIN2 (_____9___36538),
       .Q (______9__36560));
  and2s1 _______498824(.DIN1 (_________36558), .DIN2 (_________36518),
       .Q (_________36559));
  or2s1 _______498825(.DIN1 (_________38583), .DIN2 (_________36519),
       .Q (_________36557));
  nnd2s1 _______498826(.DIN1 (_________36513), .DIN2 (_________36474),
       .Q (______9__36603));
  nnd2s1 ____09_498827(.DIN1 (______0__36516), .DIN2 (_________36556),
       .Q (_________36610));
  xnr2s1 ____0__498828(.DIN1 (___009___39979), .DIN2 (_________36500),
       .Q (______0__36614));
  nnd2s1 _______498829(.DIN1 (_________36510), .DIN2 (_________36554),
       .Q (_________36555));
  nnd2s1 _______498830(.DIN1 (_________36552), .DIN2 (_________36414),
       .Q (_________36553));
  nnd2s1 _______498831(.DIN1 (____0____40802), .DIN2 (____09___35375),
       .Q (______0__36551));
  xor2s1 _____0_498832(.DIN1 (_____0___36549), .DIN2 (_________38385),
       .Q (_____0___36550));
  and2s1 _______498833(.DIN1 (____0____40804), .DIN2 (_________35073),
       .Q (______9__36597));
  nnd2s1 _______498834(.DIN1 (_____0___36548), .DIN2 (_____0___36547),
       .Q (_________37552));
  nor2s1 _______498835(.DIN1 (____09___34472), .DIN2 (_____0___36546),
       .Q (_________36599));
  nnd2s1 _______498836(.DIN1 (______0__36508), .DIN2 (_____0___36460),
       .Q (______0__37325));
  dffacs1 _______________________________________________498837(.CLRB
       (reset), .CLK (clk), .DIN (_________36506), .QN
       (______0__22040));
  nor2s1 ______498838(.DIN1 (__9__9__30047), .DIN2 (______0__36491), .Q
       (_____0___36545));
  or2s1 ____0_498839(.DIN1 (____9_9__37052), .DIN2 (_________36503), .Q
       (_____00__36544));
  and2s1 ____0_498840(.DIN1 (_________36288), .DIN2 (_________36502),
       .Q (_____99__36543));
  nor2s1 ____00_498841(.DIN1 (____0____36262), .DIN2 (_________36505),
       .Q (_____9___36542));
  or2s1 _____498842(.DIN1 (_____9___36540), .DIN2 (_________36517), .Q
       (_____9___36541));
  and2s1 _______498843(.DIN1 (_____9___36538), .DIN2 (_________35682),
       .Q (_____9___36539));
  nnd2s1 _______498844(.DIN1 (______9__36498), .DIN2 (___000___30551),
       .Q (_____9___36537));
  nor2s1 _______498845(.DIN1 (_________36497), .DIN2 (______0__36561),
       .Q (_____9___36536));
  and2s1 _______498846(.DIN1 (_________36486), .DIN2 (____9____37049),
       .Q (_____90__36535));
  nor2s1 ______498847(.DIN1 (_____9__22488), .DIN2 (_________36533), .Q
       (______9__36534));
  nnd2s1 ____09_498848(.DIN1 (______9__36515), .DIN2
       (___________9___22071), .Q (_________36609));
  xor2s1 _______498849(.DIN1 (_________36469), .DIN2 (_________38242),
       .Q (_________36585));
  xor2s1 _______498850(.DIN1 (_________36464), .DIN2 (_________36856),
       .Q (_________37494));
  and2s1 _____9_498851(.DIN1 (_________36531), .DIN2 (_________36523),
       .Q (_________36532));
  and2s1 _____9_498852(.DIN1 (_________36485), .DIN2 (_________38262),
       .Q (_________36530));
  xor2s1 _____0_498853(.DIN1 (____0____34445), .DIN2 (_____0___36456),
       .Q (_________36529));
  xor2s1 _____0_498854(.DIN1 (_____0___36457), .DIN2 (_________36527),
       .Q (_________36528));
  xor2s1 _____498855(.DIN1 (_____0___36461), .DIN2 (____9____38007), .Q
       (______0__36526));
  nor2s1 _______498856(.DIN1 (_____9___37656), .DIN2 (_________36492),
       .Q (______9__36525));
  or2s1 _____9_498857(.DIN1 (_________36523), .DIN2 (_________36531),
       .Q (_________36524));
  nor2s1 ______498858(.DIN1 (_________36521), .DIN2 (_________36484),
       .Q (_________36522));
  nnd2s1 _______498859(.DIN1 (_________36520), .DIN2 (___0_____40483),
       .Q (_________36565));
  dffacs1 ____________________________________0_498860(.CLRB (reset),
       .CLK (clk), .DIN (_________36504), .Q (___0_9___40454));
  or2s1 ______498861(.DIN1 (___0_____40483), .DIN2 (_________36520), .Q
       (_________36566));
  nor2s1 _______498862(.DIN1 (___0_0___40566), .DIN2 (_________36520),
       .Q (_________36567));
  xor2s1 _______498863(.DIN1 (_____0___36455), .DIN2 (_____9___36003),
       .Q (______0__36589));
  dffacs1 _______________________________________________498864(.CLRB
       (reset), .CLK (clk), .DIN (_________36478), .QN
       (_____________________________________________21781));
  xor2s1 _____0_498865(.DIN1 (_________36436), .DIN2 (____0____40808),
       .Q (_________36519));
  hi1s1 _______498866(.DIN (_________36517), .Q (_________36518));
  hi1s1 _______498867(.DIN (______9__36515), .Q (______0__36516));
  xor2s1 ______498868(.DIN1 (_________36443), .DIN2 (____9____38909),
       .Q (_________36514));
  or2s1 ______498869(.DIN1
       (______________________________________0______21886), .DIN2
       (______0__36473), .Q (_________36513));
  xor2s1 _____0_498870(.DIN1 (_________36445), .DIN2 (_________41341),
       .Q (_________36510));
  xor2s1 ____0__498871(.DIN1 (___0____22339), .DIN2
       (_________________________________________0___21968), .Q
       (_________36509));
  nnd2s1 _____498872(.DIN1 (____9_0__36140), .DIN2 (_____99__36454), .Q
       (______0__36508));
  nor2s1 _______498873(.DIN1 (______9__36447), .DIN2 (_________36523),
       .Q (______9__36507));
  nnd2s1 _______498874(.DIN1 (_________36467), .DIN2 (____0____37147),
       .Q (_________36506));
  nor2s1 _______498875(.DIN1 (____0____34418), .DIN2 (_________36466),
       .Q (_____0___36546));
  nor2s1 _______498876(.DIN1 (_________36314), .DIN2 (______0__36463),
       .Q (_________36552));
  nnd2s1 _______498877(.DIN1 (_________37735), .DIN2 (________22669),
       .Q (_____0___36547));
  nor2s1 _______498878(.DIN1 (_________36883), .DIN2 (_________36477),
       .Q (_________36568));
  xor2s1 _______498879(.DIN1 (___________________), .DIN2
       (_________36476), .Q (_________37341));
  nnd2s1 ____0__498880(.DIN1 (_____9___36450), .DIN2 (____0____36256),
       .Q (_________36505));
  nnd2s1 _____0_498881(.DIN1 (________23899), .DIN2
       (_________________________________________0___21968), .Q
       (_________36504));
  xor2s1 _______498882(.DIN1 (_________36423), .DIN2 (_____9___36448),
       .Q (_________36503));
  nnd2s1 _______498883(.DIN1 (___09____40675), .DIN2 (inData[2]), .Q
       (_________36502));
  nor2s1 _______498884(.DIN1 (_________36442), .DIN2 (____9____37049),
       .Q (_________36501));
  nor2s1 ______498885(.DIN1
       (_____________________________________________21953), .DIN2
       (_________36495), .Q (_________36500));
  xor2s1 ______498886(.DIN1 (_________36406), .DIN2 (___0_____40537),
       .Q (______0__36499));
  or2s1 _____9_498887(.DIN1 (______0__36766), .DIN2 (_________36444),
       .Q (______9__36498));
  and2s1 ______498888(.DIN1 (_________36493), .DIN2 (___0_____40472),
       .Q (_________36497));
  xor2s1 _______498889(.DIN1 (____0____40806), .DIN2 (___99_9__39836),
       .Q (_____9___36538));
  nor2s1 _______498890(.DIN1 (_________36494), .DIN2 (_________36495),
       .Q (_________36517));
  nnd2s1 _______498891(.DIN1 (_____9___36449), .DIN2 (______0__36404),
       .Q (______9__36515));
  nnd2s1 _______498892(.DIN1 (_________36495), .DIN2 (_________36494),
       .Q (_________36558));
  nnd2s1 _______498893(.DIN1 (_________36495), .DIN2
       (_____________________________________________21953), .Q
       (_________36616));
  nor2s1 ______498894(.DIN1 (___0_____40472), .DIN2 (_________36493),
       .Q (______0__36561));
  xor2s1 ______498895(.DIN1 (____9____36141), .DIN2 (_____0___36459),
       .Q (_________36492));
  nor2s1 ______498896(.DIN1 (_________36482), .DIN2 (__9_____30046), .Q
       (______0__36491));
  nnd2s1 _______498897(.DIN1 (_________36435), .DIN2 (_________38576),
       .Q (______9__36490));
  and2s1 _______498898(.DIN1 (_____9___36451), .DIN2 (____9_0__37080),
       .Q (_________36489));
  or2s1 _______498899(.DIN1 (________23907), .DIN2 (_________36487), .Q
       (_________36488));
  xor2s1 _______498900(.DIN1 (____0____34420), .DIN2 (_________36465),
       .Q (_________36486));
  xor2s1 ______498901(.DIN1 (______0__36410), .DIN2 (_________36432),
       .Q (_________36485));
  xor2s1 _______498902(.DIN1 (_________36407), .DIN2 (___9_____39542),
       .Q (_________36484));
  and2s1 _______498903(.DIN1
       (______________________________________0______21886), .DIN2
       (_________36482), .Q (_________36483));
  nor2s1 _______498904(.DIN1 (_________37687), .DIN2 (_________36430),
       .Q (______0__36481));
  nnd2s1 ______498905(.DIN1 (_________36431), .DIN2 (____0___24459), .Q
       (_________36478));
  nor2s1 ______498906(.DIN1 (______9__36384), .DIN2 (_________36433),
       .Q (_____0___36549));
  nnd2s1 _______498907(.DIN1 (_____9___36452), .DIN2 (__________22059),
       .Q (_____0___36548));
  nor2s1 _______498908(.DIN1 (_________36391), .DIN2 (_________36440),
       .Q (_________36533));
  hi1s1 _____9_498909(.DIN (_________36477), .Q (_________36520));
  nor2s1 _______498910(.DIN1 (_________36418), .DIN2 (_________36476),
       .Q (_________36531));
  nnd2s1 ______498911(.DIN1 (_________36415), .DIN2 (_________36417),
       .Q (_________36475));
  or2s1 ______498912(.DIN1
       (______________________________________0__0_), .DIN2
       (______________________________________0______21885), .Q
       (_________36474));
  nnd2s1 _______498913(.DIN1
       (______________________________________0______21885), .DIN2
       (______________________________________0__0_), .Q
       (______0__36473));
  nor2s1 _______498914(.DIN1 (_________36471), .DIN2 (_________36470),
       .Q (______9__36472));
  nnd2s1 ______498915(.DIN1 (_________36421), .DIN2 (_________35038),
       .Q (_________36469));
  nor2s1 _______498916(.DIN1 (_________36439), .DIN2 (______9__36419),
       .Q (_________36468));
  nor2s1 _______498917(.DIN1 (_________36411), .DIN2 (_________35662),
       .Q (_________36467));
  nor2s1 _______498918(.DIN1 (____0____34419), .DIN2 (_________36465),
       .Q (_________36466));
  xor2s1 _______498919(.DIN1 (____090__40810), .DIN2 (_____9___36363),
       .Q (_________36464));
  and2s1 ______498920(.DIN1 (____0____40808), .DIN2 (_________36298),
       .Q (______0__36463));
  and2s1 _______498921(.DIN1 (_____0___36462), .DIN2 (_________36397),
       .Q (_________36511));
  nnd2s1 ____0_498922(.DIN1 (_________36425), .DIN2 (____0____36264),
       .Q (_________36688));
  xor2s1 _______498923(.DIN1 (_________36378), .DIN2 (_____9___36725),
       .Q (_____0___36461));
  nnd2s1 _______498924(.DIN1 (_____0___36459), .DIN2 (___0_____40519),
       .Q (_____0___36460));
  xor2s1 ______498925(.DIN1 (_________36386), .DIN2 (___9_____39554),
       .Q (_____0___36458));
  xor2s1 _______498926(.DIN1 (______9__36437), .DIN2 (___0_0___40567),
       .Q (_____0___36457));
  xor2s1 _______498927(.DIN1 (_________36426), .DIN2 (_____9___41303),
       .Q (_____0___36456));
  xor2s1 _______498928(.DIN1 (_________36377), .DIN2 (________27618),
       .Q (_____0___36455));
  or2s1 ______498929(.DIN1 (___0_____40519), .DIN2 (_____0___36459), .Q
       (_____99__36454));
  xor2s1 _______498930(.DIN1 (_________36379), .DIN2 (_________37789),
       .Q (_________36477));
  hi1s1 _____9_498931(.DIN (_____9___36453), .Q (_________36523));
  hi1s1 _____9_498932(.DIN (_____9___36452), .Q (_________37735));
  xor2s1 _____498933(.DIN1 (_________36353), .DIN2 (_________36356), .Q
       (_____9___36451));
  xor2s1 _______498934(.DIN1 (____0____36261), .DIN2 (_________36424),
       .Q (_____9___36450));
  or2s1 _______498935(.DIN1 (______9__36403), .DIN2 (_____9___36448),
       .Q (_____9___36449));
  nor2s1 _____9_498936(.DIN1 (______9__36427), .DIN2 (_________36446),
       .Q (______9__36447));
  nnd2s1 _______498937(.DIN1 (_________36434), .DIN2 (_____9___36359),
       .Q (_________36445));
  xor2s1 _______498938(.DIN1 (_________35052), .DIN2 (_________36420),
       .Q (_________36444));
  nor2s1 _______498939(.DIN1 (_____0___36371), .DIN2 (_________36399),
       .Q (_________36443));
  nor2s1 _______498940(.DIN1 (___9_0__29602), .DIN2 (_________36392),
       .Q (_________36442));
  hi1s1 ______498941(.DIN (_________36554), .Q (_________36441));
  nor2s1 _______498942(.DIN1 (______0__34897), .DIN2 (_________36395),
       .Q (_________36440));
  nnd2s1 _______498943(.DIN1 (_________36396), .DIN2 (_________36439),
       .Q (_________36496));
  hi1s1 ______498944(.DIN
       (______________________________________0______21885), .Q
       (_________36482));
  dffacs1 _____________________________________________0_498945(.CLRB
       (reset), .CLK (clk), .DIN (_________36393), .Q
       (_________________________________________0___21968));
  xor2s1 _______498946(.DIN1 (_____0___36367), .DIN2 (___9_____39511),
       .Q (_________36495));
  dffacs1 _______________________________________________498947(.CLRB
       (reset), .CLK (clk), .DIN (_________36400), .Q (___0_____40472));
  nnd2s1 _______498948(.DIN1 (______9__36437), .DIN2 (___0_____40484),
       .Q (______0__36438));
  xor2s1 _______498949(.DIN1 (_________36350), .DIN2 (___0_0___40568),
       .Q (_________36436));
  xor2s1 _____0_498950(.DIN1 (____0____36243), .DIN2 (______0__36348),
       .Q (_________36435));
  dffacs1 ________________498951(.CLRB (reset), .CLK (clk), .DIN
       (_________36434), .Q (outData[11]));
  nor2s1 _______498952(.DIN1 (_________36383), .DIN2 (_________36432),
       .Q (_________36433));
  nnd2s1 _______498953(.DIN1 (_________36380), .DIN2 (_________38576),
       .Q (_________36431));
  or2s1 _______498954(.DIN1 (___0_____40484), .DIN2 (______9__36437),
       .Q (_________36430));
  and2s1 _____0_498955(.DIN1 (_________36434), .DIN2 (______0__36428),
       .Q (_________36429));
  nor2s1 _______498956(.DIN1 (_________36416), .DIN2 (_________36434),
       .Q (_________36699));
  nnd2s1 _______498957(.DIN1 (_________36446), .DIN2 (______9__36427),
       .Q (_____9___36453));
  xor2s1 _______498958(.DIN1 (______9__36347), .DIN2 (________27618),
       .Q (_____9___36452));
  xor2s1 ______498959(.DIN1 (___0_____40484), .DIN2 (_________36413),
       .Q (_________36487));
  nnd2s1 _______498960(.DIN1 (_________36426), .DIN2 (____0____34416),
       .Q (_________36479));
  nor2s1 _______498961(.DIN1 (_________37937), .DIN2 (_________36434),
       .Q (_________36476));
  dffacs1 _______________________________________________498962(.CLRB
       (reset), .CLK (clk), .DIN (_________36381), .Q
       (_____________________________________________21839));
  dffacs1 _______________________________________________498963(.CLRB
       (reset), .CLK (clk), .DIN (_____0___36373), .QN
       (_____________________________________________21825));
  nnd2s1 _______498964(.DIN1 (_________36424), .DIN2 (______0__36338),
       .Q (_________36425));
  xor2s1 _____0_498965(.DIN1
       (_________________________________________________________________________________________22091),
       .DIN2 (___0_____40473), .Q (_________36423));
  nnd2s1 _______498966(.DIN1 (_____9___36362), .DIN2 (_________36670),
       .Q (_________36422));
  or2s1 _______498967(.DIN1 (_________35042), .DIN2 (_________36420),
       .Q (_________36421));
  xor2s1 _____0_498968(.DIN1 (_________________0_), .DIN2
       (_________36323), .Q (______9__36419));
  nor2s1 _____0_498969(.DIN1 (_________36439), .DIN2 (______9__36903),
       .Q (_________36418));
  nnd2s1 _____0_498970(.DIN1 (______9__36903), .DIN2 (_________36416),
       .Q (_________36417));
  or2s1 _____498971(.DIN1 (______0__36428), .DIN2 (______9__36903), .Q
       (_________36415));
  and2s1 _______498972(.DIN1 (______9__36903), .DIN2
       (_____________________________________________21900), .Q
       (_________36470));
  nor2s1 _______498973(.DIN1
       (_____________________________________________21900), .DIN2
       (______9__36903), .Q (_________36471));
  dffacs1 __________________________________________0____498974(.CLRB
       (reset), .CLK (clk), .DIN (_____9___36365), .QN
       (______________________________________0______21885));
  nnd2s1 _______498975(.DIN1 (______9__36903), .DIN2 (_____9___36358),
       .Q (_________36554));
  or2s1 _______498976(.DIN1 (___0_0___40567), .DIN2 (_________36413),
       .Q (_________36414));
  nnd2s1 ______498977(.DIN1 (_________36413), .DIN2 (___0_0___40567),
       .Q (_________36412));
  nor2s1 _______498978(.DIN1 (_________36355), .DIN2 (____9____37049),
       .Q (_________36411));
  xor2s1 _______498979(.DIN1
       (_____________________________________________21780), .DIN2
       (____000__36182), .Q (______0__36410));
  xor2s1 _______498980(.DIN1 (_________36653), .DIN2 (_________36320),
       .Q (_________36407));
  xor2s1 _____498981(.DIN1 (______0__37507), .DIN2 (_________36858), .Q
       (_________36406));
  nnd2s1 _______498982(.DIN1 (_____9___36361), .DIN2 (____0____36202),
       .Q (_____0___36462));
  nor2s1 _______498983(.DIN1 (_________36352), .DIN2 (______9__36357),
       .Q (_________36465));
  nnd2s1 _______498984(.DIN1 (_________36343), .DIN2 (______0__36302),
       .Q (_____0___36459));
  xor2s1 _______498985(.DIN1 (____0___27033), .DIN2 (_____09__36374),
       .Q (_________36405));
  nnd2s1 _______498986(.DIN1 (_________36402), .DIN2 (___0_____40473),
       .Q (______0__36404));
  nor2s1 _______498987(.DIN1 (___0_____40473), .DIN2 (_________36402),
       .Q (______9__36403));
  or2s1 _______498988(.DIN1 (______0__36766), .DIN2 (_________36334),
       .Q (_________36401));
  nnd2s1 _______498989(.DIN1 (_________36336), .DIN2 (_________36643),
       .Q (_________36400));
  nor2s1 _____9_498990(.DIN1 (_____0___36368), .DIN2 (_________36398),
       .Q (_________36399));
  nnd2s1 _____0_498991(.DIN1 (_________36398), .DIN2 (_____0___36370),
       .Q (_________36397));
  xor2s1 _____0_498992(.DIN1 (_________36303), .DIN2
       (___________________), .Q (_________36396));
  nor2s1 _______498993(.DIN1 (________26208), .DIN2 (_________36332),
       .Q (_________36395));
  nnd2s1 _______498994(.DIN1 (______0__37507), .DIN2 (______22120), .Q
       (______0__36394));
  nnd2s1 _______498995(.DIN1 (_________36333), .DIN2 (___9____29563),
       .Q (_________36393));
  xnr2s1 _______498996(.DIN1 (_________36354), .DIN2 (______0__22040),
       .Q (_________36392));
  nor2s1 _______498997(.DIN1 (___9_____39627), .DIN2 (______9__36318),
       .Q (_________36391));
  hi1s1 ______498998(.DIN (_________36390), .Q (_________36446));
  hi1s1 _______498999(.DIN (______9__36903), .Q (_________36434));
  nnd2s1 ______499000(.DIN1 (_________36387), .DIN2 (___0_____40536),
       .Q (_________36389));
  nor2s1 _____9_499001(.DIN1 (___0_____40516), .DIN2 (_________36387),
       .Q (_________36388));
  nor2s1 _____0_499002(.DIN1 (______0__36385), .DIN2 (_________36344),
       .Q (_________36386));
  and2s1 _______499003(.DIN1 (_________36382), .DIN2
       (_____________________________________________21780), .Q
       (______9__36384));
  nor2s1 _______499004(.DIN1
       (_____________________________________________21780), .DIN2
       (_________36382), .Q (_________36383));
  nnd2s1 _______499005(.DIN1 (_________36322), .DIN2 (___9____25040),
       .Q (_________36381));
  xor2s1 _______499006(.DIN1 (______0__34949), .DIN2 (_________36342),
       .Q (_________36380));
  xor2s1 _______499007(.DIN1 (_________36341), .DIN2 (_____9___36002),
       .Q (_________36379));
  nnd2s1 _______499008(.DIN1 (_________36376), .DIN2 (____09___36273),
       .Q (_________36378));
  nnd2s1 _______499009(.DIN1 (_________36376), .DIN2 (______0__36319),
       .Q (_________36377));
  xor2s1 ______499010(.DIN1 (___0_____40516), .DIN2 (_____09__36374),
       .Q (______0__36375));
  nnd2s1 _______499011(.DIN1 (_________36326), .DIN2 (________24664),
       .Q (_____0___36373));
  xor2s1 _______499012(.DIN1 (_____________________21677), .DIN2
       (_________36294), .Q (_________36426));
  dffacs1 _______________________________________________499013(.CLRB
       (reset), .CLK (clk), .DIN (_________36330), .Q
       (_____________________________________________21838));
  dffacs1 _______________________________________________499014(.CLRB
       (reset), .CLK (clk), .DIN (_________36321), .Q
       (_____________________________________________21836));
  hi1s1 _____499015(.DIN (_________36413), .Q (______9__36437));
  nnd2s1 _______499016(.DIN1 (_____09__36374), .DIN2 (________25838),
       .Q (_____0___36372));
  nor2s1 _______499017(.DIN1 (_____0___36370), .DIN2 (_________37352),
       .Q (_____0___36371));
  nnd2s1 _____9_499018(.DIN1 (_________37352), .DIN2 (_____0___36368),
       .Q (_____0___36369));
  xor2s1 _______499019(.DIN1 (_____09__36286), .DIN2 (_____0___36279),
       .Q (_____0___36367));
  nnd2s1 _______499020(.DIN1 (_________36327), .DIN2 (___0_____40537),
       .Q (_____99__36366));
  nnd2s1 ______499021(.DIN1 (_________36311), .DIN2 (_____9__25009), .Q
       (_____9___36365));
  xnr2s1 ______499022(.DIN1
       (_____________________________________________21899), .DIN2
       (_____9___36363), .Q (_____9___36364));
  xor2s1 ______499023(.DIN1 (_________36316), .DIN2 (_____9___36363),
       .Q (_____9___36362));
  xor2s1 _______499024(.DIN1 (_____0___36280), .DIN2 (_____9___36360),
       .Q (_____9___36361));
  nnd2s1 _______499025(.DIN1 (_________36312), .DIN2 (____00___36187),
       .Q (_________36424));
  nor2s1 _______499026(.DIN1 (______0__36309), .DIN2 (_________36304),
       .Q (_________36416));
  xnr2s1 _______499027(.DIN1 (______9__36337), .DIN2 (_____9___36363),
       .Q (_________36390));
  nnd2s1 _______499028(.DIN1 (_________36306), .DIN2 (____99___36177),
       .Q (_________36420));
  xnr2s1 _______499029(.DIN1 (_________36317), .DIN2 (_________36331),
       .Q (______9__36903));
  hi1s1 _____0_499030(.DIN (_____9___36358), .Q (_____9___36359));
  nor2s1 _______499031(.DIN1 (_________36351), .DIN2 (_________36356),
       .Q (______9__36357));
  nor2s1 _______499032(.DIN1 (_________36293), .DIN2 (_________36354),
       .Q (_________36355));
  nor2s1 _______499033(.DIN1 (_________36352), .DIN2 (_________36351),
       .Q (_________36353));
  xor2s1 ______499034(.DIN1 (_________36315), .DIN2 (_________36349),
       .Q (_________36350));
  xor2s1 ______499035(.DIN1 (____09___36270), .DIN2 (___9_____39784),
       .Q (______0__36348));
  xor2s1 _______499036(.DIN1 (____090__36268), .DIN2 (____9____36135),
       .Q (______9__36347));
  nor2s1 _____9_499037(.DIN1 (______22146), .DIN2 (_____09__36374), .Q
       (_________36346));
  hi1s1 _______499038(.DIN (_________36344), .Q (_________36345));
  or2s1 _______499039(.DIN1 (_________36653), .DIN2 (_________36296),
       .Q (_________36343));
  or2s1 ______499040(.DIN1 (_____9___34925), .DIN2 (_________36342), .Q
       (_________36409));
  or2s1 _______499041(.DIN1 (_________35991), .DIN2 (_________36341),
       .Q (_________36408));
  dffacs1 _______________________________________________499042(.CLRB
       (reset), .CLK (clk), .DIN (_________36299), .Q (___0_90__40551));
  xor2s1 _______499043(.DIN1 (____09___36271), .DIN2 (_________36340),
       .Q (_________36413));
  dffacs1 _______________________________________________499044(.CLRB
       (reset), .CLK (clk), .DIN (_________36313), .Q (___0_____40523));
  xnr2s1 _______499045(.DIN1 (______0__36598), .DIN2 (____0____36259),
       .Q (_________36339));
  xor2s1 _____9_499046(.DIN1 (____0____36255), .DIN2 (______9__36337),
       .Q (______0__36338));
  nor2s1 _______499047(.DIN1 (___000___30549), .DIN2 (_________36289),
       .Q (_________36336));
  dffacs1 ______________0_499048(.CLRB (reset), .CLK (clk), .DIN
       (_____9___36363), .Q (outData[10]));
  and2s1 _______499049(.DIN1 (______0__36287), .DIN2 (_________37317),
       .Q (_________36335));
  xor2s1 ______499050(.DIN1 (____999__36181), .DIN2 (_________36305),
       .Q (_________36334));
  nnd2s1 ______499051(.DIN1 (_____0___36283), .DIN2 (___0_____40100),
       .Q (_________36333));
  and2s1 ______499052(.DIN1 (_________36331), .DIN2 (________26161), .Q
       (_________36332));
  nnd2s1 _____9_499053(.DIN1 (_____00__36278), .DIN2 (__9_9___30365),
       .Q (_________36330));
  or2s1 _____0_499054(.DIN1 (____9____36128), .DIN2 (______9__36328),
       .Q (______0__36329));
  hi1s1 ______499055(.DIN (_________37352), .Q (_________36398));
  dffacs1 _______________________________________________499056(.CLRB
       (reset), .CLK (clk), .DIN (_________36290), .Q (___0_____40473));
  hi1s1 _____0_499057(.DIN (_________36327), .Q (______0__37507));
  nnd2s1 _____9_499058(.DIN1 (____099__36277), .DIN2 (_____9___37752),
       .Q (_________36326));
  and2s1 _______499059(.DIN1 (______9__36328), .DIN2 (____9____36133),
       .Q (_________36325));
  xor2s1 _______499060(.DIN1 (____0____36246), .DIN2 (___0_____40517),
       .Q (_________36324));
  nor2s1 _______499061(.DIN1 (____0____36230), .DIN2 (_____9___36363),
       .Q (_________36323));
  nnd2s1 _______499062(.DIN1 (____09___36272), .DIN2 (_________37223),
       .Q (_________36322));
  nnd2s1 _______499063(.DIN1 (_________35681), .DIN2 (_____0___36281),
       .Q (_________36321));
  xnr2s1 _______499064(.DIN1
       (_____________________________________________21811), .DIN2
       (____09___40812), .Q (_________36320));
  nnd2s1 _______499065(.DIN1 (____09___36274), .DIN2 (_________36340),
       .Q (______0__36319));
  or2s1 _______499066(.DIN1 (_________36317), .DIN2 (_________36331),
       .Q (______9__36318));
  nor2s1 _______499067(.DIN1 (_________36316), .DIN2 (_____9___36363),
       .Q (_____9___36358));
  hi1s1 _______499068(.DIN (_____09__36374), .Q (_________36387));
  and2s1 _______499069(.DIN1 (_________36315), .DIN2
       (_____________________________________________21859), .Q
       (______0__36385));
  nor2s1 _______499070(.DIN1 (____0____36223), .DIN2 (____09___36275),
       .Q (_________36376));
  nor2s1 ______499071(.DIN1
       (_____________________________________________21859), .DIN2
       (_________36315), .Q (_________36344));
  dffacs1 _______________________________________________499072(.CLRB
       (reset), .CLK (clk), .DIN (____09___36276), .Q
       (_____________________________________________21780));
  nor2s1 _______499073(.DIN1 (___0_0___40568), .DIN2 (_________36297),
       .Q (_________36314));
  nnd2s1 _______499074(.DIN1 (____0_9__36257), .DIN2 (_____9___36996),
       .Q (_________36313));
  nor2s1 _______499075(.DIN1 (____00___36190), .DIN2 (____0____36263),
       .Q (_________36312));
  nnd2s1 _______499076(.DIN1 (____0____36251), .DIN2 (_________36670),
       .Q (_________36311));
  or2s1 _______499077(.DIN1
       (_____________________________________________21899), .DIN2
       (______0__36309), .Q (_________36310));
  and2s1 _______499078(.DIN1 (______0__36309), .DIN2
       (_____________________________________________21899), .Q
       (______9__36308));
  nnd2s1 _____9_499079(.DIN1 (____9_9__36171), .DIN2 (_________36305),
       .Q (_________36306));
  xor2s1 ______499080(.DIN1 (____0____36234), .DIN2 (_________38869),
       .Q (_________36304));
  nor2s1 _______499081(.DIN1 (____0____36233), .DIN2 (______0__36309),
       .Q (_________36303));
  xor2s1 ______499082(.DIN1 (____0____36227), .DIN2 (________27618), .Q
       (_________36327));
  nnd2s1 ______499083(.DIN1 (______0__36309), .DIN2 (____0_9__36208),
       .Q (______0__36428));
  xor2s1 _______499084(.DIN1 (____0_0__36239), .DIN2 (_____9___38412),
       .Q (_________37352));
  or2s1 _______499085(.DIN1
       (_____________________________________________21811), .DIN2
       (____09___40812), .Q (______0__36302));
  nnd2s1 _______499086(.DIN1 (____0____36247), .DIN2 (_________38262),
       .Q (_________36299));
  nnd2s1 _______499087(.DIN1 (_________36297), .DIN2 (___0_0___40568),
       .Q (_________36298));
  and2s1 _______499088(.DIN1 (____09___40812), .DIN2
       (_____________________________________________21811), .Q
       (_________36296));
  nor2s1 _____0_499089(.DIN1 (____0____34397), .DIN2 (____0____36250),
       .Q (_________36294));
  nor2s1 _______499090(.DIN1 (___0_____40485), .DIN2 (___0_____40499),
       .Q (_________36293));
  and2s1 ______499091(.DIN1 (_________36292), .DIN2 (___0_____40499),
       .Q (_________36352));
  and2s1 _______499092(.DIN1 (___0_____40499), .DIN2 (___0_____40485),
       .Q (_________36354));
  nor2s1 _____499093(.DIN1 (_________35845), .DIN2 (____0_0__36249), .Q
       (_________36341));
  nor2s1 ______499094(.DIN1 (____0____36195), .DIN2 (____0____36244),
       .Q (_________36342));
  nor2s1 _______499095(.DIN1 (___0_____40499), .DIN2 (_________36292),
       .Q (_________36351));
  xor2s1 _____499096(.DIN1 (____0____36224), .DIN2 (_____9___35730), .Q
       (_____09__36374));
  nnd2s1 ______499097(.DIN1 (____0____36237), .DIN2 (_________36643),
       .Q (_________36290));
  nor2s1 _______499098(.DIN1 (_________36288), .DIN2 (____0____36241),
       .Q (_________36289));
  xor2s1 _______499099(.DIN1 (______9__35536), .DIN2 (____0____36252),
       .Q (______0__36287));
  xor2s1 _______499100(.DIN1 (____0____36203), .DIN2 (_____0___36285),
       .Q (_____09__36286));
  xor2s1 _______499101(.DIN1
       (_____________________________________________21801), .DIN2
       (_____9___36629), .Q (_____0___36284));
  xor2s1 _____0_499102(.DIN1 (____0_0__36209), .DIN2 (___900___38985),
       .Q (_____0___36283));
  nnd2s1 ______499103(.DIN1 (____0____36242), .DIN2 (inData[6]), .Q
       (_____0___36281));
  or2s1 ______499104(.DIN1 (____9____36167), .DIN2 (_____0___36279), .Q
       (_____0___36280));
  nnd2s1 _______499105(.DIN1 (____0____36232), .DIN2 (_________37414),
       .Q (_____00__36278));
  hi1s1 _______499106(.DIN (______0__36309), .Q (_____9___36363));
  xor2s1 _______499107(.DIN1 (____0____36196), .DIN2 (_________41343),
       .Q (____099__36277));
  nor2s1 _____9_499108(.DIN1 (____0____38117), .DIN2 (____0____36222),
       .Q (____09___36276));
  nor2s1 _______499109(.DIN1 (_________38280), .DIN2 (____0_9__36218),
       .Q (____09___36275));
  nnd2s1 _______499110(.DIN1 (____09___36273), .DIN2 (_________38280),
       .Q (____09___36274));
  xor2s1 ______499111(.DIN1 (____0____34429), .DIN2 (____09___40814),
       .Q (____09___36272));
  xor2s1 _______499112(.DIN1 (____0_9__36248), .DIN2 (_________35844),
       .Q (____09___36271));
  or2s1 _______499113(.DIN1 (____0_0__36229), .DIN2 (____09___36269),
       .Q (____09___36270));
  xor2s1 ______499114(.DIN1 (____0_0__36192), .DIN2 (____0_9__36267),
       .Q (____090__36268));
  nnd2s1 _____0_499115(.DIN1 (____0____36266), .DIN2 (____0____36265),
       .Q (______9__36295));
  nnd2s1 ______499116(.DIN1 (______0__36985), .DIN2 (____0____36236),
       .Q (______9__36328));
  hi1s1 _______499117(.DIN (_________36297), .Q (_________36315));
  xor2s1 _______499118(.DIN1 (____0____36197), .DIN2 (___9_9___39790),
       .Q (_________36331));
  dffacs1 _____________________________________________0_499119(.CLRB
       (reset), .CLK (clk), .DIN (____0_9__36238), .Q
       (_________________________________________0_));
  nnd2s1 _____9_499120(.DIN1 (____0____36254), .DIN2 (____0____36260),
       .Q (____0____36264));
  nor2s1 _______499121(.DIN1 (____0____36210), .DIN2 (____0____36213),
       .Q (____0____36263));
  nnd2s1 _______499122(.DIN1 (____0____36214), .DIN2 (_________33291),
       .Q (____0____36262));
  xor2s1 _______499123(.DIN1 (___09____40677), .DIN2 (____0____36260),
       .Q (____0____36261));
  nor2s1 _______499124(.DIN1 (____0_0__36258), .DIN2 (_____9___36629),
       .Q (____0____36259));
  nor2s1 _______499125(.DIN1 (________27367), .DIN2 (____0____36207),
       .Q (____0_9__36257));
  nor2s1 _______499126(.DIN1 (______0__33292), .DIN2 (____0____36212),
       .Q (____0____36256));
  nor2s1 _____0_499127(.DIN1 (____0____36260), .DIN2 (____0____36254),
       .Q (____0____36255));
  nnd2s1 _______499128(.DIN1 (_____9___36629), .DIN2 (____0_0__36258),
       .Q (____0____36253));
  nor2s1 _____0_499129(.DIN1 (____9____36147), .DIN2 (____0____36206),
       .Q (_________36748));
  or2s1 _______499130(.DIN1 (_________35510), .DIN2 (____0____36252),
       .Q (_________36307));
  xor2s1 _______499131(.DIN1 (____00___36188), .DIN2 (_____0___36285),
       .Q (______9__36613));
  xor2s1 _______499132(.DIN1 (____0____36231), .DIN2 (_________37937),
       .Q (____0____36251));
  nor2s1 _______499133(.DIN1 (____009__34395), .DIN2 (____09___40814),
       .Q (____0____36250));
  nor2s1 _______499134(.DIN1 (_____0___35841), .DIN2 (____0_9__36248),
       .Q (____0_0__36249));
  xor2s1 _______499135(.DIN1 (____00___36183), .DIN2 (___9__9__39731),
       .Q (____0____36247));
  xor2s1 _______499136(.DIN1 (____0____36225), .DIN2 (____0____36245),
       .Q (____0____36246));
  nor2s1 ______499137(.DIN1 (_________36680), .DIN2 (____0_9__36200),
       .Q (____0____36244));
  nnd2s1 _______499138(.DIN1 (____0____36204), .DIN2 (_________34942),
       .Q (_________36305));
  nnd2s1 ______499139(.DIN1 (____0_9__36228), .DIN2 (____0____36243),
       .Q (_________36300));
  xor2s1 _______499140(.DIN1 (____99___36175), .DIN2 (______9__37429),
       .Q (_________36297));
  dffacs1 _______________________________________________499141(.CLRB
       (reset), .CLK (clk), .DIN (____0____36198), .QN
       (___0_____40499));
  xor2s1 _____9_499142(.DIN1 (____99___36180), .DIN2 (__________0_), .Q
       (______0__36309));
  nor2s1 _____499143(.DIN1 (____009__36191), .DIN2 (____9___24640), .Q
       (____0____36242));
  xor2s1 ______499144(.DIN1 (_________34944), .DIN2 (____09___40818),
       .Q (____0____36241));
  nor2s1 _______499145(.DIN1 (_________41090), .DIN2 (____00___36185),
       .Q (____0____36240));
  xor2s1 _______499146(.DIN1 (_____0___40822), .DIN2 (_________36439),
       .Q (____0_0__36239));
  nnd2s1 _____9_499147(.DIN1 (____00___36184), .DIN2 (____9___27734),
       .Q (____0_9__36238));
  nor2s1 ______499148(.DIN1 (_________35954), .DIN2 (____00___36189),
       .Q (____0____36237));
  nnd2s1 _____499149(.DIN1 (_________37937), .DIN2 (____0____36235), .Q
       (____0____36236));
  nor2s1 _____0_499150(.DIN1 (____0____36233), .DIN2 (_________37937),
       .Q (____0____36234));
  xor2s1 _______499151(.DIN1 (____9____36157), .DIN2 (_____9___37851),
       .Q (____0____36232));
  or2s1 _____0_499152(.DIN1 (____0____36231), .DIN2 (_________37937),
       .Q (_________36316));
  and2s1 _____0_499153(.DIN1 (_________37937), .DIN2 (____0____36230),
       .Q (_____0___36282));
  hi1s1 _______499154(.DIN (____0_9__36228), .Q (____0_0__36229));
  xor2s1 _______499155(.DIN1 (____9____36159), .DIN2 (_____9___38512),
       .Q (____0____36227));
  dffacs1 _____________9_(.CLRB (reset), .CLK (clk), .DIN
       (_________37937), .Q (outData[9]));
  nor2s1 _______499156(.DIN1 (________22524), .DIN2 (____0____36225),
       .Q (____0____36226));
  or2s1 _______499157(.DIN1 (____0____36223), .DIN2 (____0____36217),
       .Q (____0____36224));
  xor2s1 _______499158(.DIN1 (_________34987), .DIN2 (____0____36199),
       .Q (____0____36222));
  xor2s1 _______499159(.DIN1 (____0____36220), .DIN2 (____0_0__36219),
       .Q (____0____36221));
  nor2s1 ______499160(.DIN1 (____0____36216), .DIN2 (____0____36217),
       .Q (____0_9__36218));
  nnd2s1 _______499161(.DIN1 (____0____36225), .DIN2
       (_____________________________________________21802), .Q
       (____0____36265));
  nnd2s1 _______499162(.DIN1 (____0____36217), .DIN2 (____0____36216),
       .Q (____09___36273));
  or2s1 ______499163(.DIN1
       (_____________________________________________21802), .DIN2
       (____0____36225), .Q (____0____36266));
  xor2s1 _______499164(.DIN1 (____09___40816), .DIN2 (____0____36215),
       .Q (_____0___36279));
  nnd2s1 _______499165(.DIN1 (____0____36213), .DIN2 (____0____36211),
       .Q (____0____36214));
  nor2s1 _______499166(.DIN1 (____0____36211), .DIN2 (____0____36213),
       .Q (____0____36212));
  xor2s1 _______499167(.DIN1 (____9____36156), .DIN2 (_________38200),
       .Q (____0____36210));
  xor2s1 _______499168(.DIN1 (____9____36151), .DIN2 (____9____36152),
       .Q (____0_0__36209));
  or2s1 _______499169(.DIN1 (____0____36230), .DIN2 (_________36439),
       .Q (____0_9__36208));
  nor2s1 _______499170(.DIN1 (____0____37165), .DIN2 (____9____36161),
       .Q (____0____36207));
  nor2s1 _______499171(.DIN1 (______9__35906), .DIN2 (____9____36166),
       .Q (____0____36206));
  nnd2s1 _____9_499172(.DIN1 (_________36439), .DIN2 (____0____36233),
       .Q (____0____36205));
  nnd2s1 _____9_499173(.DIN1 (_________34943), .DIN2 (____09___40818),
       .Q (____0____36204));
  nnd2s1 _____0_499174(.DIN1 (____9____36168), .DIN2 (____0____36202),
       .Q (____0____36203));
  nor2s1 _______499175(.DIN1 (______9__35440), .DIN2 (____9____36170),
       .Q (____0____36252));
  hi1s1 _______499176(.DIN (___09____40677), .Q (____0____36254));
  nnd2s1 _______499177(.DIN1 (_________36439), .DIN2 (____0_0__36201),
       .Q (______0__36985));
  nor2s1 _______499178(.DIN1 (____0____36194), .DIN2 (____0____36199),
       .Q (____0_9__36200));
  nnd2s1 _______499179(.DIN1 (____9____36163), .DIN2 (____0____37147),
       .Q (____0____36198));
  nor2s1 _______499180(.DIN1 (________28039), .DIN2 (____9____36165),
       .Q (____0____36197));
  xor2s1 _______499181(.DIN1 (____9____36138), .DIN2 (___0_____40652),
       .Q (____0____36196));
  and2s1 ______499182(.DIN1 (____0____36199), .DIN2 (____0____36194),
       .Q (____0____36195));
  nor2s1 _______499183(.DIN1 (___0_____40517), .DIN2 (____990__36172),
       .Q (____0____36193));
  nor2s1 _____0_499184(.DIN1 (_____00__40820), .DIN2 (____9____36160),
       .Q (____0_0__36192));
  nnd2s1 _______499185(.DIN1 (____0_0__36219), .DIN2 (___0_0___40569),
       .Q (____0_9__36228));
  xor2s1 _______499186(.DIN1 (____9____36134), .DIN2 (_____0___36285),
       .Q (____0_9__36248));
  nor2s1 _______499187(.DIN1 (___0_0___40569), .DIN2 (____0_0__36219),
       .Q (____09___36269));
  dffacs1 _______________________________________________499188(.CLRB
       (reset), .CLK (clk), .DIN (____9_0__36162), .QN
       (_____________________________________________21799));
  xnr2s1 _______499189(.DIN1 (_________38280), .DIN2 (____9_9__36139),
       .Q (_____9___36629));
  xor2s1 _______499190(.DIN1
       (_____________________________________________21854), .DIN2
       (_____________________________________0______21757), .Q
       (____009__36191));
  nor2s1 _____499191(.DIN1 (_________41341), .DIN2 (____00___36186), .Q
       (____00___36190));
  nor2s1 _______499192(.DIN1 (_________36288), .DIN2 (____9_9__36148),
       .Q (____00___36189));
  nnd2s1 _______499193(.DIN1 (____9____36153), .DIN2 (____9_0__36149),
       .Q (____00___36188));
  nnd2s1 _____9_499194(.DIN1 (____00___36186), .DIN2 (_________41341),
       .Q (____00___36187));
  xor2s1 _______499195(.DIN1 (_____9___35558), .DIN2 (____9____36169),
       .Q (____00___36185));
  nor2s1 _______499196(.DIN1 (____9___28106), .DIN2 (____9____36145),
       .Q (____00___36184));
  hi1s1 _______499197(.DIN (_________36439), .Q (_________37937));
  xor2s1 _____499198(.DIN1 (____9____36119), .DIN2 (____000__36182), .Q
       (____00___36183));
  xor2s1 _______499199(.DIN1
       (_____________________________________________21854), .DIN2
       (____99___36176), .Q (____999__36181));
  xor2s1 ______499200(.DIN1 (___0__9__40590), .DIN2 (____9____36164),
       .Q (____99___36180));
  nnd2s1 ______499201(.DIN1 (____99___36178), .DIN2 (_________35946),
       .Q (____99___36179));
  nnd2s1 _____9_499202(.DIN1 (____99___36176), .DIN2 (____9____36137),
       .Q (____99___36177));
  xor2s1 _____0_499203(.DIN1 (____9____36116), .DIN2 (____99___36174),
       .Q (____99___36175));
  or2s1 _______499204(.DIN1 (______9__35941), .DIN2 (____99___36178),
       .Q (____99___36173));
  nnd2s1 _______499205(.DIN1 (____9____36136), .DIN2 (____900__36097),
       .Q (____0____36217));
  hi1s1 _____9_499206(.DIN (____990__36172), .Q (____0____36225));
  nnd2s1 _____9_499207(.DIN1 (_________35063), .DIN2
       (_____________________________________________21854), .Q
       (____9_9__36171));
  nor2s1 ______499208(.DIN1 (_________35445), .DIN2 (____9____36169),
       .Q (____9____36170));
  hi1s1 _______499209(.DIN (____9____36167), .Q (____9____36168));
  xor2s1 ______499210(.DIN1 (____9____36113), .DIN2 (_________36854),
       .Q (____9____36166));
  nor2s1 ______499211(.DIN1 (_____9__28461), .DIN2 (____9____36164), .Q
       (____9____36165));
  nor2s1 _______499212(.DIN1 (__9_0___29901), .DIN2 (____9____36126),
       .Q (____9____36163));
  nnd2s1 _______499213(.DIN1 (____9_0__36131), .DIN2 (_____9___41202),
       .Q (____9_0__36162));
  xor2s1 _______499214(.DIN1 (____0_9__35349), .DIN2 (____9____36112),
       .Q (____9____36161));
  xor2s1 _______499215(.DIN1 (____9____36154), .DIN2 (____9____36155),
       .Q (____0____36211));
  xnr2s1 _______499216(.DIN1 (_________9_), .DIN2 (____90___36103), .Q
       (_________36439));
  nor2s1 _______499217(.DIN1 (_________41367), .DIN2 (____9____36123),
       .Q (____9____36160));
  xor2s1 _____0_499218(.DIN1 (____90___36100), .DIN2 (______0__35481),
       .Q (____9____36159));
  xor2s1 _____0_499219(.DIN1 (____90___36099), .DIN2 (_________36292),
       .Q (____9____36157));
  xor2s1 _______499220(.DIN1 (_________35632), .DIN2 (_____9___36096),
       .Q (____990__36172));
  dffacs1 _______________________________________________499221(.CLRB
       (reset), .CLK (clk), .DIN (____9_9__36121), .Q (___0_9___40557));
  nnd2s1 _______499222(.DIN1 (____9____36132), .DIN2 (____9____36117),
       .Q (____0____36199));
  xor2s1 _______499223(.DIN1 (____90___36098), .DIN2 (____0____37113),
       .Q (____0_0__36219));
  dffacs1 ______________________________________499224(.CLRB (reset),
       .CLK (clk), .DIN (____9____36129), .QN (___________));
  nor2s1 _______499225(.DIN1 (____9____36155), .DIN2 (____9____36154),
       .Q (____9____36156));
  nnd2s1 _____9_499226(.DIN1 (____9____36150), .DIN2 (____9____36152),
       .Q (____9____36153));
  and2s1 _____0_499227(.DIN1 (____9____36150), .DIN2 (____9_0__36149),
       .Q (____9____36151));
  xor2s1 _______499228(.DIN1 (_____90__36089), .DIN2 (_________36054),
       .Q (____9_9__36148));
  nor2s1 _______499229(.DIN1 (_________36854), .DIN2 (____9____36111),
       .Q (____9____36147));
  nnd2s1 _______499230(.DIN1 (____9____36109), .DIN2 (_________37744),
       .Q (____9____36146));
  xor2s1 ______499231(.DIN1 (_________36083), .DIN2 (___9_____39582),
       .Q (____9____36167));
  xor2s1 _______499232(.DIN1 (_____9___36090), .DIN2 (_____00__35736),
       .Q (____0____36202));
  nnd2s1 _______499233(.DIN1 (____9____36154), .DIN2 (____9____36155),
       .Q (____00___36186));
  nor2s1 _______499234(.DIN1 (____0_0__37159), .DIN2 (____9____36108),
       .Q (____9____36145));
  or2s1 ______499235(.DIN1 (____9____36143), .DIN2 (____9____36142), .Q
       (____9____36144));
  xor2s1 _____0_499236(.DIN1 (____9_0__36140), .DIN2 (___9____26008),
       .Q (____9____36141));
  xor2s1 _______499237(.DIN1 (_________36073), .DIN2 (____0____38106),
       .Q (____9_9__36139));
  xnr2s1 _______499238(.DIN1 (___0__9__40520), .DIN2 (_____0___40824),
       .Q (____9____36138));
  hi1s1 _______499239(.DIN
       (_____________________________________________21854), .Q
       (____9____36137));
  or2s1 _______499240(.DIN1 (____9____36135), .DIN2 (____9_0__36122),
       .Q (____9____36136));
  nnd2s1 ______499241(.DIN1 (____90___36102), .DIN2 (_________35714),
       .Q (____9____36134));
  nnd2s1 _______499242(.DIN1 (____9____36133), .DIN2 (______0__36081),
       .Q (____99___36178));
  nnd2s1 _______499243(.DIN1 (____9____36118), .DIN2 (_________36382),
       .Q (____9____36132));
  or2s1 _______499244(.DIN1 (____0_0__37159), .DIN2 (_________36075),
       .Q (____9_0__36131));
  xor2s1 _______499245(.DIN1 (_________31912), .DIN2 (____9____36152),
       .Q (____9_9__36130));
  nnd2s1 _______499246(.DIN1 (_________35990), .DIN2 (______9__36088),
       .Q (____9____36129));
  nor2s1 _______499247(.DIN1 (___9_____39274), .DIN2 (____9____36127),
       .Q (____9____36128));
  and2s1 ______499248(.DIN1 (_________36078), .DIN2 (____9____37049),
       .Q (____9____36126));
  xor2s1 _______499249(.DIN1 (____9____36124), .DIN2 (_________38463),
       .Q (____9____36125));
  nor2s1 _____9_499250(.DIN1 (____9____35277), .DIN2 (_________36085),
       .Q (____9____36169));
  nor2s1 _______499251(.DIN1 (_______22231), .DIN2 (_____9___36093), .Q
       (____9____36164));
  hi1s1 _______499252(.DIN (____9_0__36122), .Q (____9____36123));
  nnd2s1 _______499253(.DIN1 (_________36077), .DIN2 (_________38262),
       .Q (____9_9__36121));
  and2s1 _______499254(.DIN1 (____9____36118), .DIN2 (____9____36117),
       .Q (____9____36119));
  xor2s1 ______499255(.DIN1 (____90___36101), .DIN2 (____0____36216),
       .Q (____9____36116));
  nor2s1 _______499256(.DIN1 (____9_9__36114), .DIN2 (_________36076),
       .Q (____9_0__36115));
  nnd2s1 _______499257(.DIN1 (_____9___35828), .DIN2 (_____0___40824),
       .Q (____9____36158));
  dffacs1 _______________________________________________499258(.CLRB
       (reset), .CLK (clk), .DIN (_____9___36091), .QN
       (_____________________________________________21854));
  dffacs1 _____________________________________________9_499259(.CLRB
       (reset), .CLK (clk), .DIN (______9__36072), .QN
       (_________22042));
  and2s1 _____499260(.DIN1 (____9____36152), .DIN2 (____9____36110), .Q
       (____9____36113));
  xor2s1 ______499261(.DIN1 (_________36084), .DIN2 (_____99__36913),
       .Q (____9____36112));
  or2s1 _______499262(.DIN1 (____9____36110), .DIN2 (____9____36152),
       .Q (____9____36111));
  and2s1 _______499263(.DIN1 (_________36069), .DIN2 (____0____36231),
       .Q (____9____36109));
  xor2s1 ______499264(.DIN1 (_________36051), .DIN2 (____9_0__36107),
       .Q (____9____36108));
  xnr2s1 _____0_499265(.DIN1 (___00____39929), .DIN2 (____099__37188),
       .Q (____909__36106));
  hi1s1 _______499266(.DIN (____9____36127), .Q (____9____36133));
  nor2s1 _______499267(.DIN1 (____0___27923), .DIN2 (______9__36427),
       .Q (____9____36142));
  nnd2s1 _______499268(.DIN1 (____90___36105), .DIN2
       (_________________________________________0___21952), .Q
       (____9____36150));
  or2s1 ______499269(.DIN1
       (_________________________________________0___21952), .DIN2
       (____90___36105), .Q (____9_0__36149));
  xor2s1 _______499270(.DIN1 (_________36058), .DIN2 (____90___36104),
       .Q (____9____36154));
  dffacs1 _____________________________________________0_499271(.CLRB
       (reset), .CLK (clk), .DIN (_________36068), .QN
       (_________________________________________0___21798));
  xor2s1 _______499272(.DIN1 (___0__0__40591), .DIN2 (_____9___36092),
       .Q (____90___36103));
  or2s1 _____0_499273(.DIN1 (_________35713), .DIN2 (____90___36101),
       .Q (____90___36102));
  nnd2s1 _____9_499274(.DIN1 (______0__36065), .DIN2 (_________35483),
       .Q (____90___36100));
  xor2s1 _____9_499275(.DIN1 (_________36071), .DIN2 (___0_____40508),
       .Q (____90___36099));
  xor2s1 _______499276(.DIN1 (_________36048), .DIN2 (_________37412),
       .Q (____90___36098));
  nnd2s1 ______499277(.DIN1 (_____9___36095), .DIN2 (________27612), .Q
       (____900__36097));
  nor2s1 _______499278(.DIN1 (_________35591), .DIN2 (_____9___36095),
       .Q (_____9___36096));
  nnd2s1 _____499279(.DIN1 (_____9___36095), .DIN2 (_____9___36094), .Q
       (____9_0__36122));
  nor2s1 _______499280(.DIN1 (_____99__33909), .DIN2 (_________36061),
       .Q (_________36356));
  nor2s1 _______499281(.DIN1 (_____0___34761), .DIN2 (_________36067),
       .Q (_________36432));
  xor2s1 _____9_499282(.DIN1 (_________36049), .DIN2 (___9_0___39619),
       .Q (____0____36243));
  dffacs1 _________________________________________9____(.CLRB (reset),
       .CLK (clk), .DIN (_________36062), .Q
       (_____________________________________9______21877));
  dffacs1 ___________________________________9_(.CLRB (reset), .CLK
       (clk), .DIN (_____0___40826), .QN (___0__0__40591));
  nor2s1 _______499283(.DIN1 (_______22179), .DIN2 (_____9___36092), .Q
       (_____9___36093));
  nnd2s1 _______499284(.DIN1 (_________36052), .DIN2 (____9___24641),
       .Q (_____9___36091));
  nor2s1 ______499285(.DIN1 (_________36082), .DIN2 (____099__37188),
       .Q (_____9___36090));
  xor2s1 _____499286(.DIN1 (_________36045), .DIN2 (_________36034), .Q
       (_____90__36089));
  nnd2s1 _______499287(.DIN1 (______9__36055), .DIN2
       (_____________________________________9_____), .Q
       (______9__36088));
  and2s1 _______499288(.DIN1 (_________36084), .DIN2 (____9____35265),
       .Q (_________36085));
  and2s1 _______499289(.DIN1 (____099__37188), .DIN2 (_________36082),
       .Q (_________36083));
  nnd2s1 _______499290(.DIN1 (______9__36080), .DIN2 (_________36079),
       .Q (______0__36081));
  nor2s1 ______499291(.DIN1
       (_____________________________________________21897), .DIN2
       (______9__36080), .Q (____9____36143));
  nor2s1 _______499292(.DIN1 (___0_____40646), .DIN2 (______9__36080),
       .Q (____9____36127));
  nor2s1 _____9_499293(.DIN1 (_________35985), .DIN2 (_________36057),
       .Q (____0____36260));
  xor2s1 _______499294(.DIN1 (_________36040), .DIN2 (_________38385),
       .Q (_________36078));
  xor2s1 ______499295(.DIN1 (_________36039), .DIN2 (_________40834),
       .Q (_________36077));
  xor2s1 _______499296(.DIN1 (_________36060), .DIN2 (______0__33946),
       .Q (_________36076));
  xor2s1 _______499297(.DIN1 (_________34786), .DIN2 (_________36066),
       .Q (_________36075));
  xor2s1 _____9_499298(.DIN1 (______9__36064), .DIN2 (_________35504),
       .Q (_________36073));
  nnd2s1 _______499299(.DIN1 (_________36050), .DIN2 (_____9___36996),
       .Q (______9__36072));
  or2s1 _______499300(.DIN1 (_________34168), .DIN2 (_________36071),
       .Q (____9____36120));
  nnd2s1 _______499301(.DIN1 (_________36070), .DIN2 (___0_9___40557),
       .Q (____9____36118));
  or2s1 _______499302(.DIN1 (___0_9___40557), .DIN2 (_________36070),
       .Q (____9____36117));
  hi1s1 _______499303(.DIN (____9____36124), .Q (____9_0__36140));
  dffacs1 ____________________________________0_499304(.CLRB (reset),
       .CLK (clk), .DIN (_________36059), .Q (___0__9__40590));
  xor2s1 ______499305(.DIN1 (_________36026), .DIN2 (_________38675),
       .Q (_________36069));
  nnd2s1 ______499306(.DIN1 (______0__36047), .DIN2 (___0____28760), .Q
       (_________36068));
  xor2s1 _____0_499307(.DIN1 (_________36033), .DIN2 (_________38200),
       .Q (____90___36105));
  xor2s1 ______499308(.DIN1 (________22381), .DIN2 (______0__36028), .Q
       (____0____36233));
  xor2s1 _______499309(.DIN1 (_________36024), .DIN2 (_____0___36015),
       .Q (____9____36152));
  dffacs1 __________________499310(.CLRB (reset), .CLK (clk), .DIN
       (_________36044), .QN
       (_________________________________________________________________________________________22095));
  nor2s1 _____499311(.DIN1 (_____0___34760), .DIN2 (_________36066), .Q
       (_________36067));
  nnd2s1 _______499312(.DIN1 (______9__36064), .DIN2 (_________35484),
       .Q (______0__36065));
  nnd2s1 _____0_499313(.DIN1 (_____9___35466), .DIN2 (_________36043),
       .Q (_________36062));
  nor2s1 _____0_499314(.DIN1 (_____00__33910), .DIN2 (_________36060),
       .Q (_________36061));
  nor2s1 ______499315(.DIN1 (_____9___35647), .DIN2 (______9__36037),
       .Q (____90___36101));
  xor2s1 _____9_499316(.DIN1 (_________36019), .DIN2 (_____9___35196),
       .Q (____9____36124));
  hi1s1 _______499317(.DIN (______9__36080), .Q (______9__36427));
  nor2s1 _______499318(.DIN1 (_________35592), .DIN2 (______9__36064),
       .Q (_____9___36095));
  or2s1 _______499319(.DIN1 (_________36032), .DIN2 (_________35705),
       .Q (_________36059));
  xor2s1 _____0_499320(.DIN1 (_____9___36008), .DIN2 (______0__36056),
       .Q (_________36058));
  nor2s1 ______499321(.DIN1 (______0__36056), .DIN2 (_________36029),
       .Q (_________36057));
  or2s1 _______499322(.DIN1 (_________36031), .DIN2 (_____9___36005),
       .Q (______9__36055));
  xor2s1 _____9_499323(.DIN1 (_____99__36009), .DIN2 (______9__34088),
       .Q (_________36084));
  nnd2s1 ______499324(.DIN1 (_________36054), .DIN2 (_________36035),
       .Q (_________36086));
  xor2s1 _____9_499325(.DIN1 (_________36053), .DIN2 (____9____37036),
       .Q (______9__36080));
  xnr2s1 _____9_499326(.DIN1 (_________36053), .DIN2 (_____0___40828),
       .Q (____099__37188));
  dffacs1 _________________________________________9_____499327(.CLRB
       (reset), .CLK (clk), .DIN (_________36021), .Q
       (_____________________________________9_____));
  nnd2s1 _____499328(.DIN1 (_____09__36017), .DIN2 (_________35680), .Q
       (_________36052));
  xor2s1 _______499329(.DIN1 (_________35995), .DIN2 (_________34791),
       .Q (_________36051));
  nor2s1 _______499330(.DIN1 (________27466), .DIN2 (_____0___36011),
       .Q (_________36050));
  nnd2s1 _______499331(.DIN1 (_____0___36012), .DIN2 (______0__35975),
       .Q (_________36049));
  xor2s1 _______499332(.DIN1 (____9____36135), .DIN2 (_________36036),
       .Q (_________36048));
  nor2s1 _______499333(.DIN1 (_____9___36004), .DIN2 (______0__36018),
       .Q (_____9___36092));
  and2s1 _______499334(.DIN1 (_____0___36013), .DIN2 (_________35978),
       .Q (_________36070));
  xor2s1 _______499335(.DIN1 (______0__35993), .DIN2 (___9_____39738),
       .Q (_________36071));
  nor2s1 _______499336(.DIN1 (_____0___36016), .DIN2 (_________36023),
       .Q (_________36074));
  or2s1 ______499337(.DIN1 (_________36521), .DIN2 (_____90__36000), .Q
       (______0__36047));
  nnd2s1 _______499338(.DIN1 (_________36053), .DIN2 (_________36020),
       .Q (_________36046));
  xor2s1 _______499339(.DIN1 (___0_____40488), .DIN2
       (___________________), .Q (_________36045));
  nnd2s1 _______499340(.DIN1 (_________36643), .DIN2 (_________35994),
       .Q (_________36044));
  nnd2s1 _______499341(.DIN1 (_____9___36001), .DIN2 (inData[2]), .Q
       (_________36043));
  nor2s1 _______499342(.DIN1 (______9__36027), .DIN2 (_________36053),
       .Q (_________36063));
  nnd2s1 _______499343(.DIN1 (_________36053), .DIN2 (_________35934),
       .Q (____0____36231));
  xor2s1 _______499344(.DIN1 (________26216), .DIN2 (_________36041),
       .Q (_________36042));
  xor2s1 _______499345(.DIN1 (_________35976), .DIN2 (______9__33945),
       .Q (_________36040));
  xor2s1 ______499346(.DIN1 (___0_09__40570), .DIN2 (_________36041),
       .Q (_________36039));
  nnd2s1 _____9_499347(.DIN1 (______9__35999), .DIN2 (______9__37314),
       .Q (______0__36038));
  nor2s1 ______499348(.DIN1 (______0__35636), .DIN2 (_________36036),
       .Q (______9__36037));
  xnr2s1 _______499349(.DIN1 (_____9___36721), .DIN2 (______0__40830),
       .Q (_________36066));
  nor2s1 _______499350(.DIN1 (_____9___33808), .DIN2 (_________35998),
       .Q (_________36060));
  nor2s1 _______499351(.DIN1 (_____9___35195), .DIN2 (_________35997),
       .Q (______9__36064));
  or2s1 _______499352(.DIN1 (___0_____40488), .DIN2 (_________36034),
       .Q (_________36035));
  nor2s1 _______499353(.DIN1 (_________32951), .DIN2 (_________35984),
       .Q (_________36033));
  nnd2s1 _____0_499354(.DIN1 (_________35989), .DIN2 (_____0__25538),
       .Q (_________36032));
  nor2s1 _____0_499355(.DIN1 (___0__9__40590), .DIN2 (_________35988),
       .Q (_________36031));
  and2s1 _______499356(.DIN1 (_________36034), .DIN2 (___0_____40488),
       .Q (_________36030));
  nor2s1 _______499357(.DIN1 (_____9___36007), .DIN2 (_________35987),
       .Q (_________36029));
  nnd2s1 _______499358(.DIN1 (_________36025), .DIN2 (______9__36027),
       .Q (______0__36028));
  nnd2s1 ______499359(.DIN1 (_________36025), .DIN2 (______0__35933),
       .Q (_________36026));
  xor2s1 ______499360(.DIN1 (_________36023), .DIN2 (_________36022),
       .Q (_________36024));
  nnd2s1 ______499361(.DIN1 (_________35981), .DIN2 (________28348), .Q
       (_________36021));
  nor2s1 _______499362(.DIN1 (_________36020), .DIN2 (_________36025),
       .Q (____0____36230));
  xor2s1 ______499363(.DIN1 (________27618), .DIN2 (_________35996), .Q
       (_________36019));
  and2s1 _______499364(.DIN1 (______0__35983), .DIN2 (_________38306),
       .Q (______0__36018));
  xor2s1 _______499365(.DIN1 (_________33835), .DIN2 (_________40832),
       .Q (_____09__36017));
  and2s1 _______499366(.DIN1 (____0____37118), .DIN2 (_____0___36015),
       .Q (_____0___36016));
  or2s1 _______499367(.DIN1 (_____0___36015), .DIN2 (____0____37118),
       .Q (_____0___36014));
  dffacs1 _______________(.CLRB (reset), .CLK (clk), .DIN
       (_________36025), .Q (outData[8]));
  nnd2s1 ______499368(.DIN1 (______0__40840), .DIN2 (_________35979),
       .Q (_____0___36013));
  nnd2s1 _______499369(.DIN1 (_________36041), .DIN2 (_________35980),
       .Q (_____0___36012));
  nor2s1 _______499370(.DIN1 (____0____37165), .DIN2 (______9__35982),
       .Q (_____0___36011));
  nnd2s1 _______499371(.DIN1 (_________35895), .DIN2 (_________35969),
       .Q (_____99__36009));
  xor2s1 _______499372(.DIN1 (_________35986), .DIN2 (_____9___36007),
       .Q (_____9___36008));
  nor2s1 _______499373(.DIN1 (_________35972), .DIN2 (_____9___36005),
       .Q (_____9___36006));
  nor2s1 ______499374(.DIN1 (_________38306), .DIN2 (_________35971),
       .Q (_____9___36004));
  xnr2s1 ____90_499375(.DIN1 (___9_____39384), .DIN2 (_____9___36002),
       .Q (_____9___36003));
  nnd2s1 _______499376(.DIN1 (_________35944), .DIN2 (______0__35965),
       .Q (_____9___36001));
  xor2s1 _______499377(.DIN1 (_________35952), .DIN2 (_________38301),
       .Q (_____90__36000));
  hi1s1 _______499378(.DIN (_________36025), .Q (_________36053));
  xor2s1 _______499379(.DIN1 (_________35704), .DIN2 (_________35973),
       .Q (______9__35999));
  nor2s1 _______499380(.DIN1 (_________33780), .DIN2 (_________40832),
       .Q (_________35998));
  nor2s1 _______499381(.DIN1 (_____9___35192), .DIN2 (_________35996),
       .Q (_________35997));
  xor2s1 _____9_499382(.DIN1 (______0__40840), .DIN2 (______0___22058),
       .Q (_________35995));
  nor2s1 _______499383(.DIN1 (_________35967), .DIN2 (__9_____30421),
       .Q (_________35994));
  nor2s1 _____0_499384(.DIN1 (_____9___33908), .DIN2 (_________35963),
       .Q (______0__35993));
  nor2s1 _______499385(.DIN1 (_________35678), .DIN2 (______9__35964),
       .Q (_________36036));
  xor2s1 _____9_499386(.DIN1 (______9__35956), .DIN2 (_________38306),
       .Q (_____9___36448));
  nor2s1 ____9__499387(.DIN1 (_________37789), .DIN2 (_____9___36002),
       .Q (______9__35992));
  and2s1 ____9__499388(.DIN1 (_____9___36002), .DIN2 (_________37789),
       .Q (_________35991));
  or2s1 _______499389(.DIN1
       (_____________________________________9___0_), .DIN2
       (________26824), .Q (_________35990));
  nnd2s1 _______499390(.DIN1 (_____9___36005), .DIN2
       (_____________________________________9___0_), .Q
       (_________35989));
  nnd2s1 _______499391(.DIN1 (___0_9__25144), .DIN2
       (_____________________________________9___0_), .Q
       (_________35988));
  nor2s1 _____0_499392(.DIN1 (_________36928), .DIN2 (_________35986),
       .Q (_________35987));
  and2s1 _____0_499393(.DIN1 (_________35986), .DIN2 (_________32307),
       .Q (_________35985));
  nnd2s1 _______499394(.DIN1 (_________35986), .DIN2 (______0__32950),
       .Q (_________35984));
  dffacs1 _______________________________________________499395(.CLRB
       (reset), .CLK (clk), .DIN (_________35959), .QN
       (___0_____40488));
  dffacs1 _______________________________________________499396(.CLRB
       (reset), .CLK (clk), .DIN (_________35960), .QN
       (_____________________________________________21853));
  dffacs1 _______________________________________________499397(.CLRB
       (reset), .CLK (clk), .DIN (_________35958), .QN
       (_____________________________________________21810));
  xor2s1 _______499398(.DIN1 (_____99__35922), .DIN2 (_________35970),
       .Q (_________36025));
  dffacs1 _______________________________________________499399(.CLRB
       (reset), .CLK (clk), .DIN (_________35951), .Q (___0__9__40500));
  nnd2s1 _______499400(.DIN1 (_________35962), .DIN2 (_____9___35921),
       .Q (______0__35983));
  xor2s1 ______499401(.DIN1 (_________35949), .DIN2 (______0__35585),
       .Q (______9__35982));
  nnd2s1 _______499402(.DIN1 (_________35953), .DIN2 (_____9___36005),
       .Q (_________35981));
  or2s1 _______499403(.DIN1 (______9__35974), .DIN2 (_________40834),
       .Q (_________35980));
  nnd2s1 _______499404(.DIN1 (_________35977), .DIN2 (______0___22058),
       .Q (_________35979));
  or2s1 _______499405(.DIN1 (______0___22058), .DIN2 (_________35977),
       .Q (_________35978));
  xor2s1 ______499406(.DIN1 (_________40836), .DIN2 (___0_____40509),
       .Q (_________35976));
  nnd2s1 _______499407(.DIN1 (_________40834), .DIN2 (______9__35974),
       .Q (______0__35975));
  or2s1 ______499408(.DIN1 (_________35973), .DIN2 (_________35669), .Q
       (_____00__36010));
  xor2s1 ______499409(.DIN1 (______9__35947), .DIN2 (_________38573),
       .Q (_________36494));
  hi1s1 _______499410(.DIN (_________36022), .Q (____0____37118));
  xor2s1 _______499411(.DIN1 (_________35950), .DIN2 (_____9___36094),
       .Q (_________36041));
  xor2s1 _______499412(.DIN1 (_________35788), .DIN2 (_____0___35926),
       .Q (_________35972));
  nnd2s1 _______499413(.DIN1 (_________35961), .DIN2 (_________35970),
       .Q (_________35971));
  nnd2s1 _______499414(.DIN1 (______0__35948), .DIN2 (_________35968),
       .Q (_________35969));
  nor2s1 _____9_499415(.DIN1 (_________35945), .DIN2 (_________35966),
       .Q (_________35967));
  xor2s1 _____9_499416(.DIN1 (_____0___35927), .DIN2 (_________38675),
       .Q (_________36022));
  dffacs1 _____________________________________________9_499417(.CLRB
       (reset), .CLK (clk), .DIN (_________35940), .QN
       (___0_____40539));
  nnd2s1 _____9_499418(.DIN1 (_________35718), .DIN2 (_________40838),
       .Q (______0__35965));
  xor2s1 _______499419(.DIN1 (_________35938), .DIN2 (_________38871),
       .Q (______9__35964));
  and2s1 _______499420(.DIN1 (_________40836), .DIN2 (______0__33918),
       .Q (_________35963));
  xnr2s1 _______499421(.DIN1 (____0_9__36267), .DIN2 (_____90__35915),
       .Q (_________35996));
  or2s1 _____499422(.DIN1 (_____0___35928), .DIN2 (_________35961), .Q
       (_________35962));
  nnd2s1 _____9_499423(.DIN1 (_____0___35925), .DIN2 (________25701),
       .Q (_________35960));
  nnd2s1 _______499424(.DIN1 (_____0___35929), .DIN2 (_________35435),
       .Q (_________35959));
  nnd2s1 _______499425(.DIN1 (_____0___35930), .DIN2 (___0_____30949),
       .Q (_________35958));
  nor2s1 ____9__499426(.DIN1 (_________35511), .DIN2 (_________35936),
       .Q (_________35973));
  dffacs1 _________________________________________9___0_499427(.CLRB
       (reset), .CLK (clk), .DIN (_____09__35932), .QN
       (_____________________________________9___0_));
  xor2s1 _______499428(.DIN1 (_________35901), .DIN2 (________22537),
       .Q (_________35986));
  xor2s1 ____9__499429(.DIN1 (_________35902), .DIN2 (______0__35957),
       .Q (_____9___36002));
  nnd2s1 _______499430(.DIN1 (_____9___35920), .DIN2 (_________35909),
       .Q (______9__35956));
  nnd2s1 _______499431(.DIN1 (_____00__35923), .DIN2 (_________36670),
       .Q (_________35955));
  nor2s1 ______499432(.DIN1 (_____0___35924), .DIN2 (_________35966),
       .Q (_________35954));
  xor2s1 _______499433(.DIN1 (_________35910), .DIN2 (_____9___35919),
       .Q (_________35953));
  xor2s1 _______499434(.DIN1 (_________35908), .DIN2
       (_________________________________________0_), .Q
       (_________35952));
  nnd2s1 ______499435(.DIN1 (_____9___35916), .DIN2 (____0____37173),
       .Q (_________35951));
  dffacs1 _____________________________________________0_499436(.CLRB
       (reset), .CLK (clk), .DIN (_________35939), .Q
       (______0___22058));
  dffacs1 _______________________________________________499437(.CLRB
       (reset), .CLK (clk), .DIN (_____0___35931), .QN
       (___0_____40524));
  xor2s1 ____499438(.DIN1 (_________35937), .DIN2
       (_______________22074), .Q (_________35950));
  xnr2s1 ____9__499439(.DIN1 (___9_0___39166), .DIN2 (_________35935),
       .Q (_________35949));
  nnd2s1 _____0_499440(.DIN1 (_________35898), .DIN2 (______0__35863),
       .Q (______0__35948));
  xor2s1 _______499441(.DIN1 (_____________22102), .DIN2
       (____________22078), .Q (_________35970));
  nor2s1 _______499442(.DIN1 (_____9___32667), .DIN2 (_________35903),
       .Q (_________36023));
  dffacs1 _______________________________________________499443(.CLRB
       (reset), .CLK (clk), .DIN (_________35914), .Q (___0_____40508));
  dffacs1 ____________________________________________9_(.CLRB (reset),
       .CLK (clk), .DIN (______0__35897), .Q (___0__9__40490));
  dffacs1 _________________(.CLRB (reset), .CLK (clk), .DIN
       (_________35899), .QN (___0_____40598));
  nnd2s1 _______499444(.DIN1 (_________35946), .DIN2 (______0__35889),
       .Q (______9__35947));
  nor2s1 _______499445(.DIN1 (_________35587), .DIN2 (_________35913),
       .Q (_________35945));
  nnd2s1 ______499446(.DIN1 (_________35857), .DIN2 (_________35943),
       .Q (_________35944));
  and2s1 _______499447(.DIN1 (_________35946), .DIN2 (_____9___36721),
       .Q (______9__35941));
  nnd2s1 _______499448(.DIN1 (_________35893), .DIN2 (______9__35683),
       .Q (_________35940));
  nnd2s1 _____499449(.DIN1 (_________35886), .DIN2 (_________38262), .Q
       (_________35939));
  and2s1 ____9__499450(.DIN1 (_________35937), .DIN2 (_________35605),
       .Q (_________35938));
  nor2s1 ____9__499451(.DIN1 (_________35521), .DIN2 (_________35935),
       .Q (_________35936));
  hi1s1 _______499452(.DIN (______0__35933), .Q (_________35934));
  nnd2s1 _____499453(.DIN1 (______0__35880), .DIN2 (____90__26857), .Q
       (_____09__35932));
  nnd2s1 _____0_499454(.DIN1 (_________35881), .DIN2 (____0____37147),
       .Q (_____0___35931));
  nnd2s1 _______499455(.DIN1 (______9__35879), .DIN2 (_________36870),
       .Q (_____0___35930));
  xor2s1 _______499456(.DIN1 (_________35877), .DIN2 (_________38155),
       .Q (_____0___35929));
  and2s1 _______499457(.DIN1 (____________22078), .DIN2
       (_____________22102), .Q (_____0___35928));
  dffacs1 _____________________________________________9_499458(.CLRB
       (reset), .CLK (clk), .DIN (_________35884), .QN
       (______0___22057));
  xor2s1 _______499459(.DIN1 (_____00__35833), .DIN2 (____0_0__36201),
       .Q (_____0___35927));
  and2s1 _______499460(.DIN1 (____________22078), .DIN2
       (___0__0__40591), .Q (_____0___35926));
  nnd2s1 _______499461(.DIN1 (_________35890), .DIN2 (_________35663),
       .Q (_____0___35925));
  xor2s1 _______499462(.DIN1 (_________35912), .DIN2
       (_________________________________________________________________________________________22095),
       .Q (_____0___35924));
  xor2s1 _______499463(.DIN1 (_________35905), .DIN2 (____0_0__36201),
       .Q (_____00__35923));
  xor2s1 _______499464(.DIN1 (_________35961), .DIN2 (________29290),
       .Q (_____99__35922));
  or2s1 _______499465(.DIN1 (_____________22102), .DIN2
       (____________22078), .Q (_____9___35921));
  or2s1 _______499466(.DIN1 (_________35892), .DIN2 (_____9___35919),
       .Q (_____9___35920));
  nor2s1 _______499467(.DIN1 (__9_____30191), .DIN2 (_________35885),
       .Q (_____9___35916));
  nnd2s1 _______499468(.DIN1 (_________35883), .DIN2 (_____9___35829),
       .Q (_____90__35915));
  nnd2s1 ____9__499469(.DIN1 (_________35866), .DIN2 (_________37322),
       .Q (_________35914));
  or2s1 _____9_499470(.DIN1 (_________35872), .DIN2 (_________35912),
       .Q (_________35913));
  nor2s1 _____9_499471(.DIN1 (____0_0__36201), .DIN2 (_________35779),
       .Q (_________35911));
  and2s1 ______499472(.DIN1 (_________35891), .DIN2 (_________35909),
       .Q (_________35910));
  xor2s1 ____90_499473(.DIN1 (_________35882), .DIN2 (_________35907),
       .Q (_________35908));
  nnd2s1 ____90_499474(.DIN1 (______0__35813), .DIN2 (____0_0__36201),
       .Q (______0__35942));
  nnd2s1 ____90_499475(.DIN1 (_________35905), .DIN2 (____0_0__36201),
       .Q (______0__35933));
  nnd2s1 ____90_499476(.DIN1 (____0_0__36201), .DIN2 (______9__35812),
       .Q (______9__36027));
  nor2s1 ____90_499477(.DIN1 (____0_0__36201), .DIN2 (_________35780),
       .Q (_________36020));
  hi1s1 ______499478(.DIN (_________35904), .Q (_________35946));
  nor2s1 _______499479(.DIN1 (_________36781), .DIN2 (_________32664),
       .Q (_________35903));
  nnd2s1 ____0__499480(.DIN1 (______9__35870), .DIN2 (_____9___35825),
       .Q (_________35902));
  xor2s1 ______499481(.DIN1 (_____90__32666), .DIN2 (_________35900),
       .Q (_________35901));
  nnd2s1 _______499482(.DIN1 (_____0___35839), .DIN2 (_________35874),
       .Q (_________35899));
  or2s1 ______499483(.DIN1 (_____00__35653), .DIN2 (_________35864), .Q
       (_________35898));
  nnd2s1 _______499484(.DIN1 (_________35869), .DIN2 (_________35795),
       .Q (______0__35897));
  nnd2s1 ____9__499485(.DIN1 (_________35865), .DIN2 (_________37317),
       .Q (______9__35896));
  or2s1 _______499486(.DIN1 (_________35968), .DIN2 (_________35876),
       .Q (_________35895));
  nor2s1 ______499487(.DIN1 (____00__26499), .DIN2 (_________35873), .Q
       (_________35893));
  hi1s1 _______499488(.DIN (____________22078), .Q (_________35943));
  hi1s1 ____9__499489(.DIN (_________35891), .Q (_________35892));
  xor2s1 _____9_499490(.DIN1 (_________33782), .DIN2 (______0__35871),
       .Q (_________35890));
  nnd2s1 _____9_499491(.DIN1 (____0____36235), .DIN2 (______9__35888),
       .Q (______0__35889));
  nnd2s1 ____90_499492(.DIN1 (_________35855), .DIN2 (_________35768),
       .Q (_________35887));
  xor2s1 ____9__499493(.DIN1 (_____9___35824), .DIN2 (_________35804),
       .Q (_________35886));
  and2s1 ____9__499494(.DIN1 (_________35849), .DIN2 (____9_0__37080),
       .Q (_________35885));
  nnd2s1 ____9__499495(.DIN1 (_________35846), .DIN2 (_____0___37283),
       .Q (_________35884));
  xnr2s1 ____9__499496(.DIN1 (______9__36337), .DIN2 (_____9___35827),
       .Q (_________35883));
  nor2s1 ____9_499497(.DIN1 (______9__35888), .DIN2 (____0____36235),
       .Q (_________35904));
  nor2s1 ____499498(.DIN1 (_________35854), .DIN2 (_____9___36540), .Q
       (______9__35906));
  nor2s1 ____9__499499(.DIN1 (_____9___34563), .DIN2 (_________35882),
       .Q (_____9___35918));
  dffacs1 _____________________________________(.CLRB (reset), .CLK
       (clk), .DIN (_________35858), .Q (____________22078));
  and2s1 _______499500(.DIN1 (_________35861), .DIN2 (__9_____30114),
       .Q (_________35881));
  nor2s1 _______499501(.DIN1 (________26855), .DIN2 (______9__35862),
       .Q (______0__35880));
  xor2s1 ______499502(.DIN1 (____9____35246), .DIN2 (_________35875),
       .Q (______9__35879));
  dffacs1 _______________499503(.CLRB (reset), .CLK (clk), .DIN
       (____0____36235), .Q (outData[7]));
  nor2s1 ____00_499504(.DIN1 (______0__35441), .DIN2 (______0__35843),
       .Q (_________35935));
  xor2s1 ____9__499505(.DIN1 (_________35820), .DIN2 (___9_____39461),
       .Q (_________35937));
  xor2s1 ____9__499506(.DIN1 (_____9___35830), .DIN2 (_________37867),
       .Q (_________36653));
  dffacs1 _______________________________________________499507(.CLRB
       (reset), .CLK (clk), .DIN (_________35851), .Q
       (_____________________________________________21837));
  dffacs1 _____________________________________499508(.CLRB (reset),
       .CLK (clk), .DIN (_________35856), .QN (___0_____40592));
  dffacs1 _________________499509(.CLRB (reset), .CLK (clk), .DIN
       (_________35850), .QN (____________));
  xor2s1 ____90_499510(.DIN1 (_________35810), .DIN2 (____00___35294),
       .Q (_________35877));
  or2s1 _____9_499511(.DIN1 (_________35875), .DIN2 (____9____35245),
       .Q (_________35876));
  nnd2s1 _____9_499512(.DIN1 (_____0___35838), .DIN2 (_____0___35834),
       .Q (_________35874));
  nor2s1 ____9__499513(.DIN1 (____99__26498), .DIN2 (_____99__35832),
       .Q (_________35873));
  nor2s1 ____9__499514(.DIN1 (___0_____40474), .DIN2
       (_________________________________________________________________________________________22094),
       .Q (_________35872));
  and2s1 ____9__499515(.DIN1
       (_________________________________________________________________________________________22094),
       .DIN2 (___0_____40474), .Q (_________35912));
  nnd2s1 ____9__499516(.DIN1 (___0__9__40412), .DIN2 (___0_____40474),
       .Q (_________35891));
  or2s1 ____9__499517(.DIN1 (___0_____40474), .DIN2 (___0__9__40412),
       .Q (_________35909));
  nor2s1 ____9__499518(.DIN1 (_________33671), .DIN2 (______0__35871),
       .Q (_________35894));
  hi1s1 _____499519(.DIN (_________35900), .Q (_________36781));
  hi1s1 ____9__499520(.DIN (____0____36235), .Q (____0_0__36201));
  nnd2s1 ____0__499521(.DIN1 (_________35818), .DIN2 (___9_____39539),
       .Q (______9__35870));
  and2s1 _______499522(.DIN1 (______0__35113), .DIN2 (_____0___35835),
       .Q (_________35869));
  and2s1 ____99_499523(.DIN1 (_________35819), .DIN2 (__9_____29757),
       .Q (_________35866));
  xor2s1 ____0__499524(.DIN1 (_________35447), .DIN2 (_____09__35842),
       .Q (_________35865));
  nor2s1 _______499525(.DIN1 (___0_____40542), .DIN2 (_________35875),
       .Q (_________35864));
  nnd2s1 _______499526(.DIN1 (_________35875), .DIN2 (___0_____40542),
       .Q (______0__35863));
  nor2s1 ____9__499527(.DIN1 (______0__35853), .DIN2 (_____0___35840),
       .Q (_________35905));
  xor2s1 ____9__499528(.DIN1 (______9__35802), .DIN2 (_____99__37662),
       .Q (_________35961));
  dffacs1 _______________________________________________499529(.CLRB
       (reset), .CLK (clk), .DIN (_____9___35831), .QN (______0_));
  dffacs1 _______________________________________________499530(.CLRB
       (reset), .CLK (clk), .DIN (_____0___35836), .QN
       (___0__9__40540));
  and2s1 _____9_499531(.DIN1 (_________35814), .DIN2 (_____9___36005),
       .Q (______9__35862));
  nnd2s1 _____9_499532(.DIN1 (_________35815), .DIN2 (____9____37049),
       .Q (_________35861));
  or2s1 ____9__499533(.DIN1 (_________35859), .DIN2 (___0_____40646),
       .Q (_________35860));
  or2s1 ____9__499534(.DIN1 (_________35857), .DIN2 (________28508), .Q
       (_________35858));
  or2s1 ____9__499535(.DIN1 (______0__35784), .DIN2 (_________35811),
       .Q (_________35856));
  nnd2s1 ____9_499536(.DIN1 (___0_____40646), .DIN2
       (_____________________________________________21896), .Q
       (_________35855));
  and2s1 ____9__499537(.DIN1 (_________36079), .DIN2 (______0__35853),
       .Q (_________35854));
  nor2s1 ____9_499538(.DIN1 (______0__35853), .DIN2 (_________36079),
       .Q (_____9___36540));
  xor2s1 ____9__499539(.DIN1 (_________35787), .DIN2 (___99_0__39864),
       .Q (_________35900));
  xnr2s1 ____9__499540(.DIN1 (_____________22101), .DIN2
       (_________35775), .Q (____0____36235));
  nnd2s1 ____9__499541(.DIN1 (_________35799), .DIN2 (___0__9__40520),
       .Q (______9__35852));
  or2s1 ____9_499542(.DIN1 (___0_____31063), .DIN2 (_________35805), .Q
       (_________35851));
  nnd2s1 _______499543(.DIN1 (________25005), .DIN2 (_________35816),
       .Q (_________35850));
  xor2s1 ____9__499544(.DIN1 (_____09__33917), .DIN2 (_________35817),
       .Q (_________35849));
  xor2s1 ____9__499545(.DIN1 (_________35847), .DIN2 (___9____27757),
       .Q (_________35848));
  nor2s1 ____9__499546(.DIN1 (_____00__41210), .DIN2 (_________35807),
       .Q (_________35846));
  and2s1 ____0__499547(.DIN1 (_________36340), .DIN2 (_________35844),
       .Q (_________35845));
  nor2s1 ____0__499548(.DIN1 (_____09__35842), .DIN2 (_________35442),
       .Q (______0__35843));
  nor2s1 ____0_499549(.DIN1 (_________35844), .DIN2 (_________36340),
       .Q (_____0___35841));
  nor2s1 ____0__499550(.DIN1 (_________35798), .DIN2 (______0__35803),
       .Q (_________35878));
  nor2s1 ____9__499551(.DIN1 (____090__34470), .DIN2 (_________35809),
       .Q (_________35882));
  nnd2s1 ____9__499552(.DIN1 (_________35777), .DIN2 (___0_____30717),
       .Q (_____0___35840));
  nor2s1 ____9_499553(.DIN1 (________25472), .DIN2 (_________35796), .Q
       (_____0___35839));
  nnd2s1 ____9__499554(.DIN1 (_________35794), .DIN2 (inData[0]), .Q
       (_____0___35838));
  nnd2s1 ____99_499555(.DIN1 (_________35847), .DIN2
       (_____________________________________________21799), .Q
       (_____0___35837));
  nnd2s1 ____9__499556(.DIN1 (_________35786), .DIN2 (____0___27303),
       .Q (_____0___35836));
  nnd2s1 ____9__499557(.DIN1 (______9__35792), .DIN2 (_____0___35834),
       .Q (_____0___35835));
  nnd2s1 ____9_499558(.DIN1 (_________35770), .DIN2 (______0__35765),
       .Q (_____00__35833));
  xor2s1 ____9_499559(.DIN1 (____09___34471), .DIN2 (_________35808),
       .Q (_____99__35832));
  or2s1 ____9__499560(.DIN1 (_____9___35559), .DIN2 (______0__35793),
       .Q (_____9___35831));
  nor2s1 ____9__499561(.DIN1 (_________33577), .DIN2 (_________35782),
       .Q (______0__35871));
  nor2s1 ____9_499562(.DIN1 (______9__35619), .DIN2 (_________35790),
       .Q (_________35875));
  dffacs1 _______________________________________________499563(.CLRB
       (reset), .CLK (clk), .DIN (______9__35783), .QN
       (___0_____40474));
  nnd2s1 ____0__499564(.DIN1 (_____9___35826), .DIN2 (_____9___35829),
       .Q (_____9___35830));
  nnd2s1 ____499565(.DIN1 (_________35847), .DIN2 (____0___28017), .Q
       (_____9___35828));
  nnd2s1 ____00_499566(.DIN1 (_____9___35826), .DIN2 (_________37867),
       .Q (_____9___35827));
  nnd2s1 _______499567(.DIN1 (______0__35774), .DIN2 (___9__9__39569),
       .Q (_____9___35825));
  xor2s1 ____0_499568(.DIN1 (______9__35822), .DIN2 (_____9__27442), .Q
       (_____9___35824));
  xor2s1 ____0_499569(.DIN1 (______9__35822), .DIN2 (_____9__26158), .Q
       (_____90__35823));
  nor2s1 ____99_499570(.DIN1
       (_____________________________________________21799), .DIN2
       (___0_____40652), .Q (_________35821));
  nnd2s1 ____0__499571(.DIN1 (_________35771), .DIN2 (_____0___35474),
       .Q (_________35820));
  nnd2s1 ____0__499572(.DIN1 (_________35778), .DIN2 (_________37223),
       .Q (_________35819));
  nnd2s1 ____499573(.DIN1 (_________35769), .DIN2 (________28232), .Q
       (_________35818));
  dffacs1 _________________________________________9____499574(.CLRB
       (reset), .CLK (clk), .DIN (_________35785), .Q (_________22033));
  or2s1 ____00_499575(.DIN1 (_________33796), .DIN2 (_________35817),
       .Q (_________35868));
  nnd2s1 ____9_499576(.DIN1 (_____0___35834), .DIN2 (_________35762),
       .Q (_________35816));
  xor2s1 ____9_499577(.DIN1 (______0__35620), .DIN2 (_________35789),
       .Q (_________35815));
  xor2s1 ____9__499578(.DIN1 (_________35752), .DIN2 (_________35747),
       .Q (_________35814));
  hi1s1 ____0__499579(.DIN (______9__35812), .Q (______0__35813));
  xor2s1 ____9__499580(.DIN1 (___0_____40627), .DIN2 (_____0___35742),
       .Q (_________35811));
  xor2s1 ____9__499581(.DIN1 (_________35781), .DIN2 (_____9___22050),
       .Q (_________35810));
  nor2s1 ____99_499582(.DIN1 (____0_9__34469), .DIN2 (_________35808),
       .Q (_________35809));
  or2s1 ____99_499583(.DIN1 (_____0__28062), .DIN2 (_________35759), .Q
       (_________35807));
  nor2s1 ____9__499584(.DIN1 (_________35766), .DIN2 (_____0___35741),
       .Q (_________35857));
  xor2s1 ____9__499585(.DIN1 (_________35776), .DIN2 (_________35806),
       .Q (_________36079));
  nor2s1 ____0__499586(.DIN1 (____9_9__36114), .DIN2 (_________35756),
       .Q (_________35805));
  xor2s1 ____0__499587(.DIN1 (______0__35803), .DIN2 (_________38871),
       .Q (_________35804));
  nor2s1 ____0__499588(.DIN1 (_______22186), .DIN2 (_________35758), .Q
       (______9__35802));
  nnd2s1 ____0__499589(.DIN1 (______9__35822), .DIN2
       (_________________________________________0___21856), .Q
       (_________35801));
  or2s1 ____0__499590(.DIN1
       (_________________________________________0___21856), .DIN2
       (______9__35822), .Q (_________35800));
  and2s1 ____0__499591(.DIN1 (______9__35822), .DIN2
       (_____________________________________0___0___21760), .Q
       (_________35798));
  or2s1 ____0__499592(.DIN1
       (_____________________________________0___0___21760), .DIN2
       (______9__35822), .Q (_________35797));
  nor2s1 ____0__499593(.DIN1 (____9____35272), .DIN2 (_________35761),
       .Q (_____09__35842));
  xor2s1 _______499594(.DIN1 (_________35772), .DIN2 (______9__35773),
       .Q (_________36340));
  nor2s1 ____9__499595(.DIN1 (_____9__23492), .DIN2 (_________35795),
       .Q (_________35796));
  and2s1 ____9__499596(.DIN1 (_________35791), .DIN2 (________22376),
       .Q (_________35794));
  nnd2s1 ____9_499597(.DIN1 (_________34999), .DIN2 (______9__35754),
       .Q (______0__35793));
  nnd2s1 ____9__499598(.DIN1 (_________35791), .DIN2 (inData[14]), .Q
       (______9__35792));
  nor2s1 ____9__499599(.DIN1 (_________35618), .DIN2 (_________35789),
       .Q (_________35790));
  xor2s1 ____9_499600(.DIN1 (___0_____40626), .DIN2
       (_____________________________________9______21877), .Q
       (_________35788));
  xor2s1 ____9__499601(.DIN1 (_________32309), .DIN2 (_________35767),
       .Q (_________35787));
  or2s1 ____0__499602(.DIN1 (____99__26498), .DIN2 (_____0___35737), .Q
       (_________35786));
  or2s1 ____499603(.DIN1 (______0__35784), .DIN2 (_________35753), .Q
       (_________35785));
  nnd2s1 ____00_499604(.DIN1 (_________35750), .DIN2 (_________36643),
       .Q (______9__35783));
  and2s1 ____00_499605(.DIN1 (_________35781), .DIN2 (______9__33584),
       .Q (_________35782));
  hi1s1 ____0_499606(.DIN (_________35779), .Q (_________35780));
  nor2s1 ____9__499607(.DIN1 (_________35751), .DIN2 (_________35749),
       .Q (_____9___35919));
  xor2s1 ____09_499608(.DIN1 (____99___35287), .DIN2 (_________35760),
       .Q (_________35778));
  nor2s1 ____0__499609(.DIN1 (_________31657), .DIN2 (_________35776),
       .Q (_________35777));
  xor2s1 ____0__499610(.DIN1 (_________35757), .DIN2 (___0_____40592),
       .Q (_________35775));
  dffacs1 _______________499611(.CLRB (reset), .CLK (clk), .DIN
       (_________35776), .Q (outData[6]));
  nor2s1 _______499612(.DIN1 (______9__35773), .DIN2 (_________35772),
       .Q (______0__35774));
  nor2s1 ____0__499613(.DIN1 (_____0___35477), .DIN2 (_____0___35743),
       .Q (_________35771));
  nnd2s1 ____0_499614(.DIN1 (______9__31939), .DIN2 (_________35776),
       .Q (_________35770));
  nnd2s1 _______499615(.DIN1 (_________35772), .DIN2 (____9___28553),
       .Q (_________35769));
  nor2s1 ____0__499616(.DIN1 (______0__33669), .DIN2 (_____0___35739),
       .Q (_________35817));
  nnd2s1 ____0__499617(.DIN1 (_________31822), .DIN2 (_________35776),
       .Q (______9__35812));
  xor2s1 ____0__499618(.DIN1 (_____9___35733), .DIN2 (_________36856),
       .Q (_____9___35826));
  dffacs1 _________________________________________0_____499619(.CLRB
       (reset), .CLK (clk), .DIN (_________35746), .QN
       (_____________________________________0_____));
  xor2s1 ____0__499620(.DIN1 (___0_____40630), .DIN2 (_________37789),
       .Q (_________35847));
  dffacs1 _______________________________________________499621(.CLRB
       (reset), .CLK (clk), .DIN (_____0___35740), .Q (___0_____40509));
  nnd2s1 ____0__499622(.DIN1 (_________35767), .DIN2 (_________35859),
       .Q (_________35768));
  nnd2s1 ____99_499623(.DIN1 (____00__28471), .DIN2 (___0_____40626),
       .Q (_________35766));
  nnd2s1 ____0__499624(.DIN1 (_________35767), .DIN2 (____0____31531),
       .Q (______0__35765));
  nor2s1 ____0__499625(.DIN1 (___0_____40626), .DIN2 (_____9__25537),
       .Q (______9__35764));
  nor2s1 ____0__499626(.DIN1
       (_____________________________________________21896), .DIN2
       (_________35767), .Q (_________35763));
  nor2s1 ____9__499627(.DIN1 (_____99__35735), .DIN2 (______0__35745),
       .Q (_________35762));
  nor2s1 ____09_499628(.DIN1 (____9____35273), .DIN2 (_________35760),
       .Q (_________35761));
  nor2s1 ____0__499629(.DIN1 (____0_0__37159), .DIN2 (_____9___35732),
       .Q (_________35759));
  and2s1 ____0__499630(.DIN1 (_________35757), .DIN2 (____9__22189), .Q
       (_________35758));
  xor2s1 ____0__499631(.DIN1 (_____0___35738), .DIN2 (_________33700),
       .Q (_________35756));
  nnd2s1 ____0__499632(.DIN1 (______9__31824), .DIN2 (_________35767),
       .Q (_________35779));
  nor2s1 ____0__499633(.DIN1 (____0____34446), .DIN2 (_____9___35734),
       .Q (_________35808));
  xor2s1 ____09_499634(.DIN1 (______0__35451), .DIN2 (_________40842),
       .Q (______9__35822));
  and2s1 ____0__499635(.DIN1 (______0__35721), .DIN2 (_________37223),
       .Q (______0__35755));
  nnd2s1 ____499636(.DIN1 (_________35448), .DIN2 (_________35729), .Q
       (______9__35754));
  nnd2s1 ____0__499637(.DIN1 (____9____35247), .DIN2 (_________35719),
       .Q (_________35753));
  nor2s1 ____00_499638(.DIN1 (_________35748), .DIN2 (_________35751),
       .Q (_________35752));
  nor2s1 ____0__499639(.DIN1 (__9999), .DIN2 (______9__35720), .Q
       (_________35750));
  nor2s1 ____99_499640(.DIN1 (_________35748), .DIN2 (_________35747),
       .Q (_________35749));
  nnd2s1 ____0_499641(.DIN1 (________25426), .DIN2 (_________35724), .Q
       (_________35746));
  nnd2s1 ____00_499642(.DIN1 (_________35722), .DIN2 (_________35727),
       .Q (_________35795));
  nor2s1 ____00_499643(.DIN1 (_________35728), .DIN2 (______0__35745),
       .Q (_________35791));
  xor2s1 ____0__499644(.DIN1 (_________35708), .DIN2 (_____09__35744),
       .Q (_________35789));
  hi1s1 ____0__499645(.DIN (_________35767), .Q (_________35776));
  nor2s1 ____09_499646(.DIN1 (_________35429), .DIN2 (_________40842),
       .Q (_____0___35743));
  nor2s1 ____0__499647(.DIN1 (_________35726), .DIN2 (_____0___35741),
       .Q (_____0___35742));
  nnd2s1 _____0_499648(.DIN1 (_________35712), .DIN2 (_________37504),
       .Q (_____0___35740));
  nor2s1 ____0__499649(.DIN1 (_________33680), .DIN2 (_____0___35738),
       .Q (_____0___35739));
  xor2s1 ____0_499650(.DIN1 (____0____34448), .DIN2 (_________40844),
       .Q (_____0___35737));
  nor2s1 ____09_499651(.DIN1 (_________35609), .DIN2 (_________35716),
       .Q (______0__35803));
  xor2s1 ____0__499652(.DIN1 (_________40846), .DIN2 (_____9___35917),
       .Q (_________35781));
  dffacs1 _______________________________________________499653(.CLRB
       (reset), .CLK (clk), .DIN (_________35725), .QN
       (___0__0__40541));
  dffacs1 _____________________________________________9_499654(.CLRB
       (reset), .CLK (clk), .DIN (_________35717), .QN
       (_________________________________________9___21779));
  dffacs1 _______________________________________________499655(.CLRB
       (reset), .CLK (clk), .DIN (_________35723), .Q
       (_____________________________________________21775));
  xor2s1 _____9_499656(.DIN1 (_________35698), .DIN2 (_____00__35736),
       .Q (_________35772));
  xor2s1 ____0__499657(.DIN1 (___0_____40475), .DIN2 (___0__9__40490),
       .Q (_____99__35735));
  nor2s1 ____0__499658(.DIN1 (____0____34447), .DIN2 (_________40844),
       .Q (_____9___35734));
  nor2s1 _____0_499659(.DIN1 (_____9___35731), .DIN2 (_________40848),
       .Q (_____9___35733));
  xor2s1 ____499660(.DIN1 (_________35640), .DIN2 (_________35715), .Q
       (_____9___35732));
  nnd2s1 ____0__499661(.DIN1 (_________35707), .DIN2 (_________35668),
       .Q (_________35757));
  nnd2s1 _____0_499662(.DIN1 (_________40848), .DIN2 (_____9___35731),
       .Q (_____9___35829));
  dffacs1 _________________________________________9__9_(.CLRB (reset),
       .CLK (clk), .DIN (_________35706), .QN (___0_____40626));
  xor2s1 ____0__499663(.DIN1 (_________35697), .DIN2
       (_____________22100), .Q (_________35767));
  xor2s1 _____9_499664(.DIN1 (____0____36216), .DIN2
       (__________________________________9__________), .Q
       (_____9___35730));
  nor2s1 _____9_499665(.DIN1
       (__________________________________9__________), .DIN2
       (_________35699), .Q (____0____36223));
  nnd2s1 _______499666(.DIN1 (____9____35221), .DIN2 (_________35700),
       .Q (_________35760));
  dffacs1 _______________________________________________499667(.CLRB
       (reset), .CLK (clk), .DIN (_________35703), .QN
       (___0_9___40558));
  dffacs1 _______________________________________________499668(.CLRB
       (reset), .CLK (clk), .DIN (______9__35710), .Q (_____9___22050));
  dffacs1 _______________________________________________499669(.CLRB
       (reset), .CLK (clk), .DIN (_________35709), .QN
       (_____________________________________________21852));
  nnd2s1 ____0_499670(.DIN1 (______9__35693), .DIN2 (inData[8]), .Q
       (_________35729));
  nor2s1 ____0_499671(.DIN1 (_________35727), .DIN2 (___0_____40475),
       .Q (_________35728));
  xor2s1 ____0__499672(.DIN1 (______9__35667), .DIN2 (_________22033),
       .Q (_________35726));
  nnd2s1 ____0__499673(.DIN1 (_________35690), .DIN2 (_____90__35555),
       .Q (_________35725));
  nnd2s1 ____0__499674(.DIN1 (______0__35694), .DIN2 (_________35692),
       .Q (_________35724));
  nnd2s1 ____0__499675(.DIN1 (_____9___35013), .DIN2 (_________35695),
       .Q (_________35723));
  and2s1 ____0__499676(.DIN1 (_____0___35834), .DIN2 (___0_____40475),
       .Q (_________35722));
  xor2s1 ____0_499677(.DIN1 (___09____40678), .DIN2 (_________35674),
       .Q (______0__35721));
  nor2s1 ____0__499678(.DIN1 (___0_____40475), .DIN2
       (_________________________________________________________________________________________22090),
       .Q (_________35751));
  and2s1 ____0__499679(.DIN1
       (_________________________________________________________________________________________22090),
       .DIN2 (___0_____40475), .Q (_________35748));
  nor2s1 ____0__499680(.DIN1 (_________36288), .DIN2 (_________35689),
       .Q (______9__35720));
  nnd2s1 ____0__499681(.DIN1 (_________35718), .DIN2 (_________35688),
       .Q (_________35719));
  nnd2s1 _______499682(.DIN1 (_________35679), .DIN2 (___0____28781),
       .Q (_________35717));
  nor2s1 _______499683(.DIN1 (_________35634), .DIN2 (_________35715),
       .Q (_________35716));
  nnd2s1 ______499684(.DIN1 (____0____36216), .DIN2 (____99___36174),
       .Q (_________35714));
  nor2s1 _____499685(.DIN1 (____99___36174), .DIN2 (____0____36216), .Q
       (_________35713));
  nor2s1 _______499686(.DIN1 (__9_____29885), .DIN2 (_________35676),
       .Q (_________35712));
  xnr2s1 _______499687(.DIN1 (______0__35711), .DIN2 (_____0___35658),
       .Q (_____0___35738));
  dffacs1 _______________________________________________499688(.CLRB
       (reset), .CLK (clk), .DIN (______0__35684), .Q
       (______0___22055));
  nnd2s1 _____0_499689(.DIN1 (_________35664), .DIN2 (________26526),
       .Q (______9__35710));
  nnd2s1 ____0__499690(.DIN1 (_________35673), .DIN2 (________24869),
       .Q (_________35709));
  nnd2s1 ____09_499691(.DIN1 (______9__35675), .DIN2 (_________35626),
       .Q (_________35708));
  nnd2s1 ____09_499692(.DIN1 (_________35696), .DIN2 (_________35670),
       .Q (_________35707));
  or2s1 ____0_499693(.DIN1 (_________35705), .DIN2 (_________35666), .Q
       (_________35706));
  xor2s1 ______499694(.DIN1 (___0__0__40521), .DIN2 (_________35685),
       .Q (_________35704));
  nnd2s1 _______499695(.DIN1 (_________35665), .DIN2 (_________36621),
       .Q (_________35703));
  nnd2s1 _______499696(.DIN1 (_____0___35656), .DIN2 (______0__35701),
       .Q (_________35702));
  nor2s1 ______499697(.DIN1 (______9__35602), .DIN2 (_____0___35654),
       .Q (_________35700));
  nor2s1 _______499698(.DIN1 (_____9___36094), .DIN2 (_____9___35651),
       .Q (_________35699));
  nor2s1 _______499699(.DIN1 (_____0__22489), .DIN2 (_____9___35649),
       .Q (_________35698));
  dffacs1 _______________________________________________499700(.CLRB
       (reset), .CLK (clk), .DIN (_____99__35652), .QN
       (___0_____40526));
  xor2s1 _______499701(.DIN1 (_________35696), .DIN2 (___0_____40593),
       .Q (_________35697));
  nnd2s1 ____0__499702(.DIN1 (______0__35694), .DIN2 (_____9___35646),
       .Q (_________35695));
  xnr2s1 ____0__499703(.DIN1
       (_____________________________________________21775), .DIN2
       (_________35691), .Q (______9__35693));
  xnr2s1 ____0_499704(.DIN1 (_________35691), .DIN2 (______0_), .Q
       (_________35692));
  and2s1 _____499705(.DIN1 (_____9___35645), .DIN2 (________26834), .Q
       (_________35690));
  xor2s1 ______499706(.DIN1 (_________35630), .DIN2
       (_____________________________________________21852), .Q
       (_________35689));
  xor2s1 _______499707(.DIN1 (___0_____40593), .DIN2 (___0_____40627),
       .Q (_________35688));
  xor2s1 ______499708(.DIN1
       (_________________________________________0___21798), .DIN2
       (_________35671), .Q (_________35687));
  dffacs1 _____________________________________________0_499709(.CLRB
       (reset), .CLK (clk), .DIN (_____90__35644), .QN
       (___0_____40475));
  nor2s1 _______499710(.DIN1
       (_________________________________________0___21798), .DIN2
       (_________35685), .Q (_________35686));
  nnd2s1 _______499711(.DIN1 (______9__35643), .DIN2 (______9__35683),
       .Q (______0__35684));
  nnd2s1 _______499712(.DIN1 (_________35685), .DIN2
       (_________________________________________0___21798), .Q
       (_________35682));
  nnd2s1 _______499713(.DIN1 (_________35642), .DIN2 (_________35680),
       .Q (_________35681));
  or2s1 ______499714(.DIN1 (_________36521), .DIN2 (_________35641), .Q
       (_________35679));
  xor2s1 _______499715(.DIN1 (_________35606), .DIN2 (_________35677),
       .Q (_________35678));
  nor2s1 _______499716(.DIN1 (_________41090), .DIN2 (_________35633),
       .Q (_________35676));
  xor2s1 _______499717(.DIN1 (______0__40850), .DIN2 (______0__35711),
       .Q (_________35715));
  xor2s1 _______499718(.DIN1 (_____0__27443), .DIN2 (_____9___35648),
       .Q (____0____36216));
  or2s1 _______499719(.DIN1 (_________35674), .DIN2 (______0__35628),
       .Q (______9__35675));
  nnd2s1 _______499720(.DIN1 (_________35625), .DIN2 (____9____35258),
       .Q (_________35673));
  and2s1 _______499721(.DIN1 (_________35671), .DIN2 (___0__0__40521),
       .Q (_________35672));
  nnd2s1 _______499722(.DIN1 (___0_____40593), .DIN2
       (_____________22100), .Q (_________35670));
  nor2s1 ______499723(.DIN1 (___0__0__40521), .DIN2 (_________35671),
       .Q (_________35669));
  or2s1 ______499724(.DIN1 (_____________22100), .DIN2
       (___0_____40593), .Q (_________35668));
  and2s1 _______499725(.DIN1 (___0_____40593), .DIN2 (___0_____40592),
       .Q (______9__35667));
  nnd2s1 ____09_499726(.DIN1 (_________35614), .DIN2 (____9___25027),
       .Q (_________35666));
  nor2s1 _______499727(.DIN1 (________27061), .DIN2 (_________35617),
       .Q (_________35665));
  nnd2s1 _______499728(.DIN1 (_________35615), .DIN2 (_________35663),
       .Q (_________35664));
  nnd2s1 ______499729(.DIN1 (_________35621), .DIN2 (_________35629),
       .Q (_________36054));
  and2s1 ______499730(.DIN1 (_________35607), .DIN2 (____9____37049),
       .Q (_________35662));
  nnd2s1 _______499731(.DIN1 (_________35613), .DIN2 (_________33588),
       .Q (_____0___35658));
  nnd2s1 ______499732(.DIN1 (____9____32436), .DIN2 (___0_____40593),
       .Q (_____0___35657));
  hi1s1 _____9_499733(.DIN (_____0___35655), .Q (_____0___35656));
  nor2s1 _____0_499734(.DIN1 (_________35604), .DIN2 (_____00__35653),
       .Q (_____0___35654));
  nnd2s1 _______499735(.DIN1 (_________35601), .DIN2 (____0____35361),
       .Q (_____99__35652));
  nnd2s1 _______499736(.DIN1 (_____9___35650), .DIN2 (____9____36135),
       .Q (_____9___35651));
  nor2s1 _____9_499737(.DIN1 (_______22221), .DIN2 (_____9___35648), .Q
       (_____9___35649));
  nor2s1 _____9_499738(.DIN1 (_______________22075), .DIN2
       (____9____36135), .Q (_____9___35647));
  dffacs1 __________________499739(.CLRB (reset), .CLK (clk), .DIN
       (_________35624), .QN (_______________22069));
  xor2s1 _______499740(.DIN1
       (_____________________________________0_____), .DIN2
       (___0_____40543), .Q (_____9___35646));
  nnd2s1 _______499741(.DIN1 (_________35596), .DIN2 (_________35394),
       .Q (_____9___35645));
  nnd2s1 _____0_499742(.DIN1 (_________35595), .DIN2 (______0__35181),
       .Q (_____90__35644));
  nor2s1 _______499743(.DIN1 (________26469), .DIN2 (______0__35594),
       .Q (______9__35643));
  xor2s1 _______499744(.DIN1 (_____9___33613), .DIN2 (______0__35612),
       .Q (_________35642));
  xor2s1 _______499745(.DIN1 (_____9___34562), .DIN2 (_________35600),
       .Q (_________35641));
  xor2s1 _____9_499746(.DIN1 (________26157), .DIN2 (_________35608),
       .Q (_________35640));
  hi1s1 _______499747(.DIN (_________35671), .Q (_________35685));
  xor2s1 ______499748(.DIN1 (_________35637), .DIN2 (___090__23301), .Q
       (_________35638));
  nor2s1 _____499749(.DIN1 (_________37412), .DIN2 (_________35597), .Q
       (______0__35636));
  nor2s1 _______499750(.DIN1 (________25534), .DIN2 (_________35631),
       .Q (_________35634));
  xor2s1 _______499751(.DIN1 (____9____35220), .DIN2 (______0__35603),
       .Q (_________35633));
  xor2s1 ______499752(.DIN1
       (__________________________________9__________), .DIN2
       (_____9___36094), .Q (_________35632));
  nnd2s1 _______499753(.DIN1 (_________35631), .DIN2
       (_________________________________________9___21855), .Q
       (______0__35701));
  nor2s1 _____0_499754(.DIN1
       (_________________________________________9___21855), .DIN2
       (_________35631), .Q (_____0___35655));
  dffacs1 _______________________________________________499755(.CLRB
       (reset), .CLK (clk), .DIN (______9__35593), .QN
       (_________22039));
  nnd2s1 _____9_499756(.DIN1 (_________35581), .DIN2 (_________35629),
       .Q (_________35630));
  nor2s1 _______499757(.DIN1 (___0_____40543), .DIN2 (______9__35627),
       .Q (______0__35628));
  nnd2s1 _______499758(.DIN1 (______9__35627), .DIN2 (___0_____40543),
       .Q (_________35626));
  xor2s1 _______499759(.DIN1 (_____0___35567), .DIN2 (_________35580),
       .Q (_________35625));
  nnd2s1 _______499760(.DIN1 (_________35588), .DIN2 (___9_9__28663),
       .Q (_________35624));
  or2s1 ______499761(.DIN1
       (_____________________________________________21852), .DIN2
       (_________35582), .Q (_________35621));
  nor2s1 _____9_499762(.DIN1 (______9__35619), .DIN2 (_________35618),
       .Q (______0__35620));
  nor2s1 _______499763(.DIN1 (_________36521), .DIN2 (_________35583),
       .Q (_________35617));
  xor2s1 _____499764(.DIN1 (_____0___35569), .DIN2 (_________40854), .Q
       (_________35615));
  nnd2s1 _______499765(.DIN1 (_________35590), .DIN2 (_____9___36005),
       .Q (_________35614));
  or2s1 ______499766(.DIN1 (___0_____40543), .DIN2
       (_____________________________________0_____), .Q
       (_________35691));
  xor2s1 _____9_499767(.DIN1 (_____0___35572), .DIN2 (_________35844),
       .Q (_________35671));
  dffacs1 _____________________________________499768(.CLRB (reset),
       .CLK (clk), .DIN (_________35586), .QN (___0_____40593));
  nnd2s1 _____0_499769(.DIN1 (______0__35612), .DIN2 (_________33567),
       .Q (_________35613));
  xor2s1 ______499770(.DIN1 (_________35610), .DIN2 (___9_0___39166),
       .Q (_________35611));
  nor2s1 _______499771(.DIN1 (___0__0__40571), .DIN2 (_________35608),
       .Q (_________35609));
  xor2s1 _______499772(.DIN1 (_____00__35565), .DIN2 (_________38395),
       .Q (_________35607));
  nnd2s1 _____0_499773(.DIN1 (_____9___36094), .DIN2 (_________37320),
       .Q (_________35606));
  or2s1 _____0_499774(.DIN1 (_________37320), .DIN2 (_____9___36094),
       .Q (_________35605));
  nor2s1 _______499775(.DIN1 (________25910), .DIN2 (______0__35603),
       .Q (_________35604));
  and2s1 _______499776(.DIN1 (______0__35603), .DIN2
       (_____________________________________________21810), .Q
       (______9__35602));
  nor2s1 _______499777(.DIN1 (_________35578), .DIN2 (_________35507),
       .Q (_________35601));
  nnd2s1 _______499778(.DIN1 (_________35600), .DIN2 (_____9___34565),
       .Q (_____0___35659));
  nor2s1 _______499779(.DIN1 (_________35598), .DIN2 (_________35599),
       .Q (_________35635));
  nor2s1 _______499780(.DIN1 (________22890), .DIN2 (_________35577),
       .Q (_____9___35648));
  nnd2s1 _______499781(.DIN1 (_________35599), .DIN2 (_________35598),
       .Q (_________35661));
  dffacs1 _______________________________________________499782(.CLRB
       (reset), .CLK (clk), .DIN (_________35589), .QN
       (_____________________________________________21809));
  hi1s1 _______499783(.DIN (_________35597), .Q (____9____36135));
  dffacs1 __________________499784(.CLRB (reset), .CLK (clk), .DIN
       (______0__35575), .QN
       (______________________________________________________________________________________0__22096));
  xor2s1 ______499785(.DIN1 (_________34246), .DIN2 (_________35579),
       .Q (_________35596));
  nor2s1 _______499786(.DIN1 (________24975), .DIN2 (_____0___35571),
       .Q (_________35595));
  nor2s1 _______499787(.DIN1 (____99__26498), .DIN2 (_____0___35568),
       .Q (______0__35594));
  nnd2s1 _______499788(.DIN1 (_____9___35563), .DIN2 (____0____37173),
       .Q (______9__35593));
  xor2s1 _______499789(.DIN1 (_________35532), .DIN2 (_________36087),
       .Q (_________35592));
  nor2s1 _______499790(.DIN1
       (__________________________________9__________), .DIN2
       (_____9___35650), .Q (_________35591));
  nor2s1 _______499791(.DIN1 (_____99__35564), .DIN2 (_____0___35573),
       .Q (_________35639));
  xor2s1 ______499792(.DIN1 (________22892), .DIN2 (_________35576), .Q
       (_________35597));
  hi1s1 _______499793(.DIN (_________35608), .Q (_________35631));
  dffacs1 _______________________________________________499794(.CLRB
       (reset), .CLK (clk), .DIN (_____0___35570), .Q (___0_____40542));
  xor2s1 _______499795(.DIN1 (_________35517), .DIN2 (_________35546),
       .Q (_________35590));
  or2s1 _____0_499796(.DIN1 (______9__35554), .DIN2 (_________35418),
       .Q (_________35589));
  or2s1 _____0_499797(.DIN1 (_________35587), .DIN2 (_________35553),
       .Q (_________35588));
  or2s1 _____0_499798(.DIN1 (______0__35784), .DIN2 (_________35551),
       .Q (_________35586));
  xor2s1 _______499799(.DIN1 (_________35516), .DIN2 (______9__35584),
       .Q (______0__35585));
  xor2s1 ______499800(.DIN1 (_________35512), .DIN2 (_________36512),
       .Q (_________35583));
  hi1s1 ______499801(.DIN (_________35581), .Q (_________35582));
  nnd2s1 _______499802(.DIN1 (_________35549), .DIN2 (_____0___34569),
       .Q (_________35629));
  or2s1 _______499803(.DIN1 (_________35550), .DIN2 (_________35580),
       .Q (_________35616));
  nor2s1 ______499804(.DIN1 (_____9___35557), .DIN2 (_________34995),
       .Q (_________35618));
  nor2s1 _______499805(.DIN1 (______0__35416), .DIN2 (_________35547),
       .Q (_________35747));
  nor2s1 _____499806(.DIN1 (_________34245), .DIN2 (_________35579), .Q
       (_________35623));
  dffacs1 _______________________________________________499807(.CLRB
       (reset), .CLK (clk), .DIN (_____9___35560), .Q (___0_____40543));
  nor2s1 _______499808(.DIN1 (_________35533), .DIN2 (_________35680),
       .Q (_________35578));
  nor2s1 _______499809(.DIN1 (________22891), .DIN2 (_________35576),
       .Q (_________35577));
  nnd2s1 _______499810(.DIN1 (_________35538), .DIN2 (_________35491),
       .Q (______0__35575));
  nor2s1 _____499811(.DIN1 (_____09__35574), .DIN2 (______0__35528), .Q
       (_________35637));
  nor2s1 _______499812(.DIN1 (_________34808), .DIN2 (_________35540),
       .Q (_________35599));
  nor2s1 _______499813(.DIN1 (_________35456), .DIN2 (_________35541),
       .Q (______0__35612));
  xor2s1 _______499814(.DIN1 (______9__35508), .DIN2 (_________36301),
       .Q (_________35600));
  nor2s1 _____499815(.DIN1 (_________34996), .DIN2 (_________35535), .Q
       (______0__35603));
  xor2s1 _______499816(.DIN1 (_________35505), .DIN2 (_____0___35573),
       .Q (_________35608));
  dffacs1 _____________________________________________0_499817(.CLRB
       (reset), .CLK (clk), .DIN (_________35543), .QN
       (___0_____40527));
  dffacs1 _______________________________________________499818(.CLRB
       (reset), .CLK (clk), .DIN (_____9___35556), .QN
       (___0_9___40559));
  dffacs1 _____________________0_499819(.CLRB (reset), .CLK (clk), .DIN
       (_________35542), .QN (_________________0_));
  xnr2s1 _______499820(.DIN1 (_________37412), .DIN2 (_________35503),
       .Q (_____9___36094));
  dffacs2 __________________499821(.CLRB (reset), .CLK (clk), .DIN
       (_________35552), .QN (_______________22070));
  xor2s1 _______499822(.DIN1 (_____9___34841), .DIN2 (_________35539),
       .Q (_____0___35572));
  nor2s1 _______499823(.DIN1 (_____0___35834), .DIN2 (_________35524),
       .Q (_____0___35571));
  nnd2s1 _______499824(.DIN1 (______9__35518), .DIN2 (_____9___35467),
       .Q (_____0___35570));
  xor2s1 ______499825(.DIN1 (_________35495), .DIN2 (_____0___35566),
       .Q (_____0___35569));
  xor2s1 _______499826(.DIN1 (____0____34456), .DIN2 (_________35492),
       .Q (_____0___35568));
  xor2s1 _______499827(.DIN1
       (_____________________________________________21835), .DIN2
       (_____0___35566), .Q (_____0___35567));
  nor2s1 ______499828(.DIN1
       (_____________________________________________21797), .DIN2
       (_________35003), .Q (______9__35619));
  nnd2s1 _______499829(.DIN1 (_________35548), .DIN2 (_________34514),
       .Q (_________35581));
  dffacs1 ________________0_(.CLRB (reset), .CLK (clk), .DIN
       (_________35515), .QN (___0__0__40413));
  xor2s1 _______499830(.DIN1 (_________35004), .DIN2 (_________35534),
       .Q (_____00__35565));
  xor2s1 _______499831(.DIN1 (_________35485), .DIN2 (_________37199),
       .Q (_____99__35564));
  nor2s1 _____499832(.DIN1 (__9_____30212), .DIN2 (_________35506), .Q
       (_____9___35563));
  nnd2s1 _____0_499833(.DIN1 (_____9___35562), .DIN2 (_____9___35561),
       .Q (_________35610));
  dffacs1 _______________________________________________499834(.CLRB
       (reset), .CLK (clk), .DIN (_________35514), .QN
       (_____________________________________________21766));
  xor2s1 _______499835(.DIN1 (_____0___35478), .DIN2 (_________38372),
       .Q (_____9___35650));
  dffacs1 _______________________________________________499836(.CLRB
       (reset), .CLK (clk), .DIN (_________35513), .Q
       (_____________________________________________21778));
  dffacs1 ______________________________________________499837(.CLRB
       (reset), .CLK (clk), .DIN (_________35522), .QN
       (____________________________________________21761));
  dffacs1 _________________________________________0____(.CLRB (reset),
       .CLK (clk), .DIN (______0__35519), .QN
       (_____________________________________0______21754));
  or2s1 _____0_499838(.DIN1 (_____9___35559), .DIN2 (_________35502),
       .Q (_____9___35560));
  xor2s1 _______499839(.DIN1 (_____9___35463), .DIN2 (___0__9__40540),
       .Q (_____9___35558));
  hi1s1 _______499840(.DIN
       (_____________________________________________21797), .Q
       (_____9___35557));
  nnd2s1 _______499841(.DIN1 (_________35501), .DIN2 (_____90__35555),
       .Q (_____9___35556));
  nor2s1 ______499842(.DIN1 (_________35493), .DIN2 (______9__35498),
       .Q (______9__35554));
  nnd2s1 _______499843(.DIN1 (_________35500), .DIN2 (______0__35537),
       .Q (_________35553));
  nnd2s1 _______499844(.DIN1 (______0__35499), .DIN2 (__9_____30228),
       .Q (_________35552));
  nnd2s1 _______499845(.DIN1 (________28532), .DIN2 (_________35494),
       .Q (_________35551));
  and2s1 _______499846(.DIN1 (______9__35544), .DIN2
       (_____________________________________________21835), .Q
       (_________35550));
  hi1s1 _______499847(.DIN (_________35548), .Q (_________35549));
  and2s1 ______499848(.DIN1 (_________35546), .DIN2 (_________35417),
       .Q (_________35547));
  or2s1 _______499849(.DIN1
       (_____________________________________________21835), .DIN2
       (______9__35544), .Q (______0__35545));
  nor2s1 ______499850(.DIN1 (_________33950), .DIN2 (_________35497),
       .Q (_________35579));
  nnd2s1 _____9_499851(.DIN1 (_________35118), .DIN2 (_________35490),
       .Q (_________35543));
  nnd2s1 _____0_499852(.DIN1 (______0__35489), .DIN2 (__9_____29834),
       .Q (_________35542));
  nor2s1 _____0_499853(.DIN1 (_____09__35480), .DIN2 (_________40854),
       .Q (_________35541));
  nor2s1 _____0_499854(.DIN1 (_________34823), .DIN2 (_________35539),
       .Q (_________35540));
  nnd2s1 _______499855(.DIN1 (_________40852), .DIN2 (______0__35537),
       .Q (_________35538));
  xor2s1 _______499856(.DIN1 (___0_____40539), .DIN2 (_________35520),
       .Q (______9__35536));
  nor2s1 ______499857(.DIN1 (_________34994), .DIN2 (_________35534),
       .Q (_________35535));
  nor2s1 _______499858(.DIN1 (____9____38963), .DIN2 (_________35486),
       .Q (_________35533));
  nor2s1 _______499859(.DIN1 (_________41367), .DIN2 (_________35482),
       .Q (_________35532));
  nor2s1 _____9_499860(.DIN1 (_________35530), .DIN2 (_________35529),
       .Q (_________35531));
  hi1s1 _______499861(.DIN (______9__35527), .Q (______0__35528));
  nor2s1 _______499862(.DIN1 (___9___22269), .DIN2 (_____0___35472), .Q
       (_________35576));
  xor2s1 _______499863(.DIN1 (_________35446), .DIN2 (_________35523),
       .Q (_________35524));
  nnd2s1 _______499864(.DIN1 (_________33977), .DIN2 (_____9___35469),
       .Q (_________35522));
  nor2s1 _______499865(.DIN1 (_________22043), .DIN2 (_________35520),
       .Q (_________35521));
  nnd2s1 ______499866(.DIN1 (_____9___35465), .DIN2 (________23994), .Q
       (______0__35519));
  xor2s1 _______499867(.DIN1 (_________33951), .DIN2 (_________35496),
       .Q (______9__35518));
  xor2s1 _______499868(.DIN1 (______0__35432), .DIN2
       (_________________________________________________________________________________________22094),
       .Q (_________35517));
  xor2s1 _______499869(.DIN1 (______9__35450), .DIN2 (_________22043),
       .Q (_________35516));
  nnd2s1 _____499870(.DIN1 (_____9___35462), .DIN2 (_________40856), .Q
       (_________35515));
  nnd2s1 _____0_499871(.DIN1 (_____90__35461), .DIN2 (___9____28661),
       .Q (_________35514));
  nnd2s1 _____0_499872(.DIN1 (_____99__35470), .DIN2 (___9____28678),
       .Q (_________35513));
  xor2s1 _______499873(.DIN1 (______0__35426), .DIN2 (_________35488),
       .Q (_________35512));
  xor2s1 _______499874(.DIN1 (_________35439), .DIN2 (___9_0___39705),
       .Q (_________35548));
  dffacs1 _______________________________________________499875(.CLRB
       (reset), .CLK (clk), .DIN (_____9___35468), .QN
       (_____________________________________________21797));
  and2s1 _______499876(.DIN1 (_________35520), .DIN2 (_________22043),
       .Q (_________35511));
  nor2s1 _______499877(.DIN1 (___0_____40539), .DIN2 (_________35520),
       .Q (_________35510));
  and2s1 _______499878(.DIN1 (_________35520), .DIN2 (___0_____40539),
       .Q (______0__35509));
  nor2s1 _______499879(.DIN1 (____0____34415), .DIN2 (_________35458),
       .Q (______9__35508));
  nnd2s1 _______499880(.DIN1 (____9____35253), .DIN2 (_________35454),
       .Q (_________35507));
  and2s1 _______499881(.DIN1 (_________35455), .DIN2 (____9_0__37080),
       .Q (_________35506));
  xor2s1 _______499882(.DIN1 (_________35504), .DIN2 (_________37321),
       .Q (_________35505));
  xor2s1 _______499883(.DIN1 (_____00__35471), .DIN2 (_________35844),
       .Q (_________35503));
  nnd2s1 _______499884(.DIN1 (_________37715), .DIN2 (__________22063),
       .Q (______9__35527));
  nnd2s1 _______499885(.DIN1 (_________37715), .DIN2 (___0_____40494),
       .Q (_____9___35561));
  or2s1 _______499886(.DIN1 (___0_____40494), .DIN2 (_________37715),
       .Q (_____9___35562));
  nor2s1 ______499887(.DIN1 (__________22063), .DIN2 (_________37715),
       .Q (_____09__35574));
  dffacs1 ____________________________________________9_499888(.CLRB
       (reset), .CLK (clk), .DIN (______9__35460), .Q
       (________________________________________9_));
  nnd2s1 ______499889(.DIN1 (_________35449), .DIN2 (________25443), .Q
       (_________35502));
  nor2s1 ______499890(.DIN1 (________27110), .DIN2 (_________35443), .Q
       (_________35501));
  nor2s1 _____9_499891(.DIN1 (_________35434), .DIN2 (____0____35363),
       .Q (_________35500));
  or2s1 _____9_499892(.DIN1 (_________35433), .DIN2 (______9__35498),
       .Q (______0__35499));
  nor2s1 _____9_499893(.DIN1 (_________33949), .DIN2 (_________35496),
       .Q (_________35497));
  xor2s1 _______499894(.DIN1 (_____9___22052), .DIN2 (___0_____40323),
       .Q (_________35495));
  nnd2s1 ______499895(.DIN1 (_________35718), .DIN2 (___0_____40627),
       .Q (_________35494));
  xnr2s1 ______499896(.DIN1 (_______________22069), .DIN2
       (_________35412), .Q (_________35493));
  xor2s1 _______499897(.DIN1 (_________35457), .DIN2 (_____99__36913),
       .Q (_________35492));
  nor2s1 _______499898(.DIN1 (________28455), .DIN2 (_________35437),
       .Q (_________35491));
  nnd2s1 _______499899(.DIN1 (_________35438), .DIN2 (________26525),
       .Q (_________35490));
  nor2s1 _______499900(.DIN1 (___9____28724), .DIN2 (______9__35431),
       .Q (______0__35489));
  xnr2s1 _______499901(.DIN1 (___0_____40323), .DIN2 (______0__35406),
       .Q (_________35539));
  xor2s1 _______499902(.DIN1 (______9__35425), .DIN2 (_________38456),
       .Q (_________35546));
  nnd2s1 ______499903(.DIN1 (_________35488), .DIN2 (_____09__35387),
       .Q (_________35525));
  dffacs1 _______________________________________________499904(.CLRB
       (reset), .CLK (clk), .DIN (_________35436), .QN
       (_____________________________________________21835));
  nnd2s1 _______499905(.DIN1 (_________35504), .DIN2 (_________37321),
       .Q (_________35487));
  nor2s1 _____9_499906(.DIN1 (_____0___35479), .DIN2 (_________35044),
       .Q (_________35486));
  nor2s1 _____9_499907(.DIN1 (_________37321), .DIN2 (_________35504),
       .Q (_________35485));
  nnd2s1 _______499908(.DIN1 (_________35504), .DIN2 (________27618),
       .Q (_________35484));
  or2s1 _______499909(.DIN1 (________27618), .DIN2 (_________35504), .Q
       (_________35483));
  and2s1 _______499910(.DIN1 (_________35504), .DIN2 (______0__35481),
       .Q (_________35482));
  nor2s1 _______499911(.DIN1 (_____0___35479), .DIN2 (_____0___35566),
       .Q (_____09__35480));
  or2s1 _______499912(.DIN1 (______0__35481), .DIN2 (_________35504),
       .Q (_____0___35478));
  nor2s1 _______499913(.DIN1 (_____9___38412), .DIN2 (_____0___35473),
       .Q (_____0___35477));
  and2s1 _______499914(.DIN1 (____00___38045), .DIN2
       (_________________________________________9_), .Q
       (_____0___35476));
  or2s1 _______499915(.DIN1
       (_________________________________________9_), .DIN2
       (____00___38045), .Q (_____0___35475));
  nnd2s1 _______499916(.DIN1 (_____0___35473), .DIN2 (_____9___38412),
       .Q (_____0___35474));
  nor2s1 _____0_499917(.DIN1 (___0_9__22333), .DIN2 (_____00__35471),
       .Q (_____0___35472));
  and2s1 ______499918(.DIN1 (_________37621), .DIN2 (___0_____40504),
       .Q (_________35530));
  nor2s1 _______499919(.DIN1 (___0_____40504), .DIN2 (_________37621),
       .Q (_________35529));
  nor2s1 _____0_499920(.DIN1 (_________34919), .DIN2 (_________35427),
       .Q (_________35534));
  or2s1 _______499921(.DIN1 (____99__26498), .DIN2 (_________35413), .Q
       (_____99__35470));
  nnd2s1 _______499922(.DIN1 (_____9___35464), .DIN2 (_________35420),
       .Q (_____9___35469));
  and2s1 _______499923(.DIN1 (_________35423), .DIN2 (_____9___35467),
       .Q (_____9___35468));
  nnd2s1 _______499924(.DIN1 (_________35422), .DIN2 (_____0___35741),
       .Q (_____9___35466));
  nnd2s1 _______499925(.DIN1 (_____9___35464), .DIN2 (_________35421),
       .Q (_____9___35465));
  xor2s1 _______499926(.DIN1 (_________35444), .DIN2 (____0____38091),
       .Q (_____9___35463));
  nor2s1 _______499927(.DIN1 (________28440), .DIN2 (______9__35415),
       .Q (_____9___35462));
  or2s1 _______499928(.DIN1 (____99__26498), .DIN2 (_________35414), .Q
       (_____90__35461));
  nnd2s1 _____0_499929(.DIN1 (______0__35171), .DIN2 (_________35424),
       .Q (______9__35460));
  nnd2s1 _______499930(.DIN1 (_________35452), .DIN2 (___0_____40495),
       .Q (_________35459));
  and2s1 _______499931(.DIN1 (_________35457), .DIN2 (____0_0__34414),
       .Q (_________35458));
  nor2s1 _______499932(.DIN1 (_____9___22052), .DIN2 (______9__35544),
       .Q (_________35456));
  xor2s1 ______499933(.DIN1 (_____0___34936), .DIN2 (_________40858),
       .Q (_________35455));
  or2s1 _____9_499934(.DIN1 (_____9___22052), .DIN2 (_________35147),
       .Q (_________35454));
  nor2s1 _______499935(.DIN1 (___0_____40495), .DIN2 (_________35452),
       .Q (_________35453));
  xor2s1 _______499936(.DIN1
       (_______________________________________________________________________________________),
       .DIN2 (______0__35481), .Q (______0__35451));
  hi1s1 _____0_499937(.DIN (______9__35450), .Q (_________35520));
  hi1s1 ______499938(.DIN (____00___38045), .Q (_________37715));
  or2s1 _______499939(.DIN1 (_________35448), .DIN2 (_________35403),
       .Q (_________35449));
  xor2s1 _______499940(.DIN1 (___0_____40522), .DIN2 (_________35390),
       .Q (_________35447));
  xor2s1 _______499941(.DIN1 (____09___35371), .DIN2 (____0____35365),
       .Q (_________35446));
  nor2s1 _______499942(.DIN1 (___0__9__40540), .DIN2 (_________35444),
       .Q (_________35445));
  nnd2s1 _______499943(.DIN1 (_________35395), .DIN2 (________26845),
       .Q (_________35443));
  nor2s1 _______499944(.DIN1 (___0_____40522), .DIN2 (_________35444),
       .Q (_________35442));
  and2s1 ______499945(.DIN1 (_________35444), .DIN2 (___0_____40522),
       .Q (______0__35441));
  and2s1 _______499946(.DIN1 (_________35444), .DIN2 (___0__9__40540),
       .Q (______9__35440));
  nor2s1 ______499947(.DIN1 (____0____35366), .DIN2 (_________35398),
       .Q (_________35439));
  nnd2s1 _____499948(.DIN1 (_________35391), .DIN2 (inData[2]), .Q
       (_________35438));
  nor2s1 _______499949(.DIN1 (_____0___32287), .DIN2 (_________40856),
       .Q (_________35437));
  and2s1 _______499950(.DIN1 (_________35393), .DIN2 (_________35435),
       .Q (_________35436));
  xor2s1 _______499951(.DIN1 (___0_____40476), .DIN2
       (_______________22070), .Q (_________35434));
  xor2s1 _______499952(.DIN1
       (_____________________________________________21809), .DIN2
       (___0_____40476), .Q (_________35433));
  xor2s1 _______499953(.DIN1 (___________________), .DIN2
       (___0_____40476), .Q (______0__35432));
  nor2s1 _______499954(.DIN1 (_____90__33805), .DIN2 (_________35400),
       .Q (_________35496));
  dffacs1 _________________________________________9____499955(.CLRB
       (reset), .CLK (clk), .DIN (_________35402), .Q (___0_____40627));
  nnd2s1 _____9_499956(.DIN1 (______0__35388), .DIN2 (________29385),
       .Q (______9__35431));
  nor2s1 ______499957(.DIN1
       (_______________________________________________________________________________________),
       .DIN2 (______0__35481), .Q (_________35429));
  xor2s1 ______499958(.DIN1 (_________37616), .DIN2 (____0____35352),
       .Q (_________35428));
  nor2s1 _______499959(.DIN1 (_________40858), .DIN2 (_________34941),
       .Q (_________35427));
  xor2s1 _______499960(.DIN1 (_________35408), .DIN2 (___0_____40572),
       .Q (______0__35426));
  nnd2s1 _____499961(.DIN1 (______0__35397), .DIN2 (____9____35214), .Q
       (_________35488));
  hi1s1 ______499962(.DIN (_____9___22052), .Q (_____0___35479));
  and2s1 _____9_499963(.DIN1 (______0__35481), .DIN2
       (_______________________________________________________________________________________),
       .Q (_____0___35473));
  nor2s1 _______499964(.DIN1 (____0____35340), .DIN2 (_________35389),
       .Q (_____00__35471));
  xor2s1 _______499965(.DIN1 (____09___35374), .DIN2
       (_______________22076), .Q (______9__35450));
  dffacs1 _______________________________________________499966(.CLRB
       (reset), .CLK (clk), .DIN (_________35401), .Q
       (_____________________________________________21777));
  nnd2s1 _____9_499967(.DIN1 (____09___35377), .DIN2 (__9_0___29997),
       .Q (____00___38045));
  hi1s1 _____0_499968(.DIN (_________35452), .Q (_________37621));
  xnr2s1 _______499969(.DIN1 (_____9___37002), .DIN2 (____0____35353),
       .Q (_________35504));
  nnd2s1 _____9_499970(.DIN1 (____0____35368), .DIN2 (____0____35330),
       .Q (______9__35425));
  nnd2s1 _______499971(.DIN1 (_____9___35464), .DIN2 (____09___35372),
       .Q (_________35424));
  xor2s1 _______499972(.DIN1 (______9__33832), .DIN2 (_________35399),
       .Q (_________35423));
  xor2s1 ______499973(.DIN1 (____0____35342), .DIN2 (____0____35367),
       .Q (_________35422));
  xor2s1 _______499974(.DIN1
       (____________________________________________21761), .DIN2
       (_________35419), .Q (_________35421));
  xnr2s1 _______499975(.DIN1
       (________________________________________9_), .DIN2
       (_________35419), .Q (_________35420));
  and2s1 _______499976(.DIN1 (____090__35370), .DIN2 (____9_0__37080),
       .Q (_________35418));
  nnd2s1 _____0_499977(.DIN1
       (_________________________________________________________________________________________22094),
       .DIN2 (___0_____40476), .Q (_________35417));
  nor2s1 _____0_499978(.DIN1 (___0_____40476), .DIN2
       (_________________________________________________________________________________________22094),
       .Q (______0__35416));
  nor2s1 _____0_499979(.DIN1 (___9____28662), .DIN2 (_________35392),
       .Q (______9__35415));
  xor2s1 _______499980(.DIN1 (____9____35236), .DIN2 (______9__35396),
       .Q (_________35414));
  xor2s1 _______499981(.DIN1
       (_____________________________________________21766), .DIN2
       (____0____35339), .Q (_________35413));
  nnd2s1 _______499982(.DIN1 (___0_____40476), .DIN2 (_________34167),
       .Q (_________35412));
  nor2s1 ______499983(.DIN1 (____0____35351), .DIN2 (_________35410),
       .Q (_________35411));
  nor2s1 _____9_499984(.DIN1 (_________22041), .DIN2 (_________35408),
       .Q (_________35409));
  xor2s1 _______499985(.DIN1 (___09___23302), .DIN2 (_____0___35386),
       .Q (_________35407));
  nor2s1 _______499986(.DIN1 (____09___35373), .DIN2 (____0_0__35360),
       .Q (______0__35406));
  and2s1 _____9_499987(.DIN1 (_________35408), .DIN2 (_________22041),
       .Q (______9__35405));
  nor2s1 _______499988(.DIN1 (____0____35321), .DIN2 (____0____35364),
       .Q (_________35457));
  xor2s1 _______499989(.DIN1 (_________37748), .DIN2 (_________35404),
       .Q (_________38154));
  xor2s1 _______499990(.DIN1
       (_____________________________________________21785), .DIN2
       (_________35404), .Q (_________35430));
  nor2s1 _______499991(.DIN1 (____999__35288), .DIN2 (____0____35354),
       .Q (_____0___35573));
  xor2s1 _______499992(.DIN1 (__9_0___29998), .DIN2 (____09___35376),
       .Q (_________35452));
  dffacs1 _______________________________________________499993(.CLRB
       (reset), .CLK (clk), .DIN (____0____35362), .Q (_____9___22052));
  dffacs1 _______________________________________________499994(.CLRB
       (reset), .CLK (clk), .DIN (____0_9__35369), .QN
       (_____________________________________________21796));
  xor2s1 ______499995(.DIN1 (____0_9__35333), .DIN2 (____9____35239),
       .Q (_________35403));
  or2s1 _______499996(.DIN1 (______0__35784), .DIN2 (____0____35348),
       .Q (_________35402));
  nnd2s1 _______499997(.DIN1 (____0____35345), .DIN2 (___0____28773),
       .Q (_________35401));
  nor2s1 ______499998(.DIN1 (_________33776), .DIN2 (_________35399),
       .Q (_________35400));
  nor2s1 _____9_499999(.DIN1 (____0____35346), .DIN2 (______0__40860),
       .Q (_________35398));
  or2s1 _______500000(.DIN1 (____9____35213), .DIN2 (______9__35396),
       .Q (______0__35397));
  nnd2s1 ______500001(.DIN1 (____0____35347), .DIN2 (_________35394),
       .Q (_________35395));
  xor2s1 ______500002(.DIN1 (____0_0__35324), .DIN2 (_________40862),
       .Q (_________35393));
  nor2s1 ______500003(.DIN1 (___09____40679), .DIN2 (________24808), .Q
       (_________35391));
  nnd2s1 _______500004(.DIN1 (____0____35344), .DIN2 (______0__34772),
       .Q (_________35674));
  hi1s1 _____0_500005(.DIN (_________35390), .Q (_________35444));
  nor2s1 _____0_500006(.DIN1 (_________38591), .DIN2 (____0____35338),
       .Q (_________35389));
  nor2s1 ______500007(.DIN1 (__909___29722), .DIN2 (____0_0__35341), .Q
       (______0__35388));
  nnd2s1 _______500008(.DIN1 (_____0___35386), .DIN2 (___0_____40572),
       .Q (_____09__35387));
  nor2s1 _______500009(.DIN1 (___0_____40572), .DIN2 (_____0___35386),
       .Q (_____0___35385));
  xor2s1 _______500010(.DIN1
       (_____________________________________________21769), .DIN2
       (_________38267), .Q (_____0___35383));
  nnd2s1 _______500011(.DIN1 (_________35404), .DIN2
       (_____________________________________________21769), .Q
       (_____0___35382));
  or2s1 _______500012(.DIN1
       (_____________________________________________21769), .DIN2
       (_________35404), .Q (_____0___35381));
  nor2s1 _______500013(.DIN1 (_________37748), .DIN2 (_________35404),
       .Q (_____0___35380));
  or2s1 _______500014(.DIN1
       (_____________________________________________21785), .DIN2
       (_________35404), .Q (_____00__35379));
  nnd2s1 _______500015(.DIN1 (_________35404), .DIN2
       (_____________________________________________21785), .Q
       (____099__35378));
  nnd2s1 _______500016(.DIN1 (____09___35376), .DIN2 (____09___35375),
       .Q (____09___35377));
  xor2s1 ______500017(.DIN1 (____0____35318), .DIN2 (____0____35302),
       .Q (______0__35481));
  or2s1 _____9_500018(.DIN1 (____09___35373), .DIN2 (____0_9__35359),
       .Q (____09___35374));
  xor2s1 _______500019(.DIN1
       (_____________________________________0______21754), .DIN2
       (___0_____40489), .Q (____09___35372));
  xor2s1 _______500020(.DIN1 (______0__40860), .DIN2 (___0_____40489),
       .Q (____09___35371));
  xor2s1 ______500021(.DIN1 (_________34777), .DIN2 (____0____35343),
       .Q (____090__35370));
  nnd2s1 _______500022(.DIN1 (____0_0__35334), .DIN2 (________26182),
       .Q (____0_9__35369));
  nnd2s1 _______500023(.DIN1 (____0____35367), .DIN2 (____0____35329),
       .Q (____0____35368));
  nor2s1 _______500024(.DIN1 (____0____35332), .DIN2 (____0____35365),
       .Q (____0____35366));
  nor2s1 _______500025(.DIN1 (____0_0__34396), .DIN2 (____0____35322),
       .Q (____0____35364));
  xor2s1 _______500026(.DIN1 (____0____35316), .DIN2 (______0__36598),
       .Q (_________35390));
  nor2s1 _______500027(.DIN1 (____0____35331), .DIN2 (____0____35363),
       .Q (_________35392));
  dffacs1 ____________________________________________9_500028(.CLRB
       (reset), .CLK (clk), .DIN (____0____35328), .QN
       (___0_____40476));
  nnd2s1 _____0_500029(.DIN1 (____0_9__35323), .DIN2 (____0____35361),
       .Q (____0____35362));
  nor2s1 _______500030(.DIN1 (____99___36174), .DIN2 (____0_9__35359),
       .Q (____0_0__35360));
  nor2s1 _______500031(.DIN1 (___0_____40505), .DIN2 (_________38267),
       .Q (____0____35358));
  nor2s1 _______500032(.DIN1 (____0____35356), .DIN2 (____0____35355),
       .Q (____0____35357));
  xnr2s1 ______500033(.DIN1 (_________38869), .DIN2 (____0____35300),
       .Q (____0____35354));
  xor2s1 ______500034(.DIN1 (____00___35297), .DIN2 (___9_9___39790),
       .Q (____0____35353));
  xnr2s1 _______500035(.DIN1 (__________22061), .DIN2 (____999__38037),
       .Q (____0____35352));
  hi1s1 _______500036(.DIN (____0_0__35350), .Q (____0____35351));
  hi1s1 _______500037(.DIN (_____0___35386), .Q (_________35408));
  dffacs1 _______________________________________________500038(.CLRB
       (reset), .CLK (clk), .DIN (____0____35326), .Q (___0_99__40560));
  dffacs1 _____________________________________________0_500039(.CLRB
       (reset), .CLK (clk), .DIN (____0____35319), .QN
       (_____90__22048));
  xor2s1 _______500040(.DIN1 (___0__0__40541), .DIN2 (____99___35285),
       .Q (____0_9__35349));
  nnd2s1 _______500041(.DIN1 (____0_9__35314), .DIN2 (________28505),
       .Q (____0____35348));
  xor2s1 _______500042(.DIN1 (____9____35215), .DIN2 (____00___35293),
       .Q (____0____35347));
  nor2s1 _______500043(.DIN1 (___0_____40489), .DIN2 (____9____34308),
       .Q (____0____35346));
  nnd2s1 _______500044(.DIN1 (____0____35311), .DIN2 (_________35394),
       .Q (____0____35345));
  or2s1 _____9_500045(.DIN1 (____0____35343), .DIN2 (_________34774),
       .Q (____0____35344));
  xor2s1 _______500046(.DIN1 (____99__25496), .DIN2 (___0_____40477),
       .Q (____0____35342));
  nnd2s1 ______500047(.DIN1 (____0____35308), .DIN2 (_____0__29235), .Q
       (____0_0__35341));
  nor2s1 _______500048(.DIN1 (______0__35161), .DIN2 (____0____35313),
       .Q (_________35399));
  nor2s1 _____9_500049(.DIN1 (____9_9__35269), .DIN2 (____0____35310),
       .Q (______9__35396));
  or2s1 ______500050(.DIN1 (___0_____40489), .DIN2
       (_____________________________________0______21754), .Q
       (_________35419));
  nor2s1 _______500051(.DIN1 (_________36291), .DIN2 (____0____35303),
       .Q (____0____35340));
  xnr2s1 ______500052(.DIN1 (_________40864), .DIN2 (____0_0__34396),
       .Q (____0____35339));
  nor2s1 _______500053(.DIN1 (________22609), .DIN2 (____0_9__35305),
       .Q (____0____35338));
  and2s1 _______500054(.DIN1 (____999__38037), .DIN2 (__________22061),
       .Q (____0____35337));
  or2s1 _______500055(.DIN1 (__________22061), .DIN2 (____999__38037),
       .Q (____0____35336));
  nnd2s1 _____500056(.DIN1 (____999__38037), .DIN2
       (_____________________________________________21784), .Q
       (____0_0__35350));
  nor2s1 _______500057(.DIN1 (____0_0__35315), .DIN2 (_________40862),
       .Q (_____0___35384));
  nor2s1 _______500058(.DIN1 (________29169), .DIN2 (____0____35307),
       .Q (____09___35376));
  nor2s1 ______500059(.DIN1
       (_____________________________________________21784), .DIN2
       (____999__38037), .Q (_________35410));
  xnr2s1 ______500060(.DIN1 (____000__35289), .DIN2 (____0____35299),
       .Q (_____0___35386));
  hi1s1 _____9_500061(.DIN (_________38267), .Q (_________35404));
  or2s1 _____500062(.DIN1 (______0__36766), .DIN2 (____00___35291), .Q
       (____0____35335));
  nnd2s1 _______500063(.DIN1 (____00___35295), .DIN2 (_________35186),
       .Q (____0_0__35334));
  xor2s1 ______500064(.DIN1 (____0____35312), .DIN2 (___90____39008),
       .Q (____0_9__35333));
  hi1s1 _______500065(.DIN (___0_____40489), .Q (____0____35332));
  nor2s1 _______500066(.DIN1 (___0_____40478), .DIN2 (___0_____40477),
       .Q (____0____35331));
  nnd2s1 _______500067(.DIN1
       (_________________________________________________________________________________________22095),
       .DIN2 (___0_____40477), .Q (____0____35330));
  or2s1 _______500068(.DIN1 (___0_____40477), .DIN2
       (_________________________________________________________________________________________22095),
       .Q (____0____35329));
  nnd2s1 _____500069(.DIN1 (____00___35296), .DIN2 (____9____35254), .Q
       (____0____35328));
  nor2s1 _____0_500070(.DIN1 (___0_____40477), .DIN2
       (______________________________________________________________________________________0__22096),
       .Q (____0____35327));
  nnd2s1 _____0_500071(.DIN1 (____00___35292), .DIN2 (_____90__35555),
       .Q (____0____35326));
  nor2s1 _______500072(.DIN1 (____9_9__36114), .DIN2 (____99___35281),
       .Q (____0____35325));
  xor2s1 _______500073(.DIN1
       (_____________________________________________21822), .DIN2
       (______0__33312), .Q (____0_0__35324));
  nor2s1 _______500074(.DIN1 (_________35078), .DIN2 (____99___35286),
       .Q (____0_9__35323));
  nor2s1 ______500075(.DIN1 (____0____35320), .DIN2 (_________40864),
       .Q (____0____35322));
  and2s1 ______500076(.DIN1 (_________40864), .DIN2 (____0____35320),
       .Q (____0____35321));
  nnd2s1 _____0_500077(.DIN1 (____00___35290), .DIN2 (____0____35361),
       .Q (____0____35319));
  xor2s1 _______500078(.DIN1 (____0____35304), .DIN2 (_________38666),
       .Q (____0____35318));
  nor2s1 _______500079(.DIN1 (___0_____40496), .DIN2 (____0____35317),
       .Q (____0____35356));
  nor2s1 _______500080(.DIN1 (______9__34523), .DIN2 (____99___35283),
       .Q (____0_9__35359));
  and2s1 _______500081(.DIN1 (____0____35317), .DIN2 (___0_____40496),
       .Q (____0____35355));
  xor2s1 ______500082(.DIN1 (__9_0___29996), .DIN2 (____0_0__35306), .Q
       (_________38267));
  xor2s1 ______500083(.DIN1 (____9_0__35262), .DIN2 (_____0___34756),
       .Q (____0____35316));
  nor2s1 _______500084(.DIN1
       (_____________________________________________21822), .DIN2
       (_________33288), .Q (____0_0__35315));
  nnd2s1 _____0_500085(.DIN1 (____9____35276), .DIN2 (_____0___35741),
       .Q (____0_9__35314));
  nor2s1 _____500086(.DIN1 (_________35163), .DIN2 (____0____35312), .Q
       (____0____35313));
  xor2s1 _______500087(.DIN1 (____9_0__35252), .DIN2 (______0__38256),
       .Q (____0____35311));
  and2s1 _______500088(.DIN1 (____9____35271), .DIN2 (____0____35309),
       .Q (____0____35310));
  and2s1 _______500089(.DIN1 (____9____35268), .DIN2 (________28960),
       .Q (____0____35308));
  nor2s1 _______500090(.DIN1 (_________34733), .DIN2 (____9____35275),
       .Q (____0____35343));
  dffacs1 _____________________________________________0_500091(.CLRB
       (reset), .CLK (clk), .DIN (____9_9__35279), .Q (___0_____40489));
  nor2s1 _______500092(.DIN1 (________29168), .DIN2 (____0_0__35306),
       .Q (____0____35307));
  and2s1 ______500093(.DIN1 (____0____35304), .DIN2 (___9____23174), .Q
       (____0_9__35305));
  or2s1 _______500094(.DIN1 (____0____35302), .DIN2 (____0____35304),
       .Q (____0____35303));
  nnd2s1 _______500095(.DIN1 (____0____35299), .DIN2 (____9____35267),
       .Q (____0____35300));
  nnd2s1 _______500096(.DIN1 (_________33288), .DIN2
       (_____________________________________________21822), .Q
       (____0_0__35298));
  xor2s1 _______500097(.DIN1 (____9____35250), .DIN2
       (_______________22075), .Q (____00___35297));
  nor2s1 _______500098(.DIN1 (_________34883), .DIN2 (____99___35282),
       .Q (____09___35373));
  hi1s1 _______500099(.DIN (____0____35317), .Q (____999__38037));
  dffacs1 _______________9_(.CLRB (reset), .CLK (clk), .DIN
       (____9____35278), .QN (__________9_));
  nor2s1 ______500100(.DIN1 (________28615), .DIN2 (____9____35257), .Q
       (____00___35296));
  xor2s1 _______500101(.DIN1 (____9____35249), .DIN2 (____00___35294),
       .Q (____00___35295));
  xor2s1 ______500102(.DIN1 (____9_0__35270), .DIN2 (___9_____39231),
       .Q (____00___35293));
  nor2s1 _______500103(.DIN1 (_____0__25721), .DIN2 (____9____35256),
       .Q (____00___35292));
  xor2s1 _______500104(.DIN1 (___0_____40632), .DIN2 (____9____35274),
       .Q (____00___35291));
  nor2s1 _______500105(.DIN1 (________24988), .DIN2 (____9____35259),
       .Q (____00___35290));
  nor2s1 _______500106(.DIN1 (___0____22304), .DIN2 (____9_9__35261),
       .Q (____0____35367));
  dffacs1 ______________________________________________500107(.CLRB
       (reset), .CLK (clk), .DIN (____9____35255), .QN
       (___0_____40477));
  nor2s1 _______500108(.DIN1 (____999__35288), .DIN2 (____9____35266),
       .Q (____000__35289));
  xor2s1 _______500109(.DIN1 (___0_____40523), .DIN2 (____99___35284),
       .Q (____99___35287));
  nnd2s1 _______500110(.DIN1 (____9_9__35251), .DIN2 (_________35080),
       .Q (____99___35286));
  xor2s1 _______500111(.DIN1 (____99___35284), .DIN2 (___090__23301),
       .Q (____99___35285));
  hi1s1 _____9_500112(.DIN (____99___35282), .Q (____99___35283));
  xor2s1 _____9_500113(.DIN1 (_________34802), .DIN2 (____9____35263),
       .Q (____99___35281));
  xor2s1 _______500114(.DIN1 (____9____35228), .DIN2 (________27618),
       .Q (____0____35317));
  xor2s1 _______500115(.DIN1 (___0_____40486), .DIN2 (____9____35211),
       .Q (____990__35280));
  nnd2s1 _______500116(.DIN1 (____9____35240), .DIN2 (________24623),
       .Q (____9_9__35279));
  nnd2s1 _______500117(.DIN1 (____0___25685), .DIN2 (____9_9__35242),
       .Q (____9____35278));
  nor2s1 _______500118(.DIN1 (____9____35264), .DIN2 (____99___35284),
       .Q (____9____35277));
  xor2s1 _______500119(.DIN1 (____0___22453), .DIN2 (____9____35260),
       .Q (____9____35276));
  nor2s1 _______500120(.DIN1 (____9____35274), .DIN2 (______9__34705),
       .Q (____9____35275));
  and2s1 _______500121(.DIN1 (____99___35284), .DIN2 (___0_____40523),
       .Q (____9____35273));
  nor2s1 _______500122(.DIN1 (___0_____40523), .DIN2 (____99___35284),
       .Q (____9____35272));
  nnd2s1 _______500123(.DIN1 (____9_0__35270), .DIN2 (___0_____40573),
       .Q (____9____35271));
  nor2s1 ______500124(.DIN1 (___0_____40573), .DIN2 (____9_0__35270),
       .Q (____9_9__35269));
  nor2s1 _______500125(.DIN1 (____9____35248), .DIN2 (____9____35244),
       .Q (____0____35312));
  nnd2s1 _____500126(.DIN1 (____9____35241), .DIN2 (________26723), .Q
       (____9____35268));
  hi1s1 _______500127(.DIN (____9____35266), .Q (____9____35267));
  nnd2s1 _______500128(.DIN1 (____99___35284), .DIN2 (____9____35264),
       .Q (____9____35265));
  nnd2s1 _______500129(.DIN1 (____9____35238), .DIN2 (_________34537),
       .Q (____99___35282));
  and2s1 ______500130(.DIN1 (____9____35263), .DIN2 (______9__34771),
       .Q (____0____35301));
  nor2s1 _______500131(.DIN1 (____9_0__35227), .DIN2 (____9_9__35226),
       .Q (____0_0__35306));
  nnd2s1 _______500132(.DIN1 (____9_9__35233), .DIN2 (________22522),
       .Q (____0____35304));
  dffacs1 _______________________________________________500133(.CLRB
       (reset), .CLK (clk), .DIN (____9_0__35234), .Q
       (_____________________________________________21822));
  dffacs1 ____________________________________________9_500134(.CLRB
       (reset), .CLK (clk), .DIN (____9____35230), .QN
       (___0_____40528));
  xor2s1 _______500135(.DIN1 (_______________22075), .DIN2
       (____9____35237), .Q (____9_0__35262));
  nor2s1 _____500136(.DIN1 (___0____22314), .DIN2 (____9____35260), .Q
       (____9_9__35261));
  and2s1 _____0_500137(.DIN1 (____9____35218), .DIN2 (____9____35258),
       .Q (____9____35259));
  nor2s1 _____0_500138(.DIN1 (______0__35537), .DIN2 (____9_0__35217),
       .Q (____9____35257));
  and2s1 _____0_500139(.DIN1 (____9_9__35216), .DIN2 (_________35394),
       .Q (____9____35256));
  nnd2s1 ______500140(.DIN1 (____9____35219), .DIN2 (____9____35254),
       .Q (____9____35255));
  nnd2s1 _____0_500141(.DIN1 (____9____35224), .DIN2 (_________35680),
       .Q (____9____35253));
  xor2s1 _______500142(.DIN1 (_____90__35191), .DIN2 (_________36292),
       .Q (____9_0__35252));
  nnd2s1 _______500143(.DIN1 (____9_0__35209), .DIN2 (_________35680),
       .Q (____9_9__35251));
  xor2s1 _______500144(.DIN1
       (_______________________________________________________________________________________),
       .DIN2 (____9____35232), .Q (____9____35250));
  nnd2s1 _______500145(.DIN1 (____9____35210), .DIN2 (_________35125),
       .Q (____0____35299));
  xnr2s1 ______500146(.DIN1 (______9__37429), .DIN2 (_____9___35197),
       .Q (____9____35266));
  dffacs1 _______________________________________________500147(.CLRB
       (reset), .CLK (clk), .DIN (____9____35222), .QN
       (_____________________________________________21795));
  dffacs1 _______________________________________________500148(.CLRB
       (reset), .CLK (clk), .DIN (____9____35223), .QN
       (___________________________________________));
  or2s1 _______500149(.DIN1 (____9_0__35243), .DIN2 (____9____35248),
       .Q (____9____35249));
  nnd2s1 _______500150(.DIN1 (____90___35207), .DIN2 (_____0___35741),
       .Q (____9____35247));
  xor2s1 _______500151(.DIN1 (____9____35245), .DIN2 (____0____36215),
       .Q (____9____35246));
  nor2s1 _______500152(.DIN1 (____00___35294), .DIN2 (____9_0__35243),
       .Q (____9____35244));
  nnd2s1 _______500153(.DIN1 (____90___35204), .DIN2 (inData[2]), .Q
       (____9_9__35242));
  nnd2s1 _______500154(.DIN1 (____909__35208), .DIN2 (________26695),
       .Q (____9____35241));
  nnd2s1 _____0_500155(.DIN1 (____90___35203), .DIN2 (______9__35170),
       .Q (____9____35240));
  xor2s1 _______500156(.DIN1 (_________35174), .DIN2 (_________35162),
       .Q (____9____35239));
  nnd2s1 ______500157(.DIN1 (____9____35237), .DIN2 (_________34540),
       .Q (____9____35238));
  nnd2s1 _______500158(.DIN1 (____90___35202), .DIN2 (____0____34425),
       .Q (____9____35274));
  xor2s1 _______500159(.DIN1
       (_____________________________________0_______21759), .DIN2
       (____9____35235), .Q (____9____35236));
  nnd2s1 _______500160(.DIN1 (____90___35206), .DIN2 (_____09__35023),
       .Q (____9_0__35234));
  nnd2s1 _______500161(.DIN1 (____9____35232), .DIN2 (__90), .Q
       (____9_9__35233));
  nnd2s1 ______500162(.DIN1 (_________35051), .DIN2 (____90___35205),
       .Q (____9____35230));
  nor2s1 ______500163(.DIN1 (____9_0__35227), .DIN2 (____9____35225),
       .Q (____9____35228));
  nor2s1 _____0_500164(.DIN1
       (__________________________________9__________), .DIN2
       (____9____35225), .Q (____9_9__35226));
  nnd2s1 _______500165(.DIN1 (_____9___35194), .DIN2 (_________34703),
       .Q (____9____35263));
  nor2s1 _______500166(.DIN1 (_________35057), .DIN2 (____90___35200),
       .Q (____9_0__35270));
  xor2s1 _______500167(.DIN1 (_________35172), .DIN2 (_________37320),
       .Q (____99___35284));
  xor2s1 ______500168(.DIN1 (____90___35201), .DIN2 (____0____34461),
       .Q (____9____35224));
  nnd2s1 _______500169(.DIN1 (______9__34676), .DIN2 (_________35185),
       .Q (____9____35223));
  nnd2s1 _____0_500170(.DIN1 (_________35187), .DIN2 (________28400),
       .Q (____9____35222));
  or2s1 _____0_500171(.DIN1 (___9_____39539), .DIN2 (____9____35220),
       .Q (____9____35221));
  nor2s1 _______500172(.DIN1 (________28429), .DIN2 (_________35175),
       .Q (____9____35219));
  xor2s1 _______500173(.DIN1 (_________35137), .DIN2 (_________35189),
       .Q (____9____35218));
  xor2s1 _______500174(.DIN1 (____9____34313), .DIN2 (_____99__35199),
       .Q (____9_0__35217));
  xor2s1 ______500175(.DIN1 (_________35089), .DIN2 (_________40866),
       .Q (____9_9__35216));
  nor2s1 _______500176(.DIN1 (______0__35132), .DIN2 (_________35184),
       .Q (____9____35260));
  nor2s1 _______500177(.DIN1 (____90___33342), .DIN2 (______9__35180),
       .Q (_________35580));
  xor2s1 _______500178(.DIN1 (____0____35309), .DIN2 (_____0__26457),
       .Q (____9____35215));
  nnd2s1 _______500179(.DIN1 (____9____35235), .DIN2
       (_____________________________________0_______21759), .Q
       (____9____35214));
  nor2s1 _______500180(.DIN1
       (_____________________________________0_______21759), .DIN2
       (____9____35235), .Q (____9____35213));
  xor2s1 _______500181(.DIN1 (____0____35309), .DIN2 (_________36512),
       .Q (____9____35211));
  xnr2s1 _____9_500182(.DIN1 (_____9___36360), .DIN2 (_________35156),
       .Q (____9____35210));
  xor2s1 _____9_500183(.DIN1 (_________34735), .DIN2 (_____9___35193),
       .Q (____9_0__35209));
  dffacs1 ______________________________________________500184(.CLRB
       (reset), .CLK (clk), .DIN (_________35188), .QN
       (____________________________________________21851));
  dffacs1 ____________________________________________9_500185(.CLRB
       (reset), .CLK (clk), .DIN (_________35173), .QN
       (_____9___22051));
  dffacs1 ______________________________________________500186(.CLRB
       (reset), .CLK (clk), .DIN (_________35182), .QN
       (___0__0__40501));
  nor2s1 _______500187(.DIN1 (_________35168), .DIN2 (____9____33367),
       .Q (____909__35208));
  xor2s1 _____500188(.DIN1 (______9__35150), .DIN2 (_________35183), .Q
       (____90___35207));
  nnd2s1 _______500189(.DIN1 (______9__35160), .DIN2 (_________35663),
       .Q (____90___35206));
  nnd2s1 _______500190(.DIN1 (_________35167), .DIN2 (______0__35050),
       .Q (____90___35205));
  nor2s1 _______500191(.DIN1 (_________35166), .DIN2 (_________33686),
       .Q (____90___35204));
  xor2s1 _______500192(.DIN1 (____9____33399), .DIN2 (_________35179),
       .Q (____90___35203));
  or2s1 _______500193(.DIN1 (____0____34433), .DIN2 (____90___35201),
       .Q (____90___35202));
  and2s1 ______500194(.DIN1 (_________40866), .DIN2 (_________35088),
       .Q (____90___35200));
  and2s1 _______500195(.DIN1 (_____9___35198), .DIN2
       (_____________________________________________21775), .Q
       (____9____35248));
  nnd2s1 _______500196(.DIN1 (_____99__35199), .DIN2 (______0__34249),
       .Q (____9____35229));
  nnd2s1 ______500197(.DIN1 (_________35165), .DIN2 (______9__35140),
       .Q (____9____35237));
  nor2s1 _______500198(.DIN1
       (_____________________________________________21775), .DIN2
       (_____9___35198), .Q (____9_0__35243));
  or2s1 _______500199(.DIN1 (___0_____40411), .DIN2 (_____9___35196),
       .Q (_____9___35197));
  and2s1 _______500200(.DIN1 (_____9___35196), .DIN2 (________27612),
       .Q (_____9___35195));
  or2s1 _____0_500201(.DIN1 (______0__34734), .DIN2 (_____9___35193),
       .Q (_____9___35194));
  nor2s1 _______500202(.DIN1 (_________41367), .DIN2 (_____9___35196),
       .Q (_____9___35192));
  xor2s1 _____9_500203(.DIN1 (___0_9___40559), .DIN2 (_________35169),
       .Q (_____90__35191));
  and2s1 ______500204(.DIN1 (_____9___35196), .DIN2 (___0_____40411),
       .Q (____999__35288));
  and2s1 ______500205(.DIN1 (______9__35190), .DIN2 (_________35844),
       .Q (____9____35225));
  nor2s1 _______500206(.DIN1 (_________35844), .DIN2 (______9__35190),
       .Q (____9_0__35227));
  xor2s1 _____0_500207(.DIN1 (______0__35141), .DIN2 (______9__37429),
       .Q (____9____35232));
  nor2s1 _____9_500208(.DIN1 (_________35136), .DIN2 (_________35189),
       .Q (____9____35231));
  dffacs1 _______________________________________________500209(.CLRB
       (reset), .CLK (clk), .DIN (_________35159), .QN
       (______0___22054));
  nnd2s1 ______500210(.DIN1 (_________35153), .DIN2 (_________34834),
       .Q (_________35188));
  nnd2s1 _______500211(.DIN1 (______0__35151), .DIN2 (_________35186),
       .Q (_________35187));
  nnd2s1 _______500212(.DIN1 (_________35154), .DIN2 (inData[10]), .Q
       (_________35185));
  nor2s1 _______500213(.DIN1 (_________35146), .DIN2 (_________35183),
       .Q (_________35184));
  nnd2s1 _______500214(.DIN1 (_________35149), .DIN2 (______0__35181),
       .Q (_________35182));
  nor2s1 _______500215(.DIN1 (____90___33341), .DIN2 (_________35179),
       .Q (______9__35180));
  xor2s1 _______500216(.DIN1
       (_____________________________________________21810), .DIN2
       (_____00__35653), .Q (____9____35220));
  xor2s1 ______500217(.DIN1 (___0_____40542), .DIN2 (_____00__35653),
       .Q (____9____35245));
  nnd2s1 ______500218(.DIN1 (_________35177), .DIN2 (_________35176),
       .Q (_________35178));
  nor2s1 _______500219(.DIN1 (______0__35537), .DIN2 (_________35144),
       .Q (_________35175));
  xor2s1 _____9_500220(.DIN1
       (_____________________________________________21776), .DIN2
       (_________38271), .Q (_________35174));
  nnd2s1 _______500221(.DIN1 (_________35148), .DIN2 (____0____35361),
       .Q (_________35173));
  and2s1 _______500222(.DIN1 (_________35139), .DIN2 (_________35164),
       .Q (_________35172));
  nnd2s1 _______500223(.DIN1 (_________35143), .DIN2 (______9__35170),
       .Q (______0__35171));
  or2s1 _______500224(.DIN1 (______9__34171), .DIN2 (_________35169),
       .Q (____9____35212));
  dffacs1 _______________________________________________500225(.CLRB
       (reset), .CLK (clk), .DIN (_________35152), .Q
       (_____________________________________________21765));
  xor2s1 _______500226(.DIN1 (_________35126), .DIN2 (_________35155),
       .Q (____9____35235));
  and2s1 _____0_500227(.DIN1 (_____0__29534), .DIN2
       (_____________________________________________21776), .Q
       (_________35168));
  nnd2s1 _____500228(.DIN1 (___0____24201), .DIN2 (_________35123), .Q
       (_________35167));
  xor2s1 _____9_500229(.DIN1 (_________35145), .DIN2
       (____________________________________________21867), .Q
       (_________35166));
  nnd2s1 _____500230(.DIN1 (_________35164), .DIN2 (_________37320), .Q
       (_________35165));
  nor2s1 ______500231(.DIN1
       (_____________________________________________21776), .DIN2
       (_________35162), .Q (_________35163));
  nnd2s1 _______500232(.DIN1 (_________35134), .DIN2 (____9____33368),
       .Q (_____9___35198));
  nnd2s1 _______500233(.DIN1 (_________35128), .DIN2 (_________34114),
       .Q (_____99__35199));
  nor2s1 _______500234(.DIN1 (_________33024), .DIN2 (______9__35131),
       .Q (_________35189));
  xor2s1 ______500235(.DIN1 (_________35114), .DIN2 (___9_0___39170),
       .Q (____90___35201));
  and2s1 _______500236(.DIN1 (_________35162), .DIN2
       (_____________________________________________21776), .Q
       (______0__35161));
  xor2s1 _______500237(.DIN1 (____0_9__34459), .DIN2 (_____0___35109),
       .Q (______9__35160));
  nnd2s1 _______500238(.DIN1 (_________35124), .DIN2 (_____9___35467),
       .Q (_________35159));
  xor2s1 _____9_500239(.DIN1 (_____9__27676), .DIN2 (_________35157),
       .Q (_________35158));
  nor2s1 _______500240(.DIN1 (_________35085), .DIN2 (_________35155),
       .Q (_________35156));
  xor2s1 _____9_500241(.DIN1 (_____9___35098), .DIN2 (_____9___41303),
       .Q (______9__35190));
  nnd2s1 _______500242(.DIN1 (______0__35122), .DIN2 (_________35091),
       .Q (_____9___35193));
  dffacs1 _______________________________________________500243(.CLRB
       (reset), .CLK (clk), .DIN (_________35129), .Q (___0_____40544));
  xor2s1 _______500244(.DIN1 (_____9___35101), .DIN2 (_________36349),
       .Q (____0____35309));
  xor2s1 _______500245(.DIN1 (_____0___35106), .DIN2
       (_______________22074), .Q (_____9___35196));
  nor2s1 ______500246(.DIN1 (_________35116), .DIN2 (________28399), .Q
       (_________35154));
  nnd2s1 _______500247(.DIN1 (_________35117), .DIN2 (_____0___34932),
       .Q (_________35153));
  and2s1 _______500248(.DIN1 (_________35115), .DIN2 (_____9___35467),
       .Q (_________35152));
  xor2s1 _____9_500249(.DIN1 (____9____33361), .DIN2 (_________35133),
       .Q (______0__35151));
  xor2s1 _____9_500250(.DIN1 (_______________22069), .DIN2
       (____________________________________________21868), .Q
       (______9__35150));
  nor2s1 _____500251(.DIN1 (________24971), .DIN2 (_____0___35110), .Q
       (_________35149));
  and2s1 _____0_500252(.DIN1 (_____09__35112), .DIN2 (_________35147),
       .Q (_________35148));
  nor2s1 _____0_500253(.DIN1 (_________35145), .DIN2
       (_______________22069), .Q (_________35146));
  xor2s1 _______500254(.DIN1 (_________34149), .DIN2 (_________35127),
       .Q (_________35144));
  xor2s1 _______500255(.DIN1 (_____0___33070), .DIN2 (_________35130),
       .Q (_________35143));
  nnd2s1 _____0_500256(.DIN1 (_________35157), .DIN2
       (_____________________________________________21826), .Q
       (_________35142));
  nnd2s1 _______500257(.DIN1 (_____9___35100), .DIN2 (_____0___35105),
       .Q (______0__35141));
  nnd2s1 _______500258(.DIN1 (_________35138), .DIN2 (_________34548),
       .Q (______9__35140));
  nnd2s1 _______500259(.DIN1 (_________35138), .DIN2 (______9__34543),
       .Q (_________35139));
  nor2s1 ______500260(.DIN1 (_________35120), .DIN2 (_________35136),
       .Q (_________35137));
  nor2s1 _______500261(.DIN1
       (_____________________________________________21826), .DIN2
       (_________35157), .Q (_________35135));
  xor2s1 _______500262(.DIN1 (_________35094), .DIN2 (_________38650),
       .Q (_________35179));
  nnd2s1 _______500263(.DIN1 (_________35157), .DIN2 (___0_____40497),
       .Q (_________35177));
  or2s1 _______500264(.DIN1 (___0_____40497), .DIN2 (_________35157),
       .Q (_________35176));
  nor2s1 _______500265(.DIN1 (_____90__33994), .DIN2 (_____0___35108),
       .Q (_________35169));
  dffacs1 ______________________________________________500266(.CLRB
       (reset), .CLK (clk), .DIN (_____0___35111), .QN
       (___0_____40478));
  or2s1 _____0_500267(.DIN1 (____9____33369), .DIN2 (_________35133),
       .Q (_________35134));
  nor2s1 _____0_500268(.DIN1
       (____________________________________________21868), .DIN2
       (_________33973), .Q (______0__35132));
  nor2s1 _______500269(.DIN1 (_________33039), .DIN2 (_________35130),
       .Q (______9__35131));
  nnd2s1 _____500270(.DIN1 (_____90__35096), .DIN2 (______0__34855), .Q
       (_________35129));
  or2s1 ______500271(.DIN1 (_________35127), .DIN2 (_________34113), .Q
       (_________35128));
  dffacs1 _______________________________________________500272(.CLRB
       (reset), .CLK (clk), .DIN (______9__35095), .Q
       (_____________________________________________21776));
  xnr2s1 _______500273(.DIN1
       (_______________________________________________________________________________________),
       .DIN2 (______0__35077), .Q (_____00__35653));
  nnd2s1 _______500274(.DIN1 (______9__35086), .DIN2 (_________35125),
       .Q (_________35126));
  xor2s1 _______500275(.DIN1 (_____0___35107), .DIN2 (_____9___33995),
       .Q (_________35124));
  xor2s1 ______500276(.DIN1
       (_________________________________________0___21821), .DIN2
       (________23052), .Q (_________35123));
  nnd2s1 _______500277(.DIN1 (_________35092), .DIN2 (____0_0__34460),
       .Q (______0__35122));
  nor2s1 _____500278(.DIN1
       (_____________________________________________21783), .DIN2
       (____9_0__37043), .Q (______9__35121));
  and2s1 _____0_500279(.DIN1 (____9_0__37043), .DIN2
       (_____________________________________________21783), .Q
       (_________35119));
  nor2s1 _______500280(.DIN1 (_________35005), .DIN2 (_________35090),
       .Q (_________35155));
  nnd2s1 _______500281(.DIN1 (_________40868), .DIN2 (_________34558),
       .Q (_________35164));
  nnd2s1 _____0_500282(.DIN1 (_________35083), .DIN2 (_________35663),
       .Q (_________35118));
  xor2s1 _______500283(.DIN1 (______0__35067), .DIN2 (_________38372),
       .Q (_________35117));
  xor2s1 _______500284(.DIN1 (___0___22204), .DIN2 (___09_9__40680), .Q
       (_________35116));
  xor2s1 _______500285(.DIN1 (_________35064), .DIN2 (_____9___37654),
       .Q (_________35115));
  nor2s1 ______500286(.DIN1 (______9__35049), .DIN2 (_________35082),
       .Q (_________35114));
  nnd2s1 _______500287(.DIN1 (______9__35076), .DIN2 (________25004),
       .Q (______0__35113));
  and2s1 _______500288(.DIN1 (______9__34714), .DIN2 (_________35081),
       .Q (_____09__35112));
  nnd2s1 _______500289(.DIN1 (_________35079), .DIN2 (____9____35254),
       .Q (_____0___35111));
  nor2s1 _______500290(.DIN1 (_____0___35834), .DIN2 (_________35075),
       .Q (_____0___35110));
  hi1s1 _______500291(.DIN
       (____________________________________________21868), .Q
       (_________35145));
  xnr2s1 _____500292(.DIN1 (___9_____39231), .DIN2 (_________41355), .Q
       (_____0___35109));
  and2s1 _______500293(.DIN1 (_____0___35107), .DIN2 (_________33943),
       .Q (_____0___35108));
  and2s1 _____9_500294(.DIN1 (_____0___35105), .DIN2 (_____9___35099),
       .Q (_____0___35106));
  or2s1 ______500295(.DIN1 (_____00__35103), .DIN2 (_____99__35102), .Q
       (_____0___35104));
  xor2s1 _____500296(.DIN1 (_________35053), .DIN2 (_________35055), .Q
       (_____9___35101));
  nnd2s1 _______500297(.DIN1 (_____9___35099), .DIN2 (_________37320),
       .Q (_____9___35100));
  nor2s1 _______500298(.DIN1 (_____9__28228), .DIN2 (_________35069),
       .Q (_____9___35098));
  and2s1 _____9_500299(.DIN1 (_________40656), .DIN2
       (_________________________________________0___21821), .Q
       (_________35136));
  hi1s1 _______500300(.DIN (_________40868), .Q (_________35138));
  nor2s1 _____9_500301(.DIN1
       (_________________________________________0___21821), .DIN2
       (_________40656), .Q (_________35120));
  hi1s1 _______500302(.DIN (____9_0__37043), .Q (_________35157));
  xor2s1 ______500303(.DIN1 (_________35046), .DIN2 (_________35065),
       .Q (_____90__35096));
  and2s1 _______500304(.DIN1 (_________35054), .DIN2 (_____9___35467),
       .Q (______9__35095));
  nnd2s1 _______500305(.DIN1 (_________35061), .DIN2 (_________33184),
       .Q (_________35094));
  xnr2s1 _____0_500306(.DIN1 (_________36087), .DIN2 (_________40870),
       .Q (_________35127));
  nor2s1 _______500307(.DIN1 (_________35030), .DIN2 (______9__35066),
       .Q (_________35133));
  dffacs1 ______________________________________________500308(.CLRB
       (reset), .CLK (clk), .DIN (_________35062), .Q
       (____________________________________________21868));
  xor2s1 ____500309(.DIN1
       (_____________________________________________21768), .DIN2
       (_________37792), .Q (_________35093));
  nnd2s1 _____0_500310(.DIN1 (_________41355), .DIN2 (___0_____40526),
       .Q (_________35092));
  or2s1 _____0_500311(.DIN1 (___0_____40526), .DIN2 (_________41355),
       .Q (_________35091));
  nnd2s1 ______500312(.DIN1 (_________35056), .DIN2 (_____9___35009),
       .Q (_________35090));
  nnd2s1 _______500313(.DIN1 (_________35088), .DIN2 (_________35058),
       .Q (_________35089));
  xor2s1 _____9_500314(.DIN1 (________23677), .DIN2 (_________37792),
       .Q (______0__35087));
  hi1s1 _______500315(.DIN (_________35085), .Q (______9__35086));
  xor2s1 _____0_500316(.DIN1 (_________35035), .DIN2 (_________35084),
       .Q (_________35130));
  xor2s1 ______500317(.DIN1 (____09__28561), .DIN2 (_________35068), .Q
       (____9_0__37043));
  xor2s1 _______500318(.DIN1 (_________35048), .DIN2 (_________35027),
       .Q (_________35083));
  nor2s1 _______500319(.DIN1 (_________35026), .DIN2 (_________35047),
       .Q (_________35082));
  nnd2s1 _______500320(.DIN1 (______9__35039), .DIN2 (_________35043),
       .Q (_________35081));
  or2s1 ______500321(.DIN1 (_____00__33066), .DIN2 (_________35147), .Q
       (_________35080));
  nor2s1 _______500322(.DIN1 (____9___28639), .DIN2 (______0__35040),
       .Q (_________35079));
  nor2s1 _______500323(.DIN1 (_________35045), .DIN2 (_________35680),
       .Q (_________35078));
  nor2s1 _______500324(.DIN1 (_________35031), .DIN2 (______0__35059),
       .Q (______0__35077));
  xor2s1 _______500325(.DIN1 (_________33226), .DIN2 (_________35060),
       .Q (______9__35076));
  xor2s1 ______500326(.DIN1 (_________32958), .DIN2 (_____0___35020),
       .Q (_________35075));
  nnd2s1 _______500327(.DIN1 (_________35033), .DIN2 (_________33777),
       .Q (_____0___35107));
  or2s1 ____90_500328(.DIN1
       (_____________________________________________21768), .DIN2
       (_________37792), .Q (_________35074));
  nnd2s1 ____90_500329(.DIN1 (_________37792), .DIN2
       (_____________________________________________21768), .Q
       (_________35073));
  and2s1 ____90_500330(.DIN1 (_________35070), .DIN2 (___0__9__40550),
       .Q (_________35072));
  nor2s1 ____500331(.DIN1 (___0__9__40550), .DIN2 (_________35070), .Q
       (_________35071));
  and2s1 _____9_500332(.DIN1 (_________35068), .DIN2 (_____0__28229),
       .Q (_________35069));
  xor2s1 _____9_500333(.DIN1 (_____0___35022), .DIN2 (_________41264),
       .Q (_________35085));
  and2s1 ____9__500334(.DIN1 (_________35070), .DIN2
       (_____________________________________________21843), .Q
       (_____00__35103));
  nor2s1 ____9__500335(.DIN1
       (_____________________________________________21843), .DIN2
       (_________35070), .Q (_____99__35102));
  nnd2s1 ____9_500336(.DIN1 (_________35037), .DIN2 (_________37321),
       .Q (_____9___35099));
  dffacs1 _____________________________________________0_500337(.CLRB
       (reset), .CLK (clk), .DIN (_________35034), .QN
       (_________________________________________0___21821));
  xor2s1 _____9_500338(.DIN1 (_____0___35019), .DIN2 (_________33006),
       .Q (______0__35067));
  and2s1 _______500339(.DIN1 (_________35065), .DIN2 (_________35029),
       .Q (______9__35066));
  xor2s1 _____9_500340(.DIN1 (_________35063), .DIN2 (_____00__35016),
       .Q (_________35064));
  nnd2s1 _______500341(.DIN1 (_________35028), .DIN2 (___9____29603),
       .Q (_________35062));
  or2s1 _______500342(.DIN1 (_________33225), .DIN2 (_________35060),
       .Q (_________35061));
  nnd2s1 _______500343(.DIN1 (_________35025), .DIN2 (_____99__35015),
       .Q (_____9___35097));
  hi1s1 _______500344(.DIN (_________35057), .Q (_________35058));
  nnd2s1 _______500345(.DIN1 (_________35055), .DIN2 (______0__34975),
       .Q (_________35056));
  xor2s1 _______500346(.DIN1 (______0__33833), .DIN2 (_________41357),
       .Q (_________35054));
  nnd2s1 _______500347(.DIN1 (_____9___35012), .DIN2 (_____0___35021),
       .Q (_________35053));
  xor2s1 _______500348(.DIN1 (________25915), .DIN2 (_________35041),
       .Q (_________35052));
  nnd2s1 ____9__500349(.DIN1 (_________35036), .DIN2
       (_______________22073), .Q (_____0___35105));
  or2s1 _______500350(.DIN1 (______0__35050), .DIN2 (_____0___35018),
       .Q (_________35051));
  nor2s1 _______500351(.DIN1
       (_________________________________________0___21794), .DIN2
       (_________35048), .Q (______9__35049));
  and2s1 _______500352(.DIN1 (_________35048), .DIN2
       (_________________________________________0___21794), .Q
       (_________35047));
  xor2s1 _____9_500353(.DIN1 (______0__33312), .DIN2 (_____99__22053),
       .Q (_________35046));
  or2s1 _____0_500354(.DIN1 (_____9___22051), .DIN2 (_________35044),
       .Q (_________35045));
  nnd2s1 _______500355(.DIN1 (_____0___35017), .DIN2 (inData[6]), .Q
       (_________35043));
  nor2s1 _______500356(.DIN1 (_________36852), .DIN2 (_________35041),
       .Q (_________35042));
  nor2s1 _______500357(.DIN1 (______0__35537), .DIN2 (_____9___35014),
       .Q (______0__35040));
  xor2s1 ______500358(.DIN1 (_________35002), .DIN2 (_________38680),
       .Q (______0__35059));
  nnd2s1 _______500359(.DIN1 (______9__35039), .DIN2 (_________35044),
       .Q (_________35147));
  nnd2s1 _______500360(.DIN1 (_________35041), .DIN2 (_________36852),
       .Q (_________35038));
  hi1s1 ____9_500361(.DIN (_________35036), .Q (_________35037));
  nor2s1 _______500362(.DIN1 (_____0___32879), .DIN2 (_____9___35011),
       .Q (_________35035));
  nnd2s1 _______500363(.DIN1 (_____9___35010), .DIN2 (____0___23693),
       .Q (_________35034));
  nnd2s1 _______500364(.DIN1 (_________41357), .DIN2 (______0__33775),
       .Q (_________35033));
  xor2s1 ____9__500365(.DIN1 (_________34986), .DIN2 (____90___36104),
       .Q (_________35068));
  nnd2s1 _______500366(.DIN1 (_________35041), .DIN2 (___0_____40574),
       .Q (_________35088));
  nor2s1 _______500367(.DIN1 (___0_____40574), .DIN2 (_________35041),
       .Q (_________35057));
  hi1s1 ____9__500368(.DIN (______0__35032), .Q (_________35070));
  nb1s1 ____9__500369(.DIN (______0__35032), .Q (_________37792));
  nor2s1 ______500370(.DIN1 (_____99__22053), .DIN2 (______0__33312),
       .Q (_________35030));
  nnd2s1 _______500371(.DIN1 (______0__33312), .DIN2 (_____99__22053),
       .Q (_________35029));
  nnd2s1 _______500372(.DIN1 (_________35001), .DIN2 (_________34877),
       .Q (_________35028));
  xnr2s1 ______500373(.DIN1
       (_________________________________________0___21794), .DIN2
       (_________35026), .Q (_________35027));
  nnd2s1 _______500374(.DIN1 (_________35063), .DIN2 (___0_____40575),
       .Q (_________35025));
  nor2s1 ______500375(.DIN1 (___0_____40575), .DIN2 (_________35063),
       .Q (______0__35024));
  nnd2s1 ______500376(.DIN1 (________25700), .DIN2 (______0__34998), .Q
       (_____09__35023));
  nor2s1 ______500377(.DIN1 (______9__33045), .DIN2 (_________34993),
       .Q (_________35060));
  nor2s1 ____9__500378(.DIN1 (_________36762), .DIN2 (_____9___35731),
       .Q (_____0___35022));
  nnd2s1 _____9_500379(.DIN1 (_________34988), .DIN2 (______0__36598),
       .Q (_____0___35021));
  xnr2s1 _______500380(.DIN1 (_________36512), .DIN2 (_________40872),
       .Q (_____0___35020));
  nnd2s1 ____9__500381(.DIN1 (_____9___35731), .DIN2 (_________36762),
       .Q (_________35125));
  xnr2s1 ____9__500382(.DIN1 (_________38385), .DIN2 (_________34977),
       .Q (_________35036));
  xor2s1 ____9_500383(.DIN1 (______9__34974), .DIN2 (_________37867),
       .Q (______0__35032));
  nnd2s1 _______500384(.DIN1 (_________34990), .DIN2 (_________34826),
       .Q (_________35055));
  dffacs1 ______________________________________________500385(.CLRB
       (reset), .CLK (clk), .DIN (_________35000), .QN
       (____________________________________________21850));
  xor2s1 _______500386(.DIN1 (___0__0__40501), .DIN2 (_________34992),
       .Q (_____0___35019));
  xor2s1 _____500387(.DIN1 (_________34968), .DIN2 (______0__40884), .Q
       (_____0___35018));
  or2s1 _______500388(.DIN1
       (_________________________________________0___21794), .DIN2
       (___0_____40526), .Q (_____0___35017));
  xnr2s1 _______500389(.DIN1 (___0_____40575), .DIN2 (_____99__35015),
       .Q (_____00__35016));
  xor2s1 _______500390(.DIN1 (______9__33794), .DIN2 (_________34966),
       .Q (_____9___35014));
  or2s1 _______500391(.DIN1 (_________35448), .DIN2 (_________34980),
       .Q (_____9___35013));
  and2s1 _______500392(.DIN1 (___0_____40526), .DIN2
       (_________________________________________0___21794), .Q
       (_________35044));
  nnd2s1 _______500393(.DIN1 (_________34978), .DIN2 (_________34961),
       .Q (_________35048));
  nnd2s1 ____9__500394(.DIN1 (_____90__35008), .DIN2 (_________33924),
       .Q (_____9___35012));
  nor2s1 _______500395(.DIN1 (_____0___32880), .DIN2 (_________40872),
       .Q (_____9___35011));
  or2s1 _____500396(.DIN1 (______0__35050), .DIN2 (_________34976), .Q
       (_____9___35010));
  nnd2s1 ____9__500397(.DIN1 (_____90__35008), .DIN2 (______0__36598),
       .Q (_____9___35009));
  nnd2s1 ____9__500398(.DIN1 (_________34984), .DIN2 (_________35006),
       .Q (______9__35007));
  nor2s1 ____9__500399(.DIN1 (______0__36598), .DIN2 (_____90__35008),
       .Q (_________35005));
  xor2s1 ____90_500400(.DIN1 (_____9___34842), .DIN2 (_________40874),
       .Q (_________35041));
  xor2s1 _______500401(.DIN1 (___0_____40524), .DIN2 (_________35003),
       .Q (_________35004));
  nnd2s1 _____9_500402(.DIN1 (______0__34982), .DIN2 (_________34983),
       .Q (_________35002));
  xor2s1 _______500403(.DIN1 (_________34957), .DIN2 (____0_0__38064),
       .Q (_________35001));
  nnd2s1 ______500404(.DIN1 (_________34971), .DIN2 (_____0__23862), .Q
       (_________35000));
  or2s1 ______500405(.DIN1 (_________35448), .DIN2 (_________34969), .Q
       (_________34999));
  xor2s1 ______500406(.DIN1 (_____9___22049), .DIN2 (______9__34997),
       .Q (______0__34998));
  and2s1 ______500407(.DIN1 (_________34995), .DIN2 (___0_____40524),
       .Q (_________34996));
  nor2s1 _______500408(.DIN1 (___0_____40524), .DIN2 (_________34995),
       .Q (_________34994));
  nor2s1 _______500409(.DIN1 (_________33040), .DIN2 (_________34992),
       .Q (_________34993));
  hi1s1 _______500410(.DIN (____99___36176), .Q (_________35063));
  dffacs1 _______________________________________________500411(.CLRB
       (reset), .CLK (clk), .DIN (_________34970), .Q (_____99__22053));
  xor2s1 ____9__500412(.DIN1 (________27450), .DIN2 (_________36680),
       .Q (_________34991));
  nnd2s1 ____90_500413(.DIN1 (_________40874), .DIN2 (______9__34827),
       .Q (_________34990));
  xor2s1 ____9__500414(.DIN1 (_________35598), .DIN2 (_________36761),
       .Q (_________34988));
  xor2s1 ____9__500415(.DIN1 (________25531), .DIN2 (_________36680),
       .Q (_________34987));
  nnd2s1 ____9__500416(.DIN1 (______0__34965), .DIN2 (_________34973),
       .Q (_________34986));
  hi1s1 ____9__500417(.DIN (_________34984), .Q (_________34985));
  nor2s1 _____500418(.DIN1 (_________34983), .DIN2 (______0__34982), .Q
       (_________35031));
  xor2s1 ___900_(.DIN1 (_________34953), .DIN2 (______9__34981), .Q
       (_____9___35731));
  dffacs1 ______________________________________________500419(.CLRB
       (reset), .CLK (clk), .DIN (_________34972), .QN
       (___0_____40502));
  dffacs1 ____0___________________(.CLRB (reset), .CLK (clk), .DIN
       (_________34963), .QN (____0_________________21725));
  xor2s1 _______500420(.DIN1 (_____99__34930), .DIN2 (_____9___33711),
       .Q (_________34980));
  nnd2s1 ______500421(.DIN1 (_________34967), .DIN2 (_________34960),
       .Q (_________34978));
  xor2s1 ____90_500422(.DIN1 (_____9___34929), .DIN2 (_________38675),
       .Q (____99___36176));
  dffacs1 _____________________________________________0_500423(.CLRB
       (reset), .CLK (clk), .DIN (_________34958), .Q
       (_________________________________________0___21794));
  nnd2s1 ___90__(.DIN1 (_________34951), .DIN2 (_________34952), .Q
       (_________34977));
  xor2s1 ____9__500424(.DIN1 (_________34962), .DIN2 (_________34255),
       .Q (_________34976));
  nnd2s1 ____9__500425(.DIN1 (_________35598), .DIN2 (_________36761),
       .Q (______0__34975));
  and2s1 ___90_0(.DIN1 (______9__34964), .DIN2 (_________34973), .Q
       (______9__34974));
  or2s1 ____9__500426(.DIN1 (_________22044), .DIN2 (_________36680),
       .Q (_________35006));
  nnd2s1 ____9__500427(.DIN1 (_________36680), .DIN2 (_________22044),
       .Q (_________34984));
  nor2s1 ____9__500428(.DIN1 (_________36761), .DIN2 (_________35598),
       .Q (_____90__35008));
  dffacs1 ______________________________________________500429(.CLRB
       (reset), .CLK (clk), .DIN (_________34959), .QN
       (___0_____40503));
  nnd2s1 ____9__500430(.DIN1 (_____0___34933), .DIN2 (________25896),
       .Q (_________34972));
  nnd2s1 _______500431(.DIN1 (_____09__34939), .DIN2 (_________34916),
       .Q (_________34971));
  nnd2s1 ______500432(.DIN1 (______0__34940), .DIN2 (__9__9__30158), .Q
       (_________34970));
  xor2s1 _____9_500433(.DIN1 (_____90__34922), .DIN2 (_____0___34934),
       .Q (_________34969));
  xor2s1 _______500434(.DIN1 (___0_____40545), .DIN2 (_________34967),
       .Q (_________34968));
  nnd2s1 ____9__500435(.DIN1 (_____0___34937), .DIN2 (_________34036),
       .Q (______0__34982));
  hi1s1 ____9__500436(.DIN (_________35003), .Q (_________34995));
  xor2s1 ____9__500437(.DIN1 (_________34945), .DIN2 (_____9___41303),
       .Q (_________34966));
  nnd2s1 ___90__500438(.DIN1 (______9__34964), .DIN2 (_________37867),
       .Q (______0__34965));
  nnd2s1 ___90__500439(.DIN1 (_____9___34927), .DIN2 (___0_____31239),
       .Q (_________34963));
  nnd2s1 ____9__500440(.DIN1 (_________34962), .DIN2 (_________34233),
       .Q (_________34989));
  nnd2s1 ____9__500441(.DIN1 (_____0___34935), .DIN2 (_________34910),
       .Q (_____99__35015));
  xor2s1 ____9__500442(.DIN1 (______0__41359), .DIN2 (___9_9___39790),
       .Q (_________34992));
  dffacs1 _______________________________________________500443(.CLRB
       (reset), .CLK (clk), .DIN (_____00__34931), .QN
       (___0_9___40552));
  or2s1 _______500444(.DIN1 (___0_____40545), .DIN2 (______0__40884),
       .Q (_________34961));
  nnd2s1 _______500445(.DIN1 (______0__40884), .DIN2 (___0_____40545),
       .Q (_________34960));
  nnd2s1 ____9_500446(.DIN1 (_________34917), .DIN2 (_____0__25806), .Q
       (_________34959));
  nnd2s1 ____90_500447(.DIN1 (_________34920), .DIN2 (_____00__41309),
       .Q (_________34958));
  xor2s1 ____9__500448(.DIN1 (______0__34905), .DIN2 (_________33683),
       .Q (_________34957));
  xor2s1 ____9_500449(.DIN1 (_________34906), .DIN2 (_________41343),
       .Q (_________35065));
  nor2s1 _______500450(.DIN1 (___9__22143), .DIN2 (___0_____40545), .Q
       (______9__34997));
  xor2s1 ____9__500451(.DIN1 (_________40876), .DIN2 (_________34062),
       .Q (_________35003));
  xnr2s1 ___90__500452(.DIN1 (___0_____40506), .DIN2 (_________34954),
       .Q (_________34955));
  nnd2s1 ___90_9(.DIN1 (_________34950), .DIN2 (_________34952), .Q
       (_________34953));
  nnd2s1 ___90__500453(.DIN1 (_________34950), .DIN2 (______9__34981),
       .Q (_________34951));
  xor2s1 ___90__500454(.DIN1 (________24571), .DIN2 (_________34954),
       .Q (______0__34949));
  or2s1 ___90_500455(.DIN1 (_________34947), .DIN2 (_________34946), .Q
       (______9__34948));
  nnd2s1 ___90__500456(.DIN1 (______9__34914), .DIN2
       (_______________22075), .Q (_________34973));
  and2s1 ____9__500457(.DIN1 (_________33789), .DIN2 (_________34945),
       .Q (_________34979));
  xor2s1 ___9009(.DIN1 (______9__34896), .DIN2 (_____0__25892), .Q
       (_________35598));
  dffacs1 ______________________________________________500458(.CLRB
       (reset), .CLK (clk), .DIN (_________34921), .QN
       (___0__0__40491));
  xnr2s1 ___90_500459(.DIN1 (_________36087), .DIN2 (_________34898),
       .Q (_________36680));
  and2s1 ____9__500460(.DIN1 (_________34943), .DIN2 (_________34942),
       .Q (_________34944));
  nor2s1 ____9__500461(.DIN1 (___0_____40525), .DIN2 (_________34902),
       .Q (_________34941));
  nnd2s1 ____9_500462(.DIN1 (_________34908), .DIN2 (_________35186),
       .Q (______0__34940));
  xor2s1 ____9__500463(.DIN1 (_________34893), .DIN2 (_____0___34938),
       .Q (_____09__34939));
  nnd2s1 ____9__500464(.DIN1 (_________40876), .DIN2 (_________34018),
       .Q (_____0___34937));
  xor2s1 _____9_500465(.DIN1 (____90__23778), .DIN2 (______9__35627),
       .Q (_____0___34936));
  nnd2s1 ____9__500466(.DIN1 (______9__34904), .DIN2 (_____0___34934),
       .Q (_____0___34935));
  nnd2s1 ____9__500467(.DIN1 (_________34900), .DIN2 (_____0___34932),
       .Q (_____0___34933));
  nnd2s1 ____9_500468(.DIN1 (_________34903), .DIN2 (___9____25986), .Q
       (_____00__34931));
  xor2s1 ____9__500469(.DIN1 (_________34911), .DIN2 (___90____39008),
       .Q (_____99__34930));
  xor2s1 ____9__500470(.DIN1 (_________34884), .DIN2 (_________36402),
       .Q (_____9___34929));
  nor2s1 ___90__500471(.DIN1 (______22148), .DIN2 (_________34954), .Q
       (_____9___34928));
  nor2s1 ___9_0_(.DIN1 (___0_0___30837), .DIN2 (_________34895), .Q
       (_____9___34927));
  and2s1 ___90_500472(.DIN1 (_________34954), .DIN2
       (_____________________________________________21782), .Q
       (_____9___34926));
  nor2s1 ___90__500473(.DIN1 (___0_9___40556), .DIN2 (_________34954),
       .Q (_____9___34925));
  and2s1 ___90__500474(.DIN1 (_________34954), .DIN2 (___0_9___40556),
       .Q (_____9___34924));
  nor2s1 ___90_500475(.DIN1
       (_____________________________________________21782), .DIN2
       (_________34954), .Q (_____9___34923));
  xnr2s1 ___900_500476(.DIN1 (___9_____39784), .DIN2 (_________40878),
       .Q (_________34962));
  nnd2s1 ___90__500477(.DIN1 (_________34913), .DIN2 (_________37412),
       .Q (______9__34964));
  dffacs1 ____________________________________________9_500478(.CLRB
       (reset), .CLK (clk), .DIN (_________34894), .QN
       (___0__0__40511));
  dffacs1 ______________________________________________500479(.CLRB
       (reset), .CLK (clk), .DIN (_________34901), .Q
       (____________________________________________21867));
  xor2s1 ____9__500480(.DIN1 (________26620), .DIN2 (_________34909),
       .Q (_____90__34922));
  nnd2s1 ____9__500481(.DIN1 (_________34892), .DIN2 (_________37722),
       .Q (_________34921));
  nnd2s1 ____9_500482(.DIN1 (_________34891), .DIN2 (_________35680),
       .Q (_________34920));
  nor2s1 ____9__500483(.DIN1 (____9___24637), .DIN2 (______9__35627),
       .Q (_________34919));
  dffacs1 ____________________________________________9_500484(.CLRB
       (reset), .CLK (clk), .DIN (_________34890), .Q (___0_____40545));
  nnd2s1 ____99_500485(.DIN1 (_________34881), .DIN2 (_________34916),
       .Q (_________34917));
  nor2s1 ___90__500486(.DIN1 (___0_____40506), .DIN2 (_________34912),
       .Q (______0__34915));
  hi1s1 ___9090(.DIN (_________34913), .Q (______9__34914));
  and2s1 ___90_500487(.DIN1 (_________34912), .DIN2 (______0___22056),
       .Q (_________34946));
  nnd2s1 ____9_500488(.DIN1 (_________34889), .DIN2 (_________33655),
       .Q (_________34945));
  nnd2s1 ___90__500489(.DIN1 (_________34886), .DIN2 (________27043),
       .Q (_________34950));
  nor2s1 ___90__500490(.DIN1 (______0___22056), .DIN2 (_________34912),
       .Q (_________34947));
  or2s1 ____9__500491(.DIN1 (_________34911), .DIN2 (_________33673),
       .Q (_________34956));
  dffacs1 ____0__________________(.CLRB (reset), .CLK (clk), .DIN
       (_________34882), .QN (____0________________21715));
  or2s1 ____99_500492(.DIN1
       (_____________________________________0_______21758), .DIN2
       (_________34909), .Q (_________34910));
  xor2s1 ____9__500493(.DIN1 (_________34867), .DIN2 (_________34907),
       .Q (_________34908));
  nnd2s1 ____9__500494(.DIN1 (______0__34880), .DIN2 (______0__33177),
       .Q (_________34906));
  xor2s1 ___900_500495(.DIN1 (___0__0__40491), .DIN2 (______0__34888),
       .Q (______0__34905));
  nnd2s1 ____99_500496(.DIN1 (_________34909), .DIN2
       (_____________________________________0_______21758), .Q
       (______9__34904));
  nnd2s1 ____99_500497(.DIN1 (_________34876), .DIN2 (_________35186),
       .Q (_________34903));
  hi1s1 ____9__500498(.DIN (______9__35627), .Q (_________34902));
  nnd2s1 ____500499(.DIN1 (_________34878), .DIN2 (________24868), .Q
       (_________34901));
  xor2s1 ___9000(.DIN1 (____0____32506), .DIN2 (______9__34887), .Q
       (_________34900));
  nnd2s1 ___900_500500(.DIN1 (_________34909), .DIN2
       (_____________________________________________21853), .Q
       (_________34943));
  or2s1 ___900_500501(.DIN1
       (_____________________________________________21853), .DIN2
       (_________34909), .Q (_________34942));
  xor2s1 ___90_500502(.DIN1 (_________34860), .DIN2 (______0__34897),
       .Q (_________34898));
  xor2s1 ___90__500503(.DIN1 (_________34861), .DIN2 (_________36762),
       .Q (______9__34896));
  nnd2s1 ___9___(.DIN1 (______9__34870), .DIN2 (__9_____30414), .Q
       (_________34895));
  nnd2s1 ___90__500504(.DIN1 (______0__34871), .DIN2 (____0____35361),
       .Q (_________34894));
  dffacs1 _______________________________________________500505(.CLRB
       (reset), .CLK (clk), .DIN (_________34879), .QN
       (___0_00__40561));
  nnd2s1 ___90__500506(.DIN1 (_________34885), .DIN2
       (_______________________________________________________________________________________),
       .Q (_________34952));
  nor2s1 ___9_0_500507(.DIN1 (___0____22290), .DIN2 (_________34873),
       .Q (_________34913));
  dffacs1 ______________________________________________500508(.CLRB
       (reset), .CLK (clk), .DIN (_________34874), .QN
       (____________________________________________21806));
  dffacs1 ______________________________________________500509(.CLRB
       (reset), .CLK (clk), .DIN (_________34875), .QN
       (____________________________________________21820));
  hi1s1 ___909_(.DIN (_________34912), .Q (_________34954));
  xor2s1 ___900_500510(.DIN1 (_____0___34853), .DIN2 (_________34626),
       .Q (_________34893));
  and2s1 ____9__500511(.DIN1 (_________34868), .DIN2 (________24574),
       .Q (_________34892));
  xor2s1 ___900_500512(.DIN1 (_________33198), .DIN2 (_________40880),
       .Q (_________34891));
  nnd2s1 ____9__500513(.DIN1 (______9__34863), .DIN2 (_________35435),
       .Q (_________34890));
  or2s1 ___90__500514(.DIN1 (______0__34888), .DIN2 (_________33654),
       .Q (_________34889));
  or2s1 ___90__500515(.DIN1 (____9____32452), .DIN2 (______9__34887),
       .Q (_________34918));
  xnr2s1 ____9__500516(.DIN1 (____90___36104), .DIN2 (_____09__34854),
       .Q (______9__35627));
  hi1s1 ___9___500517(.DIN (_________34885), .Q (_________34886));
  xor2s1 ___90__500518(.DIN1 (_________34869), .DIN2 (_________34883),
       .Q (_________34884));
  nnd2s1 ___9_0_500519(.DIN1 (_________34862), .DIN2 (_____9___34752),
       .Q (_________34882));
  xor2s1 ___90__500520(.DIN1
       (____________________________________________21819), .DIN2
       (_____9___34845), .Q (_________34881));
  nor2s1 ___90__500521(.DIN1 (_________33592), .DIN2 (_________34866),
       .Q (_________34911));
  xor2s1 ___9_0_500522(.DIN1 (________27672), .DIN2 (_________34872),
       .Q (_________34912));
  dffacs1 _____________________0_500523(.CLRB (reset), .CLK (clk), .DIN
       (_________34859), .QN (_________________0___21687));
  dffacs1 ____0__________________500524(.CLRB (reset), .CLK (clk), .DIN
       (_________34858), .QN (____0______________));
  nnd2s1 ___90__500525(.DIN1 (_________40880), .DIN2 (_________33190),
       .Q (______0__34880));
  or2s1 ___90__500526(.DIN1 (_____9___35559), .DIN2 (_____0___34850),
       .Q (_________34879));
  nnd2s1 ___90__500527(.DIN1 (_____0___34852), .DIN2 (_________34877),
       .Q (_________34878));
  xor2s1 ___90__500528(.DIN1 (_____9___33614), .DIN2 (_________34865),
       .Q (_________34876));
  nnd2s1 ___90__500529(.DIN1 (_____0___34851), .DIN2 (_________34262),
       .Q (_________34875));
  xor2s1 ___90_500530(.DIN1 (_________34832), .DIN2 (_________34907),
       .Q (_________34909));
  nnd2s1 ___90__500531(.DIN1 (_________34064), .DIN2 (_____0___34848),
       .Q (_________34874));
  nor2s1 ___9__9(.DIN1 (________22474), .DIN2 (_________34872), .Q
       (_________34873));
  nor2s1 ___90__500532(.DIN1 (___9____25059), .DIN2 (_____99__34846),
       .Q (______0__34871));
  nnd2s1 ___9__0(.DIN1 (_____9___34843), .DIN2 (____9____32424), .Q
       (______9__34870));
  nnd2s1 ___90__500533(.DIN1 (_________34869), .DIN2 (_________34579),
       .Q (_________34899));
  nnd2s1 ___9___500534(.DIN1 (_____9___34839), .DIN2 (_____9__22498),
       .Q (_________34885));
  dffacs1 _____________________________________________0_500535(.CLRB
       (reset), .CLK (clk), .DIN (_________34856), .Q (___0_9___40553));
  dffacs1 ______________________________________________500536(.CLRB
       (reset), .CLK (clk), .DIN (_________34857), .QN
       (____________________________________________21866));
  nnd2s1 ___90_500537(.DIN1 (______9__34837), .DIN2 (_________34796),
       .Q (_________34868));
  xor2s1 ___90__500538(.DIN1 (_________34812), .DIN2 (_____0___35566),
       .Q (_________34867));
  and2s1 ___90__500539(.DIN1 (_________33600), .DIN2 (_________34865),
       .Q (_________34866));
  xor2s1 ___900_500540(.DIN1 (_________34816), .DIN2 (___9_____39231),
       .Q (______9__34863));
  nor2s1 ___90__500541(.DIN1 (_________33544), .DIN2 (_________34836),
       .Q (______0__34888));
  nor2s1 ___9___500542(.DIN1 (___0_0___31123), .DIN2 (______0__34828),
       .Q (_________34862));
  xor2s1 ___9___500543(.DIN1 (_____9___34838), .DIN2 (_________37321),
       .Q (_________34861));
  xor2s1 ___9___500544(.DIN1 (_________34805), .DIN2 (_________35844),
       .Q (_________34860));
  nnd2s1 ___9___500545(.DIN1 (_________34821), .DIN2 (______0__32744),
       .Q (_________34859));
  nnd2s1 ___9__500546(.DIN1 (_________34820), .DIN2 (_________34576),
       .Q (_________34858));
  nor2s1 ___90__500547(.DIN1 (_____9___34844), .DIN2 (_________34831),
       .Q (______9__34887));
  dffacs1 ______________________________________________500548(.CLRB
       (reset), .CLK (clk), .DIN (_________34833), .QN
       (____________________________________________21834));
  nnd2s1 ___90__500549(.DIN1 (______9__34818), .DIN2 (_________34146),
       .Q (_________34857));
  nnd2s1 ___90__500550(.DIN1 (_________34817), .DIN2 (______0__34855),
       .Q (_________34856));
  xor2s1 ___90__500551(.DIN1 (_________34801), .DIN2 (______9__34981),
       .Q (_____09__34854));
  xor2s1 ___90__500552(.DIN1 (___0_____40502), .DIN2 (_________34829),
       .Q (_____0___34853));
  xor2s1 ___90_500553(.DIN1 (______0__33566), .DIN2 (_________34835),
       .Q (_____0___34852));
  nnd2s1 ___90__500554(.DIN1 (_________34813), .DIN2 (______9__35170),
       .Q (_____0___34851));
  nnd2s1 ___90__500555(.DIN1 (_________34814), .DIN2 (________25431),
       .Q (_____0___34850));
  or2s1 ___90__500556(.DIN1 (_____00__34847), .DIN2 (_________34815),
       .Q (_____0___34848));
  and2s1 ___909_500557(.DIN1 (______0__34810), .DIN2 (____9____35258),
       .Q (_____99__34846));
  nor2s1 ___909_500558(.DIN1 (_________34830), .DIN2 (_____9___34844),
       .Q (_____9___34845));
  nor2s1 ___9___500559(.DIN1 (_________41273), .DIN2 (______9__34809),
       .Q (_____9___34843));
  xor2s1 ___9__500560(.DIN1 (___________9___22071), .DIN2
       (_____9___34840), .Q (_____9___34842));
  xor2s1 ___9___500561(.DIN1 (_____9___34840), .DIN2 (_________35867),
       .Q (_____9___34841));
  or2s1 ___9___500562(.DIN1 (___0____22337), .DIN2 (_____9___34838), .Q
       (_____9___34839));
  nor2s1 ___9___500563(.DIN1 (_________34804), .DIN2 (_________34806),
       .Q (_________34872));
  xor2s1 ___9_0_500564(.DIN1 (_________34795), .DIN2 (___99_9__39836),
       .Q (_________34869));
  dffacs1 ______________________________________________500565(.CLRB
       (reset), .CLK (clk), .DIN (_________34811), .QN
       (____________________________________________21793));
  xor2s1 ___90__500566(.DIN1 (_________34763), .DIN2 (______0__34897),
       .Q (______9__34837));
  nor2s1 ___90_500567(.DIN1 (_________34835), .DIN2 (_________33563),
       .Q (_________34836));
  nnd2s1 ___90_500568(.DIN1 (______0__34800), .DIN2 (inData[0]), .Q
       (_________34834));
  nnd2s1 ___90__500569(.DIN1 (_________34797), .DIN2 (___9____23189),
       .Q (_________34833));
  xor2s1 ___9_0_500570(.DIN1 (_____0___34757), .DIN2 (___0__9__40412),
       .Q (_________34832));
  nor2s1 ___909_500571(.DIN1
       (____________________________________________21819), .DIN2
       (_________34830), .Q (_________34831));
  nnd2s1 ___90__500572(.DIN1 (______9__34799), .DIN2 (____9____33352),
       .Q (_________34865));
  or2s1 ___90__500573(.DIN1 (_________32910), .DIN2 (_________34829),
       .Q (_________34864));
  nnd2s1 ___9__500574(.DIN1 (_________34782), .DIN2 (___0_0___31124),
       .Q (______0__34828));
  or2s1 ___9___500575(.DIN1 (_________36556), .DIN2 (_____9___34840),
       .Q (______9__34827));
  nnd2s1 ___9___500576(.DIN1 (_____9___34840), .DIN2 (_________36556),
       .Q (_________34826));
  nor2s1 ___9___500577(.DIN1 (_________34824), .DIN2 (______0__34790),
       .Q (_________34825));
  nor2s1 ___9___500578(.DIN1 (_______________22077), .DIN2
       (_____9___34840), .Q (_________34823));
  xor2s1 ___9___500579(.DIN1 (_________34737), .DIN2
       (_____________________________________________21841), .Q
       (_________34822));
  nor2s1 ___9___500580(.DIN1 (___09____31428), .DIN2 (_________34783),
       .Q (_________34821));
  nor2s1 ___9__500581(.DIN1 (_________33769), .DIN2 (_________34784),
       .Q (_________34820));
  nnd2s1 ___90__500582(.DIN1 (_________34778), .DIN2 (_________34916),
       .Q (______9__34818));
  xor2s1 ___90__500583(.DIN1 (_____9___34748), .DIN2 (_________34718),
       .Q (_________34817));
  xor2s1 ___90__500584(.DIN1 (_____9___34747), .DIN2 (_________33006),
       .Q (_________34816));
  nnd2s1 ___9___500585(.DIN1 (___9_9___39339), .DIN2 (______0__34762),
       .Q (_________34815));
  or2s1 ___909_500586(.DIN1 (_________35448), .DIN2 (_________34768),
       .Q (_________34814));
  xor2s1 ___909_500587(.DIN1 (______9__34743), .DIN2 (____0____37113),
       .Q (_________34813));
  xor2s1 ___9099(.DIN1 (___________________________________________),
       .DIN2 (_________34798), .Q (_________34812));
  nnd2s1 ___9_0_500588(.DIN1 (_____9___34751), .DIN2 (________24048),
       .Q (_________34811));
  nnd2s1 ___90__500589(.DIN1 (_________34765), .DIN2 (______9__34981),
       .Q (_____0___34849));
  xor2s1 ___9___500590(.DIN1 (_____90__34181), .DIN2 (_________34794),
       .Q (______0__34810));
  nnd2s1 ___9___500591(.DIN1 (_____00__34754), .DIN2 (_________31778),
       .Q (______9__34809));
  nor2s1 ___9___500592(.DIN1 (_________35844), .DIN2 (_________34781),
       .Q (_________34808));
  xor2s1 ___9___500593(.DIN1 (___0_____40507), .DIN2 (____000__36182),
       .Q (_________34807));
  nor2s1 ___9_0_500594(.DIN1 (_________35844), .DIN2 (_________34803),
       .Q (_________34806));
  nor2s1 ___9___500595(.DIN1 (_________34804), .DIN2 (_________34803),
       .Q (_________34805));
  nor2s1 ___9___500596(.DIN1 (_________34722), .DIN2 (_____0___34755),
       .Q (_____9___34838));
  nor2s1 ___9___500597(.DIN1 (_____9___34281), .DIN2 (______0__34780),
       .Q (_____9___34844));
  dffacs1 ______________________________________________500598(.CLRB
       (reset), .CLK (clk), .DIN (_________34769), .QN
       (____________________________________________21830));
  dffacs1 ____0__________________500599(.CLRB (reset), .CLK (clk), .DIN
       (_____99__34753), .QN (____0________________21720));
  xor2s1 ___9_00(.DIN1 (_________34773), .DIN2 (________27451), .Q
       (_________34802));
  xor2s1 ___9_0_500600(.DIN1 (_________33872), .DIN2 (_________34766),
       .Q (_________34801));
  and2s1 ___9___500601(.DIN1 (___9_9___39339), .DIN2 (_____9___34749),
       .Q (______0__34800));
  nnd2s1 ___9___500602(.DIN1 (_________34798), .DIN2 (____90___33343),
       .Q (______9__34799));
  nnd2s1 ___909_500603(.DIN1 (_____90__34744), .DIN2 (_________34796),
       .Q (_________34797));
  nnd2s1 ___9___500604(.DIN1 (_________34741), .DIN2 (_________34545),
       .Q (_________34795));
  nor2s1 ___9___500605(.DIN1 (____9____34309), .DIN2 (______9__34779),
       .Q (_________34830));
  xor2s1 ___9__500606(.DIN1 (______0__34725), .DIN2 (_________35677),
       .Q (_________34835));
  xor2s1 ___9___500607(.DIN1 (_________34732), .DIN2 (_____9___37002),
       .Q (_________34829));
  nnd2s1 ___9__500608(.DIN1 (_________34067), .DIN2 (_________34794),
       .Q (______0__34819));
  nnd2s1 ___9___500609(.DIN1 (_____9___34746), .DIN2 (_________34607),
       .Q (_____0___34934));
  nor2s1 ___9___500610(.DIN1 (___0_____40507), .DIN2 (_________36382),
       .Q (_________34793));
  xor2s1 ___9___500611(.DIN1 (_________34791), .DIN2
       (_____________________________________________21825), .Q
       (_________34792));
  hi1s1 ___9__500612(.DIN (______9__34789), .Q (______0__34790));
  nor2s1 ___9___500613(.DIN1
       (_____________________________________________21841), .DIN2
       (_________36382), .Q (_________34788));
  nnd2s1 ___9___500614(.DIN1 (_________36382), .DIN2
       (_____________________________________________21841), .Q
       (_________34787));
  xor2s1 ___9___500615(.DIN1 (___0_90__40551), .DIN2 (_________35977),
       .Q (_________34786));
  and2s1 ___9___500616(.DIN1 (_________36382), .DIN2 (___0_____40507),
       .Q (_________34785));
  nnd2s1 ___9___500617(.DIN1 (_________34739), .DIN2 (_____0___34487),
       .Q (_________34784));
  nnd2s1 ___9_9_(.DIN1 (_________34742), .DIN2 (___0__9__31012), .Q
       (_________34783));
  nor2s1 ___9___500618(.DIN1 (________28912), .DIN2 (_________34738),
       .Q (_________34782));
  hi1s1 ___9_0_500619(.DIN (_________34781), .Q (_____9___34840));
  hi1s1 ___9__500620(.DIN (______9__34779), .Q (______0__34780));
  xor2s1 ___909_500621(.DIN1 (_________34717), .DIN2 (_____0___34663),
       .Q (_________34778));
  xor2s1 ___9_0_500622(.DIN1
       (_____________________________________________21796), .DIN2
       (_________34727), .Q (_________34777));
  and2s1 ___9___500623(.DIN1 (_________34773), .DIN2
       (_____________________________________________21796), .Q
       (_________34774));
  or2s1 ___9___500624(.DIN1
       (_____________________________________________21796), .DIN2
       (_________34773), .Q (______0__34772));
  nnd2s1 ___9___500625(.DIN1 (_________34773), .DIN2
       (_____________________________________________21809), .Q
       (______9__34771));
  or2s1 ___9___500626(.DIN1
       (_____________________________________________21809), .DIN2
       (_________34773), .Q (_________34770));
  nnd2s1 ___9__500627(.DIN1 (____99___34381), .DIN2 (_________34729),
       .Q (_________34769));
  xor2s1 ___9___500628(.DIN1 (_________34618), .DIN2 (_____9___34745),
       .Q (_________34768));
  nor2s1 ___9___500629(.DIN1 (_________34764), .DIN2 (_________34766),
       .Q (_________34767));
  nnd2s1 ___9___500630(.DIN1 (_________34766), .DIN2 (_________34764),
       .Q (_________34765));
  xor2s1 ___9__500631(.DIN1 (_________34716), .DIN2 (____0____32505),
       .Q (_________34763));
  nnd2s1 ___9___500632(.DIN1 (_________34731), .DIN2 (_________34691),
       .Q (______0__34762));
  nor2s1 ___9___500633(.DIN1 (___0_90__40551), .DIN2 (_________35977),
       .Q (_____0___34761));
  and2s1 ___9___500634(.DIN1 (_________35977), .DIN2 (___0_90__40551),
       .Q (_____0___34760));
  and2s1 ___9___500635(.DIN1 (_________35977), .DIN2
       (_____________________________________________21825), .Q
       (_____0___34759));
  nor2s1 ___9__500636(.DIN1
       (_____________________________________________21825), .DIN2
       (_________35977), .Q (_____0___34758));
  xor2s1 ___9___500637(.DIN1 (_____0___34756), .DIN2 (_________34740),
       .Q (_____0___34757));
  nor2s1 ___9___500638(.DIN1 (_________36480), .DIN2 (_________34721),
       .Q (_____0___34755));
  nor2s1 ___9_9_500639(.DIN1 (_________33123), .DIN2 (______9__34724),
       .Q (_____00__34754));
  nnd2s1 ___9_9_500640(.DIN1 (_________34723), .DIN2 (_____9___34752),
       .Q (_____99__34753));
  or2s1 ___9___500641(.DIN1 (______0__35050), .DIN2 (_________34726),
       .Q (_____9___34751));
  nnd2s1 ___9_9_500642(.DIN1 (_________35977), .DIN2
       (_________________________________________0___21840), .Q
       (______9__34789));
  nor2s1 ___9_9_500643(.DIN1
       (_________________________________________0___21840), .DIN2
       (_________35977), .Q (_________34824));
  xor2s1 ___9___500644(.DIN1 (_________34684), .DIN2 (_________34708),
       .Q (_________34781));
  and2s1 ___9___500645(.DIN1 (_____9___34750), .DIN2
       (_______________________________________________________________________________________),
       .Q (_________34803));
  nor2s1 ___9___500646(.DIN1
       (_______________________________________________________________________________________),
       .DIN2 (_____9___34750), .Q (_________34804));
  dffacs1 ______________________________________________500647(.CLRB
       (reset), .CLK (clk), .DIN (_________34736), .QN
       (___0_____40512));
  xnr2s1 ___9___500648(.DIN1 (_________34730), .DIN2
       (____________________________________________21806), .Q
       (_____9___34749));
  xor2s1 ___9___500649(.DIN1 (______9__34696), .DIN2 (______0__33312),
       .Q (_____9___34748));
  xor2s1 ___9___500650(.DIN1 (_____9___22051), .DIN2 (_________34728),
       .Q (_____9___34747));
  or2s1 ___9___500651(.DIN1 (_________34602), .DIN2 (_____9___34745),
       .Q (_____9___34746));
  xor2s1 ___9__500652(.DIN1 (______0__34697), .DIN2 (_________34712),
       .Q (_____90__34744));
  xor2s1 ___9___500653(.DIN1 (_________34690), .DIN2 (_________34709),
       .Q (______9__34743));
  nnd2s1 ___9___500654(.DIN1 (_________34719), .DIN2 (_________34681),
       .Q (_________34798));
  nnd2s1 ___9__500655(.DIN1 (_________34713), .DIN2 (_________34674),
       .Q (______9__34779));
  nor2s1 ___9__500656(.DIN1 (___0_____30812), .DIN2 (_________34706),
       .Q (_________34742));
  nnd2s1 ___9_0_500657(.DIN1 (_________34740), .DIN2 (_________34542),
       .Q (_________34741));
  nor2s1 ___9___500658(.DIN1 (___0_____31186), .DIN2 (_________34707),
       .Q (_________34739));
  nnd2s1 ___9___500659(.DIN1 (_________34711), .DIN2 (__9_____30022),
       .Q (_________34738));
  nnd2s1 ___9_9_500660(.DIN1 (_________34710), .DIN2 (_________34672),
       .Q (_________34794));
  hi1s1 ___9___500661(.DIN (_________34737), .Q (____000__36182));
  dffacs1 ______________________________________________500662(.CLRB
       (reset), .CLK (clk), .DIN (______0__34715), .QN
       (___0_____40492));
  nb1s1 ___9___500663(.DIN (_________34737), .Q (_________36382));
  nnd2s1 ___9_0_500664(.DIN1 (_________34695), .DIN2 (______0__35181),
       .Q (_________34736));
  nor2s1 ___9__500665(.DIN1 (_________34704), .DIN2 (______0__34734),
       .Q (_________34735));
  nnd2s1 ___9_90(.DIN1 (_________34702), .DIN2 (____9____32458), .Q
       (_________34732));
  nnd2s1 ___9___500666(.DIN1 (_________34730), .DIN2 (_____0___33161),
       .Q (_________34731));
  nnd2s1 ___9___500667(.DIN1 (_________34145), .DIN2 (_________34698),
       .Q (_________34729));
  or2s1 ___9___500668(.DIN1 (_________33042), .DIN2 (_________34728),
       .Q (_________34776));
  nor2s1 ___9___500669(.DIN1 (_____9___33806), .DIN2 (_________34700),
       .Q (_________34766));
  hi1s1 ___9__500670(.DIN (_________34727), .Q (_________34773));
  xor2s1 ___9___500671(.DIN1 (_____9___22049), .DIN2 (_________34669),
       .Q (_________34726));
  nor2s1 ___9__500672(.DIN1 (_____0___34664), .DIN2 (_________34693),
       .Q (______0__34725));
  nnd2s1 ___9___500673(.DIN1 (_________34683), .DIN2 (________27526),
       .Q (______9__34724));
  nor2s1 ___9___500674(.DIN1 (___0_____31229), .DIN2 (_________34688),
       .Q (_________34723));
  nor2s1 ___9___500675(.DIN1 (_________37452), .DIN2 (_________34685),
       .Q (_________34722));
  nor2s1 ___9___500676(.DIN1 (________22564), .DIN2 (______0__34687),
       .Q (_________34721));
  xor2s1 ___9__500677(.DIN1 (______0__34668), .DIN2 (____9____38944),
       .Q (_________34737));
  nor2s1 ___9___500678(.DIN1 (_________34689), .DIN2 (_________34694),
       .Q (_____9___34750));
  hi1s1 ___9__500679(.DIN (_________34720), .Q (_________34791));
  nb1s1 ___9___500680(.DIN (_________34720), .Q (_________35977));
  nnd2s1 ___9___500681(.DIN1 (______0__34677), .DIN2 (_________34718),
       .Q (_________34719));
  xor2s1 ___9__500682(.DIN1 (_____0___34659), .DIN2 (_________34692),
       .Q (_________34717));
  xor2s1 ___9___500683(.DIN1 (___0_____40503), .DIN2 (_________34701),
       .Q (_________34716));
  nnd2s1 ___9_09(.DIN1 (_________34673), .DIN2 (____0____34453), .Q
       (______0__34715));
  nnd2s1 ___9___500684(.DIN1 (_________34679), .DIN2 (_________35680),
       .Q (______9__34714));
  or2s1 ___9___500685(.DIN1 (_________34682), .DIN2 (_________34712),
       .Q (_________34713));
  xor2s1 ___9___500686(.DIN1 (_____00__34658), .DIN2 (_________36512),
       .Q (_____9___34745));
  xor2s1 ___9___500687(.DIN1 (_________34699), .DIN2 (_____9___33807),
       .Q (_________34727));
  nnd2s1 ___9___500688(.DIN1 (_____0___34665), .DIN2 (____9____32424),
       .Q (_________34711));
  or2s1 ___9___500689(.DIN1 (_________34670), .DIN2 (_________34709),
       .Q (_________34710));
  xor2s1 ___9_500690(.DIN1 (______9__34686), .DIN2 (____0____38091), .Q
       (_________34708));
  nnd2s1 ___9___500691(.DIN1 (_____09__34667), .DIN2 (___09_9__31426),
       .Q (_________34707));
  nor2s1 ___9___500692(.DIN1 (____0____32541), .DIN2 (_____0___34666),
       .Q (_________34706));
  xnr2s1 ___9___500693(.DIN1 (_________36527), .DIN2 (_____9___34653),
       .Q (_________34740));
  xor2s1 ___9__500694(.DIN1 (_____9___34652), .DIN2 (_________38155),
       .Q (_________34720));
  dffacs1 ______________________________________________500695(.CLRB
       (reset), .CLK (clk), .DIN (_________34678), .QN
       (____________________________________________21832));
  dffacs1 ______________________________________________500696(.CLRB
       (reset), .CLK (clk), .DIN (_________34680), .QN
       (____________________________________________21833));
  hi1s1 ___9__500697(.DIN (_________34703), .Q (_________34704));
  or2s1 ___9___500698(.DIN1 (____9____32457), .DIN2 (_________34701),
       .Q (_________34702));
  and2s1 ___9_0_500699(.DIN1 (_________34699), .DIN2 (_________33749),
       .Q (_________34700));
  xor2s1 ___9___500700(.DIN1 (___0_____40503), .DIN2 (___0_____40513),
       .Q (_________34698));
  xor2s1 ___9___500701(.DIN1 (___0_____40513), .DIN2 (_________34034),
       .Q (______0__34697));
  xor2s1 ___9__500702(.DIN1 (___0_0___40562), .DIN2 (_________38842),
       .Q (______9__34696));
  nor2s1 ___9__500703(.DIN1 (________24917), .DIN2 (_____0___34662), .Q
       (_________34695));
  nor2s1 ___9_9_500704(.DIN1 (_________34636), .DIN2 (_____0___34661),
       .Q (_________34728));
  nor2s1 ___9___500705(.DIN1 (_________37321), .DIN2 (_____9___34651),
       .Q (_________34694));
  and2s1 ___9___500706(.DIN1 (_____9___34656), .DIN2 (_________34692),
       .Q (_________34693));
  or2s1 ___9__500707(.DIN1
       (____________________________________________21819), .DIN2
       (________22441), .Q (_________34691));
  xor2s1 ___9___500708(.DIN1
       (____________________________________________21807), .DIN2
       (_________34671), .Q (_________34690));
  nor2s1 ___9_9_500709(.DIN1 (____99___36174), .DIN2 (_________40882),
       .Q (_________34689));
  nnd2s1 ___9___500710(.DIN1 (_____9___34654), .DIN2 (___0____28761),
       .Q (_________34688));
  and2s1 ___9___500711(.DIN1 (______9__34686), .DIN2 (____0___23043),
       .Q (______0__34687));
  or2s1 ___9__500712(.DIN1 (_________34684), .DIN2 (______9__34686), .Q
       (_________34685));
  nor2s1 ___9__500713(.DIN1 (________29508), .DIN2 (______9__34648), .Q
       (_________34683));
  and2s1 ___9___500714(.DIN1 (___0_____40502), .DIN2
       (____________________________________________21819), .Q
       (_________34730));
  dffacs1 ____0________________0_(.CLRB (reset), .CLK (clk), .DIN
       (_____90__34649), .QN (____0____________0___21713));
  nor2s1 ___9___500715(.DIN1 (___0_____40513), .DIN2 (___0_____31295),
       .Q (_________34682));
  or2s1 ___9__500716(.DIN1 (___0_0___40562), .DIN2 (______0__33312), .Q
       (_________34681));
  nnd2s1 ___9_0_500717(.DIN1 (_________34645), .DIN2 (____9____34339),
       .Q (_________34680));
  xor2s1 ___9___500718(.DIN1 (___09____40682), .DIN2 (___0_0___40563),
       .Q (_________34679));
  nnd2s1 ___9___500719(.DIN1 (_________34522), .DIN2 (_________34643),
       .Q (_________34678));
  nnd2s1 ___9___500720(.DIN1 (______0__33312), .DIN2 (___0_0___40562),
       .Q (______0__34677));
  nnd2s1 ___9___500721(.DIN1 (_________34646), .DIN2 (_________35186),
       .Q (______9__34676));
  nor2s1 ___9_9_500722(.DIN1
       (_____________________________________________21808), .DIN2
       (_________34675), .Q (______0__34734));
  nnd2s1 ___9_9_500723(.DIN1 (_________34675), .DIN2
       (_____________________________________________21808), .Q
       (_________34703));
  nnd2s1 ___9___500724(.DIN1 (___0_____31295), .DIN2 (___0_____40513),
       .Q (_________34674));
  nnd2s1 ___9___500725(.DIN1 (_________34642), .DIN2 (_________34644),
       .Q (_________34673));
  or2s1 ___9___500726(.DIN1
       (____________________________________________21807), .DIN2
       (_________34671), .Q (_________34672));
  and2s1 ___9___500727(.DIN1 (_________34671), .DIN2
       (____________________________________________21807), .Q
       (_________34670));
  nnd2s1 ___9___500728(.DIN1 (_________34637), .DIN2 (_____0___34660),
       .Q (_________34669));
  xnr2s1 ___9___500729(.DIN1 (_____9___34650), .DIN2 (____00__27031),
       .Q (______0__34668));
  nor2s1 ___9___500730(.DIN1 (____9____34365), .DIN2 (_________34641),
       .Q (_____09__34667));
  nnd2s1 ___9_0_500731(.DIN1 (______0__34639), .DIN2 (________29108),
       .Q (_____0___34666));
  nor2s1 ___9_500732(.DIN1 (_________32058), .DIN2 (______9__34638), .Q
       (_____0___34665));
  dffacs1 ________________________(.CLRB (reset), .CLK (clk), .DIN
       (_________34640), .QN (______________________21700));
  nor2s1 ___9___500733(.DIN1 (_____9___34655), .DIN2 (_____0___34663),
       .Q (_____0___34664));
  nor2s1 ___9___500734(.DIN1 (_____0___35834), .DIN2 (______9__34630),
       .Q (_____0___34662));
  and2s1 ___9___500735(.DIN1 (_____0___34660), .DIN2 (_____9___22049),
       .Q (_____0___34661));
  xor2s1 ___9___500736(.DIN1
       (____________________________________________21849), .DIN2
       (_________37614), .Q (_____0___34659));
  nnd2s1 ___9___500737(.DIN1 (_________34633), .DIN2 (_________34515),
       .Q (_____00__34658));
  nor2s1 ___9_9_500738(.DIN1
       (_____________________________________________21795), .DIN2
       (_____99__34657), .Q (_________34733));
  xor2s1 ___9___500739(.DIN1 (_________40886), .DIN2 (___9_____39123),
       .Q (_________34699));
  and2s1 ___9_9_500740(.DIN1 (_____99__34657), .DIN2
       (_____________________________________________21795), .Q
       (______9__34705));
  dffacs1 ______________________________________________500741(.CLRB
       (reset), .CLK (clk), .DIN (_________34635), .QN
       (____________________________________________21819));
  nnd2s1 ___9___500742(.DIN1 (_____0___34663), .DIN2 (_____9___34655),
       .Q (_____9___34656));
  nor2s1 ___9_9_500743(.DIN1 (___0_____31008), .DIN2 (_________34627),
       .Q (_____9___34654));
  nor2s1 ___9___500744(.DIN1 (______0__34544), .DIN2 (_________34629),
       .Q (_____9___34653));
  xor2s1 ___9___500745(.DIN1 (______9__34621), .DIN2 (_________37412),
       .Q (_____9___34652));
  nor2s1 ___9___500746(.DIN1 (_____9__25519), .DIN2 (_____9___34650),
       .Q (_____9___34651));
  nnd2s1 ___9_9_500747(.DIN1 (______0__34631), .DIN2 (_________33193),
       .Q (_____90__34649));
  nnd2s1 ___9___500748(.DIN1 (_________34628), .DIN2 (_________32692),
       .Q (______9__34648));
  nor2s1 ___9_9_500749(.DIN1 (_____0___32096), .DIN2 (_________34634),
       .Q (_________34701));
  xor2s1 ___9___500750(.DIN1 (_________34615), .DIN2 (_________34647),
       .Q (______9__34686));
  xor2s1 ___9___500751(.DIN1 (_____0___34570), .DIN2 (_________34632),
       .Q (_________34646));
  nnd2s1 ___9___500752(.DIN1 (_________34624), .DIN2 (_________34644),
       .Q (_________34645));
  or2s1 ___9___500753(.DIN1
       (____________________________________________21849), .DIN2
       (____9____34338), .Q (_________34643));
  xor2s1 ___9___500754(.DIN1 (_________32169), .DIN2 (_________40888),
       .Q (_________34642));
  nnd2s1 ___9___500755(.DIN1 (_________34623), .DIN2 (______0__33186),
       .Q (_________34718));
  hi1s1 ___9__500756(.DIN (_____99__34657), .Q (_________34675));
  dffacs1 _____________________________________________0_500757(.CLRB
       (reset), .CLK (clk), .DIN (_________34619), .Q (___0_0___40562));
  dffacs1 ______________________________________________500758(.CLRB
       (reset), .CLK (clk), .DIN (_________34620), .QN
       (___0_____40513));
  dffacs1 _______________________(.CLRB (reset), .CLK (clk), .DIN
       (______9__34612), .QN (_____________________21678));
  nnd2s1 ___9___500759(.DIN1 (_________34610), .DIN2 (____9____34322),
       .Q (_________34641));
  nnd2s1 ___9___500760(.DIN1 (_________34614), .DIN2 (______9__33037),
       .Q (_________34640));
  nor2s1 ___9___500761(.DIN1 (__9_____30142), .DIN2 (_________34611),
       .Q (______0__34639));
  nnd2s1 ___9__500762(.DIN1 (______0__34613), .DIN2 (_________32296),
       .Q (______9__34638));
  hi1s1 ___9_9_500763(.DIN (_________34636), .Q (_________34637));
  nor2s1 ___9_0_500764(.DIN1 (_____00__33622), .DIN2 (_________34617),
       .Q (_________34671));
  dffacs1 ______________________________________________500765(.CLRB
       (reset), .CLK (clk), .DIN (_________34625), .QN
       (____________________________________________21807));
  dffacs1 ____0________________0_500766(.CLRB (reset), .CLK (clk), .DIN
       (_________34608), .QN (____0____________0_));
  dffacs1 _______________________500767(.CLRB (reset), .CLK (clk), .DIN
       (_________34609), .QN (_____________________21695));
  nnd2s1 ___9_0_500768(.DIN1 (_________34595), .DIN2 (____0___23973),
       .Q (_________34635));
  nor2s1 ___9_500769(.DIN1 (_____0___32094), .DIN2 (_________40888), .Q
       (_________34634));
  or2s1 ___9_99(.DIN1 (_________34513), .DIN2 (_________34632), .Q
       (_________34633));
  hi1s1 ___9_9_500770(.DIN
       (____________________________________________21849), .Q
       (_____9___34655));
  nor2s1 ___9__500771(.DIN1 (___0_____30722), .DIN2 (_________34606),
       .Q (_________34712));
  xor2s1 ___9___500772(.DIN1 (_________34591), .DIN2 (_____9___33617),
       .Q (_____99__34657));
  dffacs1 ______________________________________________500773(.CLRB
       (reset), .CLK (clk), .DIN (______0__34604), .QN
       (_____9___22049));
  nor2s1 ___9___500774(.DIN1 (___0_____30910), .DIN2 (_________34599),
       .Q (______0__34631));
  xor2s1 ___9__500775(.DIN1 (_________34616), .DIN2 (_____0___33623),
       .Q (______9__34630));
  nor2s1 ___9__500776(.DIN1 (______0__34499), .DIN2 (_________34598),
       .Q (_________34629));
  nor2s1 ___9__500777(.DIN1 (_________32602), .DIN2 (______0__34594),
       .Q (_________34628));
  nnd2s1 ___9___500778(.DIN1 (_________34600), .DIN2 (___0__9__31060),
       .Q (_________34627));
  nor2s1 ___9_0_500779(.DIN1 (_________34626), .DIN2 (_________40890),
       .Q (_________34636));
  nnd2s1 ___9_0_500780(.DIN1 (_________40890), .DIN2 (_________34626),
       .Q (_____0___34660));
  nnd2s1 ___9___500781(.DIN1 (_________34597), .DIN2 (________22467),
       .Q (_____9___34650));
  dffacs1 ______________________________________________500782(.CLRB
       (reset), .CLK (clk), .DIN (______9__34603), .QN
       (____________________________________________21831));
  nnd2s1 ___9___500783(.DIN1 (_________34592), .DIN2 (________24972),
       .Q (_________34625));
  xor2s1 ___9___500784(.DIN1 (___0_____30887), .DIN2 (_________34605),
       .Q (_________34624));
  nnd2s1 ___9_9_500785(.DIN1 (______0__34622), .DIN2 (_________33183),
       .Q (_________34623));
  xor2s1 ___9___500786(.DIN1 (___0_____40411), .DIN2 (_________34596),
       .Q (______9__34621));
  nnd2s1 ___9__500787(.DIN1 (______9__34593), .DIN2 (_____0__26466), .Q
       (_________34620));
  nnd2s1 ___9___500788(.DIN1 (_________34586), .DIN2 (______0__34855),
       .Q (_________34619));
  xor2s1 ___9___500789(.DIN1 (_____0__25425), .DIN2 (_________36034),
       .Q (_________34618));
  and2s1 ___9___500790(.DIN1 (_________33564), .DIN2 (_________34616),
       .Q (_________34617));
  dffacs1 ______________________________________________500791(.CLRB
       (reset), .CLK (clk), .DIN (_________34587), .QN
       (____________________________________________21849));
  nnd2s1 ___9___500792(.DIN1 (______9__34584), .DIN2 (_________34536),
       .Q (_________34615));
  nor2s1 ___9___500793(.DIN1 (_________33143), .DIN2 (_________34578),
       .Q (_________34614));
  nor2s1 ___9___500794(.DIN1 (________29529), .DIN2 (_________34581),
       .Q (______0__34613));
  nnd2s1 ___9___500795(.DIN1 (_________34582), .DIN2 (______0__31680),
       .Q (______9__34612));
  nnd2s1 ___9___500796(.DIN1 (_________34580), .DIN2 (________29331),
       .Q (_________34611));
  nor2s1 ___9___500797(.DIN1 (______9__34266), .DIN2 (_________34583),
       .Q (_________34610));
  or2s1 ___9___500798(.DIN1 (_________33175), .DIN2 (______0__34585),
       .Q (_________34609));
  nnd2s1 ___9___500799(.DIN1 (_________34577), .DIN2 (_________34154),
       .Q (_________34608));
  dffacs1 _______________________500800(.CLRB (reset), .CLK (clk), .DIN
       (______0__34575), .QN (_____________________21680));
  dffacs1 ______________________________________________500801(.CLRB
       (reset), .CLK (clk), .DIN (_________34589), .QN
       (____________________________________________21792));
  nnd2s1 ___9___500802(.DIN1 (_________36034), .DIN2 (_________34601),
       .Q (_________34607));
  and2s1 ___9_0_500803(.DIN1 (_________34605), .DIN2 (___0__0__30721),
       .Q (_________34606));
  nnd2s1 ___9___500804(.DIN1 (_____0___34571), .DIN2 (_________35435),
       .Q (______0__34604));
  nnd2s1 ___9___500805(.DIN1 (_____09__34574), .DIN2 (____00__23502),
       .Q (______9__34603));
  nor2s1 ___9___500806(.DIN1 (_________34601), .DIN2 (_________36034),
       .Q (_________34602));
  nor2s1 ___9___500807(.DIN1 (___00____30576), .DIN2 (_____9___34561),
       .Q (_________34600));
  nnd2s1 ___9__500808(.DIN1 (_____90__34560), .DIN2 (_____9__28905), .Q
       (_________34599));
  xor2s1 ___9__500809(.DIN1 (_________34539), .DIN2 (___0_____40323),
       .Q (_________34598));
  nnd2s1 ___9___500810(.DIN1 (_________34596), .DIN2 (___9___22266), .Q
       (_________34597));
  nnd2s1 ___9___500811(.DIN1 (_____9___34567), .DIN2 (_____0___34932),
       .Q (_________34595));
  nnd2s1 ___9__500812(.DIN1 (_________34559), .DIN2 (________29056), .Q
       (______0__34594));
  nor2s1 ___9___500813(.DIN1 (____0____34426), .DIN2 (_____99__34568),
       .Q (_________34632));
  dffacs1 ______________________________________________500814(.CLRB
       (reset), .CLK (clk), .DIN (_____0___34572), .QN
       (____________________________________________21848));
  nnd2s1 ___9___500815(.DIN1 (_________34557), .DIN2 (_________34916),
       .Q (______9__34593));
  nnd2s1 ___9___500816(.DIN1 (_________34551), .DIN2 (____9____35258),
       .Q (_________34592));
  xor2s1 ___9___500817(.DIN1 (_________34519), .DIN2 (____9____38944),
       .Q (_________34591));
  nor2s1 ___9___500818(.DIN1 (_________36402), .DIN2 (_________34883),
       .Q (_________34590));
  nnd2s1 ___9___500819(.DIN1 (_________34554), .DIN2 (_________41323),
       .Q (_________34589));
  xor2s1 ___9__500820(.DIN1
       (_________________________________________0___21824), .DIN2
       (_________35907), .Q (_________34588));
  nnd2s1 ___9___500821(.DIN1 (_________34552), .DIN2 (________26478),
       .Q (_________34587));
  xor2s1 ___9__500822(.DIN1 (____0____34428), .DIN2 (_________40892),
       .Q (_________34586));
  nnd2s1 ___9___500823(.DIN1 (_________34550), .DIN2 (____9____33379),
       .Q (_________34616));
  nnd2s1 ___9__500824(.DIN1 (_________34556), .DIN2 (_________33082),
       .Q (______0__34622));
  dffacs1 ______________________________________________500825(.CLRB
       (reset), .CLK (clk), .DIN (_________34555), .QN
       (____________________________________________21791));
  nnd2s1 ___9__500826(.DIN1 (_________34527), .DIN2 (_________34531),
       .Q (______0__34585));
  or2s1 ___9___500827(.DIN1 (_________38271), .DIN2 (_________34535),
       .Q (______9__34584));
  nnd2s1 ___9__500828(.DIN1 (______9__34533), .DIN2 (____999__33432),
       .Q (_________34583));
  nnd2s1 ___9__500829(.DIN1 (_________34528), .DIN2 (______0__34524),
       .Q (_________34582));
  nnd2s1 ___9___500830(.DIN1 (_________34541), .DIN2 (________29259),
       .Q (_________34581));
  nor2s1 ___9___500831(.DIN1 (___0_____30669), .DIN2 (______0__34534),
       .Q (_________34580));
  nnd2s1 ___9___500832(.DIN1 (_________34883), .DIN2 (_________36402),
       .Q (_________34579));
  nnd2s1 ___9___500833(.DIN1 (_________34530), .DIN2 (________28482),
       .Q (_________34578));
  and2s1 ___9___500834(.DIN1 (_________34529), .DIN2 (_________34576),
       .Q (_________34577));
  nnd2s1 ___9___500835(.DIN1 (_________34525), .DIN2 (_________31917),
       .Q (______0__34575));
  dffacs1 _______________________500836(.CLRB (reset), .CLK (clk), .DIN
       (_________34532), .QN (_____________________21692));
  dffacs1 ____0__________________500837(.CLRB (reset), .CLK (clk), .DIN
       (_________34526), .QN (____0________________21663));
  nnd2s1 ___9___500838(.DIN1 (_________34518), .DIN2 (_____0___34932),
       .Q (_____09__34574));
  nnd2s1 ___9___500839(.DIN1 (_________34520), .DIN2 (____0___23884),
       .Q (_____0___34572));
  xor2s1 ___9___500840(.DIN1 (______0__33084), .DIN2 (______0__40894),
       .Q (_____0___34571));
  xor2s1 ___9___500841(.DIN1 (_____0___34569), .DIN2 (___0_____40576),
       .Q (_____0___34570));
  nor2s1 ___9___500842(.DIN1 (____0____34427), .DIN2 (_________40892),
       .Q (_____99__34568));
  xor2s1 ___9__500843(.DIN1 (____9_9__33384), .DIN2 (_________34549),
       .Q (_____9___34567));
  xor2s1 ___9___500844(.DIN1 (_________34501), .DIN2 (_________38214),
       .Q (_________34605));
  dffacs1 _____________________9_(.CLRB (reset), .CLK (clk), .DIN
       (_________34505), .QN (_________________9___21685));
  nnd2s1 ___9___500845(.DIN1 (_________35907), .DIN2
       (_________________________________________0_), .Q
       (_____9___34566));
  or2s1 ___9___500846(.DIN1 (______0___22057), .DIN2 (_________35907),
       .Q (_____9___34565));
  and2s1 ___9__500847(.DIN1 (_________35907), .DIN2 (______0___22057),
       .Q (_____9___34564));
  nor2s1 ___9___500848(.DIN1
       (_________________________________________0_), .DIN2
       (_________35907), .Q (_____9___34563));
  xor2s1 ___9__500849(.DIN1 (___9____25991), .DIN2 (_________36778), .Q
       (_____9___34562));
  nor2s1 ___9__500850(.DIN1 (___0____25136), .DIN2 (______9__34507), .Q
       (_____9___34561));
  nnd2s1 ___9___500851(.DIN1 (_________34510), .DIN2 (____9____32424),
       .Q (_____90__34560));
  nor2s1 ___9___500852(.DIN1 (________25361), .DIN2 (_________34506),
       .Q (_________34559));
  nnd2s1 ___9___500853(.DIN1 (_________34509), .DIN2 (________27108),
       .Q (_________34596));
  dffacs1 ______________________________________________500854(.CLRB
       (reset), .CLK (clk), .DIN (_________34521), .QN
       (____________________________________________21818));
  xor2s1 ___9___500855(.DIN1 (_________34558), .DIN2 (_________34500),
       .Q (_________36034));
  dffacs1 ____0__________________500856(.CLRB (reset), .CLK (clk), .DIN
       (______0__34508), .QN (____0________________21662));
  xor2s1 ___9___500857(.DIN1 (_____00__34480), .DIN2 (_________41343),
       .Q (_________34557));
  nnd2s1 ___9__500858(.DIN1 (______0__40894), .DIN2 (______9__33083),
       .Q (_________34556));
  nnd2s1 ___9___500859(.DIN1 (_________34502), .DIN2 (____0___25869),
       .Q (_________34555));
  nnd2s1 ___9___500860(.DIN1 (_________34504), .DIN2 (____9____35258),
       .Q (_________34554));
  nnd2s1 ___9___500861(.DIN1 (_________34503), .DIN2 (_________34644),
       .Q (_________34552));
  xor2s1 ___9___500862(.DIN1 (_________34511), .DIN2 (_________33781),
       .Q (_________34551));
  or2s1 ___9_9_500863(.DIN1 (_________34549), .DIN2 (____9____33377),
       .Q (_________34550));
  xor2s1 ___9___500864(.DIN1 (_________34558), .DIN2 (_________35968),
       .Q (_________34548));
  or2s1 ___9___500865(.DIN1
       (_________________________________________0___21824), .DIN2
       (_________36778), .Q (_________34547));
  nnd2s1 ___9___500866(.DIN1 (_________36778), .DIN2
       (_________________________________________0___21824), .Q
       (_________34546));
  or2s1 ___9__500867(.DIN1 (_________36493), .DIN2 (_____0___34756), .Q
       (_________34545));
  nor2s1 ___9___500868(.DIN1 (_________34538), .DIN2 (______9__34543),
       .Q (______0__34544));
  nnd2s1 ___9___500869(.DIN1 (_____0___34756), .DIN2 (_________36493),
       .Q (_________34542));
  nor2s1 ___9___500870(.DIN1 (___0____27851), .DIN2 (_________34492),
       .Q (_________34541));
  or2s1 ___9___500871(.DIN1 (_________37412), .DIN2 (_____0___34756),
       .Q (_________34540));
  nnd2s1 ___9__500872(.DIN1 (______9__34543), .DIN2 (_________34538),
       .Q (_________34539));
  nnd2s1 ___9___500873(.DIN1 (_____0___34756), .DIN2 (_________37412),
       .Q (_________34537));
  nnd2s1 ___9_500874(.DIN1 (______9__34498), .DIN2 (_________38271), .Q
       (_________34536));
  nor2s1 ___9_0_500875(.DIN1 (________22581), .DIN2 (_________34495),
       .Q (_________34535));
  nnd2s1 ___9___500876(.DIN1 (_________34491), .DIN2 (___09____31461),
       .Q (______0__34534));
  and2s1 ___9__500877(.DIN1 (_____0___34486), .DIN2 (___0_____31164),
       .Q (______9__34533));
  nnd2s1 ___9___500878(.DIN1 (_________34490), .DIN2 (_________34531),
       .Q (_________34532));
  nor2s1 ___9___500879(.DIN1 (___0_____31293), .DIN2 (______0__34489),
       .Q (_________34530));
  nor2s1 ___9_0_500880(.DIN1 (____0_0__32518), .DIN2 (_________34494),
       .Q (_________34529));
  nor2s1 ___9_0_500881(.DIN1 (_________32311), .DIN2 (_____0___34484),
       .Q (_________34528));
  nor2s1 ___9_0_500882(.DIN1 (___0_____31064), .DIN2 (_________34493),
       .Q (_________34527));
  nnd2s1 ___9_0_500883(.DIN1 (_____09__34488), .DIN2 (___9____27773),
       .Q (_________34526));
  nnd2s1 ___9___500884(.DIN1 (_____0___34485), .DIN2 (______0__34524),
       .Q (_________34525));
  hi1s1 ___9_9_500885(.DIN (______9__34523), .Q (_________34883));
  nnd2s1 ___9___500886(.DIN1 (_____0___34482), .DIN2 (_________34644),
       .Q (_________34522));
  nnd2s1 ___9__500887(.DIN1 (____099__34479), .DIN2 (_____90__33707),
       .Q (_________34521));
  nnd2s1 ___9___500888(.DIN1 (_____0___34483), .DIN2 (_________34916),
       .Q (_________34520));
  xor2s1 ___9___500889(.DIN1 (_________34496), .DIN2 (_________36761),
       .Q (_________34519));
  xor2s1 ___9___500890(.DIN1 (____0____34458), .DIN2 (______0__37673),
       .Q (_________34518));
  or2s1 ___9_9_500891(.DIN1 (___0_____40576), .DIN2 (_________34514),
       .Q (_________34515));
  and2s1 ___9_9_500892(.DIN1 (_________34514), .DIN2 (___0_____40576),
       .Q (_________34513));
  nor2s1 ___9___500893(.DIN1 (_________34511), .DIN2 (_________33761),
       .Q (_____0___34573));
  nor2s1 ___9___500894(.DIN1 (____00___31509), .DIN2 (____0____34465),
       .Q (_________34510));
  nor2s1 ___9___500895(.DIN1 (___0____27001), .DIN2 (____0____34468),
       .Q (_________34509));
  nnd2s1 ___9___500896(.DIN1 (____0____34462), .DIN2 (_________34576),
       .Q (______0__34508));
  or2s1 ___9___500897(.DIN1 (_________41273), .DIN2 (____0____34464),
       .Q (______9__34507));
  nnd2s1 ___9__500898(.DIN1 (____0____34463), .DIN2 (__9_____30325), .Q
       (_________34506));
  nnd2s1 ___9___500899(.DIN1 (____0____34466), .DIN2 (_____9___32377),
       .Q (_________34505));
  xor2s1 ___9___500900(.DIN1 (________25536), .DIN2 (_________34497),
       .Q (______9__34523));
  dffacs1 ______________________________________________500901(.CLRB
       (reset), .CLK (clk), .DIN (____09___34478), .QN
       (___0_____40529));
  dffacs1 ______________________________________________500902(.CLRB
       (reset), .CLK (clk), .DIN (_____0___34481), .Q
       (____________________________________________21805));
  dffacs1 _______________________500903(.CLRB (reset), .CLK (clk), .DIN
       (____09___34475), .QN (_____________________21710));
  hi1s1 ___9_9_500904(.DIN (_________36778), .Q (_________35907));
  xor2s1 ___9_0_500905(.DIN1 (____0____32504), .DIN2 (____09___34476),
       .Q (_________34504));
  xor2s1 ___9_0_500906(.DIN1 (_________31627), .DIN2 (____09___34477),
       .Q (_________34503));
  nnd2s1 ___9_0_500907(.DIN1 (____0____34455), .DIN2 (_________33843),
       .Q (_________34502));
  nnd2s1 ___9___500908(.DIN1 (____0____34452), .DIN2 (_________34253),
       .Q (_________34501));
  xnr2s1 ___9__500909(.DIN1
       (_________________________________________________________________________________________22090),
       .DIN2 (______0__34499), .Q (_________34500));
  nor2s1 ___9___500910(.DIN1 (________25535), .DIN2 (_________34497),
       .Q (______9__34498));
  nor2s1 ___9___500911(.DIN1 (_________33260), .DIN2 (____0_9__34450),
       .Q (_________34549));
  hi1s1 ___9___500912(.DIN (_________34514), .Q (_____0___34569));
  nnd2s1 ___9_9_500913(.DIN1 (_________34496), .DIN2 (____09___33522),
       .Q (______9__34553));
  hi1s1 ___9_9_500914(.DIN (_________34558), .Q (______9__34543));
  xor2s1 ___9___500915(.DIN1 (____0____34411), .DIN2 (_________36858),
       .Q (_____0___34756));
  xor2s1 ___9___500916(.DIN1 (________28130), .DIN2 (____0____34467),
       .Q (_________36778));
  and2s1 ___9___500917(.DIN1 (_________34497), .DIN2 (___9____23171),
       .Q (_________34495));
  nnd2s1 ___9___500918(.DIN1 (____0____34434), .DIN2 (______0__33736),
       .Q (_________34494));
  nnd2s1 ___9___500919(.DIN1 (____0____34437), .DIN2 (____0___29370),
       .Q (_________34493));
  nnd2s1 ___9__500920(.DIN1 (____0____34439), .DIN2 (________29043), .Q
       (_________34492));
  nor2s1 ___9___500921(.DIN1 (________28857), .DIN2 (____0____34442),
       .Q (_________34491));
  and2s1 ___9___500922(.DIN1 (____0____34438), .DIN2 (__9_09__30281),
       .Q (_________34490));
  nnd2s1 ___9___500923(.DIN1 (____0_0__34441), .DIN2 (__99____30484),
       .Q (______0__34489));
  and2s1 ___9__500924(.DIN1 (____0_9__34440), .DIN2 (_____0___34487),
       .Q (_____09__34488));
  nor2s1 ___9___500925(.DIN1 (___0_____31242), .DIN2 (____0____34436),
       .Q (_____0___34486));
  nor2s1 ___9___500926(.DIN1 (_________33742), .DIN2 (____0____34435),
       .Q (_____0___34485));
  nnd2s1 ___9___500927(.DIN1 (____0____34443), .DIN2 (_________33692),
       .Q (_____0___34484));
  dffacs1 ____________________________________________9_500928(.CLRB
       (reset), .CLK (clk), .DIN (____0____34454), .Q (___0_0___40563));
  dffacs1 _____________________________________500929(.CLRB (reset),
       .CLK (clk), .DIN (____0____34457), .QN (___0_____40594));
  xor2s1 ___9___500930(.DIN1 (____0____34399), .DIN2
       (____________________________________________21832), .Q
       (_____0___34483));
  xor2s1 ___9___500931(.DIN1 (_____9___34284), .DIN2 (____0_0__34451),
       .Q (_____0___34482));
  nnd2s1 ___9___500932(.DIN1 (______9__33594), .DIN2 (____0____34430),
       .Q (_____0___34481));
  xor2s1 ___9___500933(.DIN1 (___0_____40636), .DIN2 (____0____34449),
       .Q (_____00__34480));
  nnd2s1 ___9___500934(.DIN1 (____0____34421), .DIN2 (_________34796),
       .Q (____099__34479));
  nnd2s1 ___9_9_500935(.DIN1 (____0_9__34431), .DIN2 (____0___24653),
       .Q (____09___34478));
  and2s1 ___9__500936(.DIN1 (____09___34477), .DIN2 (____0____31535),
       .Q (______9__34516));
  nor2s1 ___9___500937(.DIN1 (____9____32456), .DIN2 (____09___34476),
       .Q (_________34512));
  xor2s1 ___9___500938(.DIN1 (____0____34400), .DIN2 (______0__34897),
       .Q (_________34511));
  dffacs1 ______________________________________________500939(.CLRB
       (reset), .CLK (clk), .DIN (____0_0__34432), .QN
       (____________________________________________21774));
  xor2s1 ___9___500940(.DIN1 (____0____34398), .DIN2 (_________34983),
       .Q (_________34514));
  nnd2s1 ___9__500941(.DIN1 (____0____34412), .DIN2 (_________34163),
       .Q (____09___34475));
  or2s1 ___9___500942(.DIN1 (____09___34473), .DIN2 (____09___34472),
       .Q (____09___34474));
  or2s1 ___9___500943(.DIN1 (____090__34470), .DIN2 (____0_9__34469),
       .Q (____09___34471));
  nor2s1 ___9___500944(.DIN1 (_____0__27463), .DIN2 (____0____34467),
       .Q (____0____34468));
  nor2s1 ___9__500945(.DIN1 (_________32002), .DIN2 (____0____34409),
       .Q (____0____34466));
  nnd2s1 ___9___500946(.DIN1 (____0____34408), .DIN2 (__9900), .Q
       (____0____34465));
  dffacs2 _______________________500947(.CLRB (reset), .CLK (clk), .DIN
       (____0____34406), .Q (_____________________21682));
  nnd2s1 ___9___500948(.DIN1 (____0____34407), .DIN2 (_________31738),
       .Q (____0____34464));
  nor2s1 ___9__500949(.DIN1 (________29321), .DIN2 (____0____34410), .Q
       (____0____34463));
  and2s1 ___9_9_500950(.DIN1 (____0____34417), .DIN2 (____9____33362),
       .Q (____0____34462));
  xor2s1 ___9___500951(.DIN1 (____999__34386), .DIN2 (___90____39001),
       .Q (_________34558));
  dffacs1 ______________________________________________500952(.CLRB
       (reset), .CLK (clk), .DIN (____0____34424), .QN
       (___0__9__40530));
  xnr2s1 ___9___500953(.DIN1 (___0_____40544), .DIN2 (____0_0__34460),
       .Q (____0____34461));
  xor2s1 ___9___500954(.DIN1 (________27228), .DIN2 (____0_0__34460),
       .Q (____0_9__34459));
  xor2s1 ___9___500955(.DIN1 (____99___34378), .DIN2 (_________34141),
       .Q (____0____34458));
  nnd2s1 ___9___500956(.DIN1 (____0____34402), .DIN2 (____9_9__34346),
       .Q (____0____34457));
  xor2s1 ___9___500957(.DIN1 (____9___23779), .DIN2 (____0____34444),
       .Q (____0____34456));
  xor2s1 ___9__500958(.DIN1 (____990__34377), .DIN2 (___0_9___40554),
       .Q (____0____34455));
  nnd2s1 ___9___500959(.DIN1 (____0____34405), .DIN2 (______0__34855),
       .Q (____0____34454));
  or2s1 ___9__500960(.DIN1 (_________34644), .DIN2 (____0____34403), .Q
       (____0____34453));
  nnd2s1 ___9___500961(.DIN1 (____0_0__34451), .DIN2 (_____9___34280),
       .Q (____0____34452));
  nor2s1 ___9___500962(.DIN1 (_________33214), .DIN2 (____0____34449),
       .Q (____0_9__34450));
  or2s1 ___9___500963(.DIN1 (____0____34447), .DIN2 (____0____34446),
       .Q (____0____34448));
  nor2s1 ___9__500964(.DIN1 (____0____34401), .DIN2 (____00___34394),
       .Q (_________34496));
  xor2s1 ___9___500965(.DIN1 (________22659), .DIN2 (____0____34444),
       .Q (____0____34445));
  nor2s1 ___9___500966(.DIN1 (_________32065), .DIN2 (____00___34388),
       .Q (____0____34443));
  nnd2s1 ___9_500967(.DIN1 (____99___34382), .DIN2 (____0___27573), .Q
       (____0____34442));
  nor2s1 ___9_9_500968(.DIN1 (__9_____30418), .DIN2 (____99___34383),
       .Q (____0_0__34441));
  nor2s1 ___9_9_500969(.DIN1 (_____0___34102), .DIN2 (____00___34391),
       .Q (____0_9__34440));
  and2s1 ___9_500970(.DIN1 (____00___34390), .DIN2 (_____9__26717), .Q
       (____0____34439));
  nor2s1 ___9_0_500971(.DIN1 (_________32834), .DIN2 (____99___34385),
       .Q (____0____34438));
  nor2s1 ___9_0_500972(.DIN1 (___0_____30763), .DIN2 (____00___34393),
       .Q (____0____34437));
  nnd2s1 ___9_0_500973(.DIN1 (____00___34389), .DIN2 (_________33934),
       .Q (____0____34436));
  nnd2s1 ___9___500974(.DIN1 (____000__34387), .DIN2 (______0__31921),
       .Q (____0____34435));
  nor2s1 ___9___500975(.DIN1 (____0____33485), .DIN2 (____99___34384),
       .Q (____0____34434));
  xor2s1 ___9___500976(.DIN1 (____9____34358), .DIN2 (____0_0__38064),
       .Q (_________34497));
  dffacs1 ____0__________________500977(.CLRB (reset), .CLK (clk), .DIN
       (____00___34392), .QN (____0________________21664));
  nor2s1 ___9___500978(.DIN1 (___0_____40544), .DIN2 (____0_0__34460),
       .Q (____0____34433));
  nnd2s1 ___9___500979(.DIN1 (____99___34380), .DIN2 (___99___24162),
       .Q (____0_0__34432));
  nnd2s1 ___9___500980(.DIN1 (____99___34379), .DIN2 (______9__35170),
       .Q (____0_9__34431));
  nnd2s1 ___9___500981(.DIN1 (____9____34371), .DIN2 (inData[20]), .Q
       (____0____34430));
  xor2s1 ___9___500982(.DIN1
       (_____________________________________________21823), .DIN2
       (____0_0__34396), .Q (____0____34429));
  or2s1 ___9___500983(.DIN1 (____0____34427), .DIN2 (____0____34426),
       .Q (____0____34428));
  nnd2s1 ___9___500984(.DIN1 (____0_0__34460), .DIN2 (___0_____40544),
       .Q (____0____34425));
  nnd2s1 ___9_9_500985(.DIN1 (____9____34369), .DIN2 (____0_0__34423),
       .Q (____0____34424));
  xor2s1 ___9_500986(.DIN1 (____9____34335), .DIN2 (___0__0__40531), .Q
       (____0____34421));
  nor2s1 ___9___500987(.DIN1 (____0____34419), .DIN2 (____0____34418),
       .Q (____0____34420));
  nor2s1 ___9__500988(.DIN1 (____9_9__34376), .DIN2 (____9____34375),
       .Q (____09___34476));
  nor2s1 ___9__500989(.DIN1 (_________34240), .DIN2 (____9____34364),
       .Q (______0__34499));
  nnd2s1 ___9___500990(.DIN1 (____9____34373), .DIN2 (___0__9__30729),
       .Q (____09___34477));
  nor2s1 ___9__500991(.DIN1 (_____9___32184), .DIN2 (____9_9__34366),
       .Q (____0____34417));
  or2s1 ___9___500992(.DIN1 (_________22042), .DIN2 (____0____34444),
       .Q (____0____34416));
  nor2s1 ___9___500993(.DIN1 (___0_9___40558), .DIN2 (____0____34444),
       .Q (____0____34415));
  nnd2s1 ___9___500994(.DIN1 (____0____34444), .DIN2 (___0_9___40558),
       .Q (____0_0__34414));
  and2s1 ___9___500995(.DIN1 (____0____34444), .DIN2 (_________22042),
       .Q (____0_9__34413));
  nor2s1 ___9__500996(.DIN1 (____0____32548), .DIN2 (____9_9__34356),
       .Q (____0____34412));
  xor2s1 ___9___500997(.DIN1 (____9____34331), .DIN2 (_________36761),
       .Q (____0____34411));
  nnd2s1 ___9___500998(.DIN1 (____9____34359), .DIN2 (__99____30482),
       .Q (____0____34410));
  nor2s1 ___9___500999(.DIN1 (_________32658), .DIN2 (____9____34355),
       .Q (____0____34409));
  nor2s1 ___9_9_501000(.DIN1 (___9____29615), .DIN2 (____9____34362),
       .Q (____0____34408));
  nor2s1 ___9__501001(.DIN1 (_____9___33155), .DIN2 (____9_0__34357),
       .Q (____0____34407));
  nnd2s1 ___9___501002(.DIN1 (____9____34354), .DIN2 (_____9___31986),
       .Q (____0____34406));
  and2s1 ___9___501003(.DIN1 (____0____34444), .DIN2
       (_____________________________________________21839), .Q
       (____09___34473));
  nor2s1 ___9___501004(.DIN1
       (_____________________________________________21839), .DIN2
       (____0____34444), .Q (____09___34472));
  nor2s1 ___9___501005(.DIN1 (____9____34361), .DIN2 (____9____34360),
       .Q (____0____34467));
  nor2s1 ___9_9_501006(.DIN1 (________22420), .DIN2 (____0____34444),
       .Q (____0_9__34469));
  xor2s1 ___9__501007(.DIN1 (_____90__34277), .DIN2 (____9_0__34367),
       .Q (____0____34405));
  nor2s1 ___9_0_501008(.DIN1 (____9____34345), .DIN2 (________25831),
       .Q (____0____34403));
  nor2s1 ___9_0_501009(.DIN1 (____9____34340), .DIN2 (_________34137),
       .Q (____0____34402));
  nor2s1 ___9_0_501010(.DIN1 (_____99__37662), .DIN2 (____9____34350),
       .Q (____0____34401));
  nor2s1 ___9___501011(.DIN1 (_________33541), .DIN2 (____9____34352),
       .Q (____0____34400));
  xor2s1 ___9___501012(.DIN1 (____9____34372), .DIN2 (___0_____30886),
       .Q (____0____34399));
  xor2s1 ___9__501013(.DIN1
       (_________________________________________________________________________________________22094),
       .DIN2 (____9____34363), .Q (____0____34398));
  and2s1 ___9___501014(.DIN1 (____0_0__34396), .DIN2
       (_____________________________________________21823), .Q
       (____0____34397));
  nor2s1 ___9___501015(.DIN1
       (_____________________________________________21823), .DIN2
       (____0_0__34396), .Q (____009__34395));
  nor2s1 ___9___501016(.DIN1 (_________36556), .DIN2 (____9____34344),
       .Q (____00___34394));
  and2s1 ___9_9_501017(.DIN1 (____0_0__34396), .DIN2 (______0___22055),
       .Q (____0____34447));
  nnd2s1 ___9__501018(.DIN1 (____9_9__34336), .DIN2 (____9____34334),
       .Q (____0____34449));
  nor2s1 ___9_501019(.DIN1 (______0___22055), .DIN2 (____0_0__34396),
       .Q (____0____34446));
  nor2s1 ___9_501020(.DIN1 (________27728), .DIN2 (____9____34349), .Q
       (____0_0__34451));
  nor2s1 ___9___501021(.DIN1 (____0____32541), .DIN2 (____9____34332),
       .Q (____00___34393));
  or2s1 ___9___501022(.DIN1 (_________34207), .DIN2 (____9_0__34327),
       .Q (____00___34392));
  or2s1 ___9___501023(.DIN1 (____0____33465), .DIN2 (____9____34323),
       .Q (____00___34391));
  nor2s1 ___9___501024(.DIN1 (________28911), .DIN2 (____9____34328),
       .Q (____00___34390));
  nor2s1 ___9___501025(.DIN1 (______0__32823), .DIN2 (____9____34320),
       .Q (____00___34389));
  nnd2s1 ___9__501026(.DIN1 (____9____34324), .DIN2 (_____9___32868),
       .Q (____00___34388));
  nor2s1 ___9___501027(.DIN1 (_________33580), .DIN2 (____9____34329),
       .Q (____000__34387));
  xor2s1 ___9___501028(.DIN1 (____9_9__34306), .DIN2 (___0_____40323),
       .Q (____999__34386));
  nnd2s1 ___9___501029(.DIN1 (____9_9__34326), .DIN2 (_________33026),
       .Q (____99___34385));
  nnd2s1 ___9___501030(.DIN1 (____9____34319), .DIN2 (____0____33459),
       .Q (____99___34384));
  nor2s1 ___9___501031(.DIN1 (____0____32541), .DIN2 (____9____34325),
       .Q (____99___34383));
  nor2s1 ___9___501032(.DIN1 (________28874), .DIN2 (____9____34321),
       .Q (____99___34382));
  dffacs1 _________________________________________9____501033(.CLRB
       (reset), .CLK (clk), .DIN (____9_0__34347), .Q (_________22032));
  nor2s1 ___9_9_501034(.DIN1
       (_________________________________________9___21779), .DIN2
       (____9____34353), .Q (____090__34470));
  dffacs1 ______________________________________________501035(.CLRB
       (reset), .CLK (clk), .DIN (____9_0__34337), .Q
       (____________________________________________21764));
  dffacs1 _______________________501036(.CLRB (reset), .CLK (clk), .DIN
       (____9____34330), .QN (_____________________21703));
  nnd2s1 ___9_0_501037(.DIN1 (____9____34314), .DIN2 (_________34916),
       .Q (____99___34381));
  or2s1 ___9_0_501038(.DIN1 (______0__35050), .DIN2 (____9____34318),
       .Q (____99___34380));
  xor2s1 ___9___501039(.DIN1 (_________33568), .DIN2 (____9____34351),
       .Q (____99___34379));
  xor2s1 ___9___501040(.DIN1 (____9____34348), .DIN2 (___0_____40515),
       .Q (____99___34378));
  or2s1 ___9___501041(.DIN1 (____9____34374), .DIN2 (____9_9__34376),
       .Q (____990__34377));
  nor2s1 ___9___501042(.DIN1 (___0_9___40554), .DIN2 (____9____34374),
       .Q (____9____34375));
  or2s1 ___9___501043(.DIN1 (____9____34372), .DIN2 (___0_____30728),
       .Q (____9____34373));
  nor2s1 ___9___501044(.DIN1 (____9_0__34317), .DIN2 (____9____34370),
       .Q (____9____34371));
  nor2s1 ___9___501045(.DIN1 (___9____24106), .DIN2 (____9_9__34316),
       .Q (____9____34369));
  nor2s1 ___9_9_501046(.DIN1
       (_____________________________________________21838), .DIN2
       (____9____34368), .Q (____0____34419));
  and2s1 ___9__501047(.DIN1 (____9____34368), .DIN2
       (_____________________________________________21838), .Q
       (____0____34418));
  nor2s1 ___9___501048(.DIN1 (_________34252), .DIN2 (____9_0__34367),
       .Q (____0____34422));
  xnr2s1 ___9___501049(.DIN1 (___________9___22071), .DIN2
       (____9____34343), .Q (____0_0__34460));
  or2s1 ___9___501050(.DIN1 (____9____34365), .DIN2 (____9_0__34297),
       .Q (____9_9__34366));
  nor2s1 ___9_0_501051(.DIN1 (_________34247), .DIN2 (____9____34363),
       .Q (____9____34364));
  nnd2s1 ___9___501052(.DIN1 (____9____34299), .DIN2 (__9__0__30216),
       .Q (____9____34362));
  nor2s1 ___9___501053(.DIN1
       (_______________________________________________________________________________________),
       .DIN2 (____9____34311), .Q (____9____34361));
  nor2s1 ___9___501054(.DIN1
       (______________________________________________________________________________________0),
       .DIN2 (____9____34300), .Q (____9____34360));
  nor2s1 ___9___501055(.DIN1 (________27670), .DIN2 (____9____34303),
       .Q (____9____34359));
  nor2s1 ___9__501056(.DIN1 (_____0__22479), .DIN2 (____9____34305), .Q
       (____9____34358));
  nnd2s1 ___9___501057(.DIN1 (____9____34301), .DIN2 (___9____27806),
       .Q (____9_0__34357));
  nnd2s1 ___9___501058(.DIN1 (____9____34302), .DIN2 (_________32738),
       .Q (____9_9__34356));
  nnd2s1 ___9___501059(.DIN1 (____9_0__34307), .DIN2 (______9__32019),
       .Q (____9____34355));
  nor2s1 ___9__501060(.DIN1 (______0__32596), .DIN2 (____9____34298),
       .Q (____9____34354));
  and2s1 ___9___501061(.DIN1 (____0____35365), .DIN2
       (_____________________________________0___0_), .Q
       (____0____34426));
  nor2s1 ___9___501062(.DIN1
       (_____________________________________0___0_), .DIN2
       (____0____35365), .Q (____0____34427));
  hi1s1 ___9___501063(.DIN (____9____34353), .Q (____0____34444));
  nor2s1 ___9___501064(.DIN1 (____9____34351), .DIN2 (_________33543),
       .Q (____9____34352));
  nor2s1 ___9__501065(.DIN1 (_____9___34282), .DIN2 (____90___34294),
       .Q (____9____34350));
  and2s1 ___9___501066(.DIN1 (____9____34348), .DIN2 (________27730),
       .Q (____9____34349));
  nnd2s1 ___9___501067(.DIN1 (_____99__34286), .DIN2 (____9_9__34346),
       .Q (____9_0__34347));
  xor2s1 ___9___501068(.DIN1 (_________34256), .DIN2
       (____________________________________________21805), .Q
       (____9____34345));
  nnd2s1 ___9___501069(.DIN1 (____9____34343), .DIN2 (_____99__37662),
       .Q (____9____34344));
  nnd2s1 ___9___501070(.DIN1 (____90___34293), .DIN2 (____9____34341),
       .Q (____9____34342));
  nor2s1 ___9___501071(.DIN1 (____90___34290), .DIN2 (_________34225),
       .Q (____9____34340));
  or2s1 ___9___501072(.DIN1 (____90___34292), .DIN2 (____9____34338),
       .Q (____9____34339));
  nnd2s1 ___9___501073(.DIN1 (____90___34291), .DIN2 (________25696),
       .Q (____9_0__34337));
  nnd2s1 ___9___501074(.DIN1 (____9____34333), .DIN2 (___0__0__40531),
       .Q (____9_9__34336));
  nnd2s1 ___9___501075(.DIN1 (____9____34334), .DIN2 (____9____34333),
       .Q (____9____34335));
  nnd2s1 ___9___501076(.DIN1 (____90___34289), .DIN2 (_____0___33913),
       .Q (____0____34404));
  dffacs1 ______________________________________________501077(.CLRB
       (reset), .CLK (clk), .DIN (____90___34295), .QN
       (_________22045));
  dffacs1 ______________________________________________501078(.CLRB
       (reset), .CLK (clk), .DIN (_____9___34285), .QN
       (___0_____40546));
  nnd2s1 ___9_501079(.DIN1 (_________34272), .DIN2 (________25545), .Q
       (____9____34332));
  xor2s1 ___9___501080(.DIN1 (____9____34304), .DIN2 (_________36402),
       .Q (____9____34331));
  nnd2s1 ___9___501081(.DIN1 (_________34273), .DIN2 (__9_____30348),
       .Q (____9____34330));
  nnd2s1 ___9_9_501082(.DIN1 (_________34268), .DIN2 (____9____33393),
       .Q (____9____34329));
  nnd2s1 ___9_0_501083(.DIN1 (_________40896), .DIN2 (__99____30536),
       .Q (____9____34328));
  nnd2s1 ___9_0_501084(.DIN1 (_________34270), .DIN2 (____9_0__32391),
       .Q (____9_0__34327));
  nor2s1 ___9_0_501085(.DIN1 (__99____30500), .DIN2 (_________34271),
       .Q (____9_9__34326));
  nnd2s1 ___9__501086(.DIN1 (_________34275), .DIN2 (________28320), .Q
       (____9____34325));
  nor2s1 ___9___501087(.DIN1 (________28057), .DIN2 (_________34274),
       .Q (____9____34324));
  nnd2s1 ___9__501088(.DIN1 (______0__34267), .DIN2 (____9____34322),
       .Q (____9____34323));
  nnd2s1 ___9___501089(.DIN1 (_________34265), .DIN2 (________27960),
       .Q (____9____34321));
  nnd2s1 ___9___501090(.DIN1 (_________34264), .DIN2 (____0____32516),
       .Q (____9____34320));
  and2s1 ___9___501091(.DIN1 (_________34269), .DIN2 (____9____34322),
       .Q (____9____34319));
  hi1s1 ___9___501092(.DIN (____9____34368), .Q (____0_0__34396));
  xnr2s1 ___9___501093(.DIN1 (____9____34310), .DIN2 (___0_____40644),
       .Q (____9____34353));
  dffacs1 _____________________________________501094(.CLRB (reset),
       .CLK (clk), .DIN (____909__34296), .QN (___0_____40595));
  xor2s1 ___9___501095(.DIN1 (_____0___33914), .DIN2
       (____________________________________________21763), .Q
       (____9____34318));
  xor2s1 ___9__501096(.DIN1
       (____________________________________________21833), .DIN2
       (_____9___34278), .Q (____9_0__34317));
  nor2s1 ___9___501097(.DIN1 (____9____34315), .DIN2 (_________34254),
       .Q (____9_9__34316));
  xor2s1 ___9__501098(.DIN1 (_________34224), .DIN2 (____9____38007),
       .Q (____9____34314));
  nor2s1 ___9___501099(.DIN1 (_________34250), .DIN2 (____9____34312),
       .Q (____9____34313));
  nor2s1 ___9_501100(.DIN1 (___9____25089), .DIN2 (____9____34310), .Q
       (____9____34311));
  nor2s1 ___9_9_501101(.DIN1 (__90____29685), .DIN2 (______9__34258),
       .Q (____9____34372));
  nor2s1 ___9___501102(.DIN1 (____9____34309), .DIN2 (_________34263),
       .Q (____9____34374));
  nor2s1 ___9_9_501103(.DIN1 (_________34204), .DIN2 (_________34261),
       .Q (____9_0__34367));
  xor2s1 ___9___501104(.DIN1 (_________34221), .DIN2 (_________37884),
       .Q (____9____34363));
  xor2s1 ___9___501105(.DIN1 (_________34220), .DIN2 (___909___39065),
       .Q (____9____34368));
  hi1s1 ___9__501106(.DIN (____9____34308), .Q (____0____35365));
  and2s1 ___9___501107(.DIN1 (_________34242), .DIN2 (________27163),
       .Q (____9_0__34307));
  xor2s1 ___9___501108(.DIN1 (___________9___22071), .DIN2
       (______0__34219), .Q (____9_9__34306));
  nor2s1 ___9___501109(.DIN1 (_____0__22423), .DIN2 (____9____34304),
       .Q (____9____34305));
  or2s1 ___9_9_501110(.DIN1 (________28610), .DIN2 (______9__34248), .Q
       (____9____34303));
  and2s1 ___9_9_501111(.DIN1 (_________34241), .DIN2 (_________32639),
       .Q (____9____34302));
  nor2s1 ___9_0_501112(.DIN1 (____0___28474), .DIN2 (______0__34239),
       .Q (____9____34301));
  nor2s1 ___9__501113(.DIN1 (________25899), .DIN2 (____9____34310), .Q
       (____9____34300));
  nor2s1 ___9___501114(.DIN1 (_____9___34186), .DIN2 (_________34237),
       .Q (____9____34299));
  nor2s1 ___9___501115(.DIN1 (_________32755), .DIN2 (______9__34238),
       .Q (____9____34298));
  nnd2s1 ___9___501116(.DIN1 (_________34236), .DIN2 (_________34243),
       .Q (____9_0__34297));
  dffacs1 ____________________________________________0_(.CLRB (reset),
       .CLK (clk), .DIN (_________34260), .QN (___0_____40493));
  dffacs1 ____0__________________501117(.CLRB (reset), .CLK (clk), .DIN
       (_________34244), .QN (____0________________21666));
  or2s1 ___9___501118(.DIN1 (______9__34228), .DIN2 (_________34013),
       .Q (____909__34296));
  or2s1 ___9___501119(.DIN1 (______0__34259), .DIN2 (_________34231),
       .Q (____90___34295));
  nor2s1 ___9___501120(.DIN1 (___________9___22071), .DIN2
       (_____9___34283), .Q (____90___34294));
  xor2s1 ___9_0_501121(.DIN1 (__9__0__29975), .DIN2 (_________34257),
       .Q (____90___34293));
  xor2s1 ___9_501122(.DIN1 (___0_____40492), .DIN2 (___0_____40514), .Q
       (____90___34292));
  nnd2s1 ___9___501123(.DIN1 (_________34235), .DIN2 (_________35663),
       .Q (____90___34291));
  xor2s1 ___9___501124(.DIN1 (_____09__34200), .DIN2 (_______22208), .Q
       (____90___34290));
  or2s1 ___9___501125(.DIN1
       (____________________________________________21763), .DIN2
       (____900__34287), .Q (____90___34289));
  and2s1 ___9___501126(.DIN1 (____900__34287), .DIN2
       (____________________________________________21763), .Q
       (____90___34288));
  nor2s1 ___9__501127(.DIN1 (_________34226), .DIN2 (_________33865),
       .Q (_____99__34286));
  nnd2s1 ___9___501128(.DIN1 (_________34234), .DIN2 (____0____35361),
       .Q (_____9___34285));
  xor2s1 ___9__501129(.DIN1 (_____9___34279), .DIN2 (___0_____40514),
       .Q (_____9___34284));
  xnr2s1 ___9__501130(.DIN1 (_________36527), .DIN2 (_________40900),
       .Q (____9____34351));
  xor2s1 ___9___501131(.DIN1 (_____0___34199), .DIN2 (___9_0___39170),
       .Q (____9____34348));
  nor2s1 ___9___501132(.DIN1 (_____9___34283), .DIN2 (_____9___34282),
       .Q (____9____34343));
  nor2s1 ___9__501133(.DIN1 (_____9___34281), .DIN2 (_________40898),
       .Q (____9_9__34376));
  dffacs1 ______________________________________________501134(.CLRB
       (reset), .CLK (clk), .DIN (_________34227), .Q
       (____________________________________________21846));
  nnd2s1 ___9___501135(.DIN1 (_____9___34279), .DIN2 (_____9___34278),
       .Q (_____9___34280));
  nnd2s1 ___9___501136(.DIN1 (______9__34276), .DIN2 (_________34251),
       .Q (_____90__34277));
  nor2s1 ___9___501137(.DIN1 (_____9___33997), .DIN2 (_________34211),
       .Q (_________34275));
  nnd2s1 ___9___501138(.DIN1 (_________34216), .DIN2 (__99____30468),
       .Q (_________34274));
  nor2s1 ___9_0_501139(.DIN1 (________28635), .DIN2 (______9__34218),
       .Q (_________34273));
  nor2s1 ___9__501140(.DIN1 (___090___31413), .DIN2 (_________34213),
       .Q (_________34272));
  nnd2s1 ___9___501141(.DIN1 (_________34212), .DIN2 (___0_____31047),
       .Q (_________34271));
  nor2s1 ___9___501142(.DIN1 (_____0___33821), .DIN2 (_________34222),
       .Q (_________34270));
  nor2s1 ___9___501143(.DIN1 (____0____31589), .DIN2 (______0__34210),
       .Q (_________34269));
  nor2s1 ___9___501144(.DIN1 (__99____30463), .DIN2 (_________34215),
       .Q (_________34268));
  nor2s1 ___9___501145(.DIN1 (______9__34266), .DIN2 (______9__34209),
       .Q (______0__34267));
  nor2s1 ___9___501146(.DIN1 (___0_____30816), .DIN2 (_________34217),
       .Q (_________34265));
  nor2s1 ___9___501147(.DIN1 (_____0__29305), .DIN2 (_________34214),
       .Q (_________34264));
  xor2s1 ___9___501148(.DIN1 (______0__34201), .DIN2 (_________34061),
       .Q (____9____34308));
  nnd2s1 ___9__501149(.DIN1 (_________34230), .DIN2 (_________33783),
       .Q (____9____34333));
  dffacs1 ____0________________9_(.CLRB (reset), .CLK (clk), .DIN
       (_________34208), .QN (____0____________9_));
  hi1s1 ___9__501150(.DIN (_________40898), .Q (_________34263));
  nnd2s1 ___9_0_501151(.DIN1 (_________34202), .DIN2 (inData[0]), .Q
       (_________34262));
  nor2s1 ___9___501152(.DIN1 (_________34148), .DIN2 (_________34206),
       .Q (_________34261));
  or2s1 ___9___501153(.DIN1 (______0__34259), .DIN2 (_________34203),
       .Q (_________34260));
  and2s1 ___9___501154(.DIN1 (__90____29690), .DIN2 (_________34257),
       .Q (______9__34258));
  or2s1 ___9___501155(.DIN1 (___0_____40514), .DIN2
       (____________________________________________21833), .Q
       (_________34256));
  xor2s1 ___9__501156(.DIN1 (________28565), .DIN2 (_________35026), .Q
       (_________34255));
  xor2s1 ___9__501157(.DIN1
       (____________________________________________21791), .DIN2
       (______0__34172), .Q (_________34254));
  nnd2s1 ___9___501158(.DIN1 (______0__33640), .DIN2 (___0_____40514),
       .Q (_________34253));
  hi1s1 ___9___501159(.DIN (_________34251), .Q (_________34252));
  hi1s1 ___9___501160(.DIN (______0__34249), .Q (_________34250));
  nnd2s1 ___9___501161(.DIN1 (______0__34229), .DIN2 (_________33840),
       .Q (____9____34334));
  nnd2s1 ___9__501162(.DIN1 (_____9___34185), .DIN2 (__9_____30229), .Q
       (______9__34248));
  nor2s1 ___9___501163(.DIN1
       (_________________________________________________________________________________________22094),
       .DIN2 (_________34983), .Q (_________34247));
  nor2s1 ___9___501164(.DIN1 (_____0___34196), .DIN2 (_________34245),
       .Q (_________34246));
  nnd2s1 ___99__(.DIN1 (_____0___34197), .DIN2 (_________34243), .Q
       (_________34244));
  nor2s1 ___9___501165(.DIN1 (__9_____30335), .DIN2 (_____0___34198),
       .Q (_________34242));
  nor2s1 ___9__501166(.DIN1 (__99____30467), .DIN2 (_____00__34191), .Q
       (_________34241));
  and2s1 ___9__501167(.DIN1 (_________34983), .DIN2
       (_________________________________________________________________________________________22094),
       .Q (_________34240));
  nnd2s1 ___9___501168(.DIN1 (_____9___34187), .DIN2 (___0_____30807),
       .Q (______0__34239));
  nnd2s1 ___9___501169(.DIN1 (_____0___34192), .DIN2 (_________33000),
       .Q (______9__34238));
  nnd2s1 ___9___501170(.DIN1 (_____9___34188), .DIN2 (________28605),
       .Q (_________34237));
  nor2s1 ___99__501171(.DIN1 (_________33986), .DIN2 (_____9___34184),
       .Q (_________34236));
  nor2s1 ___9___501172(.DIN1 (_______22177), .DIN2 (_____0___34194), .Q
       (____9____34304));
  nnd2s1 ___9___501173(.DIN1 (_________34131), .DIN2 (_____99__34190),
       .Q (____9____34310));
  xor2s1 ___9___501174(.DIN1 (_________34205), .DIN2 (_________34139),
       .Q (_________34235));
  nor2s1 ___9__501175(.DIN1 (_____9__24496), .DIN2 (_____9___34182), .Q
       (_________34234));
  or2s1 ___9___501176(.DIN1 (___0_____40527), .DIN2 (_________35026),
       .Q (_________34233));
  and2s1 ___9___501177(.DIN1 (_________35026), .DIN2 (___0_____40527),
       .Q (_________34232));
  nnd2s1 ___9___501178(.DIN1 (____90___33344), .DIN2 (______9__34180),
       .Q (_________34231));
  hi1s1 ___9___501179(.DIN (______0__34229), .Q (_________34230));
  nnd2s1 ___9_9_501180(.DIN1 (_________34174), .DIN2 (__9_9___29797),
       .Q (______9__34228));
  nnd2s1 ___9___501181(.DIN1 (_________34176), .DIN2 (________26531),
       .Q (_________34227));
  nor2s1 ___9___501182(.DIN1 (_________34175), .DIN2 (_________34225),
       .Q (_________34226));
  xor2s1 ___9__501183(.DIN1 (_________34144), .DIN2 (_________34054),
       .Q (_________34224));
  nor2s1 ___9_501184(.DIN1 (___0__9__40490), .DIN2 (_________34223), .Q
       (____9____34312));
  hi1s1 ___9__501185(.DIN (___0_____40514), .Q (_____9___34278));
  nor2s1 ___9___501186(.DIN1 (_________33586), .DIN2 (_________34179),
       .Q (_____9___34283));
  nnd2s1 ___9_0_501187(.DIN1 (_________34223), .DIN2 (___0__9__40490),
       .Q (______0__34249));
  or2s1 ___9___501188(.DIN1 (___0_____40577), .DIN2 (_________34223),
       .Q (______9__34276));
  dffacs1 ______________________________________________501189(.CLRB
       (reset), .CLK (clk), .DIN (_________34177), .Q
       (____________________________________________21763));
  dffacs1 ______________________0_(.CLRB (reset), .CLK (clk), .DIN
       (_________34164), .QN (__________________0___21712));
  nnd2s1 ___99__501190(.DIN1 (______9__34161), .DIN2 (____9____34322),
       .Q (_________34222));
  nnd2s1 ___9___501191(.DIN1 (_________34170), .DIN2 (_________34032),
       .Q (_________34221));
  xor2s1 ___9___501192(.DIN1 (_________34130), .DIN2 (____9_9__38931),
       .Q (_________34220));
  xor2s1 ___9___501193(.DIN1 (_____0___34193), .DIN2 (_________36493),
       .Q (______0__34219));
  or2s1 ___9___501194(.DIN1 (__9_____29817), .DIN2 (_________34158), .Q
       (______9__34218));
  nnd2s1 ___990_(.DIN1 (_________34160), .DIN2 (______0__41062), .Q
       (_________34217));
  nor2s1 ___99_0(.DIN1 (___0_09__31127), .DIN2 (______0__34162), .Q
       (_________34216));
  or2s1 ___99__501195(.DIN1 (_________32748), .DIN2 (_________34159),
       .Q (_________34215));
  nnd2s1 ___99__501196(.DIN1 (_________34157), .DIN2 (________29253),
       .Q (_________34214));
  nnd2s1 ___99__501197(.DIN1 (______9__34152), .DIN2 (____09___31598),
       .Q (_________34213));
  nor2s1 ___99__501198(.DIN1 (__9__9__29915), .DIN2 (_________34150),
       .Q (_________34212));
  nnd2s1 ___99__501199(.DIN1 (_________34166), .DIN2 (_________33931),
       .Q (_________34211));
  nnd2s1 ___99__501200(.DIN1 (______0__34153), .DIN2 (______0__41319),
       .Q (______0__34210));
  nnd2s1 ___99_501201(.DIN1 (_________34151), .DIN2 (_____90__33327),
       .Q (______9__34209));
  or2s1 ___99__501202(.DIN1 (_________34207), .DIN2 (_________34155),
       .Q (_________34208));
  nnd2s1 ___9__501203(.DIN1 (_________34223), .DIN2 (___0_____40577),
       .Q (_________34251));
  dffacs1 _____________________0_501204(.CLRB (reset), .CLK (clk), .DIN
       (_________34165), .QN (_________________0___21702));
  nor2s1 ___9_9_501205(.DIN1
       (_____________________________________0______21757), .DIN2
       (_________34205), .Q (_________34206));
  and2s1 ___9_9_501206(.DIN1 (_________34205), .DIN2
       (_____________________________________0______21757), .Q
       (_________34204));
  nnd2s1 ___9_0_501207(.DIN1 (_________34138), .DIN2 (________24495),
       .Q (_________34203));
  and2s1 ___9___501208(.DIN1 (_____9___35464), .DIN2 (_________34147),
       .Q (_________34202));
  xor2s1 ___9___501209(.DIN1 (_________34169), .DIN2
       (_________________________________________________________________________________________22095),
       .Q (______0__34201));
  xor2s1 ___9___501210(.DIN1 (_________34173), .DIN2 (_________22032),
       .Q (_____09__34200));
  nnd2s1 ___9___501211(.DIN1 (_________34135), .DIN2 (_________34081),
       .Q (_____0___34199));
  nor2s1 ___9___501212(.DIN1 (_____0___33255), .DIN2 (_________34178),
       .Q (_____9___34282));
  xnr2s1 ___9___501213(.DIN1 (_________38242), .DIN2 (_________40902),
       .Q (______0__34229));
  nnd2s1 ___9__501214(.DIN1 (_________34142), .DIN2 (_________34087),
       .Q (_________34257));
  dffacs1 ______________________________________________501215(.CLRB
       (reset), .CLK (clk), .DIN (_________34140), .Q (___0_____40514));
  nnd2s1 ___99__501216(.DIN1 (______0__34125), .DIN2 (___99___29629),
       .Q (_____0___34198));
  nor2s1 ___999_(.DIN1 (______0__32892), .DIN2 (_________34128), .Q
       (_____0___34197));
  hi1s1 ___9___501217(.DIN (_____0___34195), .Q (_____0___34196));
  nor2s1 ___9___501218(.DIN1 (___0____22303), .DIN2 (_____0___34193),
       .Q (_____0___34194));
  nor2s1 ___99__501219(.DIN1 (___0_____30882), .DIN2 (_________34127),
       .Q (_____0___34192));
  nnd2s1 ___99__501220(.DIN1 (______0__34134), .DIN2 (________28959),
       .Q (_____00__34191));
  nnd2s1 ___9___501221(.DIN1 (_________34132), .DIN2 (_____9___34189),
       .Q (_____99__34190));
  nor2s1 ___99__501222(.DIN1 (________28225), .DIN2 (______9__34124),
       .Q (_____9___34188));
  nor2s1 ___99__501223(.DIN1 (_____9___34186), .DIN2 (_________34123),
       .Q (_____9___34187));
  nor2s1 ___99_501224(.DIN1 (___0_0___30933), .DIN2 (_________34156),
       .Q (_____9___34185));
  nnd2s1 ___99__501225(.DIN1 (_________34121), .DIN2 (__9_____30239),
       .Q (_____9___34184));
  xor2s1 ___9___501226(.DIN1 (_________34120), .DIN2
       (_________________________________________________________________________________________22091),
       .Q (_________34983));
  and2s1 ___9___501227(.DIN1 (_________36292), .DIN2 (___0_9___40559),
       .Q (_____9___34183));
  nor2s1 ___9___501228(.DIN1 (_________33596), .DIN2 (_________34115),
       .Q (_____9___34182));
  xor2s1 ___9___501229(.DIN1 (___0_____40528), .DIN2 (_____90__34089),
       .Q (_____90__34181));
  nnd2s1 ___9_9_501230(.DIN1 (________24500), .DIN2 (_________34119),
       .Q (______9__34180));
  hi1s1 ___9___501231(.DIN (_________34178), .Q (_________34179));
  and2s1 ___9___501232(.DIN1 (______9__34116), .DIN2 (_________35435),
       .Q (_________34177));
  nnd2s1 ___9___501233(.DIN1 (_________34118), .DIN2 (____9____34341),
       .Q (_________34176));
  xor2s1 ___9___501234(.DIN1 (___0_____40595), .DIN2
       (_____________________________________9______21876), .Q
       (_________34175));
  nnd2s1 ___9__501235(.DIN1 (_________34136), .DIN2 (_________34173),
       .Q (_________34174));
  nnd2s1 ___9_9_501236(.DIN1 (_________34126), .DIN2 (______9__34143),
       .Q (______0__34172));
  nor2s1 ___9___501237(.DIN1 (___0_9___40559), .DIN2 (_________36292),
       .Q (______9__34171));
  or2s1 ___9___501238(.DIN1 (_________34027), .DIN2 (_________34169),
       .Q (_________34170));
  nor2s1 ___9___501239(.DIN1 (___0_____30948), .DIN2 (_________36292),
       .Q (_________34168));
  xor2s1 ___9_9_501240(.DIN1 (_________34077), .DIN2 (_________34167),
       .Q (_________34223));
  xnr2s1 ___9___501241(.DIN1
       (_________________________________________________________________________________________22091),
       .DIN2 (_____9___34092), .Q (_________35026));
  nor2s1 ___99__501242(.DIN1 (__9_9___29892), .DIN2 (_____99__34097),
       .Q (_________34166));
  or2s1 ___99__501243(.DIN1 (__90_9__29659), .DIN2 (_________34109), .Q
       (_________34165));
  nnd2s1 ___99__501244(.DIN1 (_________34110), .DIN2 (_________34163),
       .Q (_________34164));
  nnd2s1 ___99__501245(.DIN1 (_____09__34107), .DIN2 (__9_____29981),
       .Q (______0__34162));
  nor2s1 ___99__501246(.DIN1 (_________33551), .DIN2 (_____0___34106),
       .Q (______9__34161));
  and2s1 ___99__501247(.DIN1 (_________34111), .DIN2 (___0_____30971),
       .Q (_________34160));
  nnd2s1 ___99_501248(.DIN1 (_____0___34100), .DIN2 (___0__9__30880),
       .Q (_________34159));
  nnd2s1 ___9909(.DIN1 (_____0___34104), .DIN2 (__9_____30108), .Q
       (_________34158));
  nor2s1 ___99__501249(.DIN1 (_________33849), .DIN2 (_____0___34101),
       .Q (_________34157));
  nnd2s1 ___99__501250(.DIN1 (_____0___34103), .DIN2 (_________34154),
       .Q (_________34155));
  nor2s1 ___99__501251(.DIN1 (____0____33491), .DIN2 (_____0___34105),
       .Q (______0__34153));
  nor2s1 ___99_9(.DIN1 (____0___29374), .DIN2 (_____0___34099), .Q
       (______9__34152));
  nor2s1 ___999_501252(.DIN1 (_________33553), .DIN2 (_____00__34098),
       .Q (_________34151));
  nor2s1 ___9999(.DIN1 (____0____32541), .DIN2 (______0__34108), .Q
       (_________34150));
  nnd2s1 ___9___501253(.DIN1 (_________36292), .DIN2
       (_____________________________________________21778), .Q
       (_____0___34195));
  nor2s1 ___9___501254(.DIN1
       (_____________________________________________21778), .DIN2
       (_________36292), .Q (_________34245));
  xor2s1 ___9__501255(.DIN1 (____9___23132), .DIN2 (_________34148), .Q
       (_________34149));
  xor2s1 ___9___501256(.DIN1 (___9_), .DIN2 (___09_0__40681), .Q
       (_________34147));
  nnd2s1 ___9___501257(.DIN1 (_________34145), .DIN2 (_____9___34094),
       .Q (_________34146));
  nnd2s1 ___9___501258(.DIN1 (_________34082), .DIN2 (_________34056),
       .Q (_________34144));
  nnd2s1 ___9___501259(.DIN1 (_________34141), .DIN2 (_________34084),
       .Q (_________34142));
  nnd2s1 ___9___501260(.DIN1 (_________34085), .DIN2 (_________38172),
       .Q (_________34140));
  xnr2s1 ___9___501261(.DIN1
       (_____________________________________0______21757), .DIN2
       (_________34148), .Q (_________34139));
  nnd2s1 ___9___501262(.DIN1 (_________34083), .DIN2 (______9__33955),
       .Q (_________34138));
  nor2s1 ___9__501263(.DIN1
       (_____________________________________9______21876), .DIN2
       (_________34136), .Q (_________34137));
  xor2s1 ___9___501264(.DIN1 (_________34055), .DIN2 (_________36349),
       .Q (_________34135));
  nnd2s1 ___9___501265(.DIN1 (_____9___34093), .DIN2 (_____9___34090),
       .Q (_________34178));
  nnd2s1 ___9___501266(.DIN1 (_____9___34096), .DIN2 (______0__33756),
       .Q (_________34205));
  dffacs1 ______________________________________________501267(.CLRB
       (reset), .CLK (clk), .DIN (_____9___34095), .Q (___0__0__40531));
  nor2s1 ___99__501268(.DIN1 (________27597), .DIN2 (_________34072),
       .Q (______0__34134));
  nor2s1 ___9___501269(.DIN1 (___0_____40508), .DIN2 (_________34112),
       .Q (______9__34133));
  nnd2s1 ___9___501270(.DIN1 (_________34080), .DIN2 (________22713),
       .Q (_________34132));
  nnd2s1 ___9__501271(.DIN1 (_________34129), .DIN2 (_____9___37851),
       .Q (_________34131));
  nor2s1 ___9_9_501272(.DIN1 (______0__34079), .DIN2 (_________34129),
       .Q (_________34130));
  nnd2s1 ___00__(.DIN1 (_________34076), .DIN2 (_________33172), .Q
       (_________34128));
  nnd2s1 ___99__501273(.DIN1 (_________34073), .DIN2 (__99____30506),
       .Q (_________34127));
  nor2s1 ___99__501274(.DIN1 (____9___29458), .DIN2 (_________34071),
       .Q (______0__34125));
  nnd2s1 ___99__501275(.DIN1 (_________34122), .DIN2 (______9__32204),
       .Q (______9__34124));
  nnd2s1 ___99_501276(.DIN1 (_________34122), .DIN2 (_________32357),
       .Q (_________34123));
  nor2s1 ___00__501277(.DIN1 (_________33609), .DIN2 (______0__34069),
       .Q (_________34121));
  nnd2s1 ___000_(.DIN1 (_________34122), .DIN2 (________28315), .Q
       (_________34156));
  nor2s1 ___99__501278(.DIN1 (________22368), .DIN2 (_________34075),
       .Q (_____0___34193));
  dffacs1 _______________________501279(.CLRB (reset), .CLK (clk), .DIN
       (_________34070), .QN (_____________________21681));
  xor2s1 ___99__501280(.DIN1 (_________34074), .DIN2 (_________34538),
       .Q (_________34120));
  nnd2s1 ___9__501281(.DIN1 (_________34063), .DIN2 (inData[30]), .Q
       (_________34119));
  xor2s1 ___9___501282(.DIN1 (_____9__29164), .DIN2 (_________34086),
       .Q (_________34118));
  xor2s1 ___9___501283(.DIN1 (_________33793), .DIN2 (_____90__40904),
       .Q (______9__34116));
  xor2s1 ___9___501284(.DIN1 (_________34035), .DIN2 (_________34052),
       .Q (_________34115));
  or2s1 ___9_501285(.DIN1
       (____________________________________________21851), .DIN2
       (_________34148), .Q (_________34114));
  and2s1 ___9_0_501286(.DIN1 (_________34148), .DIN2
       (____________________________________________21851), .Q
       (_________34113));
  nnd2s1 ___9___501287(.DIN1 (____9____33383), .DIN2 (_________34058),
       .Q (_________34126));
  hi1s1 ___9_9_501288(.DIN
       (_____________________________________9______21876), .Q
       (_________34173));
  nor2s1 ___990_501289(.DIN1 (_________33826), .DIN2 (______0__34060),
       .Q (_________34169));
  hi1s1 ___99__501290(.DIN (_________34112), .Q (_________36292));
  nor2s1 ___00_0(.DIN1 (__9__9__29984), .DIN2 (_________34047), .Q
       (_________34111));
  nor2s1 ___99__501291(.DIN1 (___0_____31092), .DIN2 (_________34043),
       .Q (_________34110));
  nnd2s1 ___99__501292(.DIN1 (_________34049), .DIN2 (__9_____30251),
       .Q (_________34109));
  nnd2s1 ___00__501293(.DIN1 (_________34037), .DIN2 (______0__32108),
       .Q (______0__34108));
  nor2s1 ___00__501294(.DIN1 (_____9__29218), .DIN2 (_________34045),
       .Q (_____09__34107));
  nnd2s1 ___00__501295(.DIN1 (______0__34051), .DIN2 (______0__33727),
       .Q (_____0___34106));
  nnd2s1 ___00_9(.DIN1 (_________34046), .DIN2 (____0_9__33489), .Q
       (_____0___34105));
  nor2s1 ___99__501296(.DIN1 (________29348), .DIN2 (_________34048),
       .Q (_____0___34104));
  nor2s1 ___00__501297(.DIN1 (_____0___34102), .DIN2 (_________34038),
       .Q (_____0___34103));
  or2s1 ___00__501298(.DIN1 (___0_____30986), .DIN2 (______0__34041),
       .Q (_____0___34101));
  nor2s1 ___00__501299(.DIN1 (________29264), .DIN2 (_________34044),
       .Q (_____0___34100));
  nnd2s1 ___00__501300(.DIN1 (______9__34040), .DIN2 (___0_____31156),
       .Q (_____0___34099));
  nnd2s1 ___00__501301(.DIN1 (_________34039), .DIN2 (______9__34050),
       .Q (_____00__34098));
  nnd2s1 ___00__501302(.DIN1 (_________34042), .DIN2 (_____9__29425),
       .Q (_____99__34097));
  dffacs1 ______________________________________________501303(.CLRB
       (reset), .CLK (clk), .DIN (_________34065), .QN
       (___0_____40547));
  nnd2s1 ___9_501304(.DIN1 (_____90__40904), .DIN2 (_________33758), .Q
       (_____9___34096));
  nnd2s1 ___9___501305(.DIN1 (_________34033), .DIN2 (_________37722),
       .Q (_____9___34095));
  xor2s1 ___9__501306(.DIN1 (___9___22191), .DIN2 (_____0___34006), .Q
       (_____9___34094));
  nnd2s1 ___9___501307(.DIN1 (_____9___34091), .DIN2 (_________36402),
       .Q (_____9___34093));
  and2s1 ___9_501308(.DIN1 (_____9___34091), .DIN2 (_____9___34090), .Q
       (_____9___34092));
  xor2s1 ___9___501309(.DIN1 (_________34967), .DIN2 (______9__34088),
       .Q (_____90__34089));
  or2s1 ___9_0_501310(.DIN1
       (____________________________________________21830), .DIN2
       (_________34086), .Q (_________34087));
  nor2s1 ___9_0_501311(.DIN1 (________25387), .DIN2 (_________34029),
       .Q (_________34085));
  nnd2s1 ___9__501312(.DIN1 (_________34086), .DIN2
       (____________________________________________21830), .Q
       (_________34084));
  nnd2s1 ___9___501313(.DIN1 (_________34086), .DIN2 (_________34028),
       .Q (_________34083));
  and2s1 ___9___501314(.DIN1 (______9__34030), .DIN2 (_________34081),
       .Q (_________34082));
  nnd2s1 ___9___501315(.DIN1 (____9____33378), .DIN2 (_________34057),
       .Q (______9__34143));
  dffacs1 _________________________________________9____501316(.CLRB
       (reset), .CLK (clk), .DIN (______0__34031), .Q
       (_____________________________________9______21876));
  dffacs1 _______________________501317(.CLRB (reset), .CLK (clk), .DIN
       (______9__34020), .QN (_____________________21677));
  nnd2s1 ___99_501318(.DIN1 (______9__34078), .DIN2 (________22712), .Q
       (_________34080));
  and2s1 ___99__501319(.DIN1 (______9__34078), .DIN2 (______9__34068),
       .Q (______0__34079));
  xor2s1 ___9_501320(.DIN1 (______9__34059), .DIN2 (_________34764), .Q
       (_________34077));
  nor2s1 ___0_0_(.DIN1 (____90__25948), .DIN2 (_________34017), .Q
       (_________34076));
  nor2s1 ___000_501321(.DIN1 (________22477), .DIN2 (_________34074),
       .Q (_________34075));
  nor2s1 ___00__501322(.DIN1 (___0_____30939), .DIN2 (_________34025),
       .Q (_________34073));
  nor2s1 ___00__501323(.DIN1 (_________31809), .DIN2 (______0__34021),
       .Q (_________34072));
  nnd2s1 ___00__501324(.DIN1 (_________34023), .DIN2 (_____0__28158),
       .Q (_________34071));
  nnd2s1 ___00__501325(.DIN1 (_________34022), .DIN2 (______0__32980),
       .Q (_________34070));
  nnd2s1 ___0_0_501326(.DIN1 (_________34024), .DIN2 (____0____33487),
       .Q (______0__34069));
  xor2s1 ___99__501327(.DIN1 (______0__34012), .DIN2 (______9__34981),
       .Q (_________34112));
  nor2s1 ___99_501328(.DIN1 (______9__34068), .DIN2 (______9__34078),
       .Q (_________34129));
  nnd2s1 ___00__501329(.DIN1 (_________34019), .DIN2 (_________31879),
       .Q (_________34122));
  dffacs1 _______________________501330(.CLRB (reset), .CLK (clk), .DIN
       (_________34016), .QN (_____________________21675));
  or2s1 ___9_0_501331(.DIN1 (___0_____40528), .DIN2 (_________34967),
       .Q (_________34067));
  and2s1 ___9_0_501332(.DIN1 (_________34967), .DIN2 (___0_____40528),
       .Q (_________34066));
  or2s1 ___9___501333(.DIN1 (______0__34259), .DIN2 (_____0___34010),
       .Q (_________34065));
  nnd2s1 ___9__501334(.DIN1 (_________34015), .DIN2 (_____0___34932),
       .Q (_________34064));
  xor2s1 ___9___501335(.DIN1
       (________________________________________0___21829), .DIN2
       (___9_0__23192), .Q (_________34063));
  xor2s1 ___99__501336(.DIN1 (_________34061), .DIN2 (_________37321),
       .Q (_________34062));
  and2s1 ___99_501337(.DIN1 (______9__34059), .DIN2 (_________33830),
       .Q (______0__34060));
  hi1s1 ___9___501338(.DIN (_________34057), .Q (_________34058));
  nnd2s1 ___9___501339(.DIN1 (_________34053), .DIN2 (___9_____39274),
       .Q (_________34056));
  nnd2s1 ___9_9_501340(.DIN1 (_________34054), .DIN2 (_________34053),
       .Q (_________34055));
  nor2s1 ___9___501341(.DIN1 (_____0___34008), .DIN2 (_________34052),
       .Q (______0__34117));
  dffacs1 ______________________________________________501342(.CLRB
       (reset), .CLK (clk), .DIN (_____0___34009), .Q
       (____________________________________________21762));
  xnr2s1 ___990_501343(.DIN1 (_________33730), .DIN2 (_________33974),
       .Q (_________34148));
  and2s1 ___0090(.DIN1 (_________33985), .DIN2 (______9__34050), .Q
       (______0__34051));
  nor2s1 ___00_501344(.DIN1 (___0_0___30644), .DIN2 (_____9___34002),
       .Q (_________34049));
  nor2s1 ___00__501345(.DIN1 (_________31809), .DIN2 (_____9___34000),
       .Q (_________34048));
  nnd2s1 ___00__501346(.DIN1 (_________33992), .DIN2 (____9___28644),
       .Q (_________34047));
  and2s1 ___00__501347(.DIN1 (_____9___33999), .DIN2 (__9__9__29849),
       .Q (_________34046));
  nnd2s1 ___00_501348(.DIN1 (_____9___33996), .DIN2 (________28447), .Q
       (_________34045));
  nnd2s1 ___00_501349(.DIN1 (_____99__34003), .DIN2 (________26742), .Q
       (_________34044));
  nnd2s1 ___00__501350(.DIN1 (_____9___34001), .DIN2 (___0__0__31241),
       .Q (_________34043));
  nor2s1 ___009_(.DIN1 (__9_____29847), .DIN2 (_________33991), .Q
       (_________34042));
  nnd2s1 ___009_501351(.DIN1 (_________33988), .DIN2 (_____9___31888),
       .Q (______0__34041));
  nor2s1 ___009_501352(.DIN1 (_________32815), .DIN2 (_____9___33998),
       .Q (______9__34040));
  nor2s1 ___0099(.DIN1 (______0__33984), .DIN2 (______9__33993), .Q
       (_________34039));
  nnd2s1 ___0_00(.DIN1 (_________33987), .DIN2 (_____0___33721), .Q
       (_________34038));
  nor2s1 ___0_09(.DIN1 (_________31836), .DIN2 (_________33989), .Q
       (_________34037));
  dffacs1 _____________________________________501353(.CLRB (reset),
       .CLK (clk), .DIN (_________34014), .QN (___0_____40596));
  nnd2s1 ___999_501354(.DIN1 (_________34061), .DIN2
       (_______________22073), .Q (_________34036));
  xor2s1 ___9__501355(.DIN1 (_________22047), .DIN2 (_________34034),
       .Q (_________34035));
  nor2s1 ___9___501356(.DIN1 (________24522), .DIN2 (_________33982),
       .Q (_________34033));
  nnd2s1 ___999_501357(.DIN1 (_________34061), .DIN2
       (_________________________________________________________________________________________22095),
       .Q (_________34032));
  nnd2s1 ___9___501358(.DIN1 (__9_____30112), .DIN2 (______9__33975),
       .Q (______0__34031));
  nnd2s1 ___9___501359(.DIN1 (_____00__34004), .DIN2 (___9_____39123),
       .Q (______9__34030));
  and2s1 ___9__501360(.DIN1 (_________33976), .DIN2 (____0_9__38073),
       .Q (_________34029));
  or2s1 ___9_9_501361(.DIN1
       (________________________________________0___21829), .DIN2
       (_________34026), .Q (_________34028));
  nor2s1 ___9990(.DIN1
       (_________________________________________________________________________________________22095),
       .DIN2 (_________34061), .Q (_________34027));
  xor2s1 ___9__501362(.DIN1 (_________33953), .DIN2 (______0__34897),
       .Q (_____9___34091));
  nnd2s1 ___9___501363(.DIN1 (_________33980), .DIN2 (_________33211),
       .Q (_________34057));
  nnd2s1 ___99_501364(.DIN1 (______9__33983), .DIN2 (_____09__34011),
       .Q (______9__34078));
  nnd2s1 ___990_501365(.DIN1 (_________34026), .DIN2
       (________________________________________0___21829), .Q
       (_________34086));
  nnd2s1 ___0_0_501366(.DIN1 (_________33963), .DIN2 (__9__9__29859),
       .Q (_________34025));
  and2s1 ___0___(.DIN1 (_________33972), .DIN2 (_____9___41206), .Q
       (_________34024));
  nor2s1 ___00__501367(.DIN1 (__9_____30016), .DIN2 (_________33968),
       .Q (_________34023));
  nor2s1 ___00__501368(.DIN1 (_________32138), .DIN2 (_________33970),
       .Q (_________34022));
  nnd2s1 ___00__501369(.DIN1 (_________33964), .DIN2 (____9___29007),
       .Q (______0__34021));
  nnd2s1 ___009_501370(.DIN1 (_________33969), .DIN2 (_________32015),
       .Q (______9__34020));
  nor2s1 ___0_0_501371(.DIN1 (_________41273), .DIN2 (_________33961),
       .Q (_________34019));
  or2s1 ___999_501372(.DIN1 (_______________22073), .DIN2
       (_________34061), .Q (_________34018));
  nnd2s1 ___0___501373(.DIN1 (_________33960), .DIN2 (_____9___41206),
       .Q (_________34017));
  or2s1 ___0__9(.DIN1 (___9____29568), .DIN2 (_________33959), .Q
       (_________34016));
  nor2s1 ___00__501374(.DIN1 (_____9___33906), .DIN2 (_________33971),
       .Q (_________34074));
  dffacs1 ______________________________________________501375(.CLRB
       (reset), .CLK (clk), .DIN (_________33981), .Q (___0_9___40554));
  dffacs1 ______________________________________________501376(.CLRB
       (reset), .CLK (clk), .DIN (_________33978), .Q (___0_____40515));
  dffacs1 _____________________9_501377(.CLRB (reset), .CLK (clk), .DIN
       (______9__33965), .QN (_________________9___21737));
  dffacs1 _______________________501378(.CLRB (reset), .CLK (clk), .DIN
       (______0__33966), .QN (_____________________21735));
  xor2s1 ___9_9_501379(.DIN1 (______9__33213), .DIN2 (_________33979),
       .Q (_________34015));
  or2s1 ___9_9_501380(.DIN1 (_________33952), .DIN2 (_________34013),
       .Q (_________34014));
  and2s1 ___00_501381(.DIN1 (_________33958), .DIN2 (_____09__34011),
       .Q (______0__34012));
  nnd2s1 ___9___501382(.DIN1 (______0__33956), .DIN2 (________24501),
       .Q (_____0___34010));
  nnd2s1 ___9__501383(.DIN1 (_________33954), .DIN2 (___9____24103), .Q
       (_____0___34009));
  nor2s1 ___9_9_501384(.DIN1 (_________22047), .DIN2 (___0_____31295),
       .Q (_____0___34008));
  nnd2s1 ___9_9_501385(.DIN1 (___0_____31295), .DIN2 (_________22047),
       .Q (_____0___34007));
  xor2s1 ___9_9_501386(.DIN1
       (____________________________________________21848), .DIN2
       (____________________________________________21817), .Q
       (_____0___34006));
  nnd2s1 ___00__501387(.DIN1 (_________33948), .DIN2 (_________33731),
       .Q (______9__34059));
  hi1s1 ___99__501388(.DIN (_____00__34004), .Q (_________34053));
  xor2s1 ___990_501389(.DIN1 (_________33919), .DIN2 (_________36871),
       .Q (_________34052));
  xor2s1 ___9___501390(.DIN1 (_________33922), .DIN2 (_________37864),
       .Q (_____9___34090));
  xor2s1 ___9_9_501391(.DIN1 (_________33926), .DIN2 (_________35084),
       .Q (_________34967));
  nor2s1 ___0___501392(.DIN1 (_________31716), .DIN2 (_________33930),
       .Q (_____99__34003));
  nnd2s1 ___00__501393(.DIN1 (_________33939), .DIN2 (____9___28104),
       .Q (_____9___34002));
  and2s1 ___00__501394(.DIN1 (_________33940), .DIN2 (__9__9__29945),
       .Q (_____9___34001));
  nor2s1 ___009_501395(.DIN1 (________28318), .DIN2 (_________33941),
       .Q (_____9___34000));
  nor2s1 ___0__501396(.DIN1 (____9____32434), .DIN2 (______9__33936),
       .Q (_____9___33999));
  or2s1 ___0__0(.DIN1 (_____9___33997), .DIN2 (_________33932), .Q
       (_____9___33998));
  nor2s1 ___0___501397(.DIN1 (____0____31519), .DIN2 (_________33929),
       .Q (_____9___33996));
  nor2s1 ___00__501398(.DIN1 (_____90__33994), .DIN2 (_________33944),
       .Q (_____9___33995));
  nnd2s1 ___0___501399(.DIN1 (_________33938), .DIN2 (___9____29597),
       .Q (______9__33993));
  nor2s1 ___0___501400(.DIN1 (__9_0___30086), .DIN2 (_________33990),
       .Q (_________33992));
  or2s1 ___0___501401(.DIN1 (___0_____30991), .DIN2 (_________33990),
       .Q (_________33991));
  nnd2s1 ___0___501402(.DIN1 (_________33933), .DIN2 (___9____27764),
       .Q (_________33989));
  nnd2s1 ___0___501403(.DIN1 (______0__33928), .DIN2 (________26723),
       .Q (_________33988));
  nor2s1 ___0___501404(.DIN1 (_________33986), .DIN2 (_________33935),
       .Q (_________33987));
  nor2s1 ___0___501405(.DIN1 (______0__33984), .DIN2 (______0__33937),
       .Q (_________33985));
  or2s1 ___00__501406(.DIN1 (___0_____40411), .DIN2 (_________33957),
       .Q (______9__33983));
  and2s1 ___9_501407(.DIN1 (_________33925), .DIN2 (_________34796), .Q
       (_________33982));
  nnd2s1 ___990_501408(.DIN1 (_________33920), .DIN2 (____0____35361),
       .Q (_________33981));
  nnd2s1 ___99__501409(.DIN1 (_________33212), .DIN2 (_________33979),
       .Q (_________33980));
  nnd2s1 ___99__501410(.DIN1 (______9__33927), .DIN2 (_________41256),
       .Q (_________33978));
  nnd2s1 ___9___501411(.DIN1 (_________33923), .DIN2 (______9__35170),
       .Q (_________33977));
  xor2s1 ___99__501412(.DIN1 (____09___32571), .DIN2 (_________33942),
       .Q (_________33976));
  nnd2s1 ___99__501413(.DIN1 (_________34225), .DIN2 (_____0___33915),
       .Q (______9__33975));
  xor2s1 ___000_501414(.DIN1 (_________33947), .DIN2 (_________33973),
       .Q (_________33974));
  nor2s1 ___99__501415(.DIN1
       (____________________________________________21817), .DIN2
       (_________34026), .Q (_____00__34004));
  nnd2s1 ___99__501416(.DIN1 (_________34026), .DIN2
       (____________________________________________21817), .Q
       (_________34081));
  dffacs1 ____________________________________________0_501417(.CLRB
       (reset), .CLK (clk), .DIN (_________33921), .Q
       (________________________________________0___21829));
  nor2s1 ___0___501418(.DIN1 (________28216), .DIN2 (_____0___33911),
       .Q (_________33972));
  nor2s1 ___0_0_501419(.DIN1 (___90____39001), .DIN2 (_____9___33907),
       .Q (_________33971));
  or2s1 ___0___501420(.DIN1 (____00___32480), .DIN2 (_____9___33904),
       .Q (_________33970));
  nor2s1 ___0___501421(.DIN1 (___0_9___31400), .DIN2 (_____90__33900),
       .Q (_________33969));
  nnd2s1 ___0___501422(.DIN1 (_________33962), .DIN2 (_____9___32375),
       .Q (_________33968));
  and2s1 ___0___501423(.DIN1 (_____9___33905), .DIN2 (_____9___32276),
       .Q (_________33967));
  nnd2s1 ___0___501424(.DIN1 (_____0___33912), .DIN2 (______9__32733),
       .Q (______0__33966));
  nnd2s1 ___0___501425(.DIN1 (_____9___33902), .DIN2 (_________33695),
       .Q (______9__33965));
  nor2s1 ___0___501426(.DIN1 (________27964), .DIN2 (_____9___33901),
       .Q (_________33964));
  and2s1 ___0___501427(.DIN1 (_________33962), .DIN2 (_____9___31985),
       .Q (_________33963));
  nnd2s1 ___0___501428(.DIN1 (______9__33899), .DIN2 (________28900),
       .Q (_________33961));
  nor2s1 ___0__501429(.DIN1 (________26382), .DIN2 (_________33898), .Q
       (_________33960));
  nnd2s1 ___0_9_(.DIN1 (_____9___33903), .DIN2 (___0_____30674), .Q
       (_________33959));
  xor2s1 ___00__501430(.DIN1 (_________33887), .DIN2 (_________33859),
       .Q (_________34061));
  hi1s1 ___00_501431(.DIN (_________33957), .Q (_________33958));
  nnd2s1 ___99__501432(.DIN1 (_________33891), .DIN2 (______9__33955),
       .Q (______0__33956));
  or2s1 ___99__501433(.DIN1 (______0__35050), .DIN2 (______0__33890),
       .Q (_________33954));
  nnd2s1 ___99__501434(.DIN1 (_________33893), .DIN2 (______9__33121),
       .Q (_________33953));
  nnd2s1 ___9___501435(.DIN1 (_________33888), .DIN2 (__9_9___29798),
       .Q (_________33952));
  or2s1 ___00__501436(.DIN1 (_________33950), .DIN2 (_________33949),
       .Q (_________33951));
  or2s1 ___00_501437(.DIN1 (_____09__33726), .DIN2 (_________33947), .Q
       (_________33948));
  xnr2s1 ___00__501438(.DIN1 (___0__9__40500), .DIN2 (______9__33945),
       .Q (______0__33946));
  hi1s1 ___00_501439(.DIN (_________33943), .Q (_________33944));
  or2s1 ___99__501440(.DIN1 (____9_9__32459), .DIN2 (_________33942),
       .Q (_____0___34005));
  nor2s1 ___99_501441(.DIN1 (_____0__22559), .DIN2 (_________33895), .Q
       (_________35183));
  dffacs1 ______________________________________________501442(.CLRB
       (reset), .CLK (clk), .DIN (______9__33889), .QN
       (_________22047));
  nor2s1 ___0__501443(.DIN1 (_________32305), .DIN2 (_________33878),
       .Q (_________33941));
  nor2s1 ___0___501444(.DIN1 (____0___29373), .DIN2 (_________33884),
       .Q (_________33940));
  nnd2s1 ___0__501445(.DIN1 (_________33883), .DIN2 (________25545), .Q
       (_________33939));
  nor2s1 ___0___501446(.DIN1 (__9__0__29841), .DIN2 (______0__33881),
       .Q (_________33938));
  nnd2s1 ___0___501447(.DIN1 (_________33877), .DIN2 (_________41198),
       .Q (______0__33937));
  nnd2s1 ___0___501448(.DIN1 (_________33882), .DIN2 (____9____32432),
       .Q (______9__33936));
  nnd2s1 ___0_9_501449(.DIN1 (_________33876), .DIN2 (_________33934),
       .Q (_________33935));
  nor2s1 ___0_99(.DIN1 (____9_0__33415), .DIN2 (______9__33880), .Q
       (_________33933));
  nnd2s1 ___0_0_501450(.DIN1 (_________33885), .DIN2 (_________33931),
       .Q (_________33932));
  nnd2s1 ___0___501451(.DIN1 (_____9___40906), .DIN2 (________27091),
       .Q (_________33930));
  nnd2s1 ___0___501452(.DIN1 (_____9___40906), .DIN2 (_________41154),
       .Q (_________33929));
  nor2s1 ___0__501453(.DIN1 (inData[31]), .DIN2 (_________33874), .Q
       (______0__33928));
  nnd2s1 ___0__501454(.DIN1 (_________33875), .DIN2 (__9_00__30177), .Q
       (_________33990));
  nnd2s1 ___0000(.DIN1 (_________33867), .DIN2 (_________34644), .Q
       (______9__33927));
  xor2s1 ___9_9_501455(.DIN1 (_________33845), .DIN2 (_________33316),
       .Q (_________33926));
  xor2s1 ___99__501456(.DIN1 (______9__33841), .DIN2 (_________33924),
       .Q (_________33925));
  xor2s1 ___99_501457(.DIN1 (______0__33842), .DIN2 (_________36512),
       .Q (_________33923));
  nnd2s1 ___99__501458(.DIN1 (_________33892), .DIN2 (____9____33347),
       .Q (_________33922));
  nnd2s1 ___99_501459(.DIN1 (_________33864), .DIN2 (___909__25037), .Q
       (_________33921));
  nor2s1 ___99__501460(.DIN1 (________24957), .DIN2 (_________33866),
       .Q (_________33920));
  nor2s1 ___99__501461(.DIN1 (___0_____30724), .DIN2 (______0__33871),
       .Q (_________33919));
  nnd2s1 ___00__501462(.DIN1 (______9__33945), .DIN2 (___0_____40509),
       .Q (______0__33918));
  xor2s1 ___00__501463(.DIN1 (_________33836), .DIN2 (______0__22040),
       .Q (_____09__33917));
  xor2s1 ___000_501464(.DIN1 (________22560), .DIN2 (_________33894),
       .Q (_____0___33915));
  xor2s1 ___000_501465(.DIN1 (_____0___33913), .DIN2 (_________34626),
       .Q (_____0___33914));
  nor2s1 ___00__501466(.DIN1 (_________36402), .DIN2 (_________33896),
       .Q (_________33957));
  nor2s1 ___00__501467(.DIN1 (___0_99__40560), .DIN2 (______9__33945),
       .Q (_____90__33994));
  xor2s1 ___00_501468(.DIN1 (_________33837), .DIN2 (_________35806),
       .Q (_________33979));
  dffacs1 ______________________________________________501469(.CLRB
       (reset), .CLK (clk), .DIN (_________33868), .Q
       (____________________________________________21817));
  dffacs1 _________________________________________9____501470(.CLRB
       (reset), .CLK (clk), .DIN (_________33869), .Q (___0_____40620));
  nor2s1 ___0_501471(.DIN1 (_________32254), .DIN2 (_________33856), .Q
       (_____0___33912));
  nnd2s1 ___0__501472(.DIN1 (_________33847), .DIN2 (_____0__27039), .Q
       (_____0___33911));
  and2s1 ___009_501473(.DIN1 (______9__33945), .DIN2 (___0__9__40500),
       .Q (_____00__33910));
  nor2s1 ___009_501474(.DIN1 (___0__9__40500), .DIN2 (______9__33945),
       .Q (_____99__33909));
  nor2s1 ___0_0_501475(.DIN1 (___0_____40509), .DIN2 (______9__33945),
       .Q (_____9___33908));
  nor2s1 ___0__501476(.DIN1 (________22873), .DIN2 (_________33862), .Q
       (_____9___33907));
  and2s1 ___0__501477(.DIN1 (______9__33860), .DIN2 (___90____39001),
       .Q (_____9___33906));
  nnd2s1 ___0___501478(.DIN1 (_________33854), .DIN2 (_________32140),
       .Q (_____9___33905));
  nor2s1 ___0___501479(.DIN1 (_________33897), .DIN2 (_________33858),
       .Q (_____9___33904));
  nor2s1 ___0___501480(.DIN1 (____0_0__31553), .DIN2 (_________33848),
       .Q (_____9___33903));
  nor2s1 ___0_0_501481(.DIN1 (___0__0__30899), .DIN2 (_________33855),
       .Q (_____9___33902));
  nnd2s1 ___0__501482(.DIN1 (______0__33852), .DIN2 (________27448), .Q
       (_____9___33901));
  nor2s1 ___0___501483(.DIN1 (_________32001), .DIN2 (______9__33851),
       .Q (_____90__33900));
  nor2s1 ___0___501484(.DIN1 (________29115), .DIN2 (_________33857),
       .Q (______9__33899));
  nnd2s1 ___0___501485(.DIN1 (_________33850), .DIN2 (_________33020),
       .Q (_________33898));
  nnd2s1 ___00__501486(.DIN1 (______9__33945), .DIN2 (___0_99__40560),
       .Q (_________33943));
  nor2s1 ___0___501487(.DIN1 (_________33897), .DIN2 (_____9___40908),
       .Q (_________33962));
  nnd2s1 ___00_501488(.DIN1 (_________33896), .DIN2 (_________36402),
       .Q (_____09__34011));
  dffacs1 _____________________________________501489(.CLRB (reset),
       .CLK (clk), .DIN (_________33873), .QN (___0_____40597));
  nor2s1 ___00__501490(.DIN1 (____09__22558), .DIN2 (_________33894),
       .Q (_________33895));
  hi1s1 ___99__501491(.DIN (_________33892), .Q (_________33893));
  xor2s1 ___99__501492(.DIN1 (___0_____31334), .DIN2 (______9__33870),
       .Q (_________33891));
  xor2s1 ___999_501493(.DIN1 (_________33684), .DIN2 (_________33863),
       .Q (______0__33890));
  nnd2s1 ___999_501494(.DIN1 (_________33844), .DIN2 (________26462),
       .Q (______9__33889));
  nnd2s1 ___99__501495(.DIN1 (_________34136), .DIN2 (_________33846),
       .Q (_________33888));
  xor2s1 ___0___501496(.DIN1 (______0__33861), .DIN2 (_________37199),
       .Q (_________33887));
  nor2s1 ___00__501497(.DIN1
       (_____________________________________________21777), .DIN2
       (_________33886), .Q (_________33949));
  xor2s1 ___0___501498(.DIN1 (_____9___40910), .DIN2 (___9_0___39619),
       .Q (_________33947));
  and2s1 ___00_501499(.DIN1 (_________33886), .DIN2
       (_____________________________________________21777), .Q
       (_________33950));
  nor2s1 ___00__501500(.DIN1 (_________32075), .DIN2 (_________33839),
       .Q (_________33942));
  and2s1 ___0___501501(.DIN1 (_________33879), .DIN2 (____00___32485),
       .Q (_________33885));
  nor2s1 ___0___501502(.DIN1 (_________31809), .DIN2 (_________33828),
       .Q (_________33884));
  nor2s1 ___0__501503(.DIN1 (___0_____31274), .DIN2 (_________33827),
       .Q (_________33883));
  nnd2s1 ___0__501504(.DIN1 (_________33831), .DIN2 (inData[31]), .Q
       (_________33882));
  nnd2s1 ___0___501505(.DIN1 (_________33824), .DIN2 (_________32696),
       .Q (______0__33881));
  nnd2s1 ___0___501506(.DIN1 (_________33879), .DIN2 (_________32122),
       .Q (______9__33880));
  nnd2s1 ___0___501507(.DIN1 (_________33829), .DIN2 (________27598),
       .Q (_________33878));
  and2s1 ___0___501508(.DIN1 (_________33825), .DIN2 (_____99__33716),
       .Q (_________33877));
  nor2s1 ___0___501509(.DIN1 (_________32701), .DIN2 (______0__33823),
       .Q (_________33876));
  and2s1 ___0___501510(.DIN1 (_________33879), .DIN2 (___0_____31078),
       .Q (_________33875));
  nnd2s1 ___0___501511(.DIN1 (_____0___33822), .DIN2 (_________34154),
       .Q (_________33874));
  nnd2s1 ___99_501512(.DIN1 (___0____28792), .DIN2 (_____0___33818), .Q
       (_________33873));
  xor2s1 ___0___501513(.DIN1 (_________34764), .DIN2 (_________35867),
       .Q (_________33872));
  nor2s1 ___00__501514(.DIN1 (___0_____30723), .DIN2 (______9__33870),
       .Q (______0__33871));
  nnd2s1 ___00__501515(.DIN1 (_____0___33815), .DIN2 (____9_9__34346),
       .Q (_________33869));
  nnd2s1 ___00__501516(.DIN1 (_____00__33814), .DIN2 (________23393),
       .Q (_________33868));
  xor2s1 ___00__501517(.DIN1 (_________32076), .DIN2 (_________33838),
       .Q (_________33867));
  and2s1 ___00__501518(.DIN1 (_____9___33810), .DIN2 (____9____35258),
       .Q (_________33866));
  nor2s1 ___00__501519(.DIN1 (_____9___33812), .DIN2 (_________34136),
       .Q (_________33865));
  nnd2s1 ___00__501520(.DIN1 (_____9___33811), .DIN2 (______9__33955),
       .Q (_________33864));
  or2s1 ___00_501521(.DIN1 (_________33653), .DIN2 (_________33863), .Q
       (_____0___33916));
  nnd2s1 ___000_501522(.DIN1 (_____0___33820), .DIN2 (______0__33046),
       .Q (_________33892));
  nnd2s1 ___0___501523(.DIN1 (_____0___33817), .DIN2 (________24985),
       .Q (_________33896));
  hi1s1 ___0___501524(.DIN (_________33886), .Q (______9__33945));
  nor2s1 ___0___501525(.DIN1 (________22874), .DIN2 (______0__33861),
       .Q (_________33862));
  and2s1 ___0___501526(.DIN1 (______0__33861), .DIN2 (_________33859),
       .Q (______9__33860));
  nnd2s1 ___0___501527(.DIN1 (_________33853), .DIN2 (_________32904),
       .Q (_________33858));
  nnd2s1 ___0___501528(.DIN1 (_________33801), .DIN2 (_________31725),
       .Q (_________33857));
  nnd2s1 ___0__501529(.DIN1 (_________33800), .DIN2 (_________32062),
       .Q (_________33856));
  nnd2s1 ___0___501530(.DIN1 (_________33803), .DIN2 (_________31643),
       .Q (_________33855));
  nor2s1 ___0___501531(.DIN1 (_________31866), .DIN2 (_________33802),
       .Q (_________33854));
  nor2s1 ___0__501532(.DIN1 (_________32982), .DIN2 (______9__33804),
       .Q (______0__33852));
  nnd2s1 ___0___501533(.DIN1 (_________33853), .DIN2 (_________32013),
       .Q (______9__33851));
  nor2s1 ___0_0_501534(.DIN1 (_________33849), .DIN2 (_________33798),
       .Q (_________33850));
  or2s1 ___0_0_501535(.DIN1 (________29243), .DIN2 (_________33797), .Q
       (_________33848));
  nor2s1 ___0___501536(.DIN1 (____9_0__33356), .DIN2 (_________33799),
       .Q (_________33847));
  xor2s1 ___999_501537(.DIN1
       (_____________________________________9____), .DIN2
       (___0_____40597), .Q (_________33846));
  xor2s1 ___0009(.DIN1 (_____0___33819), .DIN2 (_________36493), .Q
       (_________33845));
  nnd2s1 ___00__501538(.DIN1 (______0__33795), .DIN2 (_________33843),
       .Q (_________33844));
  xor2s1 ___00__501539(.DIN1 (______9__33755), .DIN2 (_________33763),
       .Q (______0__33842));
  xor2s1 ___00__501540(.DIN1 (_________33760), .DIN2 (_________33840),
       .Q (______9__33841));
  nor2s1 ___00__501541(.DIN1 (_________32074), .DIN2 (_________33838),
       .Q (_________33839));
  nnd2s1 ___00__501542(.DIN1 (______9__33784), .DIN2 (_________33733),
       .Q (_________33837));
  xor2s1 ___0___501543(.DIN1 (______0__41339), .DIN2 (_________33834),
       .Q (_________33836));
  xor2s1 ___0__501544(.DIN1
       (_____________________________________________21837), .DIN2
       (_________33834), .Q (_________33835));
  xor2s1 ___0___501545(.DIN1 (________25247), .DIN2 (_________33834),
       .Q (______0__33833));
  xor2s1 ___0___501546(.DIN1 (______0___22054), .DIN2 (_________33834),
       .Q (______9__33832));
  nnd2s1 ___00__501547(.DIN1 (_________33786), .DIN2 (____0____32565),
       .Q (_____0___33913));
  nor2s1 ___00__501548(.DIN1 (________22415), .DIN2 (_________33791),
       .Q (_________33894));
  or2s1 ___0_9_501549(.DIN1 (____9___25855), .DIN2 (_________33771), .Q
       (_________33831));
  nnd2s1 ___0___501550(.DIN1 (_________34764), .DIN2
       (_______________22070), .Q (_________33830));
  nor2s1 ___0__501551(.DIN1 (________29068), .DIN2 (_________33773), .Q
       (_________33829));
  nnd2s1 ___0__501552(.DIN1 (______9__33774), .DIN2 (__90_9__29688), .Q
       (_________33828));
  nnd2s1 ___0___501553(.DIN1 (_________33772), .DIN2 (___0_____31094),
       .Q (_________33827));
  nor2s1 ___0___501554(.DIN1 (_______________22070), .DIN2
       (_________34764), .Q (_________33826));
  nor2s1 ___0_501555(.DIN1 (_________33664), .DIN2 (______0__33765), .Q
       (_________33825));
  nor2s1 ___0_0_501556(.DIN1 (_________31647), .DIN2 (_________33770),
       .Q (_________33824));
  nnd2s1 ___0_501557(.DIN1 (_________33768), .DIN2 (________26292), .Q
       (______0__33823));
  nor2s1 ___0___501558(.DIN1 (_____0___33821), .DIN2 (_________33766),
       .Q (_____0___33822));
  xor2s1 ___0___501559(.DIN1 (________26189), .DIN2 (_____0___33816),
       .Q (_________33886));
  nnd2s1 ___0___501560(.DIN1 (_________33767), .DIN2 (________25545),
       .Q (_________33879));
  or2s1 ___00_501561(.DIN1 (_________33047), .DIN2 (_____0___33819), .Q
       (_____0___33820));
  nnd2s1 ___00_501562(.DIN1 (_________33650), .DIN2
       (_____________________________________9____), .Q
       (_____0___33818));
  nnd2s1 ___0_9_501563(.DIN1 (_____0___33816), .DIN2 (________26188),
       .Q (_____0___33817));
  nor2s1 ___009_501564(.DIN1 (__9_____29733), .DIN2 (_________33752),
       .Q (_____0___33815));
  nnd2s1 ___0_0_501565(.DIN1 (_________33757), .DIN2 (_____0___34932),
       .Q (_____00__33814));
  nnd2s1 ___0_0_501566(.DIN1 (_________33759), .DIN2 (_________37717),
       .Q (_____99__33813));
  xor2s1 ___0__501567(.DIN1 (____0___22645), .DIN2 (_________33790), .Q
       (_____9___33812));
  xor2s1 ___0___501568(.DIN1
       (________________________________________0___21816), .DIN2
       (_________33778), .Q (_____9___33811));
  xor2s1 ___0___501569(.DIN1 (______0__33785), .DIN2 (____0_9__32566),
       .Q (_____9___33810));
  nor2s1 ___0___501570(.DIN1 (______22150), .DIN2 (_________33834), .Q
       (_____9___33809));
  nor2s1 ___0__501571(.DIN1 (________22561), .DIN2 (_________33834), .Q
       (_____9___33808));
  xor2s1 ___0___501572(.DIN1 (_________33732), .DIN2 (______0__41289),
       .Q (______9__33870));
  nor2s1 ___00__501573(.DIN1 (_________33753), .DIN2 (______9__33764),
       .Q (_________33863));
  nor2s1 ___0___501574(.DIN1 (_________33750), .DIN2 (_____9___33806),
       .Q (_____9___33807));
  nor2s1 ___0_9_501575(.DIN1 (____9___22636), .DIN2 (_________33834),
       .Q (_____90__33805));
  nnd2s1 ___0_0_501576(.DIN1 (______0__33746), .DIN2 (_________31655),
       .Q (______9__33804));
  nnd2s1 ___0_0_501577(.DIN1 (_________33744), .DIN2 (_____90__32080),
       .Q (_________33803));
  nnd2s1 ___0___501578(.DIN1 (______9__33745), .DIN2 (_____9__26727),
       .Q (_________33802));
  nor2s1 ___0___501579(.DIN1 (________27217), .DIN2 (_________33751),
       .Q (_________33801));
  nnd2s1 ___0__501580(.DIN1 (_________33740), .DIN2 (______9__32753),
       .Q (_________33800));
  nnd2s1 ___0___501581(.DIN1 (_________33739), .DIN2 (___0____26079),
       .Q (_________33799));
  nnd2s1 ___0___501582(.DIN1 (_________33738), .DIN2 (___9____27787),
       .Q (_________33798));
  nor2s1 ___0___501583(.DIN1 (___0900), .DIN2 (_________33741), .Q
       (_________33797));
  nor2s1 ___0_9_501584(.DIN1 (________22377), .DIN2 (_________33748),
       .Q (______0__33861));
  nnd2s1 ___0__501585(.DIN1 (_________33743), .DIN2 (________27613), .Q
       (_________33853));
  dffacs1 ____0__________________501586(.CLRB (reset), .CLK (clk), .DIN
       (_________33737), .QN (____0________________21668));
  nor2s1 ___0___501587(.DIN1 (______0__22040), .DIN2 (_________33779),
       .Q (_________33796));
  xor2s1 ___0___501588(.DIN1 (_________33705), .DIN2 (___9_____39384),
       .Q (______0__33795));
  xor2s1 ___0___501589(.DIN1 (_____9__24515), .DIN2 (_________33792),
       .Q (______9__33794));
  xor2s1 ___0___501590(.DIN1
       (_____________________________________0______21756), .DIN2
       (_________33792), .Q (_________33793));
  nor2s1 ___0___501591(.DIN1 (_____9__22508), .DIN2 (_________33790),
       .Q (_________33791));
  nnd2s1 ___0__501592(.DIN1 (_________33787), .DIN2
       (____________________________________________21850), .Q
       (_________33789));
  nor2s1 ___0___501593(.DIN1
       (____________________________________________21850), .DIN2
       (_________33787), .Q (_________33788));
  nnd2s1 ___0___501594(.DIN1 (______0__33785), .DIN2 (____0____32564),
       .Q (_________33786));
  nnd2s1 ___0__501595(.DIN1 (_________33783), .DIN2 (_________33734),
       .Q (______9__33784));
  xor2s1 ___0___501596(.DIN1
       (_____________________________________________21836), .DIN2
       (_____9___33713), .Q (_________33782));
  xnr2s1 ___00__501597(.DIN1
       (____________________________________________21793), .DIN2
       (_________34709), .Q (_________33781));
  nor2s1 ___0__501598(.DIN1
       (_____________________________________________21837), .DIN2
       (_________33779), .Q (_________33780));
  xor2s1 ___0___501599(.DIN1 (_____9___33710), .DIN2 (___009___39979),
       .Q (_________33838));
  nor2s1 ___0___501600(.DIN1
       (________________________________________0___21816), .DIN2
       (_________33778), .Q (_________34054));
  nnd2s1 ___0_9_501601(.DIN1 (_________33779), .DIN2
       (_____________________________________________21765), .Q
       (_________33777));
  nor2s1 ___0_9_501602(.DIN1 (______0___22054), .DIN2 (_________33779),
       .Q (_________33776));
  or2s1 ___0_90(.DIN1
       (_____________________________________________21765), .DIN2
       (_________33779), .Q (______0__33775));
  nor2s1 ___0_9_501603(.DIN1 (________29088), .DIN2 (_____0___33724),
       .Q (______9__33774));
  or2s1 ___0_501604(.DIN1 (____9___26676), .DIN2 (_____0___33725), .Q
       (_________33773));
  nor2s1 ___0___501605(.DIN1 (____0___26782), .DIN2 (_____0___33723),
       .Q (_________33772));
  nor2s1 ___0___501606(.DIN1 (_________34207), .DIN2 (_________33728),
       .Q (_________33771));
  nor2s1 ___0___501607(.DIN1 (_________33769), .DIN2 (_____0___33719),
       .Q (_________33770));
  nor2s1 ___0___501608(.DIN1 (________29500), .DIN2 (_____00__33717),
       .Q (_________33768));
  nor2s1 ___0___501609(.DIN1 (____0____32521), .DIN2 (_____0___33718),
       .Q (_________33767));
  nnd2s1 ___0__501610(.DIN1 (_____0___33722), .DIN2 (_________32114),
       .Q (_________33766));
  nnd2s1 ___0___501611(.DIN1 (_____0___33720), .DIN2 (___0____26110),
       .Q (______0__33765));
  xor2s1 ___0_9_501612(.DIN1 (________23775), .DIN2 (_________33747),
       .Q (_________34764));
  dffacs1 _________________501613(.CLRB (reset), .CLK (clk), .DIN
       (______9__33735), .QN (______________22067));
  nor2s1 ___0__501614(.DIN1 (_________33763), .DIN2 (_________33754),
       .Q (______9__33764));
  or2s1 ___00__501615(.DIN1
       (____________________________________________21793), .DIN2
       (_________34709), .Q (_________33762));
  and2s1 ___00__501616(.DIN1 (_________34709), .DIN2
       (____________________________________________21793), .Q
       (_________33761));
  xor2s1 ___0__501617(.DIN1 (___0_____40547), .DIN2 (_____9___40912),
       .Q (_________33760));
  xor2s1 ___0___501618(.DIN1 (_________33675), .DIN2 (_________33676),
       .Q (_________33759));
  or2s1 ___0___501619(.DIN1
       (_____________________________________0______21756), .DIN2
       (_________33792), .Q (_________33758));
  xor2s1 ___0___501620(.DIN1 (_________33674), .DIN2 (_________38463),
       .Q (_________33757));
  nnd2s1 ___0___501621(.DIN1 (_________33792), .DIN2
       (_____________________________________0______21756), .Q
       (______0__33756));
  nor2s1 ___0___501622(.DIN1 (_________33754), .DIN2 (_________33753),
       .Q (______9__33755));
  nor2s1 ___0___501623(.DIN1 (_____9___33709), .DIN2 (_________34136),
       .Q (_________33752));
  dffacs1 _________________________________________9____501624(.CLRB
       (reset), .CLK (clk), .DIN (_____9___33714), .QN
       (_____________________________________9____));
  xor2s1 ___0___501625(.DIN1 (_________33685), .DIN2 (_____9___38611),
       .Q (_____0___33819));
  dffacs1 ______________________________________________501626(.CLRB
       (reset), .CLK (clk), .DIN (_____9___33715), .Q (___0_0___40564));
  dffacs1 ______________________________________________501627(.CLRB
       (reset), .CLK (clk), .DIN (_____9___33708), .QN
       (__________________________________________));
  nnd2s1 ___0___501628(.DIN1 (_________33694), .DIN2 (__9_____30024),
       .Q (_________33751));
  hi1s1 ___0_9_501629(.DIN (_________33749), .Q (_________33750));
  and2s1 ___0___501630(.DIN1 (_________33747), .DIN2 (________22466),
       .Q (_________33748));
  nor2s1 ___0__501631(.DIN1 (________28334), .DIN2 (______9__33698), .Q
       (______0__33746));
  nor2s1 ___0___501632(.DIN1 (_____0__27932), .DIN2 (______0__33699),
       .Q (______9__33745));
  nor2s1 ___0__501633(.DIN1 (____00___33437), .DIN2 (_________33697),
       .Q (_________33744));
  nor2s1 ___0___501634(.DIN1 (_________33742), .DIN2 (_________33693),
       .Q (_________33743));
  nnd2s1 ___0___501635(.DIN1 (_________33690), .DIN2 (___0_____30958),
       .Q (_________33741));
  nor2s1 ___0___501636(.DIN1 (_________31955), .DIN2 (_________33691),
       .Q (_________33740));
  nor2s1 ___0_0_501637(.DIN1 (_________31813), .DIN2 (______9__33688),
       .Q (_________33739));
  and2s1 ___0__501638(.DIN1 (_________33703), .DIN2 (____9___26582), .Q
       (_________33738));
  nnd2s1 ___0___501639(.DIN1 (______0__33689), .DIN2 (______0__33736),
       .Q (_________33737));
  nor2s1 ___0___501640(.DIN1 (_____0__28424), .DIN2 (_________33701),
       .Q (_____0___33816));
  dffacs1 _____________________________________501641(.CLRB (reset),
       .CLK (clk), .DIN (_____9___33712), .QN (__________));
  hi1s1 ___0___501642(.DIN (_________33779), .Q (_________33834));
  dffacs1 _______________________501643(.CLRB (reset), .CLK (clk), .DIN
       (_________33696), .QN (_____________________21732));
  nnd2s1 ___0___501644(.DIN1 (____0___25686), .DIN2 (_________33687),
       .Q (______9__33735));
  or2s1 ___0_9_501645(.DIN1 (___0_____40547), .DIN2 (_____9___40912),
       .Q (_________33734));
  nnd2s1 ___0_9_501646(.DIN1 (_____9___40912), .DIN2 (___0_____40547),
       .Q (_________33733));
  nor2s1 ___0___501647(.DIN1 (_________33642), .DIN2 (_________33677),
       .Q (_________33732));
  or2s1 ___0_9_501648(.DIN1 (_______________22069), .DIN2
       (_________33730), .Q (_________33731));
  hi1s1 ___0_0_501649(.DIN (_________33792), .Q (_________33787));
  nor2s1 ___0_0_501650(.DIN1 (________22589), .DIN2 (_________33682),
       .Q (_________33790));
  xor2s1 ___0___501651(.DIN1 (______9__33658), .DIN2 (_________33729),
       .Q (______0__33785));
  nnd2s1 ___0___501652(.DIN1 (_________33730), .DIN2 (_________36762),
       .Q (_________33749));
  dffacs1 ____________________________________________0_501653(.CLRB
       (reset), .CLK (clk), .DIN (______9__33678), .QN
       (________________________________________0___21816));
  xor2s1 ___0_9_501654(.DIN1 (______9__33639), .DIN2 (_________36291),
       .Q (_________33779));
  nnd2s1 ___0_0_501655(.DIN1 (_________33661), .DIN2 (______0__33727),
       .Q (_________33728));
  and2s1 ___0___501656(.DIN1 (_________33730), .DIN2
       (_______________22069), .Q (_____09__33726));
  nnd2s1 ___0___501657(.DIN1 (______9__33668), .DIN2 (________26744),
       .Q (_____0___33725));
  nnd2s1 ___0__501658(.DIN1 (_________33667), .DIN2 (___90___28650), .Q
       (_____0___33724));
  nnd2s1 ___0___501659(.DIN1 (_________33666), .DIN2 (_____9__28100),
       .Q (_____0___33723));
  and2s1 ___0_0_501660(.DIN1 (_________33663), .DIN2 (_____0___33721),
       .Q (_____0___33722));
  nor2s1 ___0___501661(.DIN1 (________25351), .DIN2 (_________33660),
       .Q (_____0___33720));
  nnd2s1 ___0_501662(.DIN1 (_________33662), .DIN2 (_________33570), .Q
       (_____0___33719));
  nnd2s1 ___0__501663(.DIN1 (______0__33659), .DIN2 (___0_____31182),
       .Q (_____0___33718));
  nnd2s1 ___0___501664(.DIN1 (_________33665), .DIN2 (_____99__33716),
       .Q (_____00__33717));
  nor2s1 ___0___501665(.DIN1 (_________36762), .DIN2 (_________33730),
       .Q (_____9___33806));
  dffacs1 ______________________________________________501666(.CLRB
       (reset), .CLK (clk), .DIN (______0__33679), .QN
       (_________22046));
  nnd2s1 ___0___501667(.DIN1 (_________33652), .DIN2 (____0____35361),
       .Q (_____9___33715));
  nnd2s1 ___0___501668(.DIN1 (___9____28682), .DIN2 (_________33646),
       .Q (_____9___33714));
  xnr2s1 ___0___501669(.DIN1 (_________38666), .DIN2 (_________35162),
       .Q (_____9___33713));
  or2s1 ___0___501670(.DIN1 (_________33651), .DIN2 (________28354), .Q
       (_____9___33712));
  xor2s1 ___0___501671(.DIN1 (________26156), .DIN2 (_________35162),
       .Q (_____9___33711));
  nor2s1 ___0___501672(.DIN1 (____9_0__32460), .DIN2 (_________33645),
       .Q (_____9___33710));
  xor2s1 ___0_501673(.DIN1 (________22591), .DIN2 (_________33681), .Q
       (_____9___33709));
  nnd2s1 ___0___501674(.DIN1 (_________33656), .DIN2 (________23553),
       .Q (_____9___33708));
  nnd2s1 ___0___501675(.DIN1 (________23552), .DIN2 (______9__33648),
       .Q (_____90__33707));
  and2s1 ___0___501676(.DIN1 (_________33647), .DIN2 (____0_9__38073),
       .Q (______9__33706));
  xor2s1 ___0___501677(.DIN1 (_____9___33615), .DIN2 (_____9___34281),
       .Q (_________33705));
  nor2s1 ___0_0_501678(.DIN1
       (_____________________________________0______21755), .DIN2
       (_________33704), .Q (_________33754));
  and2s1 ___0_0_501679(.DIN1 (_________33704), .DIN2
       (_____________________________________0______21755), .Q
       (_________33753));
  xnr2s1 ___0___501680(.DIN1
       (_________________________________________________________________________________________22090),
       .DIN2 (_____0___33626), .Q (_________34709));
  xor2s1 ___0___501681(.DIN1 (_____9___33618), .DIN2 (____0___28555),
       .Q (_________33792));
  nor2s1 ___0__501682(.DIN1 (_____9___31792), .DIN2 (_________33643),
       .Q (_________33703));
  xnr2s1 ___0___501683(.DIN1 (_________38395), .DIN2 (_________33602),
       .Q (_________33701));
  xor2s1 ___0_501684(.DIN1 (________23051), .DIN2 (_________35162), .Q
       (_________33700));
  nnd2s1 ___0___501685(.DIN1 (_________33636), .DIN2 (___0__9__31280),
       .Q (______0__33699));
  nnd2s1 ___0___501686(.DIN1 (_________33635), .DIN2 (___09____31438),
       .Q (______9__33698));
  nnd2s1 ___0___501687(.DIN1 (_________33634), .DIN2 (______9__33575),
       .Q (_________33697));
  nnd2s1 ___0___501688(.DIN1 (_________33638), .DIN2 (_________33695),
       .Q (_________33696));
  nor2s1 ___0___501689(.DIN1 (________27158), .DIN2 (_________33633),
       .Q (_________33694));
  nnd2s1 ___0___501690(.DIN1 (_________33637), .DIN2 (_________33692),
       .Q (_________33693));
  nnd2s1 ___0___501691(.DIN1 (_________33632), .DIN2 (_________32078),
       .Q (_________33691));
  nor2s1 ___0___501692(.DIN1 (______0__31903), .DIN2 (_________33631),
       .Q (_________33690));
  and2s1 ___0___501693(.DIN1 (______0__33630), .DIN2 (____0____33493),
       .Q (______0__33689));
  and2s1 ___0___501694(.DIN1 (_____0___33629), .DIN2 (_____0___34487),
       .Q (______9__33688));
  xor2s1 ___0_9_501695(.DIN1 (_________33611), .DIN2 (_________36928),
       .Q (_________33747));
  or2s1 ___0___501696(.DIN1 (_____0___33628), .DIN2 (_________33686),
       .Q (_________33687));
  nnd2s1 ___0___501697(.DIN1 (_____0___33627), .DIN2 (_____0___33625),
       .Q (_________33685));
  xor2s1 ___0___501698(.DIN1 (___0_____40578), .DIN2 (_________33683),
       .Q (_________33684));
  nor2s1 ___0___501699(.DIN1 (________22590), .DIN2 (_________33681),
       .Q (_________33682));
  nor2s1 ___0___501700(.DIN1 (_________22039), .DIN2 (_________35162),
       .Q (_________33680));
  nnd2s1 ___0___501701(.DIN1 (_____9___33620), .DIN2 (____0____35361),
       .Q (______0__33679));
  nor2s1 ___0___501702(.DIN1 (____0____33482), .DIN2 (_____99__33621),
       .Q (______9__33678));
  nor2s1 ___0___501703(.DIN1 (_____9___33619), .DIN2 (_________33676),
       .Q (_________33677));
  xor2s1 ___0___501704(.DIN1 (_________33641), .DIN2 (_____9___34279),
       .Q (_________33675));
  xor2s1 ___0_9_501705(.DIN1 (____9____32461), .DIN2 (_________33644),
       .Q (_________33674));
  nor2s1 ___0_0_501706(.DIN1 (______0_), .DIN2 (_________35162), .Q
       (_________33673));
  and2s1 ___0_0_501707(.DIN1 (_________35162), .DIN2 (______0_), .Q
       (_________33672));
  nor2s1 ___0___501708(.DIN1
       (_____________________________________________21836), .DIN2
       (_________35162), .Q (_________33671));
  nnd2s1 ___0___501709(.DIN1 (_________35162), .DIN2
       (_____________________________________________21836), .Q
       (_________33670));
  and2s1 ___0___501710(.DIN1 (_________35162), .DIN2 (_________22039),
       .Q (______0__33669));
  nor2s1 ___0_0_501711(.DIN1 (______9__33267), .DIN2 (_____90__33612),
       .Q (______9__33668));
  nor2s1 ___0_0_501712(.DIN1 (_________33030), .DIN2 (_____00__40914),
       .Q (_________33667));
  nor2s1 ___0___501713(.DIN1 (___9_0__28655), .DIN2 (_____0___40916),
       .Q (_________33666));
  nor2s1 ___0___501714(.DIN1 (_________33664), .DIN2 (_________33607),
       .Q (_________33665));
  nor2s1 ___0__501715(.DIN1 (___00____30625), .DIN2 (_________33605),
       .Q (_________33663));
  nor2s1 ___0___501716(.DIN1 (_________33106), .DIN2 (_________33608),
       .Q (_________33662));
  nor2s1 ___0___501717(.DIN1 (_________33549), .DIN2 (_________33610),
       .Q (_________33661));
  nnd2s1 ___0__501718(.DIN1 (_________33603), .DIN2 (_________32160),
       .Q (_________33660));
  nor2s1 ___0___501719(.DIN1 (________28600), .DIN2 (______9__33604),
       .Q (______0__33659));
  xor2s1 ___0_501720(.DIN1 (_________33583), .DIN2
       (_________________________________________________________________________________________22094),
       .Q (_________33730));
  dffacs1 ____0_________________0_(.CLRB (reset), .CLK (clk), .DIN
       (_________33606), .QN (____0_____________0_));
  nnd2s1 ___0__501721(.DIN1 (_________33590), .DIN2 (_____09__32097),
       .Q (______9__33658));
  and2s1 ___0___501722(.DIN1 (_________33598), .DIN2 (____0_9__38073),
       .Q (_________33657));
  nnd2s1 ___0___501723(.DIN1 (_________33599), .DIN2 (_________34796),
       .Q (_________33656));
  nnd2s1 ___0___501724(.DIN1 (_________33683), .DIN2 (___0__0__40491),
       .Q (_________33655));
  nor2s1 ___0___501725(.DIN1 (___0__0__40491), .DIN2 (_________33683),
       .Q (_________33654));
  nor2s1 ___0___501726(.DIN1 (___0_____40578), .DIN2 (_________33683),
       .Q (_________33653));
  nor2s1 ___0__501727(.DIN1 (________24579), .DIN2 (_________33597), .Q
       (_________33652));
  nor2s1 ___0__501728(.DIN1 (______0__33595), .DIN2 (_________33650),
       .Q (_________33651));
  and2s1 ___0___501729(.DIN1 (_________33683), .DIN2 (___0_____40578),
       .Q (______0__33649));
  xor2s1 ___0___501730(.DIN1 (________22427), .DIN2
       (____________________________________________21773), .Q
       (______9__33648));
  xor2s1 ___0___501731(.DIN1 (_________32618), .DIN2 (_____0___33624),
       .Q (_________33647));
  nnd2s1 ___0__501732(.DIN1 (_________33650), .DIN2 (_________33593),
       .Q (_________33646));
  nor2s1 ___0__501733(.DIN1 (_________33644), .DIN2 (_________32318),
       .Q (_________33645));
  xor2s1 ___0__501734(.DIN1 (_________33561), .DIN2 (_________36301),
       .Q (_________33704));
  nor2s1 ___0___501735(.DIN1 (___0900), .DIN2 (_________33572), .Q
       (_________33643));
  nor2s1 ___0__501736(.DIN1 (_________33641), .DIN2 (______0__33640),
       .Q (_________33642));
  xor2s1 ___0_9_501737(.DIN1 (_________33601), .DIN2 (________28425),
       .Q (______9__33639));
  nor2s1 ___0___501738(.DIN1 (_________32268), .DIN2 (_________33579),
       .Q (_________33638));
  nor2s1 ___0__501739(.DIN1 (_________31906), .DIN2 (_________33581),
       .Q (_________33637));
  nor2s1 ___0___501740(.DIN1 (___0_____31088), .DIN2 (_________33582),
       .Q (_________33636));
  nor2s1 ___0___501741(.DIN1 (_________32836), .DIN2 (_____0___40918),
       .Q (_________33635));
  nor2s1 ___0___501742(.DIN1 (_____9___33059), .DIN2 (_________33578),
       .Q (_________33634));
  nnd2s1 ___0___501743(.DIN1 (______0__33585), .DIN2 (___9____27784),
       .Q (_________33633));
  nor2s1 ___0___501744(.DIN1 (______9__32852), .DIN2 (______0__33576),
       .Q (_________33632));
  nnd2s1 ___0_0_501745(.DIN1 (_________33573), .DIN2 (________29090),
       .Q (_________33631));
  and2s1 ___0___501746(.DIN1 (_________33574), .DIN2 (_________41198),
       .Q (______0__33630));
  nor2s1 ___0__501747(.DIN1 (________26605), .DIN2 (_________33571), .Q
       (_____0___33629));
  nor2s1 ___0_9_501748(.DIN1 (_________33587), .DIN2 (_____9___33616),
       .Q (_________33702));
  xor2s1 ___0___501749(.DIN1 (______0__33538), .DIN2 (________22410),
       .Q (_____0___33628));
  xor2s1 ___0___501750(.DIN1 (_________33540), .DIN2 (________22381),
       .Q (_____0___33627));
  nnd2s1 ___0___501751(.DIN1 (_________33569), .DIN2 (_____0___33625),
       .Q (_____0___33626));
  nor2s1 ___0___501752(.DIN1 (_____00__33622), .DIN2 (______9__33565),
       .Q (_____0___33623));
  xor2s1 ___0__501753(.DIN1 (___0_____40533), .DIN2 (____9____33371),
       .Q (_____99__33621));
  nor2s1 ___0___501754(.DIN1 (________24583), .DIN2 (_________33559),
       .Q (_____9___33620));
  nor2s1 ___0__501755(.DIN1
       (____________________________________________21773), .DIN2
       (_____9___34279), .Q (_____9___33619));
  xor2s1 ___0___501756(.DIN1 (_____9___33617), .DIN2 (_____9___33616),
       .Q (_____9___33618));
  xor2s1 ___0___501757(.DIN1
       (____________________________________________21761), .DIN2
       (_________33589), .Q (_____9___33615));
  xor2s1 ___0___501758(.DIN1 (___0_00__40561), .DIN2 (____00___35294),
       .Q (_____9___33614));
  nor2s1 ___0___501759(.DIN1 (____0_0__33480), .DIN2 (_________33560),
       .Q (_________33681));
  xnr2s1 ___0_0_501760(.DIN1 (_________36556), .DIN2 (_____0___33532),
       .Q (_________35162));
  xor2s1 ___0__501761(.DIN1 (___9____23141), .DIN2 (____00___35294), .Q
       (_____9___33613));
  nnd2s1 ___0___501762(.DIN1 (_________33557), .DIN2 (____9___27296),
       .Q (_____90__33612));
  nor2s1 ___0__501763(.DIN1 (____9___22448), .DIN2 (______9__33556), .Q
       (_________33611));
  or2s1 ___0_9_501764(.DIN1 (_________33609), .DIN2 (_________33554),
       .Q (_________33610));
  nnd2s1 ___0_501765(.DIN1 (_________33550), .DIN2 (______0__33727), .Q
       (_________33608));
  or2s1 ___0_0_501766(.DIN1 (________26290), .DIN2 (_________33558), .Q
       (_________33607));
  nnd2s1 ___0__501767(.DIN1 (_________33552), .DIN2 (___0_____31034),
       .Q (_________33606));
  nnd2s1 ___0__501768(.DIN1 (______0__33548), .DIN2 (______0__41319),
       .Q (_________33605));
  nnd2s1 ___0___501769(.DIN1 (_________33546), .DIN2 (_________31811),
       .Q (______9__33604));
  nnd2s1 ___0___501770(.DIN1 (______9__33547), .DIN2 (_________33016),
       .Q (_________33603));
  nor2s1 ___0___501771(.DIN1 (_____9__28423), .DIN2 (_________33601),
       .Q (_________33602));
  dffacs1 ___________________________________0_(.CLRB (reset), .CLK
       (clk), .DIN (_________33562), .QN (_______________0));
  nnd2s1 ___0___501772(.DIN1 (____00___35294), .DIN2 (_________33591),
       .Q (_________33600));
  xor2s1 ___0__501773(.DIN1 (____0_9__33519), .DIN2 (_________36871),
       .Q (_________33599));
  xor2s1 ___0___501774(.DIN1 (____090__33520), .DIN2 (____9____37036),
       .Q (_________33598));
  nor2s1 ___0___501775(.DIN1 (_________33596), .DIN2 (_____09__33537),
       .Q (_________33597));
  nnd2s1 ___0___501776(.DIN1 (________27054), .DIN2 (_____0___33535),
       .Q (______0__33595));
  nnd2s1 ___0___501777(.DIN1 (_____0___33536), .DIN2 (____0_9__38073),
       .Q (______9__33594));
  xor2s1 ___0__501778(.DIN1 (____09___33521), .DIN2 (___0_____40308),
       .Q (_________33593));
  nor2s1 ___0___501779(.DIN1 (_________33591), .DIN2 (____00___35294),
       .Q (_________33592));
  or2s1 ___0___501780(.DIN1 (______0__32098), .DIN2 (_________33589),
       .Q (_________33590));
  nnd2s1 ___0___501781(.DIN1 (____00___35294), .DIN2 (___9____23140),
       .Q (_________33588));
  xnr2s1 ___0___501782(.DIN1 (_________38533), .DIN2 (____0____33504),
       .Q (_________33587));
  nnd2s1 ___0_501783(.DIN1 (____9____33400), .DIN2 (___0_____40533), .Q
       (_________33644));
  hi1s1 ___0___501784(.DIN
       (____________________________________________21773), .Q
       (_________33641));
  xor2s1 ___0__501785(.DIN1 (____0____33508), .DIN2 (_________33586),
       .Q (_________33683));
  nor2s1 ___0___501786(.DIN1 (______0__32214), .DIN2 (____09___33526),
       .Q (______0__33585));
  nnd2s1 ___0___501787(.DIN1 (____00___35294), .DIN2 (_____9___22050),
       .Q (______9__33584));
  xor2s1 ___0_501788(.DIN1 (_________33555), .DIN2 (_________34167), .Q
       (_________33583));
  nnd2s1 ___0_9_501789(.DIN1 (_____0___33530), .DIN2 (________28876),
       .Q (_________33582));
  or2s1 ___0_0_501790(.DIN1 (_________33580), .DIN2 (____09___33528),
       .Q (_________33581));
  nnd2s1 ___0_501791(.DIN1 (____09___33527), .DIN2 (______0__32754), .Q
       (_________33579));
  nnd2s1 ___0___501792(.DIN1 (_____0___40920), .DIN2 (___0__9__31299),
       .Q (_________33578));
  nor2s1 ___0__501793(.DIN1 (_____9___22050), .DIN2 (____00___35294),
       .Q (_________33577));
  nnd2s1 ___0__501794(.DIN1 (_____00__33529), .DIN2 (______9__33575),
       .Q (______0__33576));
  nor2s1 ___0___501795(.DIN1 (_____0__29262), .DIN2 (____09___33524),
       .Q (_________33574));
  nor2s1 ___0__501796(.DIN1 (___0__0__31061), .DIN2 (____09___33525),
       .Q (_________33573));
  nnd2s1 ___0___501797(.DIN1 (_____0___33531), .DIN2 (____0____31527),
       .Q (_________33572));
  nnd2s1 ___0__501798(.DIN1 (_____0___33533), .DIN2 (_________33570),
       .Q (_________33571));
  dffacs1 ______________________________________________501799(.CLRB
       (reset), .CLK (clk), .DIN (_________33545), .QN
       (____________________________________________21804));
  xnr2s1 ___0___501800(.DIN1 (_________38842), .DIN2 (_________33539),
       .Q (_________33569));
  xor2s1 ___0___501801(.DIN1 (_________33542), .DIN2 (___0____23284),
       .Q (_________33568));
  nnd2s1 ___0__501802(.DIN1 (____09___33523), .DIN2 (___0__9__40510),
       .Q (_________33567));
  xor2s1 ___0___501803(.DIN1 (___0_____40492), .DIN2 (_________33763),
       .Q (______0__33566));
  hi1s1 ___0___501804(.DIN (_________33564), .Q (______9__33565));
  nor2s1 ___0___501805(.DIN1 (___0_____40492), .DIN2 (____0____33514),
       .Q (_________33563));
  nnd2s1 ___0___501806(.DIN1 (___0____28819), .DIN2 (____0____33513),
       .Q (_________33562));
  nnd2s1 ___0__501807(.DIN1 (____0____33518), .DIN2 (____9____33382),
       .Q (_________33561));
  nor2s1 ___0___501808(.DIN1 (____0_0__33510), .DIN2 (_________33322),
       .Q (_________33560));
  nor2s1 ___0___501809(.DIN1 (_________33596), .DIN2 (____0____33511),
       .Q (_________33559));
  nor2s1 ___0___501810(.DIN1 (_________32033), .DIN2 (____0____33516),
       .Q (_____0___33624));
  xor2s1 ___0___501811(.DIN1 (____0____33484), .DIN2 (_________36871),
       .Q (_____0___33625));
  dffacs1 ______________________________________________501812(.CLRB
       (reset), .CLK (clk), .DIN (____0____33512), .Q
       (____________________________________________21773));
  nnd2s1 ___0___501813(.DIN1 (____0____33497), .DIN2 (_________32354),
       .Q (_________33558));
  nor2s1 ___0_9_501814(.DIN1 (_________32750), .DIN2 (____0____33502),
       .Q (_________33557));
  nor2s1 ___0_0_501815(.DIN1 (__9___22169), .DIN2 (_________33555), .Q
       (______9__33556));
  or2s1 ___0__501816(.DIN1 (_________33553), .DIN2 (____0____33488), .Q
       (_________33554));
  or2s1 ___0___501817(.DIN1 (_________33551), .DIN2 (____0____33494),
       .Q (_________33552));
  nor2s1 ___0___501818(.DIN1 (_________33549), .DIN2 (____0_0__33490),
       .Q (_________33550));
  nor2s1 ___0___501819(.DIN1 (___0_9___31401), .DIN2 (____0____33492),
       .Q (______0__33548));
  nor2s1 ___0___501820(.DIN1 (____0____33496), .DIN2 (____0____33486),
       .Q (______9__33547));
  nor2s1 ___0___501821(.DIN1 (______9__32117), .DIN2 (____0____33495),
       .Q (_________33546));
  nnd2s1 ___0_9_501822(.DIN1 (____0_9__33499), .DIN2 (________22426),
       .Q (_________33601));
  dffacs1 _________________________________________9____501823(.CLRB
       (reset), .CLK (clk), .DIN (____0____33506), .Q (___0_99__40460));
  nnd2s1 ___0___501824(.DIN1 (____0____33481), .DIN2 (________27137),
       .Q (_________33545));
  nor2s1 ___0___501825(.DIN1 (_____22118), .DIN2 (_________33763), .Q
       (_________33544));
  and2s1 ___0___501826(.DIN1 (_________33542), .DIN2
       (____________________________________________21792), .Q
       (_________33543));
  nor2s1 ___0___501827(.DIN1
       (____________________________________________21792), .DIN2
       (_________33542), .Q (_________33541));
  nor2s1 ___0__501828(.DIN1
       (_________________________________________________________________________________________22090),
       .DIN2 (_________33539), .Q (_________33540));
  xor2s1 ___0_9_501829(.DIN1 (____0_9__33509), .DIN2 (___0_____40479),
       .Q (______0__33538));
  xor2s1 ___0_9_501830(.DIN1 (____0____33517), .DIN2 (____9_0__33405),
       .Q (_____09__33537));
  xor2s1 ___0__501831(.DIN1 (_________32102), .DIN2 (____0____33515),
       .Q (_____0___33536));
  xor2s1 ___0_501832(.DIN1 (___0__9__40628), .DIN2 (_______________0),
       .Q (_____0___33535));
  nnd2s1 ___0__501833(.DIN1 (____0____33477), .DIN2 (_________31720),
       .Q (_________33589));
  dffacs1 ____________________________________________0_501834(.CLRB
       (reset), .CLK (clk), .DIN (____0____33483), .QN
       (___0_____40533));
  nnd2s1 ___0___501835(.DIN1 (_________33542), .DIN2 (_____0___33534),
       .Q (_________33564));
  nor2s1 ___0___501836(.DIN1 (_____0___33534), .DIN2 (_________33542),
       .Q (_____00__33622));
  nor2s1 ___0___501837(.DIN1 (_________31958), .DIN2 (____0____33468),
       .Q (_____0___33533));
  xor2s1 ___0___501838(.DIN1 (____0____33498), .DIN2
       (_________________________________________________________________________________________22094),
       .Q (_____0___33532));
  and2s1 ___0_0_501839(.DIN1 (____0____33466), .DIN2 (_____0___33721),
       .Q (_____0___33531));
  nor2s1 ___0___501840(.DIN1 (________28875), .DIN2 (____0____33469),
       .Q (_____0___33530));
  nor2s1 ___0___501841(.DIN1 (_________32931), .DIN2 (____0_0__33471),
       .Q (_____00__33529));
  nnd2s1 ___0__501842(.DIN1 (____0____33473), .DIN2 (_________32239),
       .Q (____09___33528));
  nnd2s1 ___0___501843(.DIN1 (____0_9__33470), .DIN2 (___9____26906),
       .Q (____09___33527));
  nnd2s1 ___0___501844(.DIN1 (____0____33472), .DIN2 (________29525),
       .Q (____09___33526));
  nnd2s1 ___0___501845(.DIN1 (____0____33464), .DIN2 (_________31933),
       .Q (____09___33525));
  or2s1 ___0_501846(.DIN1 (___90___29559), .DIN2 (____0____33467), .Q
       (____09___33524));
  nor2s1 ___0___501847(.DIN1 (_________33266), .DIN2 (____0_9__33479),
       .Q (_____9___33616));
  hi1s1 ___0___501848(.DIN (____09___33523), .Q (____00___35294));
  or2s1 ___0___501849(.DIN1 (_________36761), .DIN2 (_____9___33617),
       .Q (____09___33522));
  xor2s1 ___0_9_501850(.DIN1 (_________33323), .DIN2
       (____________________________________________21865), .Q
       (____09___33521));
  xor2s1 ___0_9_501851(.DIN1 (____0____33444), .DIN2 (_________34141),
       .Q (____090__33520));
  xor2s1 ___0_9_501852(.DIN1 (____0____33445), .DIN2 (_____0___33257),
       .Q (____0_9__33519));
  or2s1 ___0_0_501853(.DIN1 (____9____33381), .DIN2 (____0____33517),
       .Q (____0____33518));
  nor2s1 ___0___501854(.DIN1 (______0__32030), .DIN2 (____0____33515),
       .Q (____0____33516));
  hi1s1 ___0___501855(.DIN (_________33763), .Q (____0____33514));
  or2s1 ___0___501856(.DIN1 (___0__9__40628), .DIN2 (____990__33424),
       .Q (____0____33513));
  nnd2s1 ___0___501857(.DIN1 (____0_0__33462), .DIN2 (___90___25036),
       .Q (____0____33512));
  xor2s1 ___0___501858(.DIN1 (_________31721), .DIN2 (____0____33476),
       .Q (____0____33511));
  nor2s1 ___0___501859(.DIN1 (____0_9__33509), .DIN2 (_________33321),
       .Q (____0_0__33510));
  xor2s1 ___0__501860(.DIN1 (___0__0__40413), .DIN2 (____0____33478),
       .Q (____0____33508));
  nnd2s1 ___0___501861(.DIN1 (_____9___33617), .DIN2 (_________36761),
       .Q (____0____33507));
  nnd2s1 ___0___501862(.DIN1 (____0____33463), .DIN2 (___09___28831),
       .Q (____0____33506));
  and2s1 ___0___501863(.DIN1 (_____9___33617), .DIN2
       (______________________________________________________________________________________0__22096),
       .Q (____0____33505));
  or2s1 ___0___501864(.DIN1
       (______________________________________________________________________________________0__22096),
       .DIN2 (_____9___33617), .Q (____0____33504));
  nnd2s1 ___0__501865(.DIN1 (____0____33501), .DIN2 (______9__31622),
       .Q (____0____33503));
  nnd2s1 ___0___501866(.DIN1 (____0____33501), .DIN2 (___0_____31383),
       .Q (____0____33502));
  nnd2s1 ___0___501867(.DIN1 (____0____33455), .DIN2 (________27709),
       .Q (____0_0__33500));
  nnd2s1 ___0___501868(.DIN1 (____0____33498), .DIN2 (________22378),
       .Q (____0_9__33499));
  or2s1 ___0___501869(.DIN1 (____0____33496), .DIN2 (____0____33457),
       .Q (____0____33497));
  nnd2s1 ___0__501870(.DIN1 (____0_9__33461), .DIN2 (________27311), .Q
       (____0____33495));
  nnd2s1 ___0_9_501871(.DIN1 (____0____33454), .DIN2 (____0____33493),
       .Q (____0____33494));
  or2s1 ___0_9_501872(.DIN1 (____0____33491), .DIN2 (____0____33453),
       .Q (____0____33492));
  nnd2s1 ___0_9_501873(.DIN1 (____0_0__33452), .DIN2 (____0_9__33489),
       .Q (____0_0__33490));
  nnd2s1 ___0_501874(.DIN1 (____0____33456), .DIN2 (____0____33487), .Q
       (____0____33488));
  or2s1 ___0_501875(.DIN1 (____0____33485), .DIN2 (____0____33460), .Q
       (____0____33486));
  xor2s1 ___0___501876(.DIN1 (____0____33450), .DIN2
       (_________________________________________________________________________________________22091),
       .Q (____09___33523));
  nor2s1 ___0___501877(.DIN1 (____9____33398), .DIN2 (____0____33458),
       .Q (_________33555));
  nnd2s1 ___0___501878(.DIN1 (____0____33474), .DIN2 (____0____33475),
       .Q (____0____33484));
  or2s1 ___0___501879(.DIN1 (____0____33482), .DIN2 (____0____33448),
       .Q (____0____33483));
  nnd2s1 ___0__501880(.DIN1 (____0____33447), .DIN2 (_________34644),
       .Q (____0____33481));
  nor2s1 ___0___501881(.DIN1
       (____________________________________________21865), .DIN2
       (______________22068), .Q (____0_0__33480));
  nor2s1 ___0___501882(.DIN1 (_____0___33256), .DIN2 (____0____33478),
       .Q (____0_9__33479));
  or2s1 ___0___501883(.DIN1 (_________31625), .DIN2 (____0____33476),
       .Q (____0____33477));
  nor2s1 ___0___501884(.DIN1 (____0____33475), .DIN2 (____0____33474),
       .Q (_________33539));
  xor2s1 ___0_9_501885(.DIN1 (____9____33420), .DIN2 (_________38456),
       .Q (____0____36213));
  xor2s1 ___0___501886(.DIN1 (____9____33421), .DIN2 (_________38203),
       .Q (_________33763));
  xor2s1 ___0___501887(.DIN1 (___0_____40634), .DIN2
       (_________________________________________________________________________________________22094),
       .Q (_________33542));
  nor2s1 ___0___501888(.DIN1 (_________32903), .DIN2 (____0____33443),
       .Q (____0____33473));
  nor2s1 ___0___501889(.DIN1 (___9____27762), .DIN2 (____009__33441),
       .Q (____0____33472));
  or2s1 ___0_9_501890(.DIN1 (_____0___31994), .DIN2 (____00___33439),
       .Q (____0_0__33471));
  nor2s1 ___0_9_501891(.DIN1 (___0_____31345), .DIN2 (____00___33438),
       .Q (____0_9__33470));
  nnd2s1 ___0_9_501892(.DIN1 (____0_0__33442), .DIN2 (____9____32398),
       .Q (____0____33469));
  nnd2s1 ___0___501893(.DIN1 (____000__33433), .DIN2 (_____9___32965),
       .Q (____0____33468));
  nnd2s1 ___0___501894(.DIN1 (____00___33436), .DIN2 (___0_____31154),
       .Q (____0____33467));
  nor2s1 ___0__501895(.DIN1 (____0____33465), .DIN2 (____00___33435),
       .Q (____0____33466));
  nor2s1 ___0___501896(.DIN1 (_________31668), .DIN2 (____00___33434),
       .Q (____0____33464));
  nor2s1 ___0_0_501897(.DIN1 (____99___33425), .DIN2 (_____0__29083),
       .Q (____0____33463));
  nnd2s1 ___0___501898(.DIN1 (____9____33422), .DIN2 (______9__33955),
       .Q (____0_0__33462));
  nor2s1 ___0___501899(.DIN1 (_________33233), .DIN2 (____99___33429),
       .Q (____0____33517));
  hi1s1 ___0___501900(.DIN
       (____________________________________________21865), .Q
       (____0_9__33509));
  nor2s1 ___0___501901(.DIN1 (____9___27737), .DIN2 (____99___33428),
       .Q (_________33676));
  nnd2s1 ___0___501902(.DIN1 (____9____33413), .DIN2 (____0____33449),
       .Q (____0____33498));
  nor2s1 ___0___501903(.DIN1 (_________32315), .DIN2 (____99___33426),
       .Q (____0____33515));
  dffacs1 _________________________________________9__0_(.CLRB (reset),
       .CLK (clk), .DIN (____99___33430), .QN (___0__9__40628));
  dffacs1 _________________501904(.CLRB (reset), .CLK (clk), .DIN
       (____99___33431), .QN
       (_________________________________________________________________________________________22092));
  dffacs1 ______________________________________________501905(.CLRB
       (reset), .CLK (clk), .DIN (____9_9__33423), .Q (___0_____40479));
  xor2s1 ___0__501906(.DIN1 (____9____33396), .DIN2 (_________38214),
       .Q (_____9___33617));
  and2s1 ___0___501907(.DIN1 (____9____33416), .DIN2 (_____9__27289),
       .Q (____0_9__33461));
  nnd2s1 ___0___501908(.DIN1 (____9____33417), .DIN2 (____0____33459),
       .Q (____0____33460));
  nor2s1 ___0___501909(.DIN1 (___9_0___39170), .DIN2 (____9____33418),
       .Q (____0____33458));
  nnd2s1 ___0__501910(.DIN1 (____9____33410), .DIN2 (____9____33353),
       .Q (____0____33457));
  nor2s1 ___0___501911(.DIN1 (___0_____31194), .DIN2 (____9____33408),
       .Q (____0____33456));
  nor2s1 ___0_9_501912(.DIN1 (_________31724), .DIN2 (____0_9__33451),
       .Q (____0____33455));
  nor2s1 ___0___501913(.DIN1 (_________32246), .DIN2 (____9____33411),
       .Q (____0____33454));
  nnd2s1 ___0__501914(.DIN1 (____9_9__33414), .DIN2 (_________32720),
       .Q (____0____33453));
  nor2s1 ___0___501915(.DIN1 (__9_9___30362), .DIN2 (____9____33409),
       .Q (____0_0__33452));
  nor2s1 ___0_0_501916(.DIN1 (________29431), .DIN2 (____0_9__33451),
       .Q (____0____33501));
  dffacs1 ____0__________________501917(.CLRB (reset), .CLK (clk), .DIN
       (____9____33419), .QN (____0________________21665));
  and2s1 ___0___501918(.DIN1 (____9____33412), .DIN2 (____0____33449),
       .Q (____0____33450));
  or2s1 ___0___501919(.DIN1 (____9____33401), .DIN2 (____0____33446),
       .Q (____0____33448));
  xor2s1 ___0___501920(.DIN1 (_________32316), .DIN2 (____0____33446),
       .Q (____0____33447));
  xor2s1 ___0___501921(.DIN1 (_________33206), .DIN2 (______0__40924),
       .Q (____0____33445));
  xor2s1 ___0__501922(.DIN1 (________), .DIN2 (____99___33427), .Q
       (____0____33444));
  nnd2s1 ___0__501923(.DIN1 (____9____33406), .DIN2 (____9____33380),
       .Q (____0____33474));
  nor2s1 ___0___501924(.DIN1 (_________33220), .DIN2 (____9____33402),
       .Q (____0____33478));
  nor2s1 ___0___501925(.DIN1 (___0_____30726), .DIN2 (____9_9__33404),
       .Q (____0____33476));
  dffacs1 ______________________________________________501926(.CLRB
       (reset), .CLK (clk), .DIN (____9____33407), .Q
       (____________________________________________21865));
  nnd2s1 ___0___501927(.DIN1 (____9_9__33394), .DIN2 (___09____31443),
       .Q (____0____33443));
  nor2s1 ___0___501928(.DIN1 (_____9___32275), .DIN2 (____00___33440),
       .Q (____0_0__33442));
  nnd2s1 ___0___501929(.DIN1 (____9____33392), .DIN2 (___0_9___31301),
       .Q (____009__33441));
  nnd2s1 ___0___501930(.DIN1 (____9____33391), .DIN2 (_________41321),
       .Q (____00___33439));
  or2s1 ___0___501931(.DIN1 (____00___33437), .DIN2 (____9_0__33395),
       .Q (____00___33438));
  nnd2s1 ___0_501932(.DIN1 (____9____33388), .DIN2 (_________32104), .Q
       (____00___33436));
  nnd2s1 ___0_0_501933(.DIN1 (____9____33387), .DIN2 (____0____33459),
       .Q (____00___33435));
  nnd2s1 ___0_0_501934(.DIN1 (____9____33390), .DIN2 (_____9___32673),
       .Q (____00___33434));
  and2s1 ___0_501935(.DIN1 (____9____33389), .DIN2 (____999__33432), .Q
       (____000__33433));
  or2s1 ___0_0_501936(.DIN1 (____9_9__33375), .DIN2 (_____9__26354), .Q
       (____99___33431));
  or2s1 ___0_9_501937(.DIN1 (____9___28286), .DIN2 (____9_0__33385), .Q
       (____99___33430));
  nor2s1 ___0_501938(.DIN1 (_________33207), .DIN2 (______0__40924), .Q
       (____99___33429));
  and2s1 ___0_0_501939(.DIN1 (____99___33427), .DIN2 (____90__27732),
       .Q (____99___33428));
  and2s1 ___0_0_501940(.DIN1 (_________32225), .DIN2 (____0____33446),
       .Q (____99___33426));
  nor2s1 ___0___501941(.DIN1 (____9_0__33376), .DIN2 (____990__33424),
       .Q (____99___33425));
  nnd2s1 ___0___501942(.DIN1 (____9____33374), .DIN2 (____00__25862),
       .Q (____9_9__33423));
  xor2s1 ___0__501943(.DIN1 (___0_____30884), .DIN2 (____9____33403),
       .Q (____9____33422));
  xor2s1 ___0___501944(.DIN1 (____9____33348), .DIN2 (__________9_), .Q
       (____9____33421));
  nnd2s1 ___0___501945(.DIN1 (____9____33372), .DIN2 (______9__33311),
       .Q (____9____33420));
  nnd2s1 ___0___501946(.DIN1 (____9____33363), .DIN2 (_____0___34487),
       .Q (____9____33419));
  nor2s1 ___0___501947(.DIN1 (_____9__22710), .DIN2 (____9_9__33365),
       .Q (____9____33418));
  and2s1 ___0___501948(.DIN1 (____9____33354), .DIN2 (______0__41319),
       .Q (____9____33417));
  nor2s1 ___0___501949(.DIN1 (____9_0__33415), .DIN2 (____9____33370),
       .Q (____9____33416));
  nor2s1 ___0__501950(.DIN1 (________25746), .DIN2 (____9____33358), .Q
       (____9_9__33414));
  nnd2s1 ___0___501951(.DIN1 (____9____33412), .DIN2 (_________36402),
       .Q (____9____33413));
  nnd2s1 ___0___501952(.DIN1 (____9_9__33355), .DIN2 (______0__31815),
       .Q (____9____33411));
  nor2s1 ___0_0_501953(.DIN1 (___0_____30977), .DIN2 (____9____33360),
       .Q (____9____33410));
  nnd2s1 ___0__501954(.DIN1 (____9____33357), .DIN2 (________26430), .Q
       (____9____33409));
  nnd2s1 ___0___501955(.DIN1 (____9____33359), .DIN2 (_____9___33329),
       .Q (____9____33408));
  nor2s1 ___0___501956(.DIN1 (___0_____30695), .DIN2 (____9_0__33366),
       .Q (____0_9__33451));
  nnd2s1 ___0_0_501957(.DIN1 (____9____33351), .DIN2 (________27626),
       .Q (____9____33407));
  xor2s1 ___0___501958(.DIN1 (_________33325), .DIN2 (_________38591),
       .Q (____9____33406));
  xnr2s1 ___0___501959(.DIN1
       (_____________________________________0______21754), .DIN2
       (_________34692), .Q (____9_0__33405));
  and2s1 ___0___501960(.DIN1 (____9____33403), .DIN2 (___0_____30725),
       .Q (____9_9__33404));
  xor2s1 ___0__501961(.DIN1 (_________33314), .DIN2 (____0_9__36267),
       .Q (____9____33402));
  nor2s1 ___0___501962(.DIN1 (____9____33349), .DIN2 (____9____33400),
       .Q (____9____33401));
  xor2s1 ___0___501963(.DIN1 (_________33288), .DIN2 (_____90__22048),
       .Q (____9____33399));
  nor2s1 ___0__501964(.DIN1 (____9____33397), .DIN2 (____9_0__33346),
       .Q (____9____33398));
  xor2s1 ___0___501965(.DIN1 (____9____33364), .DIN2 (____909__33345),
       .Q (____9____33396));
  nnd2s1 ___0___501966(.DIN1 (____90___33340), .DIN2 (_________33117),
       .Q (____0____33449));
  nnd2s1 ___0___501967(.DIN1 (_____9___33334), .DIN2 (___0_____30771),
       .Q (____9_0__33395));
  and2s1 ___0___501968(.DIN1 (_____9___33333), .DIN2 (____9____33393),
       .Q (____9_9__33394));
  nor2s1 ___0___501969(.DIN1 (________29251), .DIN2 (_________40926),
       .Q (____9____33392));
  nor2s1 ___0__501970(.DIN1 (___0__0__31080), .DIN2 (_____99__33336),
       .Q (____9____33391));
  nor2s1 ___0__501971(.DIN1 (____0___28472), .DIN2 (_____9___33331), .Q
       (____9____33390));
  nor2s1 ___0___501972(.DIN1 (___0____28779), .DIN2 (_____9___33332),
       .Q (____9____33389));
  nor2s1 ___0___501973(.DIN1 (____0____33491), .DIN2 (_____9___33330),
       .Q (____9____33388));
  nor2s1 ___0___501974(.DIN1 (_________33217), .DIN2 (_____9___33328),
       .Q (____9____33387));
  or2s1 ___0_9_501975(.DIN1 (____9____33386), .DIN2 (____900__33337),
       .Q (____00___33440));
  dffacs1 ____0________________9_501976(.CLRB (reset), .CLK (clk), .DIN
       (____90___33338), .QN (____0____________9___21722));
  nnd2s1 ___0___501977(.DIN1 (___9_0__28673), .DIN2 (______9__33326),
       .Q (____9_0__33385));
  xor2s1 ___0___501978(.DIN1 (____9____33383), .DIN2 (___0__9__40530),
       .Q (____9_9__33384));
  or2s1 ___0___501979(.DIN1
       (_____________________________________0______21754), .DIN2
       (_________34692), .Q (____9____33382));
  and2s1 ___0___501980(.DIN1 (_________34692), .DIN2
       (_____________________________________0______21754), .Q
       (____9____33381));
  nnd2s1 ___0___501981(.DIN1 (____9____33378), .DIN2 (___0__9__40530),
       .Q (____9____33379));
  nor2s1 ___0___501982(.DIN1 (___0__9__40530), .DIN2 (____9____33378),
       .Q (____9____33377));
  xor2s1 ___0___501983(.DIN1 (_________33294), .DIN2 (____9____38944),
       .Q (____9_0__33376));
  nor2s1 ___0___501984(.DIN1 (_________40928), .DIN2 (____9____33350),
       .Q (____9_9__33375));
  nnd2s1 ___0__501985(.DIN1 (_________33319), .DIN2 (_________34877),
       .Q (____9____33374));
  nnd2s1 ___0___501986(.DIN1 (_________33320), .DIN2 (_________37717),
       .Q (____9____33373));
  nor2s1 ___0___501987(.DIN1 (_________33219), .DIN2 (_________33324),
       .Q (____9____33372));
  xor2s1 ___0___501988(.DIN1 (_________33297), .DIN2 (_____99__37662),
       .Q (____99___33427));
  nor2s1 ___0__501989(.DIN1
       (________________________________________0___21788), .DIN2
       (____9____33371), .Q (____0____33446));
  nnd2s1 ___0___501990(.DIN1 (_________33305), .DIN2 (___9____29590),
       .Q (____9____33370));
  nor2s1 ___0___501991(.DIN1 (___0_9___40552), .DIN2 (_____0___35566),
       .Q (____9____33369));
  nnd2s1 ___0___501992(.DIN1 (_____0___35566), .DIN2 (___0_9___40552),
       .Q (____9____33368));
  nor2s1 ___0_0_501993(.DIN1 (____0___29283), .DIN2 (_________33315),
       .Q (____9____33367));
  nnd2s1 ___0__501994(.DIN1 (_________33308), .DIN2 (__9_9___30267), .Q
       (____9_0__33366));
  and2s1 ___0___501995(.DIN1 (____9____33364), .DIN2 (________22531),
       .Q (____9_9__33365));
  and2s1 ___0__501996(.DIN1 (_________33307), .DIN2 (____9____33362),
       .Q (____9____33363));
  xor2s1 ___0___501997(.DIN1 (___0_9___40552), .DIN2 (______9__35544),
       .Q (____9____33361));
  or2s1 ___0___501998(.DIN1 (_________33609), .DIN2 (______0__33302),
       .Q (____9____33360));
  nor2s1 ___0___501999(.DIN1 (________26444), .DIN2 (_________33309),
       .Q (____9____33359));
  nnd2s1 ___0__502000(.DIN1 (_________33304), .DIN2 (________25602), .Q
       (____9____33358));
  nor2s1 ___0___502001(.DIN1 (____9_0__33356), .DIN2 (_________33306),
       .Q (____9____33357));
  nor2s1 ___0___502002(.DIN1 (___0____27906), .DIN2 (______9__33301),
       .Q (____9_9__33355));
  and2s1 ___0___502003(.DIN1 (_________33299), .DIN2 (____9____33353),
       .Q (____9____33354));
  nnd2s1 ___0___502004(.DIN1 (____90___33339), .DIN2
       (_________________________________________________________________________________________22095),
       .Q (____9____33412));
  or2s1 ___0__502005(.DIN1
       (___________________________________________), .DIN2
       (______9__35544), .Q (____9____33352));
  nnd2s1 ___0___502006(.DIN1 (_________33296), .DIN2 (____9____33350),
       .Q (____9____33351));
  hi1s1 ___0___502007(.DIN
       (________________________________________0___21788), .Q
       (____9____33349));
  xor2s1 ___0___502008(.DIN1 (____9____33347), .DIN2 (_________33313),
       .Q (____9____33348));
  nnd2s1 ___0___502009(.DIN1 (_________33298), .DIN2 (____909__33345),
       .Q (____9_0__33346));
  nnd2s1 ___0___502010(.DIN1 (_________33295), .DIN2 (______9__33955),
       .Q (____90___33344));
  nnd2s1 ___0__502011(.DIN1 (______9__35544), .DIN2
       (___________________________________________), .Q
       (____90___33343));
  and2s1 ___0___502012(.DIN1 (_________33288), .DIN2 (_____90__22048),
       .Q (____90___33342));
  nor2s1 ___0___502013(.DIN1 (_____90__22048), .DIN2 (_________33288),
       .Q (____90___33341));
  hi1s1 ___0_502014(.DIN (____90___33339), .Q (____90___33340));
  xor2s1 ___0___502015(.DIN1 (_________33273), .DIN2 (___090__23301),
       .Q (____9____33403));
  nnd2s1 ___0___502016(.DIN1 (_________33287), .DIN2 (_____9___34752),
       .Q (____90___33338));
  nnd2s1 ___0___502017(.DIN1 (_____9___33335), .DIN2 (________26239),
       .Q (____900__33337));
  nnd2s1 ___0___502018(.DIN1 (_____9___33335), .DIN2 (_________32821),
       .Q (_____99__33336));
  and2s1 ___0___502019(.DIN1 (_____9___33335), .DIN2 (_____0___32972),
       .Q (_____9___33334));
  and2s1 ___0__502020(.DIN1 (_________33285), .DIN2 (___0_00__31216),
       .Q (_____9___33333));
  nnd2s1 ___0__502021(.DIN1 (_________33280), .DIN2 (_________33934),
       .Q (_____9___33332));
  nnd2s1 ___0___502022(.DIN1 (_________33281), .DIN2 (________28162),
       .Q (_____9___33331));
  nnd2s1 ___0___502023(.DIN1 (______9__33283), .DIN2 (_____9___33329),
       .Q (_____9___33330));
  nnd2s1 ___0_0_502024(.DIN1 (_________33286), .DIN2 (_____90__33327),
       .Q (_____9___33328));
  dffacs1 ____0___________________502025(.CLRB (reset), .CLK (clk),
       .DIN (______0__33284), .QN (____0_________________21724));
  nnd2s1 ___0___502026(.DIN1 (_________33650), .DIN2 (_________33274),
       .Q (______9__33326));
  nnd2s1 ___0_502027(.DIN1 (_________33318), .DIN2 (____9___22447), .Q
       (_________33325));
  and2s1 ___0___502028(.DIN1 (_________33310), .DIN2 (___9_____39332),
       .Q (_________33324));
  xor2s1 ___0___502029(.DIN1 (_________33322), .DIN2 (_________33321),
       .Q (_________33323));
  xor2s1 ___0__502030(.DIN1 (___0_____30705), .DIN2 (______0__33259),
       .Q (_________33320));
  xor2s1 ___0_0_502031(.DIN1 (_____09__33258), .DIN2 (______0__33277),
       .Q (_________33319));
  nnd2s1 ___0___502032(.DIN1 (_________33275), .DIN2 (____0_9__38073),
       .Q (_________33317));
  dffacs1 ____________________________________________0_502033(.CLRB
       (reset), .CLK (clk), .DIN (______9__33276), .QN
       (________________________________________0___21788));
  nnd2s1 ___0_0_502034(.DIN1 (_________33278), .DIN2 (______9__33230),
       .Q (_____0___34663));
  hi1s1 ___0_0_502035(.DIN (____9____33383), .Q (____9____33378));
  xnr2s1 ___0__502036(.DIN1 (_________33316), .DIN2 (_________33261),
       .Q (_________34692));
  nnd2s1 ___0___502037(.DIN1 (_________33271), .DIN2 (________29384),
       .Q (_________33315));
  nor2s1 ___0___502038(.DIN1 (_____0___33160), .DIN2 (_________33313),
       .Q (_________33314));
  or2s1 ___0__502039(.DIN1 (___0_____40650), .DIN2 (_________33310), .Q
       (______9__33311));
  or2s1 ___0_0_502040(.DIN1 (____9____32433), .DIN2 (_________33303),
       .Q (_________33309));
  nor2s1 ___0___502041(.DIN1 (________27704), .DIN2 (______0__33268),
       .Q (_________33308));
  nor2s1 ___0_0_502042(.DIN1 (___0__9__31147), .DIN2 (_________33265),
       .Q (_________33307));
  nnd2s1 ___0___502043(.DIN1 (_________33300), .DIN2 (_____9___31983),
       .Q (_________33306));
  nor2s1 ___0___502044(.DIN1 (________29026), .DIN2 (_________33264),
       .Q (_________33305));
  nor2s1 ___0___502045(.DIN1 (_____0___31802), .DIN2 (_________33303),
       .Q (_________33304));
  or2s1 ___0___502046(.DIN1 (_________33553), .DIN2 (_________33272),
       .Q (______0__33302));
  nnd2s1 ___0___502047(.DIN1 (_________33300), .DIN2 (____0____31560),
       .Q (______9__33301));
  nor2s1 ___0_502048(.DIN1 (____09___32572), .DIN2 (_________33303), .Q
       (_________33299));
  hi1s1 ___0___502049(.DIN (_________33298), .Q (____9____33364));
  nor2s1 ___0___502050(.DIN1 (________23116), .DIN2 (_________33270),
       .Q (____90___33339));
  hi1s1 ___0_0_502051(.DIN (______9__35544), .Q (_____0___35566));
  nnd2s1 ___0__502052(.DIN1 (_________33263), .DIN2 (________26550), .Q
       (_________33297));
  xor2s1 ___0___502053(.DIN1 (_________33235), .DIN2 (______0__40934),
       .Q (_________33296));
  xor2s1 ___0__502054(.DIN1 (_________33238), .DIN2 (_________33228),
       .Q (_________33295));
  xor2s1 ___0___502055(.DIN1 (_________33239), .DIN2 (_________33293),
       .Q (_________33294));
  nor2s1 ___0___502056(.DIN1 (_________33289), .DIN2 (_________33290),
       .Q (______0__33292));
  nnd2s1 ___0___502057(.DIN1 (_________33290), .DIN2 (_________33289),
       .Q (_________33291));
  xor2s1 ___0___502058(.DIN1 (_____9___33246), .DIN2
       (_________________________________________________________________________________________22095),
       .Q (____9____33383));
  hi1s1 ___0_0_502059(.DIN (_________33288), .Q (______0__33312));
  nor2s1 ___0__502060(.DIN1 (_____00__33249), .DIN2 (_____0___33252),
       .Q (_________33287));
  nor2s1 ___0___502061(.DIN1 (____0_9__32546), .DIN2 (_________33282),
       .Q (_________33286));
  nor2s1 ___0___502062(.DIN1 (___0__9__30813), .DIN2 (_____99__33248),
       .Q (_________33285));
  nnd2s1 ___0___502063(.DIN1 (_____0___33250), .DIN2 (_________33128),
       .Q (______0__33284));
  nor2s1 ___0__502064(.DIN1 (_____9___32280), .DIN2 (_________33282),
       .Q (______9__33283));
  nor2s1 ___0___502065(.DIN1 (________29415), .DIN2 (_____0___33254),
       .Q (_________33281));
  nor2s1 ___0___502066(.DIN1 (_________32697), .DIN2 (_________33282),
       .Q (_________33280));
  xor2s1 ___0___502067(.DIN1 (_________33223), .DIN2 (_________37864),
       .Q (_________33298));
  nnd2s1 ___0_9_502068(.DIN1 (_____0___33253), .DIN2 (__9__0__30196),
       .Q (_____9___33335));
  xor2s1 ___0__502069(.DIN1 (____0___25868), .DIN2 (_________33269), .Q
       (______9__35544));
  or2s1 ___0__502070(.DIN1 (_________33229), .DIN2 (______0__33277), .Q
       (_________33278));
  nor2s1 ___0___502071(.DIN1 (____0____33482), .DIN2 (_____9___33242),
       .Q (______9__33276));
  xor2s1 ___0___502072(.DIN1 (___9____27759), .DIN2 (_________33262),
       .Q (_________33275));
  xor2s1 ___0___502073(.DIN1 (______0__33204), .DIN2 (___9_____39372),
       .Q (_________33274));
  nnd2s1 ___0_9_502074(.DIN1 (_________33232), .DIN2 (__90____29697),
       .Q (_________33273));
  nor2s1 ___0___502075(.DIN1 (_________33289), .DIN2 (_____9___33245),
       .Q (_________33310));
  xnr2s1 ___0___502076(.DIN1 (____0_9__36267), .DIN2 (_________33205),
       .Q (_________33318));
  nnd2s1 ___0___502077(.DIN1 (_____9___33247), .DIN2 (_________32620),
       .Q (_________33272));
  nor2s1 ___0___502078(.DIN1 (________26300), .DIN2 (_________40930),
       .Q (_________33271));
  nor2s1 ___0___502079(.DIN1 (_____0__24576), .DIN2 (_________33269),
       .Q (_________33270));
  or2s1 ___0___502080(.DIN1 (______9__33267), .DIN2 (_________33224),
       .Q (______0__33268));
  nor2s1 ___0_0_502081(.DIN1 (______9__32959), .DIN2 (_________33586),
       .Q (_________33266));
  nnd2s1 ___0___502082(.DIN1 (_________33218), .DIN2 (______0__33727),
       .Q (_________33265));
  nnd2s1 ___0__502083(.DIN1 (_________33216), .DIN2 (_____0___31895),
       .Q (_________33264));
  nor2s1 ___0___502084(.DIN1 (_________33036), .DIN2 (_________33237),
       .Q (_________33313));
  nor2s1 ___0___502085(.DIN1 (_________33170), .DIN2 (______0__33222),
       .Q (_________33300));
  xor2s1 ___0___502086(.DIN1 (_________33199), .DIN2 (____9____38909),
       .Q (_________33288));
  nnd2s1 ___0___502087(.DIN1 (_________33227), .DIN2 (_________32811),
       .Q (_________33303));
  nnd2s1 ___0___502088(.DIN1 (_________33262), .DIN2 (________26551),
       .Q (_________33263));
  xor2s1 ___0__502089(.DIN1 (_________33236), .DIN2
       (______________22068), .Q (_________33261));
  xor2s1 ___0___502090(.DIN1 (______0__33231), .DIN2 (_________37202),
       .Q (______0__33259));
  xor2s1 ___0___502091(.DIN1 (________23837), .DIN2 (_____0___33257),
       .Q (_____09__33258));
  nor2s1 ___0_0_502092(.DIN1 (___0__0__40413), .DIN2 (_____0___33255),
       .Q (_____0___33256));
  nor2s1 ___0_9_502093(.DIN1 (_____9__22412), .DIN2 (_________33210),
       .Q (_________33322));
  xor2s1 ___0___502094(.DIN1 (_____9___33243), .DIN2 (_____9___33244),
       .Q (_________33290));
  nnd2s1 ___0___502095(.DIN1 (_________33197), .DIN2 (___0____27013),
       .Q (_____0___33254));
  nor2s1 ___0__502096(.DIN1 (_____90__41299), .DIN2 (_________33200),
       .Q (_____0___33253));
  nnd2s1 ___0___502097(.DIN1 (_________33192), .DIN2 (_________33096),
       .Q (_____0___33252));
  nnd2s1 ___0___502098(.DIN1 (______0__33195), .DIN2 (________28445),
       .Q (_____0___33251));
  nor2s1 ___0__502099(.DIN1 (_____00__33249), .DIN2 (______9__33194),
       .Q (_____0___33250));
  nnd2s1 ___0___502100(.DIN1 (_________33196), .DIN2 (_____9__26737),
       .Q (_____99__33248));
  dffacs1 _______________________________________________502101(.CLRB
       (reset), .CLK (clk), .DIN (_________33208), .Q
       (_____________________________________________21907));
  hi1s1 ___0___502102(.DIN (_____9___33247), .Q (_________33282));
  dffacs1 ______________________________________________502103(.CLRB
       (reset), .CLK (clk), .DIN (______9__33203), .QN
       (____________________________________________21772));
  xor2s1 ___0___502104(.DIN1 (_________33169), .DIN2 (_____99__36913),
       .Q (_____9___33246));
  and2s1 ___0__502105(.DIN1 (_____9___33244), .DIN2 (_____9___33243),
       .Q (_____9___33245));
  xor2s1 ___0___502106(.DIN1 (_________33778), .DIN2
       (________________________________________0___21771), .Q
       (_____9___33242));
  xnr2s1 ___0___502107(.DIN1 (_________33209), .DIN2
       (______________22067), .Q (_________33239));
  xor2s1 ___0__502108(.DIN1 (_________33187), .DIN2 (_________33234),
       .Q (_________33238));
  and2s1 ___0___502109(.DIN1 (_________33236), .DIN2 (_________33035),
       .Q (_________33237));
  xor2s1 ___0___502110(.DIN1 (_________33234), .DIN2
       (____________________________________________21847), .Q
       (_________33235));
  nor2s1 ___0___502111(.DIN1
       (_____________________________________0____), .DIN2
       (_____0___33257), .Q (_________33233));
  or2s1 ___0__502112(.DIN1 (__90____29696), .DIN2 (______0__33231), .Q
       (_________33232));
  or2s1 ___0___502113(.DIN1
       (____________________________________________21848), .DIN2
       (_____0___33257), .Q (______9__33230));
  and2s1 ___0___502114(.DIN1 (_____0___33257), .DIN2
       (____________________________________________21848), .Q
       (_________33229));
  nnd2s1 ___0_9_502115(.DIN1 (_________33189), .DIN2 (_________33228),
       .Q (_________33279));
  nor2s1 ___0_9_502116(.DIN1 (_________33147), .DIN2 (_________33191),
       .Q (______0__33277));
  nor2s1 ___0___502117(.DIN1 (________27374), .DIN2 (______9__33221),
       .Q (_________33227));
  nor2s1 ___0_9_502118(.DIN1 (______9__33185), .DIN2 (_________33225),
       .Q (_________33226));
  or2s1 ___0___502119(.DIN1 (_________41351), .DIN2 (_________33179),
       .Q (_________33224));
  nor2s1 ___0___502120(.DIN1 (_______22188), .DIN2 (_________33181), .Q
       (_________33223));
  or2s1 ___0___502121(.DIN1 (____9___28008), .DIN2 (______9__33221), .Q
       (______0__33222));
  xnr2s1 ___0___502122(.DIN1 (_________38155), .DIN2 (_____99__33158),
       .Q (_________33220));
  nor2s1 ___0___502123(.DIN1 (_____9___33243), .DIN2 (_____9___33244),
       .Q (_________33219));
  nor2s1 ___0___502124(.DIN1 (_________33217), .DIN2 (_________33173),
       .Q (_________33218));
  nor2s1 ___0__502125(.DIN1 (____0___28930), .DIN2 (_________33174), .Q
       (_________33216));
  nor2s1 ___0__502126(.DIN1 (inData[31]), .DIN2 (______9__33221), .Q
       (_____9___33247));
  nor2s1 ___0___502127(.DIN1 (___9____26880), .DIN2 (_________33171),
       .Q (_________33269));
  hi1s1 ___0___502128(.DIN (_____0___33255), .Q (_________33586));
  dffacs1 ________________________502129(.CLRB (reset), .CLK (clk),
       .DIN (______9__33176), .QN (______________________21699));
  dffacs2 _______________________502130(.CLRB (reset), .CLK (clk), .DIN
       (_________33178), .QN (_____________________21691));
  nnd2s1 ___0___502131(.DIN1 (_________33234), .DIN2 (___0_____40579),
       .Q (_________33215));
  and2s1 ___0_9_502132(.DIN1 (_________33212), .DIN2 (_________33211),
       .Q (______9__33213));
  and2s1 ___0___502133(.DIN1 (_________33209), .DIN2 (____0___22361),
       .Q (_________33210));
  or2s1 ___0___502134(.DIN1 (_____0___33166), .DIN2 (____0____32515),
       .Q (_________33208));
  nor2s1 ___0___502135(.DIN1 (_________33206), .DIN2 (_________33182),
       .Q (_________33207));
  nor2s1 ___0___502136(.DIN1 (_________33201), .DIN2 (_________33202),
       .Q (_________33205));
  and2s1 ___0___502137(.DIN1 (_____0___33164), .DIN2 (_________33209),
       .Q (______0__33204));
  nnd2s1 ___0___502138(.DIN1 (______0__33168), .DIN2 (________26342),
       .Q (______9__33203));
  nnd2s1 ___0__502139(.DIN1 (_________33202), .DIN2 (_________33201),
       .Q (____9____33380));
  nnd2s1 ___0___502140(.DIN1 (_____9___33151), .DIN2 (_____09__31612),
       .Q (_________33200));
  xor2s1 ___0_502141(.DIN1 (____09__28117), .DIN2 (_________40932), .Q
       (_________33199));
  xor2s1 ___0__502142(.DIN1 (_________40656), .DIN2 (__9__9__29974), .Q
       (_________33198));
  nor2s1 ___0_9_502143(.DIN1 (________29256), .DIN2 (_____00__33159),
       .Q (_________33197));
  nor2s1 ___0__502144(.DIN1 (__900_), .DIN2 (_____9___33154), .Q
       (_________33196));
  nor2s1 ___0__502145(.DIN1 (____0___28473), .DIN2 (_____9___33156), .Q
       (______0__33195));
  nnd2s1 ___0___502146(.DIN1 (_____9___33152), .DIN2 (_________33193),
       .Q (______9__33194));
  nor2s1 ___0___502147(.DIN1 (________28963), .DIN2 (_____9___33153),
       .Q (_________33192));
  and2s1 ___0___502148(.DIN1 (___0____27010), .DIN2
       (________________________________________0___21771), .Q
       (_________33262));
  xor2s1 ___0___502149(.DIN1 (___909__26872), .DIN2 (_________33180),
       .Q (_____0___33255));
  dffacs1 ______________________________________________502150(.CLRB
       (reset), .CLK (clk), .DIN (_____09__33167), .QN
       (___0_0___40565));
  nor2s1 ___0___502151(.DIN1 (______9__33148), .DIN2 (_________33188),
       .Q (_________33191));
  nnd2s1 ___0___502152(.DIN1 (_________40656), .DIN2 (___0_9___40553),
       .Q (_________33190));
  nnd2s1 ___0___502153(.DIN1 (_________33188), .DIN2 (_________33187),
       .Q (_________33189));
  or2s1 ___0___502154(.DIN1 (___0_0___40563), .DIN2 (_________40656),
       .Q (______0__33186));
  hi1s1 ___0___502155(.DIN (_________33184), .Q (______9__33185));
  nnd2s1 ___0__502156(.DIN1 (_________40656), .DIN2 (___0_0___40563),
       .Q (_________33183));
  nor2s1 ___0_9_502157(.DIN1 (_________33114), .DIN2 (_________33146),
       .Q (______0__33231));
  nnd2s1 ___0___502158(.DIN1 (_____90__33149), .DIN2 (_________33010),
       .Q (_________33236));
  xor2s1 ___0___502159(.DIN1
       (________________________________________0___21863), .DIN2
       (_________32611), .Q (______9__33240));
  xnr2s1 ___0___502160(.DIN1 (_________38666), .DIN2 (_________33134),
       .Q (_____9___33244));
  hi1s1 ___0_9_502161(.DIN (_________33182), .Q (_____0___33257));
  and2s1 ___0___502162(.DIN1 (_________33180), .DIN2 (_______22181), .Q
       (_________33181));
  nnd2s1 ___0___502163(.DIN1 (______9__33140), .DIN2 (________28040),
       .Q (_________33179));
  nnd2s1 ___0_9_502164(.DIN1 (_________33142), .DIN2 (_________33137),
       .Q (_________33178));
  or2s1 ___0___502165(.DIN1 (___0_9___40553), .DIN2 (_________40656),
       .Q (______0__33177));
  or2s1 ___090_(.DIN1 (_________33175), .DIN2 (_________33138), .Q
       (______9__33176));
  nnd2s1 ___0909(.DIN1 (______0__33141), .DIN2 (________28602), .Q
       (_________33174));
  nnd2s1 ___09__(.DIN1 (_________33145), .DIN2 (_________33172), .Q
       (_________33173));
  and2s1 ___0___502166(.DIN1 (_________40932), .DIN2 (____0___28116),
       .Q (_________33171));
  nor2s1 ___090_502167(.DIN1 (_________33170), .DIN2 (_________33139),
       .Q (______9__33221));
  dffacs1 _______________________502168(.CLRB (reset), .CLK (clk), .DIN
       (_________33144), .QN (_____________________21689));
  nnd2s1 ___0_502169(.DIN1 (_____0___33163), .DIN2 (_________33118), .Q
       (_________33169));
  nnd2s1 ___0_0_502170(.DIN1 (______0__33132), .DIN2 (_________38177),
       .Q (______0__33168));
  nnd2s1 ___0___502171(.DIN1 (_________33133), .DIN2 (___9_9__25094),
       .Q (_____09__33167));
  nor2s1 ___0___502172(.DIN1 (______9__33131), .DIN2 (_____0___33165),
       .Q (_____0___33166));
  or2s1 ___0_502173(.DIN1
       (________________________________________0___21863), .DIN2
       (______________22066), .Q (_____0___33164));
  nnd2s1 ___0___502174(.DIN1 (_____0___33162), .DIN2 (___0_____40546),
       .Q (_________33211));
  nnd2s1 ___0_9_502175(.DIN1 (_____0___33163), .DIN2 (_________33119),
       .Q (_________33202));
  dffacs1 ____________________________________________0_502176(.CLRB
       (reset), .CLK (clk), .DIN (_________33135), .Q
       (________________________________________0___21771));
  or2s1 ___0___502177(.DIN1 (___0_____40546), .DIN2 (_____0___33162),
       .Q (_________33212));
  hi1s1 ___0_9_502178(.DIN (_________33188), .Q (_________33234));
  nnd2s1 ___0___502179(.DIN1 (______________22066), .DIN2
       (________________________________________0___21863), .Q
       (_________33209));
  nor2s1 ___0___502180(.DIN1 (_____0___33161), .DIN2 (_____0___33162),
       .Q (_________33214));
  nor2s1 ___090_502181(.DIN1 (_____9___33157), .DIN2 (____9____33347),
       .Q (_____0___33160));
  nnd2s1 ___09__502182(.DIN1 (_________33136), .DIN2 (____0____31574),
       .Q (_____00__33159));
  nnd2s1 ___09__502183(.DIN1 (____9____33347), .DIN2 (_____9___33157),
       .Q (_____99__33158));
  or2s1 ___0_9_502184(.DIN1 (_____9___33155), .DIN2 (_________33124),
       .Q (_____9___33156));
  nnd2s1 ___0_9_502185(.DIN1 (_________33126), .DIN2 (________29158),
       .Q (_____9___33154));
  nnd2s1 ___0_502186(.DIN1 (_________33125), .DIN2 (__9_____30027), .Q
       (_____9___33153));
  nor2s1 ___09__502187(.DIN1 (_____9__27533), .DIN2 (_________33127),
       .Q (_____9___33152));
  nor2s1 ___09_0(.DIN1 (___9____28679), .DIN2 (______0__33122), .Q
       (_____9___33151));
  nor2s1 ___0___502188(.DIN1
       (________________________________________9_), .DIN2
       (_____9___33150), .Q (_________33225));
  xor2s1 ___0___502189(.DIN1 (_________33113), .DIN2
       (______________22067), .Q (_________33182));
  nnd2s1 ___0___502190(.DIN1 (_____9___33150), .DIN2
       (________________________________________9_), .Q
       (_________33184));
  dffacs1 ____0__________________502191(.CLRB (reset), .CLK (clk), .DIN
       (_________33129), .QN (____0________________21714));
  xor2s1 ___0__502192(.DIN1 (_________33100), .DIN2 (_____0___36285),
       .Q (_____90__33149));
  and2s1 ___0__502193(.DIN1 (______0__40934), .DIN2
       (____________________________________________21847), .Q
       (______9__33148));
  nor2s1 ___0___502194(.DIN1
       (____________________________________________21847), .DIN2
       (______0__40934), .Q (_________33147));
  and2s1 ___0___502195(.DIN1 (_________34141), .DIN2 (_________33116),
       .Q (_________33146));
  nor2s1 ___0__502196(.DIN1
       (____________________________________________21806), .DIN2
       (_________33130), .Q (_________33260));
  xor2s1 ___0___502197(.DIN1 (_________33101), .DIN2
       (______________22066), .Q (_________33188));
  hi1s1 ___0___502198(.DIN (_____9___33150), .Q (_________40656));
  nor2s1 ___09_502199(.DIN1 (__99____30487), .DIN2 (_________33111), .Q
       (_________33145));
  or2s1 ___0_9_502200(.DIN1 (_________33143), .DIN2 (_________33108),
       .Q (_________33144));
  nor2s1 ___09_502201(.DIN1 (_________32688), .DIN2 (_________33110),
       .Q (_________33142));
  nor2s1 ___09__502202(.DIN1 (____9____32449), .DIN2 (______9__33112),
       .Q (______0__33141));
  nor2s1 ___0_9_502203(.DIN1 (___0_____30798), .DIN2 (_________33120),
       .Q (______9__33140));
  nnd2s1 ___09__502204(.DIN1 (_________33107), .DIN2 (_________34243),
       .Q (_________33139));
  nnd2s1 ___09__502205(.DIN1 (_________33109), .DIN2 (_________33137),
       .Q (_________33138));
  xnr2s1 ___09_9(.DIN1 (____0____38091), .DIN2 (_________33091), .Q
       (_________33180));
  nor2s1 ___0___502206(.DIN1 (____0____33482), .DIN2 (______0__33103),
       .Q (_________33135));
  nor2s1 ___0___502207(.DIN1 (_________32708), .DIN2 (_________33098),
       .Q (_________33134));
  nnd2s1 ___0_0_502208(.DIN1 (_________33095), .DIN2 (_________37717),
       .Q (_________33133));
  xor2s1 ___0___502209(.DIN1 (________28119), .DIN2 (_________33115),
       .Q (______0__33132));
  xor2s1 ___0__502210(.DIN1 (_________33086), .DIN2 (___0_9__22316), .Q
       (______9__33131));
  xor2s1 ___0___502211(.DIN1 (_________33087), .DIN2 (_________35968),
       .Q (_____0___33163));
  hi1s1 ___0_9_502212(.DIN (_________33130), .Q (_____0___33162));
  dffacs1 ____________________________________________0_502213(.CLRB
       (reset), .CLK (clk), .DIN (_________33104), .Q
       (________________________________________0___21863));
  nnd2s1 ___090_502214(.DIN1 (_________33097), .DIN2 (_________33128),
       .Q (_________33129));
  nnd2s1 ___09__502215(.DIN1 (_________33089), .DIN2 (________28302),
       .Q (_________33127));
  nor2s1 ___09__502216(.DIN1 (____0_0__32557), .DIN2 (______9__33092),
       .Q (_________33126));
  nor2s1 ___09__502217(.DIN1 (_____0___32777), .DIN2 (______0__33093),
       .Q (_________33125));
  or2s1 ___09__502218(.DIN1 (_________33123), .DIN2 (_________33090),
       .Q (_________33124));
  nnd2s1 ___09__502219(.DIN1 (_________33105), .DIN2 (___0_____31035),
       .Q (______0__33122));
  nnd2s1 ___09__502220(.DIN1 (_________33094), .DIN2 (_____0__28538),
       .Q (_________33136));
  hi1s1 ___09_502221(.DIN (______9__33121), .Q (____9____33347));
  xor2s1 ___0_502222(.DIN1 (_________33081), .DIN2 (___9_____39384), .Q
       (_____9___33150));
  nnd2s1 ___09__502223(.DIN1 (_________33088), .DIN2 (_____9__29455),
       .Q (_________33120));
  nnd2s1 ___0__502224(.DIN1 (_________33118), .DIN2 (_________33117),
       .Q (_________33119));
  or2s1 ___0___502225(.DIN1 (___0_0___40565), .DIN2 (_________33115),
       .Q (_________33116));
  and2s1 ___0___502226(.DIN1 (_________33115), .DIN2 (___0_0___40565),
       .Q (_________33114));
  xor2s1 ___0___502227(.DIN1 (____0____33475), .DIN2 (_________33099),
       .Q (_________33113));
  xor2s1 ___0___502228(.DIN1 (_____0___33073), .DIN2 (_____0___32286),
       .Q (_________33130));
  nnd2s1 ___09__502229(.DIN1 (______0__33075), .DIN2 (________29311),
       .Q (______9__33112));
  nnd2s1 ___099_(.DIN1 (_____09__33074), .DIN2 (__90____29672), .Q
       (_________33111));
  nnd2s1 ___09__502230(.DIN1 (_________33076), .DIN2 (__9_9___30446),
       .Q (_________33110));
  nor2s1 ___09__502231(.DIN1 (________28886), .DIN2 (_________33078),
       .Q (_________33109));
  nnd2s1 ___09_502232(.DIN1 (_________33085), .DIN2 (_____9___32968),
       .Q (_________33108));
  nor2s1 ___09_502233(.DIN1 (_________33106), .DIN2 (_________33077),
       .Q (_________33107));
  xor2s1 ___09__502234(.DIN1 (______9__33055), .DIN2 (_________33973),
       .Q (______9__33121));
  dffacs1 ______________________0_502235(.CLRB (reset), .CLK (clk),
       .DIN (_________33079), .QN (__________________0___21750));
  nor2s1 ___09_502236(.DIN1 (____0_0__31523), .DIN2 (_____9___33060),
       .Q (_________33105));
  nnd2s1 ___0___502237(.DIN1 (_____0___33072), .DIN2 (____9___27652),
       .Q (_________33104));
  xor2s1 ___0___502238(.DIN1
       (________________________________________0_), .DIN2
       (_________34026), .Q (______0__33103));
  nor2s1 ___0___502239(.DIN1 (_________38833), .DIN2 (_____0___33068),
       .Q (______9__33102));
  xor2s1 ___0___502240(.DIN1 (_________33043), .DIN2 (___90____39001),
       .Q (_________33101));
  nor2s1 ___090_502241(.DIN1 (_________32919), .DIN2 (_________33099),
       .Q (_________33100));
  nor2s1 ___09__502242(.DIN1 (________24760), .DIN2 (_____0___33071),
       .Q (_________33098));
  and2s1 ___09__502243(.DIN1 (_____9___33063), .DIN2 (_________33096),
       .Q (_________33097));
  xor2s1 ___0__502244(.DIN1 (_________33048), .DIN2 (_________37616),
       .Q (_________33095));
  nor2s1 ____0__502245(.DIN1 (___9_0__26930), .DIN2 (_________33051),
       .Q (_________33094));
  nnd2s1 ___09__502246(.DIN1 (_____90__33056), .DIN2 (__99____30497),
       .Q (______0__33093));
  nnd2s1 ___0990(.DIN1 (_____9___33058), .DIN2 (________29393), .Q
       (______9__33092));
  nnd2s1 ____00_502247(.DIN1 (_____9___33057), .DIN2 (_________33053),
       .Q (_________33091));
  nnd2s1 ___09__502248(.DIN1 (_____9___33062), .DIN2 (___09____31469),
       .Q (_________33090));
  nor2s1 ___09__502249(.DIN1 (______0__33008), .DIN2 (_____0___33069),
       .Q (_________33089));
  dffacs1 ____0___________________502250(.CLRB (reset), .CLK (clk),
       .DIN (_________33052), .QN (____0_________________21726));
  dffacs1 _______________________502251(.CLRB (reset), .CLK (clk), .DIN
       (_________33050), .QN (_____________________21674));
  dffacs1 ________________________502252(.CLRB (reset), .CLK (clk),
       .DIN (_____9___33061), .QN (____________________));
  nor2s1 ___09__502253(.DIN1 (________27042), .DIN2 (_________33031),
       .Q (_________33088));
  nor2s1 ___090_502254(.DIN1 (_________33080), .DIN2 (_________40936),
       .Q (_________33087));
  xor2s1 ___0___502255(.DIN1 (___0_____40613), .DIN2
       (__________________________________________________________________21989),
       .Q (_________33086));
  nor2s1 ___09__502256(.DIN1 (_____0___32775), .DIN2 (______9__33027),
       .Q (_________33085));
  and2s1 ___09__502257(.DIN1 (______9__33083), .DIN2 (_________33082),
       .Q (______0__33084));
  xor2s1 ___09__502258(.DIN1 (________28129), .DIN2 (_____9___33064),
       .Q (_________33081));
  nnd2s1 ___090_502259(.DIN1 (_________40936), .DIN2 (_________33080),
       .Q (_________33118));
  nor2s1 ___09_502260(.DIN1
       (________________________________________0_), .DIN2
       (___9____27758), .Q (_________33115));
  dffacs1 _______________________502261(.CLRB (reset), .CLK (clk), .DIN
       (______0__33038), .QN (_____________________21688));
  nnd2s1 ____0_502262(.DIN1 (______0__33018), .DIN2 (_________33032),
       .Q (_________33079));
  nnd2s1 ____0__502263(.DIN1 (_________33023), .DIN2 (________28214),
       .Q (_________33078));
  nnd2s1 ____0_502264(.DIN1 (_________33022), .DIN2 (___0090__30632),
       .Q (_________33077));
  nor2s1 ____0__502265(.DIN1 (_____9__28432), .DIN2 (_________33019),
       .Q (_________33076));
  nor2s1 ____0_502266(.DIN1 (___09____31478), .DIN2 (_________33034),
       .Q (______0__33075));
  nor2s1 ____0__502267(.DIN1 (_____9__26812), .DIN2 (_________33021),
       .Q (_____09__33074));
  dffacs1 ______________________0_502268(.CLRB (reset), .CLK (clk),
       .DIN (_________33029), .QN (__________________0___21697));
  dffacs1 ____0_________________0_502269(.CLRB (reset), .CLK (clk),
       .DIN (_________33025), .Q (____0_____________0___21723));
  dffacs1 _______________________502270(.CLRB (reset), .CLK (clk), .DIN
       (_________33041), .QN (_____________________21684));
  dffacs1 _______________________502271(.CLRB (reset), .CLK (clk), .DIN
       (_________33033), .QN (_____________________21744));
  xor2s1 ___0___502272(.DIN1 (_________32992), .DIN2 (_________41248),
       .Q (_____0___33073));
  nnd2s1 ___09__502273(.DIN1 (_________33015), .DIN2 (____9____33350),
       .Q (_____0___33072));
  nnd2s1 ___09__502274(.DIN1 (_________33013), .DIN2 (_________32795),
       .Q (_____0___33071));
  xor2s1 ___09__502275(.DIN1 (________24428), .DIN2 (_________33006),
       .Q (_____0___33070));
  nnd2s1 ____0__502276(.DIN1 (_________33003), .DIN2 (______9__32998),
       .Q (_____0___33069));
  xor2s1 ___09__502277(.DIN1 (_________32986), .DIN2 (_____0___32977),
       .Q (_____0___33068));
  nor2s1 ___09__502278(.DIN1 (_____00__33066), .DIN2 (_____0___32976),
       .Q (_____0___33067));
  nnd2s1 ___09_502279(.DIN1 (_____9___33064), .DIN2 (_____0__28128), .Q
       (_____99__33065));
  nor2s1 ___099_502280(.DIN1 (_________33002), .DIN2 (______9__33007),
       .Q (_____9___33063));
  nor2s1 ____0_502281(.DIN1 (________28268), .DIN2 (_________32993), .Q
       (_____9___33062));
  xnr2s1 ___09__502282(.DIN1 (____9_9__37984), .DIN2 (_________32984),
       .Q (_________33099));
  nor2s1 ___09__502283(.DIN1 (_________32988), .DIN2 (_________33012),
       .Q (____9____36155));
  nnd2s1 ____0__502284(.DIN1 (_________32995), .DIN2 (______0__33028),
       .Q (_____9___33061));
  or2s1 ____0__502285(.DIN1 (_____9___33059), .DIN2 (_________33004),
       .Q (_____9___33060));
  nor2s1 ____0__502286(.DIN1 (________27141), .DIN2 (_________33001),
       .Q (_____9___33058));
  nnd2s1 ____0__502287(.DIN1 (_________33054), .DIN2 (_________33973),
       .Q (_____9___33057));
  nor2s1 ____0__502288(.DIN1 (____0___28560), .DIN2 (_________33009),
       .Q (_____90__33056));
  and2s1 ____0__502289(.DIN1 (_________33054), .DIN2 (_________33053),
       .Q (______9__33055));
  nnd2s1 ____0__502290(.DIN1 (_________33005), .DIN2 (_________33128),
       .Q (_________33052));
  nnd2s1 ____0__502291(.DIN1 (_________32996), .DIN2 (___99___28731),
       .Q (_________33051));
  nnd2s1 _____502292(.DIN1 (_________32994), .DIN2 (_____0___32577), .Q
       (_________33050));
  dffacs1 ____0__________________502293(.CLRB (reset), .CLK (clk), .DIN
       (______9__33017), .QN (____0________________21667));
  dffacs1 ____0__________________502294(.CLRB (reset), .CLK (clk), .DIN
       (______0__32999), .QN (____0________________21719));
  dffacs1 _______________________502295(.CLRB (reset), .CLK (clk), .DIN
       (_________32997), .QN (_____________________21670));
  hi1s1 ___0_9_502296(.DIN
       (__________________________________________________________________21989),
       .Q (_________33049));
  xor2s1 ___09__502297(.DIN1 (_________32954), .DIN2 (______0__32990),
       .Q (_________33048));
  nor2s1 ___099_502298(.DIN1 (_________36493), .DIN2 (_________33316),
       .Q (_________33047));
  nnd2s1 ___099_502299(.DIN1 (_________33316), .DIN2 (_________36493),
       .Q (______0__33046));
  and2s1 ___09__502300(.DIN1 (_________33006), .DIN2 (___0__0__40501),
       .Q (______9__33045));
  xor2s1 ___09_502301(.DIN1 (_________32946), .DIN2 (_________33201),
       .Q (_________33043));
  nor2s1 ___09__502302(.DIN1 (_____9___22051), .DIN2 (_________33006),
       .Q (_________33042));
  or2s1 ___09__502303(.DIN1 (_________32128), .DIN2 (_________32981),
       .Q (_________33041));
  nor2s1 ___09__502304(.DIN1 (___0__0__40501), .DIN2 (_________33006),
       .Q (_________33040));
  nor2s1 ___09__502305(.DIN1 (___0__0__40511), .DIN2 (_________33006),
       .Q (_________33039));
  nnd2s1 ___09__502306(.DIN1 (_________32991), .DIN2 (_________32922),
       .Q (_________33228));
  nnd2s1 ___09__502307(.DIN1 (_________33006), .DIN2
       (____________________________________________21764), .Q
       (_________33082));
  or2s1 ___09__502308(.DIN1
       (____________________________________________21764), .DIN2
       (_________33006), .Q (______9__33083));
  dffacs1 ____________________________________________0_502309(.CLRB
       (reset), .CLK (clk), .DIN (______9__32989), .QN
       (________________________________________0_));
  nnd2s1 ____0_502310(.DIN1 (_____0___32974), .DIN2 (______9__33037),
       .Q (______0__33038));
  and2s1 ____00_502311(.DIN1 (_________33316), .DIN2
       (______________22068), .Q (_________33036));
  or2s1 ____00_502312(.DIN1 (______________22068), .DIN2
       (_________33316), .Q (_________33035));
  nnd2s1 _____0_502313(.DIN1 (_____9___32964), .DIN2 (_________31935),
       .Q (_________33034));
  nnd2s1 ____0__502314(.DIN1 (_____00__32970), .DIN2 (_________33032),
       .Q (_________33033));
  or2s1 ____0__502315(.DIN1 (_________33030), .DIN2 (_________32983),
       .Q (_________33031));
  nnd2s1 ____0__502316(.DIN1 (_____99__32969), .DIN2 (______0__33028),
       .Q (_________33029));
  nnd2s1 ____0__502317(.DIN1 (_____0___32973), .DIN2 (_________33026),
       .Q (______9__33027));
  nnd2s1 ____0__502318(.DIN1 (_____9___32967), .DIN2 (_________32808),
       .Q (_________33025));
  and2s1 ___099_502319(.DIN1 (_________33006), .DIN2 (___0__0__40511),
       .Q (_________33024));
  and2s1 ____0__502320(.DIN1 (_____9___32963), .DIN2 (_________34531),
       .Q (_________33023));
  and2s1 ____0_502321(.DIN1 (_____9___32966), .DIN2 (____9____32417),
       .Q (_________33022));
  nnd2s1 ____0_502322(.DIN1 (_____0___32975), .DIN2 (_________33020),
       .Q (_________33021));
  nnd2s1 ____0__502323(.DIN1 (_____9___32961), .DIN2 (___90___29558),
       .Q (_________33019));
  and2s1 ____502324(.DIN1 (_____9___32962), .DIN2 (_________32898), .Q
       (______0__33018));
  nnd2s1 ____00_502325(.DIN1 (_________33011), .DIN2 (_____09__32979),
       .Q (_____9___33243));
  dffacs1 ____0___________________502326(.CLRB (reset), .CLK (clk),
       .DIN (_____0___32971), .QN (____0_________________21727));
  dffacs1 ______________________0_502327(.CLRB (reset), .CLK (clk),
       .DIN (_____90__32960), .QN (__________________0___21686));
  nnd2s1 ____502328(.DIN1 (_________32943), .DIN2 (_________33016), .Q
       (______9__33017));
  xor2s1 ___09__502329(.DIN1 (_________32915), .DIN2 (_____99__36913),
       .Q (_________33015));
  xor2s1 ___09__502330(.DIN1 (_________32913), .DIN2 (_________32761),
       .Q (_________33014));
  nor2s1 ___099_502331(.DIN1 (_________31928), .DIN2 (_________32952),
       .Q (_________33013));
  nor2s1 ___099_502332(.DIN1 (____9_9__38931), .DIN2 (_________33011),
       .Q (_________33012));
  xor2s1 ____502333(.DIN1 (_________32920), .DIN2 (_________38242), .Q
       (_________33010));
  or2s1 ____0__502334(.DIN1 (______0__33008), .DIN2 (_________32937),
       .Q (_________33009));
  nnd2s1 ____0__502335(.DIN1 (_________32944), .DIN2 (____99___32478),
       .Q (______9__33007));
  nor2s1 ____0__502336(.DIN1 (_____0___32875), .DIN2 (_________32945),
       .Q (_____9___33064));
  dffacs1 ________________________________________________502337(.CLRB
       (reset), .CLK (clk), .DIN (_________32957), .QN
       (__________________________________________________________________21989));
  dffacs1 ____0__________________502338(.CLRB (reset), .CLK (clk), .DIN
       (_________32935), .QN (____0________________21718));
  dffacs1 ____0__________________502339(.CLRB (reset), .CLK (clk), .DIN
       (_________32936), .QN (____0________________21716));
  nor2s1 ____0__502340(.DIN1 (_________32598), .DIN2 (_________32941),
       .Q (_________33005));
  nnd2s1 ____0__502341(.DIN1 (_________32932), .DIN2 (_________31831),
       .Q (_________33004));
  nor2s1 _____0_502342(.DIN1 (_________33002), .DIN2 (______9__32939),
       .Q (_________33003));
  nnd2s1 _____0_502343(.DIN1 (_________32933), .DIN2 (_________33000),
       .Q (_________33001));
  nnd2s1 _____0_502344(.DIN1 (_________32942), .DIN2 (______9__32998),
       .Q (______0__32999));
  nnd2s1 ____0__502345(.DIN1 (_________32953), .DIN2 (____0____32534),
       .Q (_________32997));
  nor2s1 _______502346(.DIN1 (________28991), .DIN2 (______9__32929),
       .Q (_________32996));
  nor2s1 _______502347(.DIN1 (__9_____29979), .DIN2 (_________32928),
       .Q (_________32995));
  nor2s1 _______502348(.DIN1 (_________32105), .DIN2 (_________32927),
       .Q (_________32994));
  nnd2s1 ____0__502349(.DIN1 (_________32938), .DIN2 (________28585),
       .Q (_________32993));
  nnd2s1 ______502350(.DIN1 (_________32948), .DIN2 (___0__0__40413),
       .Q (_________33054));
  dffacs1 _______________________502351(.CLRB (reset), .CLK (clk), .DIN
       (_________32934), .QN (_____________________21694));
  dffacs1 ________________________502352(.CLRB (reset), .CLK (clk),
       .DIN (______0__32930), .QN (______________________21698));
  dffacs1 _____________________0_502353(.CLRB (reset), .CLK (clk), .DIN
       (_________32955), .QN (_________________0___21740));
  xor2s1 ___09_502354(.DIN1 (_____09__32881), .DIN2 (_________34167),
       .Q (_________32992));
  or2s1 ___09_502355(.DIN1 (______0__32990), .DIN2 (_________32924), .Q
       (_________32991));
  nor2s1 ___099_502356(.DIN1 (____0____33482), .DIN2 (_________32916),
       .Q (______9__32989));
  nor2s1 ___0999(.DIN1 (_________32987), .DIN2 (_________32917), .Q
       (_________32988));
  nnd2s1 ____00_502357(.DIN1 (_________32985), .DIN2 (_____0___32978),
       .Q (_________32986));
  nor2s1 ____0__502358(.DIN1 (______0__32606), .DIN2 (______0__32912),
       .Q (_________32984));
  or2s1 ____0__502359(.DIN1 (_________32982), .DIN2 (_________32905),
       .Q (_________32983));
  nnd2s1 ____0__502360(.DIN1 (_________32906), .DIN2 (______0__32980),
       .Q (_________32981));
  nnd2s1 ____0__502361(.DIN1 (_________32909), .DIN2 (_________31617),
       .Q (_____09__32979));
  hi1s1 ___09__502362(.DIN (_________33840), .Q (_________33783));
  and2s1 ____00_502363(.DIN1 (_____0___32978), .DIN2 (_____0___32977),
       .Q (_________33044));
  xor2s1 ____0__502364(.DIN1 (_____0___32876), .DIN2
       (______________________________________________________________________________________0__22096),
       .Q (_________33316));
  hi1s1 ____0__502365(.DIN (_____0___32976), .Q (_________33006));
  nor2s1 _______502366(.DIN1 (_____09__31999), .DIN2 (_________32894),
       .Q (_____0___32975));
  and2s1 ____0__502367(.DIN1 (_________32896), .DIN2 (______0__33028),
       .Q (_____0___32974));
  nor2s1 ____0__502368(.DIN1 (__9_____30292), .DIN2 (______9__32901),
       .Q (_____0___32973));
  nor2s1 _____0_502369(.DIN1 (________26614), .DIN2 (_________32926),
       .Q (_____0___32972));
  or2s1 ______502370(.DIN1 (______0__33008), .DIN2 (_________32897), .Q
       (_____0___32971));
  nor2s1 _______502371(.DIN1 (_________32818), .DIN2 (_________32900),
       .Q (_____00__32970));
  and2s1 ____0__502372(.DIN1 (_________32925), .DIN2 (_____9___32968),
       .Q (_____99__32969));
  nor2s1 ____0__502373(.DIN1 (______9__32703), .DIN2 (______0__32902),
       .Q (_____9___32967));
  and2s1 _______502374(.DIN1 (_________32893), .DIN2 (_____9___32965),
       .Q (_____9___32966));
  nor2s1 _______502375(.DIN1 (___0__9__31347), .DIN2 (______9__32891),
       .Q (_____9___32964));
  nor2s1 _______502376(.DIN1 (_________32854), .DIN2 (_________32890),
       .Q (_____9___32963));
  nor2s1 _______502377(.DIN1 (_________31665), .DIN2 (_________32889),
       .Q (_____9___32962));
  nor2s1 _______502378(.DIN1 (____9____32439), .DIN2 (_________32895),
       .Q (_____9___32961));
  nnd2s1 ______502379(.DIN1 (_________32888), .DIN2 (______0__32980),
       .Q (_____90__32960));
  nnd2s1 _______502380(.DIN1 (_________32947), .DIN2 (______9__32959),
       .Q (_________33053));
  dffacs1 ________________________502381(.CLRB (reset), .CLK (clk),
       .DIN (_________32899), .QN (______________________21751));
  xor2s1 ____0__502382(.DIN1 (_____0__26159), .DIN2 (____900__34287),
       .Q (_________32958));
  or2s1 ___09__502383(.DIN1 (_________32886), .DIN2 (_________32956),
       .Q (_________32957));
  nnd2s1 ______502384(.DIN1 (_________32860), .DIN2 (_____9___41208),
       .Q (_________32955));
  xor2s1 ____00_502385(.DIN1 (________24494), .DIN2 (_________32923),
       .Q (_________32954));
  and2s1 _______502386(.DIN1 (_____9___32866), .DIN2 (_________31944),
       .Q (_________32953));
  and2s1 ____0_502387(.DIN1 (_________32887), .DIN2 (_________32951),
       .Q (_________32952));
  and2s1 ____0__502388(.DIN1 (_____0___32878), .DIN2 (______9__32949),
       .Q (______0__32950));
  hi1s1 _______502389(.DIN (_________32947), .Q (_________32948));
  xor2s1 ____0_502390(.DIN1 (______9__32911), .DIN2 (_________37687),
       .Q (_________32946));
  nor2s1 _______502391(.DIN1 (______0__34897), .DIN2 (_____00__32872),
       .Q (_________32945));
  nor2s1 ____09_502392(.DIN1 (_____0___32780), .DIN2 (_____0___32873),
       .Q (_________32944));
  and2s1 ____0__502393(.DIN1 (_____0___32874), .DIN2 (____9____34322),
       .Q (_________32943));
  xor2s1 ____0__502394(.DIN1 (______0__32793), .DIN2 (______9__32832),
       .Q (_____0___32976));
  nnd2s1 ____0__502395(.DIN1 (_________32908), .DIN2 (______0__32843),
       .Q (_________33011));
  xor2s1 ___09__502396(.DIN1 (_________32845), .DIN2 (___0_____40308),
       .Q (_________33840));
  nor2s1 ____00_502397(.DIN1 (_________32762), .DIN2 (_________32883),
       .Q (_________33289));
  dffacs1 _____________________________________________0_502398(.CLRB
       (reset), .CLK (clk), .DIN (_________32884), .QN
       (_______________________________________________________________0));
  dffacs1 ________________________________________________502399(.CLRB
       (reset), .CLK (clk), .DIN (_________32885), .QN
       (______________________________________________21906));
  and2s1 _______502400(.DIN1 (_________32859), .DIN2 (______0__32940),
       .Q (_________32942));
  nnd2s1 _______502401(.DIN1 (_________32857), .DIN2 (______0__32940),
       .Q (_________32941));
  nnd2s1 ______502402(.DIN1 (_____9___32863), .DIN2 (______9__32615),
       .Q (______9__32939));
  nor2s1 _______502403(.DIN1 (____0_9__31542), .DIN2 (_____9___32867),
       .Q (_________32938));
  nnd2s1 _______502404(.DIN1 (_____9___32864), .DIN2 (____0____32499),
       .Q (_________32937));
  or2s1 _______502405(.DIN1 (______0__33008), .DIN2 (_____9___32865),
       .Q (_________32936));
  nnd2s1 _______502406(.DIN1 (_________32858), .DIN2 (_____9___34752),
       .Q (_________32935));
  nnd2s1 _______502407(.DIN1 (_________32855), .DIN2 (_____9__28157),
       .Q (_________32934));
  nor2s1 _______502408(.DIN1 (______0__31950), .DIN2 (_____9___32869),
       .Q (_________32933));
  nor2s1 _______502409(.DIN1 (_________32931), .DIN2 (______0__32853),
       .Q (_________32932));
  or2s1 _______502410(.DIN1 (_________33175), .DIN2 (______9__32861),
       .Q (______0__32930));
  nnd2s1 _____0_502411(.DIN1 (_________32851), .DIN2 (__9__0__30003),
       .Q (______9__32929));
  nnd2s1 ______502412(.DIN1 (_________32849), .DIN2 (_________32797),
       .Q (_________32928));
  nnd2s1 _______502413(.DIN1 (_________32850), .DIN2 (_________31873),
       .Q (_________32927));
  dffacs1 _____________________9_502414(.CLRB (reset), .CLK (clk), .DIN
       (_____0___32877), .QN (_________________9___21696));
  dffacs1 _______________________502415(.CLRB (reset), .CLK (clk), .DIN
       (_____9___32870), .QN (_____________________21747));
  dffacs1 _______________________502416(.CLRB (reset), .CLK (clk), .DIN
       (_____90__32862), .QN (_____________________21690));
  dffacs1 _____________________9_502417(.CLRB (reset), .CLK (clk), .DIN
       (_________32856), .QN (_________________9___21749));
  nnd2s1 ______502418(.DIN1 (_________32829), .DIN2 (________29023), .Q
       (_________32926));
  and2s1 _______502419(.DIN1 (_________32835), .DIN2 (_________32347),
       .Q (_________32925));
  nor2s1 ____0__502420(.DIN1 (___0__9__40580), .DIN2 (_________32923),
       .Q (_________32924));
  nnd2s1 ____0__502421(.DIN1 (_________32923), .DIN2 (___0__9__40580),
       .Q (_________32922));
  nnd2s1 _______502422(.DIN1 (____0____33475), .DIN2 (_________32918),
       .Q (_________32920));
  nor2s1 _______502423(.DIN1 (_________32918), .DIN2 (____0____33475),
       .Q (_________32919));
  nor2s1 ____0__502424(.DIN1 (_____99__32871), .DIN2 (_________32844),
       .Q (_________32917));
  xor2s1 ____0__502425(.DIN1 (___0__0__40581), .DIN2 (_________32914),
       .Q (_________32916));
  xor2s1 ____0__502426(.DIN1 (___0_____40493), .DIN2 (_________32914),
       .Q (_________32915));
  xor2s1 ____0__502427(.DIN1 (_________32800), .DIN2 (______0__32882),
       .Q (_________32913));
  nor2s1 ____0__502428(.DIN1 (______9__32605), .DIN2 (______9__32911),
       .Q (______0__32912));
  nor2s1 ____0__502429(.DIN1 (___0_____40502), .DIN2 (____900__34287),
       .Q (_________32910));
  hi1s1 ____09_502430(.DIN (_________32908), .Q (_________32909));
  and2s1 ____09_502431(.DIN1 (____900__34287), .DIN2 (___0_____40502),
       .Q (_________32907));
  nor2s1 _____0_502432(.DIN1 (___0_____30683), .DIN2 (______0__32833),
       .Q (_________32906));
  nnd2s1 ____0_502433(.DIN1 (_________32923), .DIN2
       (____________________________________________21846), .Q
       (_________32985));
  or2s1 ____0_502434(.DIN1
       (____________________________________________21846), .DIN2
       (_________32923), .Q (_____0___32978));
  dffacs2 _______________________502435(.CLRB (reset), .CLK (clk), .DIN
       (_________32839), .Q (_____________________21742));
  dffacs1 ________________________502436(.CLRB (reset), .CLK (clk),
       .DIN (_________32827), .QN (______________________21752));
  or2s1 _______502437(.DIN1 (_____9__29074), .DIN2 (_________32837), .Q
       (_________32905));
  nor2s1 _______502438(.DIN1 (_________32903), .DIN2 (_________32838),
       .Q (_________32904));
  nnd2s1 ______502439(.DIN1 (_________32828), .DIN2 (__990___30456), .Q
       (______0__32902));
  nnd2s1 _______502440(.DIN1 (_________32848), .DIN2 (___0_____30675),
       .Q (______9__32901));
  nnd2s1 _______502441(.DIN1 (_________32847), .DIN2 (___0_____31160),
       .Q (_________32900));
  nnd2s1 _______502442(.DIN1 (_________32826), .DIN2 (_________32898),
       .Q (_________32899));
  nnd2s1 ______502443(.DIN1 (_________32809), .DIN2 (_________33193),
       .Q (_________32897));
  nor2s1 _______502444(.DIN1 (__9_____30053), .DIN2 (_________32846),
       .Q (_________32896));
  nnd2s1 _____9_502445(.DIN1 (_________32817), .DIN2 (_____0__28881),
       .Q (_________32895));
  or2s1 ______502446(.DIN1 (_________33849), .DIN2 (_________32824), .Q
       (_________32894));
  nor2s1 _______502447(.DIN1 (______0__32892), .DIN2 (______9__32812),
       .Q (_________32893));
  nnd2s1 _______502448(.DIN1 (_________32816), .DIN2 (___0_____30676),
       .Q (______9__32891));
  nnd2s1 _______502449(.DIN1 (_________32814), .DIN2 (___0_____30752),
       .Q (_________32890));
  nnd2s1 _______502450(.DIN1 (_________32810), .DIN2 (_____0___32284),
       .Q (_________32889));
  nor2s1 _______502451(.DIN1 (___0_____30967), .DIN2 (______0__32813),
       .Q (_________32888));
  nnd2s1 _______502452(.DIN1 (_________32841), .DIN2 (__9___22167), .Q
       (_________32947));
  dffacs1 ______________________0_502453(.CLRB (reset), .CLK (clk),
       .DIN (______9__32822), .QN (__________________0___21738));
  dffacs1 _____________________9_502454(.CLRB (reset), .CLK (clk), .DIN
       (_________32830), .QN (_________________9___21711));
  dffacs1 ________________________502455(.CLRB (reset), .CLK (clk),
       .DIN (_________32825), .QN (______________________21753));
  dffacs1 ______________________0_502456(.CLRB (reset), .CLK (clk),
       .DIN (_________32820), .QN (__________________0_));
  dffacs1 _______________________502457(.CLRB (reset), .CLK (clk), .DIN
       (_________32819), .QN (_____________________21743));
  nnd2s1 _______502458(.DIN1 (_________32796), .DIN2 (____0_9__32507),
       .Q (_________32887));
  nnd2s1 ___09__502459(.DIN1 (________24331), .DIN2 (_________32804),
       .Q (_________32886));
  nnd2s1 ____0__502460(.DIN1 (______9__32802), .DIN2 (________24432),
       .Q (_________32885));
  nnd2s1 ____0_502461(.DIN1 (_________32799), .DIN2 (________27094), .Q
       (_________32884));
  nor2s1 ____0__502462(.DIN1 (_________32801), .DIN2 (______0__32882),
       .Q (_________32883));
  xor2s1 ____0_502463(.DIN1 (_________32831), .DIN2 (______0__37673),
       .Q (_____09__32881));
  nor2s1 ____0_502464(.DIN1
       (____________________________________________21820), .DIN2
       (_________34626), .Q (_____0___32880));
  and2s1 ____0_502465(.DIN1 (_________34626), .DIN2
       (____________________________________________21820), .Q
       (_____0___32879));
  nor2s1 _______502466(.DIN1 (_____99__31989), .DIN2 (_________32807),
       .Q (_____0___32878));
  nnd2s1 _____9_502467(.DIN1 (_____0___32776), .DIN2 (_________32649),
       .Q (_____0___32877));
  xor2s1 _______502468(.DIN1 (_________32840), .DIN2 (_____9___33157),
       .Q (_____0___32876));
  nor2s1 _______502469(.DIN1 (___9_____39627), .DIN2 (_________32794),
       .Q (_____0___32875));
  and2s1 _______502470(.DIN1 (_________32791), .DIN2 (____0____32524),
       .Q (_____0___32874));
  nnd2s1 _______502471(.DIN1 (_________32789), .DIN2 (________29058),
       .Q (_____0___32873));
  nor2s1 _______502472(.DIN1 (___0____22291), .DIN2 (_________32790),
       .Q (_____00__32872));
  nor2s1 _______502473(.DIN1 (________22394), .DIN2 (_________32914),
       .Q (_____0___32977));
  nor2s1 _______502474(.DIN1 (_____99__32871), .DIN2 (______9__32842),
       .Q (_________32908));
  dffacs1 _______________________502475(.CLRB (reset), .CLK (clk), .DIN
       (_____9___32769), .QN (_____________________21748));
  nnd2s1 _______502476(.DIN1 (_________40938), .DIN2 (_________32898),
       .Q (_____9___32870));
  nnd2s1 _____502477(.DIN1 (_________32785), .DIN2 (_____9___32868), .Q
       (_____9___32869));
  nnd2s1 _____0_502478(.DIN1 (_________32784), .DIN2 (________29246),
       .Q (_____9___32867));
  nor2s1 _____502479(.DIN1 (_____9___31690), .DIN2 (______0__32783), .Q
       (_____9___32866));
  nnd2s1 _______502480(.DIN1 (_____0___32781), .DIN2 (______9__32998),
       .Q (_____9___32865));
  nor2s1 _______502481(.DIN1 (________28161), .DIN2 (_____0___32779),
       .Q (_____9___32864));
  nor2s1 _______502482(.DIN1 (___0_____31010), .DIN2 (_____0___32778),
       .Q (_____9___32863));
  nnd2s1 ______502483(.DIN1 (_________32805), .DIN2 (_____0__29107), .Q
       (_____90__32862));
  nnd2s1 ______502484(.DIN1 (_____99__32773), .DIN2 (__99____30490), .Q
       (______9__32861));
  and2s1 _____9_502485(.DIN1 (_____0___32774), .DIN2 (___0_____31075),
       .Q (_________32860));
  nor2s1 _______502486(.DIN1 (___0_____31100), .DIN2 (_____9___32770),
       .Q (_________32859));
  nor2s1 ______502487(.DIN1 (_____00__33249), .DIN2 (_____9___32767),
       .Q (_________32858));
  nor2s1 _______502488(.DIN1 (_________32218), .DIN2 (_____09__32782),
       .Q (_________32857));
  nnd2s1 _______502489(.DIN1 (_____9___32772), .DIN2 (_____9___41208),
       .Q (_________32856));
  nor2s1 ______502490(.DIN1 (_________32854), .DIN2 (_________32798),
       .Q (_________32855));
  or2s1 _______502491(.DIN1 (______9__32852), .DIN2 (_____9___32768),
       .Q (______0__32853));
  nor2s1 _______502492(.DIN1 (________28573), .DIN2 (_____9___32765),
       .Q (_________32851));
  nor2s1 _______502493(.DIN1 (__9_00), .DIN2 (_____9___32766), .Q
       (_________32850));
  nor2s1 _______502494(.DIN1 (__9_____30247), .DIN2 (_____90__32764),
       .Q (_________32849));
  nor2s1 _______502495(.DIN1 (__9_____30409), .DIN2 (_________32760),
       .Q (_________32848));
  nor2s1 _______502496(.DIN1 (_____9___31793), .DIN2 (_________32736),
       .Q (_________32847));
  nnd2s1 _______502497(.DIN1 (_________32752), .DIN2 (____0___28019),
       .Q (_________32846));
  xor2s1 ____0__502498(.DIN1 (_________32710), .DIN2
       (_______________22069), .Q (_________32845));
  nor2s1 _______502499(.DIN1 (______0__32843), .DIN2 (______9__32842),
       .Q (_________32844));
  nnd2s1 _____0_502500(.DIN1 (_________32840), .DIN2 (________22515),
       .Q (_________32841));
  nnd2s1 _____0_502501(.DIN1 (_________32747), .DIN2 (_________33032),
       .Q (_________32839));
  nnd2s1 _____0_502502(.DIN1 (_________32749), .DIN2 (____9____33393),
       .Q (_________32838));
  or2s1 _____502503(.DIN1 (_________32836), .DIN2 (_________32751), .Q
       (_________32837));
  nor2s1 _____9_502504(.DIN1 (_________32834), .DIN2 (_________32737),
       .Q (_________32835));
  nor2s1 _______502505(.DIN1 (_________33897), .DIN2 (_________32756),
       .Q (______0__32833));
  xor2s1 _______502506(.DIN1 (______9__32792), .DIN2 (_________38306),
       .Q (______9__32832));
  nor2s1 ______502507(.DIN1 (____0____32503), .DIN2 (_________32757),
       .Q (______9__32911));
  nnd2s1 _______502508(.DIN1 (_________32786), .DIN2 (___0__0__40581),
       .Q (______0__32990));
  nnd2s1 ______502509(.DIN1 (_________32831), .DIN2 (_____9___32278),
       .Q (______9__32921));
  xor2s1 _______502510(.DIN1 (_________33080), .DIN2 (_________32706),
       .Q (_________32923));
  hi1s1 _______502511(.DIN (_________34626), .Q (____900__34287));
  dffacs1 _______________________502512(.CLRB (reset), .CLK (clk), .DIN
       (_________32730), .QN (_____________________21671));
  xor2s1 _____9_502513(.DIN1 (_________32699), .DIN2 (___0__0__40413),
       .Q (____0____33475));
  dffacs1 ________________________502514(.CLRB (reset), .CLK (clk),
       .DIN (_________32745), .QN (______________________21701));
  dffacs1 _______________________502515(.CLRB (reset), .CLK (clk), .DIN
       (______9__32743), .QN (_____________________21745));
  nnd2s1 _______502516(.DIN1 (_________32739), .DIN2 (_________34163),
       .Q (_________32830));
  nor2s1 _______502517(.DIN1 (_____0__29028), .DIN2 (_________32741),
       .Q (_________32829));
  nor2s1 _______502518(.DIN1 (__9_____30252), .DIN2 (_________32735),
       .Q (_________32828));
  nnd2s1 _______502519(.DIN1 (_________32758), .DIN2 (_____9___41208),
       .Q (_________32827));
  nor2s1 _______502520(.DIN1 (_________32746), .DIN2 (_________32742),
       .Q (_________32826));
  nnd2s1 _______502521(.DIN1 (_________32759), .DIN2 (________28869),
       .Q (_________32825));
  or2s1 _______502522(.DIN1 (______0__32823), .DIN2 (_________32731),
       .Q (_________32824));
  nnd2s1 _______502523(.DIN1 (_________32729), .DIN2 (______0__32646),
       .Q (______9__32822));
  nor2s1 _______502524(.DIN1 (________26296), .DIN2 (_________32728),
       .Q (_________32821));
  nnd2s1 ______502525(.DIN1 (_________32726), .DIN2 (_____0___32676),
       .Q (_________32820));
  or2s1 _______502526(.DIN1 (_________32818), .DIN2 (_________32718),
       .Q (_________32819));
  nor2s1 _______502527(.DIN1 (________27550), .DIN2 (_________32727),
       .Q (_________32817));
  nor2s1 _______502528(.DIN1 (_________32815), .DIN2 (______0__32724),
       .Q (_________32816));
  nor2s1 _____502529(.DIN1 (__9_____30067), .DIN2 (_________32722), .Q
       (_________32814));
  nnd2s1 _______502530(.DIN1 (_________32725), .DIN2 (_________32018),
       .Q (______0__32813));
  nnd2s1 _______502531(.DIN1 (_________32721), .DIN2 (_________32811),
       .Q (______9__32812));
  nnd2s1 _______502532(.DIN1 (_________32719), .DIN2 (____0____32543),
       .Q (_________32810));
  and2s1 _______502533(.DIN1 (______9__32763), .DIN2 (_________32808),
       .Q (_________32809));
  dffacs1 ________________________502534(.CLRB (reset), .CLK (clk),
       .DIN (______0__32734), .QN (______________________21739));
  dffacs1 _______________________502535(.CLRB (reset), .CLK (clk), .DIN
       (______9__32723), .QN (_____________________21746));
  dffacs1 _______________________502536(.CLRB (reset), .CLK (clk), .DIN
       (_________32732), .QN (_____________________21683));
  or2s1 _______502537(.DIN1 (_________32806), .DIN2 (_________32788),
       .Q (_________32807));
  and2s1 _______502538(.DIN1 (_________32691), .DIN2 (________29482),
       .Q (_________32805));
  nnd2s1 ____0__502539(.DIN1 (______0__32803), .DIN2 (_________32716),
       .Q (_________32804));
  nnd2s1 ____0__502540(.DIN1 (_________32715), .DIN2 (inData[26]), .Q
       (______9__32802));
  nor2s1 _____0_502541(.DIN1 (_________32800), .DIN2 (______0__32714),
       .Q (_________32801));
  nor2s1 _____0_502542(.DIN1 (____90__25398), .DIN2 (______9__32713),
       .Q (_________32799));
  nnd2s1 _______502543(.DIN1 (_________32689), .DIN2 (_________32797),
       .Q (_________32798));
  nnd2s1 ______502544(.DIN1 (_________32707), .DIN2 (_________32613),
       .Q (_________32796));
  nnd2s1 ______502545(.DIN1 (_________32787), .DIN2 (___9_____39582),
       .Q (_________32795));
  or2s1 _______502546(.DIN1 (______0__32793), .DIN2 (______9__32792),
       .Q (_________32794));
  and2s1 _______502547(.DIN1 (_________32702), .DIN2 (_____9___41206),
       .Q (_________32791));
  and2s1 _______502548(.DIN1 (______9__32792), .DIN2 (________22709),
       .Q (_________32790));
  and2s1 _____0_502549(.DIN1 (______0__32704), .DIN2 (___9____28726),
       .Q (_________32789));
  nor2s1 _______502550(.DIN1 (___0_9___31211), .DIN2 (_________32788),
       .Q (_____99__32871));
  nor2s1 ______502551(.DIN1 (______9__32665), .DIN2 (_________32787),
       .Q (______0__32882));
  dffacs2 ____0___________________502552(.CLRB (reset), .CLK (clk),
       .DIN (_________32698), .Q (____0_______________));
  hi1s1 ______502553(.DIN (_________32786), .Q (_________32914));
  xnr2s1 _____9_502554(.DIN1 (_______________22070), .DIN2
       (_________32657), .Q (_________34626));
  dffacs1 _______________________502555(.CLRB (reset), .CLK (clk), .DIN
       (_________32700), .QN (_____________________21709));
  and2s1 ______502556(.DIN1 (_____9___32672), .DIN2 (__99____30473), .Q
       (_________32785));
  nor2s1 _______502557(.DIN1 (__9_9___30449), .DIN2 (______9__32693),
       .Q (_________32784));
  nnd2s1 _______502558(.DIN1 (_________32705), .DIN2 (__9__0__29789),
       .Q (______0__32783));
  nnd2s1 _______502559(.DIN1 (_____0___32683), .DIN2 (___0_____30854),
       .Q (_____09__32782));
  nor2s1 _______502560(.DIN1 (_____0___32780), .DIN2 (_________32709),
       .Q (_____0___32781));
  nnd2s1 _______502561(.DIN1 (_________32717), .DIN2 (________27233),
       .Q (_____0___32779));
  or2s1 _____0_502562(.DIN1 (_____0___32777), .DIN2 (_____0___32680),
       .Q (_____0___32778));
  nor2s1 _____0_502563(.DIN1 (_____0___32775), .DIN2 (_____0___32682),
       .Q (_____0___32776));
  nor2s1 _____0_502564(.DIN1 (_____09__32684), .DIN2 (____0_9__32526),
       .Q (_____0___32774));
  nor2s1 _______502565(.DIN1 (__9_____30415), .DIN2 (______0__32685),
       .Q (_____99__32773));
  nor2s1 _______502566(.DIN1 (_____9___32771), .DIN2 (_________32687),
       .Q (_____9___32772));
  nnd2s1 _______502567(.DIN1 (_____0___32681), .DIN2 (____0____32512),
       .Q (_____9___32770));
  nnd2s1 _______502568(.DIN1 (_____0___32678), .DIN2 (_________32055),
       .Q (_____9___32769));
  nnd2s1 _______502569(.DIN1 (_________32686), .DIN2 (________27633),
       .Q (_____9___32768));
  nnd2s1 _______502570(.DIN1 (_____0___32679), .DIN2 (___00____30578),
       .Q (_____9___32767));
  nnd2s1 _______502571(.DIN1 (_____0___32677), .DIN2 (____0___28838),
       .Q (_____9___32766));
  nnd2s1 _______502572(.DIN1 (_____99__32674), .DIN2 (________29309),
       .Q (_____9___32765));
  nnd2s1 ______502573(.DIN1 (_____00__32675), .DIN2 (___9____28684), .Q
       (_____90__32764));
  dffacs1 _______________________502574(.CLRB (reset), .CLK (clk), .DIN
       (_________32690), .QN (_____________________21730));
  nor2s1 _______502575(.DIN1 (__9_____30137), .DIN2 (_________32651),
       .Q (______9__32763));
  nor2s1 _______502576(.DIN1 (______0__32361), .DIN2 (_________32761),
       .Q (_________32762));
  nnd2s1 _______502577(.DIN1 (_________32648), .DIN2 (________29358),
       .Q (_________32760));
  nor2s1 _______502578(.DIN1 (____9____32404), .DIN2 (_________32622),
       .Q (_________32759));
  nor2s1 ______502579(.DIN1 (_________32308), .DIN2 (_________32643),
       .Q (_________32758));
  nnd2s1 _____0_502580(.DIN1 (_________32661), .DIN2 (____0____32502),
       .Q (_________32757));
  nor2s1 _____0_502581(.DIN1 (_________32755), .DIN2 (_________32659),
       .Q (_________32756));
  nnd2s1 ______502582(.DIN1 (_________32740), .DIN2 (______9__32753),
       .Q (______0__32754));
  and2s1 _______502583(.DIN1 (_________32650), .DIN2 (__9_____30354),
       .Q (_________32752));
  or2s1 _______502584(.DIN1 (_________32750), .DIN2 (_________32654),
       .Q (_________32751));
  nor2s1 _______502585(.DIN1 (_________32748), .DIN2 (_________32653),
       .Q (_________32749));
  nor2s1 ______502586(.DIN1 (_________32746), .DIN2 (______0__32656),
       .Q (_________32747));
  nnd2s1 _______502587(.DIN1 (_________32632), .DIN2 (______0__32744),
       .Q (_________32745));
  nnd2s1 _______502588(.DIN1 (_________32662), .DIN2 (____0____32532),
       .Q (______9__32743));
  nnd2s1 _______502589(.DIN1 (_________32652), .DIN2 (____0____32550),
       .Q (_________32742));
  or2s1 _______502590(.DIN1 (_________32267), .DIN2 (_________32740),
       .Q (_________32741));
  and2s1 ______502591(.DIN1 (_________32640), .DIN2 (_________32738),
       .Q (_________32739));
  nor2s1 _______502592(.DIN1 (___0__0__30842), .DIN2 (______0__32694),
       .Q (______9__32842));
  xor2s1 _____9_502593(.DIN1 (_________32612), .DIN2 (____0____37113),
       .Q (_________32786));
  nor2s1 ______502594(.DIN1 (______0__32010), .DIN2 (_____9___32668),
       .Q (_________32831));
  dffacs1 _______________________502595(.CLRB (reset), .CLK (clk), .DIN
       (_________32641), .QN (_____________________21729));
  nnd2s1 ______502596(.DIN1 (______9__32655), .DIN2 (____0___29100), .Q
       (_________32737));
  nor2s1 _______502597(.DIN1 (____0____32539), .DIN2 (_____9___32669),
       .Q (_________32736));
  nnd2s1 ______502598(.DIN1 (_________32642), .DIN2 (_________33096),
       .Q (_________32735));
  nnd2s1 _______502599(.DIN1 (_________32624), .DIN2 (______9__32733),
       .Q (______0__32734));
  nnd2s1 _______502600(.DIN1 (_________32637), .DIN2 (_________31626),
       .Q (_________32732));
  or2s1 ______502601(.DIN1 (______9__32009), .DIN2 (_________32631), .Q
       (_________32731));
  nnd2s1 _______502602(.DIN1 (______0__32636), .DIN2 (____9____32413),
       .Q (_________32730));
  nor2s1 _______502603(.DIN1 (_________32112), .DIN2 (_________32634),
       .Q (_________32729));
  nnd2s1 _______502604(.DIN1 (______9__32625), .DIN2 (__9_____29758),
       .Q (_________32728));
  nnd2s1 _______502605(.DIN1 (_________32627), .DIN2 (__9_____30218),
       .Q (_________32727));
  nor2s1 _______502606(.DIN1 (_________32364), .DIN2 (_________32623),
       .Q (_________32726));
  nnd2s1 _______502607(.DIN1 (_________32628), .DIN2 (______0__34524),
       .Q (_________32725));
  nnd2s1 _____9_502608(.DIN1 (_________32644), .DIN2 (__9_____30322),
       .Q (______0__32724));
  nnd2s1 _____9_502609(.DIN1 (_________32630), .DIN2 (_____9___41208),
       .Q (______9__32723));
  nnd2s1 _____9_502610(.DIN1 (______0__32626), .DIN2 (________28363),
       .Q (_________32722));
  and2s1 _____9_502611(.DIN1 (_________32629), .DIN2 (_________32720),
       .Q (_________32721));
  nnd2s1 _____0_502612(.DIN1 (_________32638), .DIN2 (_____0___41313),
       .Q (_________32719));
  nnd2s1 _____0_502613(.DIN1 (______9__32635), .DIN2 (___0_____31045),
       .Q (_________32718));
  nnd2s1 _______502614(.DIN1 (_____9___32671), .DIN2 (________28222),
       .Q (_________32840));
  dffacs1 _______________________502615(.CLRB (reset), .CLK (clk), .DIN
       (_________32647), .Q (_____________________21733));
  dffacs1 _______________________502616(.CLRB (reset), .CLK (clk), .DIN
       (_________32633), .QN (_____________________21741));
  nor2s1 _______502617(.DIN1 (_____0__29436), .DIN2 (______0__32586),
       .Q (_________32717));
  xor2s1 _____502618(.DIN1
       (______________________________________________21906), .DIN2
       (___0_____40613), .Q (_________32716));
  nor2s1 _______502619(.DIN1 (_________32711), .DIN2 (_____0___33165),
       .Q (_________32715));
  hi1s1 ______502620(.DIN (_________32761), .Q (______0__32714));
  and2s1 _______502621(.DIN1 (_________32712), .DIN2 (_________32711),
       .Q (______9__32713));
  xor2s1 _______502622(.DIN1 (_________32099), .DIN2 (_________40940),
       .Q (_________32710));
  nnd2s1 ______502623(.DIN1 (_________32600), .DIN2 (_________32349),
       .Q (_________32709));
  nor2s1 ______502624(.DIN1 (______9__36337), .DIN2 (_________32614),
       .Q (_________32708));
  nnd2s1 _______502625(.DIN1 (_________32695), .DIN2 (___9_____39582),
       .Q (_________32707));
  xnr2s1 ______502626(.DIN1
       (_________________________________________________________________________________________22092),
       .DIN2 (_________32660), .Q (_________32706));
  nor2s1 _______502627(.DIN1 (__9_____30095), .DIN2 (_________32601),
       .Q (_________32705));
  nor2s1 _______502628(.DIN1 (______9__32703), .DIN2 (_________32610),
       .Q (______0__32704));
  nor2s1 _______502629(.DIN1 (_________32701), .DIN2 (_________32607),
       .Q (_________32702));
  nnd2s1 _______502630(.DIN1 (_________32587), .DIN2 (__9_____30436),
       .Q (_________32700));
  xor2s1 ______502631(.DIN1 (_____9___32670), .DIN2
       (______________22068), .Q (_________32699));
  nnd2s1 _______502632(.DIN1 (_________32599), .DIN2 (_________33128),
       .Q (_________32698));
  nnd2s1 ______502633(.DIN1 (_________32589), .DIN2 (_________32696),
       .Q (_________32697));
  nor2s1 _______502634(.DIN1 (_________31710), .DIN2 (_________32695),
       .Q (_________32787));
  hi1s1 ______502635(.DIN (______0__32694), .Q (_________32788));
  nnd2s1 _____9_502636(.DIN1 (_________32609), .DIN2 (_______22230), .Q
       (______9__32792));
  dffacs2 _______________________502637(.CLRB (reset), .CLK (clk), .DIN
       (_____0___32584), .Q (_____________________21736));
  nnd2s1 _____0_502638(.DIN1 (_________32603), .DIN2 (_________32692),
       .Q (______9__32693));
  nor2s1 _______502639(.DIN1 (__9_____29830), .DIN2 (_________32619),
       .Q (_________32691));
  or2s1 _______502640(.DIN1 (_____0___32583), .DIN2 (_________32592),
       .Q (_________32690));
  nor2s1 _______502641(.DIN1 (_________32688), .DIN2 (_________32621),
       .Q (_________32689));
  nnd2s1 ______502642(.DIN1 (_________32591), .DIN2 (___0_____30941),
       .Q (_________32687));
  nor2s1 _____9_502643(.DIN1 (_________32130), .DIN2 (_________32590),
       .Q (_________32686));
  nnd2s1 _____502644(.DIN1 (_________32593), .DIN2 (____0___27574), .Q
       (______0__32685));
  nor2s1 _____502645(.DIN1 (___99___25116), .DIN2 (_________32594), .Q
       (_____09__32684));
  nor2s1 _______502646(.DIN1 (___0____27909), .DIN2 (______0__32616),
       .Q (_____0___32683));
  nnd2s1 _____0_502647(.DIN1 (_____09__32585), .DIN2 (__9_9___30358),
       .Q (_____0___32682));
  nor2s1 _______502648(.DIN1 (____09__29287), .DIN2 (_____0___32582),
       .Q (_____0___32681));
  nnd2s1 _______502649(.DIN1 (_____0___32581), .DIN2 (__9_____30248),
       .Q (_____0___32680));
  nor2s1 _______502650(.DIN1 (________27992), .DIN2 (_____0___32580),
       .Q (_____0___32679));
  nor2s1 ______502651(.DIN1 (_____0___32190), .DIN2 (_____0___32579),
       .Q (_____0___32678));
  and2s1 _______502652(.DIN1 (_____00__32576), .DIN2 (_____0___32676),
       .Q (_____0___32677));
  nor2s1 _______502653(.DIN1 (________29489), .DIN2 (____099__32575),
       .Q (_____00__32675));
  and2s1 _____0_502654(.DIN1 (____09___32574), .DIN2 (_____9___32673),
       .Q (_____99__32674));
  nor2s1 _______502655(.DIN1 (__9_____29883), .DIN2 (______9__32595),
       .Q (_____9___32672));
  dffacs2 _______________________502656(.CLRB (reset), .CLK (clk), .DIN
       (_____0___32578), .QN (___________________));
  dffacs1 ____0__________________502657(.CLRB (reset), .CLK (clk), .DIN
       (_________32588), .QN (____0________________21721));
  nnd2s1 _____9_502658(.DIN1 (_____9___32670), .DIN2 (________28142),
       .Q (_____9___32671));
  nor2s1 _____502659(.DIN1 (________29229), .DIN2 (____0_9__32556), .Q
       (_____9___32669));
  nor2s1 ______502660(.DIN1 (_________32011), .DIN2 (_________40940),
       .Q (_____9___32668));
  nor2s1 _______502661(.DIN1 (_________32663), .DIN2 (_____90__32666),
       .Q (_____9___32667));
  nor2s1 _______502662(.DIN1 (_________31630), .DIN2 (_________32597),
       .Q (______9__32665));
  and2s1 _______502663(.DIN1 (_____90__32666), .DIN2 (_________32663),
       .Q (_________32664));
  nor2s1 _______502664(.DIN1 (________29293), .DIN2 (____0____32561),
       .Q (_________32662));
  nnd2s1 ______502665(.DIN1 (_________32660), .DIN2 (_____9___32378),
       .Q (_________32661));
  or2s1 _______502666(.DIN1 (_________32658), .DIN2 (____0____32563),
       .Q (_________32659));
  xor2s1 _______502667(.DIN1 (_________32608), .DIN2 (_____9___33157),
       .Q (_________32657));
  or2s1 _______502668(.DIN1 (_____9___32771), .DIN2 (____09___32568),
       .Q (______0__32656));
  nor2s1 _______502669(.DIN1 (____0___29201), .DIN2 (____090__32567),
       .Q (______9__32655));
  nnd2s1 ______502670(.DIN1 (____0____32560), .DIN2 (___0_____31258),
       .Q (_________32654));
  nnd2s1 _______502671(.DIN1 (____0____32558), .DIN2 (___0_____31376),
       .Q (_________32653));
  nor2s1 _______502672(.DIN1 (___0_0___30930), .DIN2 (____0____32545),
       .Q (_________32652));
  nnd2s1 ______502673(.DIN1 (____0____32554), .DIN2 (___0_____30970),
       .Q (_________32651));
  and2s1 ______502674(.DIN1 (____0____32553), .DIN2 (_________32649),
       .Q (_________32650));
  nor2s1 _______502675(.DIN1 (___0____28753), .DIN2 (____0____32552),
       .Q (_________32648));
  nnd2s1 _______502676(.DIN1 (____0____32562), .DIN2 (______0__32646),
       .Q (_________32647));
  nnd2s1 _______502677(.DIN1 (_____90__32666), .DIN2 (____90___32385),
       .Q (______0__32694));
  nnd2s1 ______502678(.DIN1 (____0____32559), .DIN2 (______0__32196),
       .Q (_________32740));
  dffacs1 _______________________502679(.CLRB (reset), .CLK (clk), .DIN
       (____0_0__32547), .Q (_____________________21734));
  nnd2s1 _____502680(.DIN1 (______9__32645), .DIN2 (___0_____31333), .Q
       (_________32761));
  and2s1 _______502681(.DIN1 (____0____32520), .DIN2 (_________33931),
       .Q (_________32644));
  nnd2s1 _____0_502682(.DIN1 (____09___32569), .DIN2 (___0__0__31232),
       .Q (_________32643));
  nor2s1 _____0_502683(.DIN1 (____0___28476), .DIN2 (____0____32531),
       .Q (_________32642));
  nnd2s1 _______502684(.DIN1 (____09___32573), .DIN2 (_________33695),
       .Q (_________32641));
  and2s1 _______502685(.DIN1 (____0____32549), .DIN2 (_________32639),
       .Q (_________32640));
  nor2s1 _______502686(.DIN1 (_____0___31604), .DIN2 (____0_9__32536),
       .Q (_________32638));
  nor2s1 _______502687(.DIN1 (____0____32490), .DIN2 (____0____32538),
       .Q (_________32637));
  nor2s1 ______502688(.DIN1 (__909___29718), .DIN2 (____0_0__32537), .Q
       (______0__32636));
  nor2s1 _______502689(.DIN1 (___0__0__30891), .DIN2 (____0____32540),
       .Q (______9__32635));
  nnd2s1 ______502690(.DIN1 (____0____32530), .DIN2 (_________32116),
       .Q (_________32634));
  or2s1 _______502691(.DIN1 (_________32746), .DIN2 (____0____32551),
       .Q (_________32633));
  nor2s1 _____9_502692(.DIN1 (________29078), .DIN2 (____0____32555),
       .Q (_________32632));
  nor2s1 _______502693(.DIN1 (inData[31]), .DIN2 (____0____32519), .Q
       (_________32631));
  nor2s1 _______502694(.DIN1 (___09___27918), .DIN2 (____0____32533),
       .Q (_________32630));
  and2s1 _______502695(.DIN1 (____0____32525), .DIN2 (_____9___33329),
       .Q (_________32629));
  nnd2s1 _____9_502696(.DIN1 (____0____32523), .DIN2 (_________31781),
       .Q (_________32628));
  nnd2s1 _____0_502697(.DIN1 (____0____32522), .DIN2 (________25544),
       .Q (_________32627));
  nor2s1 _____0_502698(.DIN1 (___0_____30901), .DIN2 (____0____32542),
       .Q (______0__32626));
  nor2s1 _____0_502699(.DIN1 (________29336), .DIN2 (____0_0__32527),
       .Q (______9__32625));
  nor2s1 _____0_502700(.DIN1 (___0_____31252), .DIN2 (____0____32528),
       .Q (_________32624));
  nnd2s1 _______502701(.DIN1 (____0____32529), .DIN2 (_________32325),
       .Q (_________32623));
  nnd2s1 _____9_502702(.DIN1 (____0____32544), .DIN2 (_________32067),
       .Q (_________32622));
  dffacs1 _______________________502703(.CLRB (reset), .CLK (clk), .DIN
       (____0____32535), .QN (_____________________21673));
  nnd2s1 _______502704(.DIN1 (____009__32487), .DIN2 (___0_____30663),
       .Q (_________32621));
  nor2s1 _______502705(.DIN1 (_____9__26294), .DIN2 (____990__32470),
       .Q (_________32620));
  nnd2s1 _______502706(.DIN1 (____0____32514), .DIN2 (__9_99__30271),
       .Q (_________32619));
  nor2s1 _______502707(.DIN1 (____09___32570), .DIN2 (_________32617),
       .Q (_________32618));
  nnd2s1 _______502708(.DIN1 (____999__32479), .DIN2 (______9__32615),
       .Q (______0__32616));
  nnd2s1 _______502709(.DIN1 (____0_0__32508), .DIN2 (_________32613),
       .Q (_________32614));
  xor2s1 ______502710(.DIN1 (____9____32445), .DIN2 (_________32611),
       .Q (_________32612));
  nnd2s1 _______502711(.DIN1 (____0_0__32498), .DIN2 (__9_____30147),
       .Q (_________32610));
  nnd2s1 _______502712(.DIN1 (_________32608), .DIN2 (___0____22349),
       .Q (_________32609));
  nnd2s1 _______502713(.DIN1 (____0_9__32517), .DIN2 (_________41238),
       .Q (_________32607));
  and2s1 _____502714(.DIN1 (_________33201), .DIN2
       (______________22066), .Q (______0__32606));
  nor2s1 ______502715(.DIN1 (______________22066), .DIN2
       (_________33201), .Q (______9__32605));
  nor2s1 _______502716(.DIN1 (___0_____31244), .DIN2 (____0____32494),
       .Q (_________32604));
  nor2s1 _______502717(.DIN1 (_________32602), .DIN2 (____0_0__32488),
       .Q (_________32603));
  nnd2s1 _______502718(.DIN1 (____0_9__32497), .DIN2 (___0_____30905),
       .Q (_________32601));
  nor2s1 _______502719(.DIN1 (____9___28370), .DIN2 (____0____32496),
       .Q (_________32600));
  nor2s1 _______502720(.DIN1 (_________32598), .DIN2 (____0____32495),
       .Q (_________32599));
  hi1s1 _____9_502721(.DIN (___0_____40613), .Q (_________32711));
  hi1s1 _____0_502722(.DIN (_________32597), .Q (_________32695));
  dffacs1 ______________________________________________9_502723(.CLRB
       (reset), .CLK (clk), .DIN (____0____32509), .Q
       (__________________________________________9_));
  dffacs1 ____0__________________502724(.CLRB (reset), .CLK (clk), .DIN
       (____0____32500), .QN (____0________________21717));
  nor2s1 _____502725(.DIN1 (_________32001), .DIN2 (____99___32471), .Q
       (______0__32596));
  nnd2s1 _______502726(.DIN1 (____0____32491), .DIN2 (___0_____30719),
       .Q (______9__32595));
  nor2s1 _______502727(.DIN1 (______0__41140), .DIN2 (____00___32486),
       .Q (_________32594));
  nor2s1 _______502728(.DIN1 (__99_0__30499), .DIN2 (____99___32474),
       .Q (_________32593));
  nnd2s1 _______502729(.DIN1 (____99___32477), .DIN2 (___0__0__31222),
       .Q (_________32592));
  nor2s1 ______502730(.DIN1 (______9__31775), .DIN2 (____00___32484),
       .Q (_________32591));
  nnd2s1 ______502731(.DIN1 (____99___32475), .DIN2 (___9_9__29627), .Q
       (_________32590));
  nor2s1 _______502732(.DIN1 (________26739), .DIN2 (____0____32493),
       .Q (_________32589));
  nnd2s1 _______502733(.DIN1 (____0____32513), .DIN2 (_________32808),
       .Q (_________32588));
  nor2s1 ______502734(.DIN1 (________28245), .DIN2 (____0____32492), .Q
       (_________32587));
  nor2s1 _____9_502735(.DIN1 (___0____25136), .DIN2 (____99___32473),
       .Q (______0__32586));
  nor2s1 ______502736(.DIN1 (___9____29591), .DIN2 (____99___32476), .Q
       (_____09__32585));
  or2s1 _____0_502737(.DIN1 (_____0___32583), .DIN2 (____00___32482),
       .Q (_____0___32584));
  nnd2s1 _____0_502738(.DIN1 (____00___32483), .DIN2 (____0___29103),
       .Q (_____0___32582));
  nor2s1 _____0_502739(.DIN1 (___0_____31337), .DIN2 (____00___32481),
       .Q (_____0___32581));
  nnd2s1 _____502740(.DIN1 (____0____32489), .DIN2 (___0_____31230), .Q
       (_____0___32580));
  nor2s1 _______502741(.DIN1 (___0__9__30890), .DIN2 (____99___32472),
       .Q (_____0___32579));
  nnd2s1 _______502742(.DIN1 (____9____32467), .DIN2 (_____0___32577),
       .Q (_____0___32578));
  and2s1 _______502743(.DIN1 (____9____32468), .DIN2 (__99____30520),
       .Q (_____00__32576));
  nnd2s1 _______502744(.DIN1 (____9____32465), .DIN2 (________29392),
       .Q (____099__32575));
  nor2s1 _______502745(.DIN1 (__9__0__30093), .DIN2 (____9_9__32469),
       .Q (____09___32574));
  dffacs1 _______________________502746(.CLRB (reset), .CLK (clk), .DIN
       (____9____32466), .QN (_____________________21672));
  nor2s1 _______502747(.DIN1 (____9_0__32451), .DIN2 (______0__32341),
       .Q (____09___32573));
  nnd2s1 _____502748(.DIN1 (____9____32435), .DIN2 (________25733), .Q
       (____09___32572));
  xor2s1 _______502749(.DIN1 (________25249), .DIN2 (____0____32510),
       .Q (____09___32571));
  nnd2s1 _______502750(.DIN1 (____9____32429), .DIN2 (________26299),
       .Q (____09___32569));
  nnd2s1 _______502751(.DIN1 (____9____32428), .DIN2 (___0_____31052),
       .Q (____09___32568));
  nnd2s1 _______502752(.DIN1 (____9____32408), .DIN2 (__9_____30070),
       .Q (____090__32567));
  nnd2s1 ______502753(.DIN1 (____0____32565), .DIN2 (____0____32564),
       .Q (____0_9__32566));
  nnd2s1 _______502754(.DIN1 (____9____32447), .DIN2 (______9__31632),
       .Q (____0____32563));
  nor2s1 _______502755(.DIN1 (_____0___31898), .DIN2 (____9____32448),
       .Q (____0____32562));
  nnd2s1 _______502756(.DIN1 (____9____32442), .DIN2 (_________31916),
       .Q (____0____32561));
  nor2s1 ______502757(.DIN1 (___0_____31198), .DIN2 (____9____32438),
       .Q (____0____32560));
  nor2s1 _______502758(.DIN1 (______9__31884), .DIN2 (____9____32463),
       .Q (____0____32559));
  nor2s1 _______502759(.DIN1 (____0_0__32557), .DIN2 (____9____32437),
       .Q (____0____32558));
  nnd2s1 ______502760(.DIN1 (____9_0__32441), .DIN2 (___0_9___31403),
       .Q (____0_9__32556));
  nnd2s1 _______502761(.DIN1 (____9_9__32440), .DIN2 (___9____29588),
       .Q (____0____32555));
  and2s1 _______502762(.DIN1 (____9____32425), .DIN2 (___0_____30800),
       .Q (____0____32554));
  and2s1 _______502763(.DIN1 (____9_0__32431), .DIN2 (______9__31910),
       .Q (____0____32553));
  nor2s1 _______502764(.DIN1 (____0____32541), .DIN2 (____9_9__32450),
       .Q (____0____32552));
  xnr2s1 _______502765(.DIN1 (_________32613), .DIN2 (_________32951),
       .Q (_________32597));
  xor2s1 ______502766(.DIN1 (____90___32388), .DIN2 (_________32613),
       .Q (______9__32645));
  nnd2s1 _______502767(.DIN1 (____9____32464), .DIN2 (____9____32443),
       .Q (_________32660));
  dffacs1 _____________________________________________0_502768(.CLRB
       (reset), .CLK (clk), .DIN (____9____32462), .QN
       (___0_____40613));
  xor2s1 _______502769(.DIN1 (____90___32383), .DIN2 (___9_____39554),
       .Q (_____90__32666));
  nnd2s1 _______502770(.DIN1 (____9____32409), .DIN2 (____0____32550),
       .Q (____0____32551));
  nor2s1 _____9_502771(.DIN1 (____0____32548), .DIN2 (____9____32427),
       .Q (____0____32549));
  nnd2s1 _____9_502772(.DIN1 (____9____32419), .DIN2 (_________31848),
       .Q (____0_0__32547));
  nnd2s1 _____502773(.DIN1 (____9____32418), .DIN2 (______0__41180), .Q
       (____0_9__32546));
  nnd2s1 _______502774(.DIN1 (_________31977), .DIN2 (____9____32416),
       .Q (____0____32545));
  nnd2s1 _______502775(.DIN1 (____9____32423), .DIN2 (____0____32543),
       .Q (____0____32544));
  nor2s1 _______502776(.DIN1 (____0____32541), .DIN2 (____9____32393),
       .Q (____0____32542));
  nor2s1 _______502777(.DIN1 (____0____32539), .DIN2 (____9_9__32430),
       .Q (____0____32540));
  nor2s1 _______502778(.DIN1 (_____9___32376), .DIN2 (____9____32397),
       .Q (____0____32538));
  nnd2s1 _______502779(.DIN1 (____9____32405), .DIN2 (_____9__29324),
       .Q (____0_0__32537));
  nnd2s1 ______502780(.DIN1 (____9____32403), .DIN2 (___0__0__31290),
       .Q (____0_9__32536));
  nnd2s1 ______502781(.DIN1 (____9____32414), .DIN2 (____0____32534),
       .Q (____0____32535));
  nnd2s1 _______502782(.DIN1 (____9____32406), .DIN2 (____0____32532),
       .Q (____0____32533));
  nnd2s1 _____9_502783(.DIN1 (____9____32426), .DIN2 (__9__9__30253),
       .Q (____0____32531));
  nnd2s1 _______502784(.DIN1 (____9_0__32411), .DIN2 (______9__32753),
       .Q (____0____32530));
  nor2s1 _______502785(.DIN1 (___00_9__30564), .DIN2 (____9____32412),
       .Q (____0____32529));
  nnd2s1 _____9_502786(.DIN1 (____9____32402), .DIN2 (____0____31550),
       .Q (____0____32528));
  nnd2s1 _____9_502787(.DIN1 (____9_9__32400), .DIN2 (____9___27564),
       .Q (____0_0__32527));
  nor2s1 _____0_502788(.DIN1 (___0__9__30890), .DIN2 (____9_0__32401),
       .Q (____0_9__32526));
  and2s1 _______502789(.DIN1 (____9____32395), .DIN2 (____0____32524),
       .Q (____0____32525));
  nor2s1 _______502790(.DIN1 (_________31762), .DIN2 (____9____32407),
       .Q (____0____32523));
  or2s1 _______502791(.DIN1 (____0____32521), .DIN2 (____9____32396),
       .Q (____0____32522));
  nor2s1 _______502792(.DIN1 (_____9__27986), .DIN2 (____9____32394),
       .Q (____0____32520));
  nor2s1 _______502793(.DIN1 (____0_0__32518), .DIN2 (____9____32392),
       .Q (____0____32519));
  nnd2s1 _______502794(.DIN1 (____9_0__32421), .DIN2 (___0_9), .Q
       (_____9___32670));
  dffacs1 _______________________502795(.CLRB (reset), .CLK (clk), .DIN
       (____9____32415), .QN (_____________________21679));
  and2s1 ______502796(.DIN1 (_____9___32373), .DIN2 (____0____32516),
       .Q (____0_9__32517));
  nor2s1 _______502797(.DIN1 (______0__32803), .DIN2 (____90___32389),
       .Q (____0____32515));
  and2s1 _______502798(.DIN1 (______9__32370), .DIN2 (_________32649),
       .Q (____0____32514));
  and2s1 _______502799(.DIN1 (____909__32390), .DIN2 (____0____32512),
       .Q (____0____32513));
  nor2s1 _______502800(.DIN1 (________25248), .DIN2 (____0____32510),
       .Q (____0____32511));
  nnd2s1 _______502801(.DIN1 (____90___32387), .DIN2 (___0____26129),
       .Q (____0____32509));
  and2s1 _______502802(.DIN1 (_________32951), .DIN2 (____0_9__32507),
       .Q (____0_0__32508));
  xor2s1 _______502803(.DIN1 (___0_____40512), .DIN2 (____0____32505),
       .Q (____0____32506));
  xor2s1 _______502804(.DIN1
       (____________________________________________21774), .DIN2
       (____0____32505), .Q (____0____32504));
  nor2s1 _______502805(.DIN1 (______9__35584), .DIN2 (____0____32501),
       .Q (____0____32503));
  nnd2s1 _______502806(.DIN1 (____0____32501), .DIN2 (______9__35584),
       .Q (____0____32502));
  nnd2s1 _______502807(.DIN1 (____90___32386), .DIN2 (____0____32499),
       .Q (____0____32500));
  nor2s1 _______502808(.DIN1 (________29057), .DIN2 (_____9___32374),
       .Q (____0_0__32498));
  nor2s1 _______502809(.DIN1 (________29052), .DIN2 (_____90__32371),
       .Q (____0_9__32497));
  nnd2s1 _______502810(.DIN1 (_____99__32380), .DIN2 (___0_____30915),
       .Q (____0____32496));
  nnd2s1 _______502811(.DIN1 (______9__32350), .DIN2 (______9__32615),
       .Q (____0____32495));
  nnd2s1 _______502812(.DIN1 (_________32338), .DIN2 (___0_____31180),
       .Q (____0____32494));
  nnd2s1 _______502813(.DIN1 (_________32367), .DIN2 (_________32298),
       .Q (____0____32493));
  nnd2s1 _______502814(.DIN1 (_________32345), .DIN2 (__90____29705),
       .Q (____0____32492));
  nor2s1 _______502815(.DIN1 (___0_9___31015), .DIN2 (_________32369),
       .Q (____0____32491));
  nor2s1 ______502816(.DIN1 (_________33897), .DIN2 (_________32362),
       .Q (____0____32490));
  nnd2s1 _______502817(.DIN1 (_____9___32372), .DIN2 (_____9___32379),
       .Q (_________32608));
  and2s1 ______502818(.DIN1 (____0____32510), .DIN2
       (____________________________________________21790), .Q
       (_________32617));
  nor2s1 _____502819(.DIN1
       (____________________________________________21790), .DIN2
       (____0____32510), .Q (____09___32570));
  xor2s1 _______502820(.DIN1 (____0___23792), .DIN2 (____9_9__32420),
       .Q (_________33201));
  dffacs1 _____________________9_502821(.CLRB (reset), .CLK (clk), .DIN
       (______0__32331), .QN (_________________9_));
  nor2s1 _____0_502822(.DIN1 (__9__9__30029), .DIN2 (_________32342),
       .Q (____0____32489));
  nnd2s1 ______502823(.DIN1 (_________32343), .DIN2 (________28537), .Q
       (____0_0__32488));
  nor2s1 _______502824(.DIN1 (________29402), .DIN2 (_________32353),
       .Q (____009__32487));
  nnd2s1 _______502825(.DIN1 (_________32346), .DIN2 (___9____26921),
       .Q (____00___32486));
  nor2s1 _______502826(.DIN1 (________27720), .DIN2 (______9__32340),
       .Q (____00___32485));
  nor2s1 _______502827(.DIN1 (___99___25116), .DIN2 (_________32352),
       .Q (____00___32484));
  nor2s1 _______502828(.DIN1 (________28950), .DIN2 (_________32363),
       .Q (____00___32483));
  nnd2s1 ______502829(.DIN1 (_________32332), .DIN2 (___009___30637),
       .Q (____00___32482));
  nnd2s1 _____9_502830(.DIN1 (_________32336), .DIN2 (__9_9___30175),
       .Q (____00___32481));
  nor2s1 _____9_502831(.DIN1 (_________32001), .DIN2 (_________32366),
       .Q (____00___32480));
  and2s1 _____502832(.DIN1 (_________32339), .DIN2 (____99___32478), .Q
       (____999__32479));
  nor2s1 _____0_502833(.DIN1 (___0_____30707), .DIN2 (_________32356),
       .Q (____99___32477));
  nnd2s1 _____0_502834(.DIN1 (_________32348), .DIN2 (__99____30491),
       .Q (____99___32476));
  nor2s1 _______502835(.DIN1 (___0_9___31111), .DIN2 (_________32355),
       .Q (____99___32475));
  nnd2s1 _____0_502836(.DIN1 (_________32337), .DIN2 (____9___29366),
       .Q (____99___32474));
  nor2s1 _______502837(.DIN1 (___099___31496), .DIN2 (_________32328),
       .Q (____99___32473));
  nor2s1 _______502838(.DIN1 (______0__32351), .DIN2 (_________32333),
       .Q (____99___32472));
  nor2s1 ______502839(.DIN1 (____9____32446), .DIN2 (_________32329),
       .Q (____99___32471));
  nnd2s1 _______502840(.DIN1 (_________32335), .DIN2 (____0____32516),
       .Q (____990__32470));
  nnd2s1 _______502841(.DIN1 (_________32327), .DIN2 (___9____27814),
       .Q (____9_9__32469));
  nor2s1 _______502842(.DIN1 (________29030), .DIN2 (_________32323),
       .Q (____9____32468));
  and2s1 ______502843(.DIN1 (_________32326), .DIN2 (____0____32534),
       .Q (____9____32467));
  nnd2s1 _______502844(.DIN1 (_________32324), .DIN2 (______9__32330),
       .Q (____9____32466));
  nor2s1 _______502845(.DIN1 (________28235), .DIN2 (_________32322),
       .Q (____9____32465));
  dffacs1 _______________________502846(.CLRB (reset), .CLK (clk), .DIN
       (_________32365), .QN (_____________________21669));
  dffacs1 _______________________502847(.CLRB (reset), .CLK (clk), .DIN
       (_________32368), .QN (_____________________21704));
  nnd2s1 _______502848(.DIN1 (____9____32444), .DIN2 (_________32611),
       .Q (____9____32464));
  nnd2s1 _______502849(.DIN1 (______0__32293), .DIN2 (______9__31688),
       .Q (____9____32463));
  or2s1 _______502850(.DIN1 (_________32956), .DIN2 (______9__32320),
       .Q (____9____32462));
  or2s1 _____9_502851(.DIN1 (____9_0__32460), .DIN2 (_________32319),
       .Q (____9____32461));
  nor2s1 _____0_502852(.DIN1 (___0_____40532), .DIN2 (_________32359),
       .Q (____9_9__32459));
  nnd2s1 _______502853(.DIN1 (____0____32505), .DIN2 (___0_____40503),
       .Q (____9____32458));
  nor2s1 _______502854(.DIN1 (___0_____40503), .DIN2 (____0____32505),
       .Q (____9____32457));
  nor2s1 ______502855(.DIN1 (____9____32454), .DIN2 (____0____32505),
       .Q (____9____32456));
  nnd2s1 ______502856(.DIN1 (____0____32505), .DIN2 (____9____32454),
       .Q (____9____32455));
  and2s1 _______502857(.DIN1 (____0____32505), .DIN2 (___0_____40512),
       .Q (____9____32453));
  nor2s1 _______502858(.DIN1 (___0_____40512), .DIN2 (____0____32505),
       .Q (____9____32452));
  nnd2s1 ______502859(.DIN1 (_________32271), .DIN2 (_________32238),
       .Q (____9_0__32451));
  nor2s1 _______502860(.DIN1 (____9____32449), .DIN2 (_________32294),
       .Q (____9_9__32450));
  nnd2s1 _______502861(.DIN1 (_____00__32283), .DIN2 (___0_____30665),
       .Q (____9____32448));
  nor2s1 _____9_502862(.DIN1 (____9____32446), .DIN2 (______9__32312),
       .Q (____9____32447));
  nnd2s1 _______502863(.DIN1 (____9____32444), .DIN2 (____9____32443),
       .Q (____9____32445));
  nnd2s1 ______502864(.DIN1 (_____0___32290), .DIN2 (____0____32543),
       .Q (____9____32442));
  and2s1 ______502865(.DIN1 (_________32310), .DIN2 (____00__27922), .Q
       (____9_0__32441));
  nor2s1 _______502866(.DIN1 (____9____32439), .DIN2 (______0__32321),
       .Q (____9_9__32440));
  nnd2s1 _______502867(.DIN1 (_________32306), .DIN2 (___00____30627),
       .Q (____9____32438));
  or2s1 _______502868(.DIN1 (____9____32436), .DIN2 (______0__32303),
       .Q (____9____32437));
  nor2s1 _______502869(.DIN1 (____9____32434), .DIN2 (_________32300),
       .Q (____9____32435));
  nnd2s1 ______502870(.DIN1 (_________32301), .DIN2 (________27309), .Q
       (____9____32433));
  nor2s1 _______502871(.DIN1 (________25840), .DIN2 (_____99__32282),
       .Q (____9____32432));
  nor2s1 _______502872(.DIN1 (___0_____31076), .DIN2 (_________32295),
       .Q (____9_0__32431));
  or2s1 ______502873(.DIN1
       (____________________________________________21762), .DIN2
       (____0____32505), .Q (____0____32564));
  nnd2s1 _______502874(.DIN1 (____0____32505), .DIN2
       (____________________________________________21762), .Q
       (____0____32565));
  dffacs1 _______________________502875(.CLRB (reset), .CLK (clk), .DIN
       (_____09__32292), .QN (_____________________21693));
  dffacs1 _______________________502876(.CLRB (reset), .CLK (clk), .DIN
       (_________32304), .QN (_____________________21707));
  dffacs1 _______________________502877(.CLRB (reset), .CLK (clk), .DIN
       (_________32317), .QN (_____________________21731));
  nor2s1 _______502878(.DIN1 (____0____31545), .DIN2 (______9__32262),
       .Q (____9_9__32430));
  nnd2s1 _______502879(.DIN1 (_____9___32277), .DIN2 (____9____32422),
       .Q (____9____32429));
  nor2s1 _____502880(.DIN1 (___00____30619), .DIN2 (_____0___32291), .Q
       (____9____32428));
  nnd2s1 _____9_502881(.DIN1 (______9__32302), .DIN2 (________28309),
       .Q (____9____32427));
  nor2s1 _____0_502882(.DIN1 (__9__9__30243), .DIN2 (______9__32242),
       .Q (____9____32426));
  nnd2s1 _____0_502883(.DIN1 (_________32297), .DIN2 (____9____32424),
       .Q (____9____32425));
  nnd2s1 _____502884(.DIN1 (_____0___32289), .DIN2 (____9____32422), .Q
       (____9____32423));
  nnd2s1 _______502885(.DIN1 (____9_9__32420), .DIN2 (___9___22270), .Q
       (____9_0__32421));
  nor2s1 _______502886(.DIN1 (_________32053), .DIN2 (_____9___32274),
       .Q (____9____32419));
  and2s1 ______502887(.DIN1 (_________32299), .DIN2 (____9____32417),
       .Q (____9____32418));
  nnd2s1 _______502888(.DIN1 (______9__32272), .DIN2 (____9_9__32410),
       .Q (____9____32416));
  nnd2s1 _______502889(.DIN1 (_________32249), .DIN2 (_________31620),
       .Q (____9____32415));
  and2s1 ______502890(.DIN1 (_________32269), .DIN2 (____9____32413),
       .Q (____9____32414));
  nnd2s1 _______502891(.DIN1 (_________32248), .DIN2 (___999__28735),
       .Q (____9____32412));
  nnd2s1 _______502892(.DIN1 (_________32264), .DIN2 (____9_9__32410),
       .Q (____9_0__32411));
  nor2s1 _______502893(.DIN1 (___0_____30856), .DIN2 (_________32256),
       .Q (____9____32409));
  nor2s1 _______502894(.DIN1 (__9_____30288), .DIN2 (______0__32313),
       .Q (____9____32408));
  nnd2s1 _______502895(.DIN1 (_________32261), .DIN2 (____0____31517),
       .Q (____9____32407));
  and2s1 _______502896(.DIN1 (_________32257), .DIN2 (_________31937),
       .Q (____9____32406));
  nor2s1 _______502897(.DIN1 (___000___30553), .DIN2 (_________32244),
       .Q (____9____32405));
  nor2s1 _____502898(.DIN1 (___0__9__30890), .DIN2 (______0__32263), .Q
       (____9____32404));
  nor2s1 _____0_502899(.DIN1 (_____0___31803), .DIN2 (_________32259),
       .Q (____9____32403));
  nnd2s1 _____0_502900(.DIN1 (_________32258), .DIN2 (______9__32753),
       .Q (____9____32402));
  nor2s1 ______502901(.DIN1 (___0_9___31405), .DIN2 (_________32255),
       .Q (____9_0__32401));
  nor2s1 _______502902(.DIN1 (________27320), .DIN2 (_________32265),
       .Q (____9_9__32400));
  nor2s1 _______502903(.DIN1 (______0__32253), .DIN2 (____9____32398),
       .Q (____9____32399));
  nor2s1 ______502904(.DIN1 (____00__25768), .DIN2 (_________32270), .Q
       (____9____32397));
  nnd2s1 ______502905(.DIN1 (_________32250), .DIN2 (________27446), .Q
       (____9____32396));
  nor2s1 _______502906(.DIN1 (___9____27790), .DIN2 (_________32247),
       .Q (____9____32395));
  nnd2s1 ______502907(.DIN1 (_________32251), .DIN2 (____0____31556),
       .Q (____9____32394));
  nor2s1 _______502908(.DIN1 (_________31817), .DIN2 (______0__32243),
       .Q (____9____32393));
  nnd2s1 _______502909(.DIN1 (_________32245), .DIN2 (____9_0__32391),
       .Q (____9____32392));
  and2s1 _______502910(.DIN1 (_________32229), .DIN2 (____0___28378),
       .Q (____909__32390));
  xor2s1 _______502911(.DIN1 (_____9___32182), .DIN2 (_____9___36360),
       .Q (____90___32389));
  xor2s1 _______502912(.DIN1 (_____9___32177), .DIN2 (_________38214),
       .Q (____90___32388));
  nnd2s1 ______502913(.DIN1 (_________32237), .DIN2 (inData[30]), .Q
       (____90___32387));
  nor2s1 _______502914(.DIN1 (_________32598), .DIN2 (_________32219),
       .Q (____90___32386));
  nnd2s1 _______502915(.DIN1 (______9__32213), .DIN2 (____90___32384),
       .Q (____90___32385));
  nnd2s1 _______502916(.DIN1 (_________32358), .DIN2 (____90___32382),
       .Q (____90___32383));
  xor2s1 ______502917(.DIN1 (____90___32382), .DIN2 (____9____38944),
       .Q (____900__32381));
  nor2s1 _______502918(.DIN1 (___0_____31011), .DIN2 (_________32221),
       .Q (_____99__32380));
  nnd2s1 _______502919(.DIN1 (_________32236), .DIN2 (_________33321),
       .Q (_____9___32379));
  nnd2s1 _______502920(.DIN1 (_________33080), .DIN2 (______9__32360),
       .Q (_____9___32378));
  or2s1 _____9_502921(.DIN1 (_____9___32376), .DIN2 (_____9___32375),
       .Q (_____9___32377));
  nnd2s1 _____9_502922(.DIN1 (_________32231), .DIN2 (__9___), .Q
       (_____9___32374));
  nor2s1 _____502923(.DIN1 (___9____26890), .DIN2 (______0__32234), .Q
       (_____9___32373));
  nnd2s1 ______502924(.DIN1 (_________32232), .DIN2
       (_______________22069), .Q (_____9___32372));
  nor2s1 _______502925(.DIN1 (___0900), .DIN2 (_________32217), .Q
       (_____90__32371));
  and2s1 _______502926(.DIN1 (_________32203), .DIN2 (________28349),
       .Q (______9__32370));
  or2s1 _______502927(.DIN1 (________27665), .DIN2 (_________32228), .Q
       (_________32369));
  or2s1 ______502928(.DIN1 (_________32344), .DIN2 (_________32227), .Q
       (_________32368));
  and2s1 _______502929(.DIN1 (______9__32223), .DIN2 (__9__9__29779),
       .Q (_________32367));
  nor2s1 _______502930(.DIN1 (____9____32446), .DIN2 (_________32240),
       .Q (_________32366));
  or2s1 _______502931(.DIN1 (_________32364), .DIN2 (_________32226),
       .Q (_________32365));
  nnd2s1 ______502932(.DIN1 (_________32200), .DIN2 (___09____31472),
       .Q (_________32363));
  nor2s1 ______502933(.DIN1 (___0_____31324), .DIN2 (_________32222),
       .Q (_________32362));
  hi1s1 _______502934(.DIN (______0__32361), .Q (_________32800));
  nor2s1 _______502935(.DIN1 (______9__32360), .DIN2 (_________33080),
       .Q (____0____32501));
  hi1s1 _______502936(.DIN (_________32359), .Q (____0____32510));
  nor2s1 _______502937(.DIN1 (_____9___32179), .DIN2 (_________32358),
       .Q (_________32951));
  nor2s1 _______502938(.DIN1 (_________41262), .DIN2 (_________32215),
       .Q (_________32357));
  nor2s1 _______502939(.DIN1 (_____90__32273), .DIN2 (_________32212),
       .Q (_________32356));
  or2s1 ______502940(.DIN1 (_________31783), .DIN2 (______9__32233), .Q
       (_________32355));
  nnd2s1 _______502941(.DIN1 (_________32334), .DIN2 (inData[31]), .Q
       (_________32354));
  nnd2s1 _______502942(.DIN1 (_________32211), .DIN2 (__9_0___29812),
       .Q (_________32353));
  nor2s1 _______502943(.DIN1 (______0__32351), .DIN2 (_________32202),
       .Q (_________32352));
  and2s1 _______502944(.DIN1 (_____0___32194), .DIN2 (_________32349),
       .Q (______9__32350));
  and2s1 ______502945(.DIN1 (_________32210), .DIN2 (_________32347),
       .Q (_________32348));
  nor2s1 ______502946(.DIN1 (_____0___31991), .DIN2 (_________32209),
       .Q (_________32346));
  nor2s1 _______502947(.DIN1 (_________32344), .DIN2 (_________32220),
       .Q (_________32345));
  nor2s1 _____0_502948(.DIN1 (_____9___31886), .DIN2 (_________32207),
       .Q (_________32343));
  nnd2s1 _____0_502949(.DIN1 (_________32216), .DIN2 (________29048),
       .Q (_________32342));
  nor2s1 _______502950(.DIN1 (____9____33386), .DIN2 (_________32197),
       .Q (______0__32341));
  nnd2s1 _______502951(.DIN1 (_____0___32191), .DIN2 (_________31953),
       .Q (______9__32340));
  nor2s1 _______502952(.DIN1 (__9_____30030), .DIN2 (_________32230),
       .Q (_________32339));
  nnd2s1 _______502953(.DIN1 (_________32206), .DIN2 (____9_9__32410),
       .Q (_________32338));
  nor2s1 ______502954(.DIN1 (_____0__28238), .DIN2 (_________32199), .Q
       (_________32337));
  nnd2s1 _______502955(.DIN1 (_________32201), .DIN2 (____9____32424),
       .Q (_________32336));
  nor2s1 _______502956(.DIN1 (______0__41150), .DIN2 (_________32334),
       .Q (_________32335));
  or2s1 _______502957(.DIN1 (_____0___32288), .DIN2 (_____0___32189),
       .Q (_________32333));
  nor2s1 _______502958(.DIN1 (___0_____30757), .DIN2 (_________32198),
       .Q (_________32332));
  nnd2s1 _______502959(.DIN1 (_____09__32195), .DIN2 (______9__32330),
       .Q (______0__32331));
  nnd2s1 _______502960(.DIN1 (_____0___32192), .DIN2 (_____0__27167),
       .Q (_________32329));
  nnd2s1 _______502961(.DIN1 (_____0___32193), .DIN2 (_____9__27551),
       .Q (_________32328));
  nor2s1 _______502962(.DIN1 (________27512), .DIN2 (_____0___32187),
       .Q (_________32327));
  and2s1 _______502963(.DIN1 (_____0___32188), .DIN2 (_________32325),
       .Q (_________32326));
  nor2s1 _______502964(.DIN1 (_________31881), .DIN2 (_____00__32186),
       .Q (_________32324));
  nor2s1 ______502965(.DIN1 (___0900), .DIN2 (_____99__32185), .Q
       (_________32323));
  nnd2s1 _______502966(.DIN1 (_________32208), .DIN2 (________28401),
       .Q (_________32322));
  nnd2s1 _____502967(.DIN1 (______0__32147), .DIN2 (____0___28477), .Q
       (______0__32321));
  nnd2s1 _______502968(.DIN1 (_____9___32183), .DIN2 (____9___24832),
       .Q (______9__32320));
  xor2s1 _____0_502969(.DIN1 (_________32318), .DIN2 (_________34647),
       .Q (_________32319));
  nnd2s1 _____0_502970(.DIN1 (_________32174), .DIN2 (___0_____31253),
       .Q (_________32317));
  nor2s1 ______502971(.DIN1 (_________32315), .DIN2 (______0__32224),
       .Q (_________32316));
  nor2s1 _____0_502972(.DIN1 (____0____32541), .DIN2 (_________32148),
       .Q (______0__32313));
  or2s1 _______502973(.DIN1 (_________32311), .DIN2 (_________32172),
       .Q (______9__32312));
  nor2s1 _____0_502974(.DIN1 (_________32042), .DIN2 (_________32170),
       .Q (_________32310));
  nnd2s1 _______502975(.DIN1 (_________32171), .DIN2 (_________31823),
       .Q (_________32309));
  nor2s1 _____502976(.DIN1 (____0____32539), .DIN2 (_________32150), .Q
       (_________32308));
  or2s1 _____502977(.DIN1 (___0_____31335), .DIN2 (_____9___36007), .Q
       (_________32307));
  nor2s1 ______502978(.DIN1 (_________32305), .DIN2 (_________32167),
       .Q (_________32306));
  nnd2s1 _______502979(.DIN1 (______0__32166), .DIN2 (_____0___31705),
       .Q (_________32304));
  or2s1 _______502980(.DIN1 (________26666), .DIN2 (______9__32165), .Q
       (______0__32303));
  nor2s1 _______502981(.DIN1 (________28572), .DIN2 (_________32164),
       .Q (______9__32302));
  nor2s1 _______502982(.DIN1 (________28525), .DIN2 (_____9___32281),
       .Q (_________32301));
  or2s1 _______502983(.DIN1 (__9_____29860), .DIN2 (_________32163), .Q
       (_________32300));
  and2s1 ______502984(.DIN1 (_________32157), .DIN2 (_________32298),
       .Q (_________32299));
  nnd2s1 _______502985(.DIN1 (______0__32156), .DIN2 (_________32296),
       .Q (_________32297));
  nnd2s1 _______502986(.DIN1 (______9__32155), .DIN2 (__9__9__30356),
       .Q (_________32295));
  or2s1 _______502987(.DIN1 (___0____27863), .DIN2 (_________32154), .Q
       (_________32294));
  nor2s1 _______502988(.DIN1 (_________32056), .DIN2 (_________32153),
       .Q (______0__32293));
  nnd2s1 _______502989(.DIN1 (_________32173), .DIN2 (__9_____30259),
       .Q (_____09__32292));
  and2s1 _______502990(.DIN1 (_________32152), .DIN2 (____0____32543),
       .Q (_____0___32291));
  nnd2s1 _______502991(.DIN1 (_________32151), .DIN2 (______0__32205),
       .Q (_____0___32290));
  nor2s1 _____9_502992(.DIN1 (_____0___32288), .DIN2 (_________32149),
       .Q (_____0___32289));
  xor2s1 _______502993(.DIN1 (_________32101), .DIN2 (_____0___32287),
       .Q (_________32359));
  nnd2s1 _____9_502994(.DIN1 (_________32162), .DIN2 (________28891),
       .Q (____9_9__32420));
  or2s1 ______502995(.DIN1 (_____0___32286), .DIN2 (_____0___32285), .Q
       (____9____32444));
  nnd2s1 _______502996(.DIN1 (_____0___32285), .DIN2 (_____0___32286),
       .Q (____9____32443));
  nor2s1 _______502997(.DIN1 (______9__32175), .DIN2 (_____9___32178),
       .Q (______0__32361));
  dffacs1 _______________________502998(.CLRB (reset), .CLK (clk), .DIN
       (_________32168), .QN (_____________________21706));
  xnr2s1 _______502999(.DIN1 (_________32235), .DIN2 (___00_9__30592),
       .Q (____0____32505));
  nnd2s1 ____9__503000(.DIN1 (_________32134), .DIN2 (________26299),
       .Q (_____0___32284));
  nnd2s1 _______503001(.DIN1 (_____9___32181), .DIN2 (______9__32753),
       .Q (_____00__32283));
  and2s1 _______503002(.DIN1 (_____9___32281), .DIN2 (_________32159),
       .Q (_____99__32282));
  nnd2s1 ______503003(.DIN1 (_________32139), .DIN2 (____0____32524),
       .Q (_____9___32280));
  nnd2s1 _______503004(.DIN1 (_____0___32286), .DIN2
       (_______________22070), .Q (_____9___32279));
  or2s1 _______503005(.DIN1 (_______________22070), .DIN2
       (_____0___32286), .Q (_____9___32278));
  nor2s1 _______503006(.DIN1 (_____0___32288), .DIN2 (_________32144),
       .Q (_____9___32277));
  nnd2s1 _______503007(.DIN1 (_____9___32275), .DIN2 (______9__32753),
       .Q (_____9___32276));
  nor2s1 _______503008(.DIN1 (_____90__32273), .DIN2 (_________32143),
       .Q (_____9___32274));
  nnd2s1 _______503009(.DIN1 (______9__32136), .DIN2 (___0_____31394),
       .Q (______9__32272));
  nnd2s1 _______503010(.DIN1 (_________32141), .DIN2 (_________32266),
       .Q (_________32271));
  or2s1 ______503011(.DIN1 (_________33580), .DIN2 (_________32129), .Q
       (_________32270));
  nor2s1 _____503012(.DIN1 (___0__0__30778), .DIN2 (_________32124), .Q
       (_________32269));
  and2s1 _____503013(.DIN1 (_________32267), .DIN2 (_________32266), .Q
       (_________32268));
  nnd2s1 _____0_503014(.DIN1 (______9__32252), .DIN2 (__9_____30096),
       .Q (_________32265));
  nor2s1 _____0_503015(.DIN1 (_________32241), .DIN2 (_________32113),
       .Q (_________32264));
  nor2s1 _____0_503016(.DIN1 (__909___29721), .DIN2 (______9__32126),
       .Q (______0__32263));
  nnd2s1 _____503017(.DIN1 (_________32121), .DIN2 (______0__31825), .Q
       (______9__32262));
  and2s1 ______503018(.DIN1 (______0__32127), .DIN2 (_________32260),
       .Q (_________32261));
  nnd2s1 _______503019(.DIN1 (_________32119), .DIN2 (____0____31581),
       .Q (_________32259));
  nnd2s1 _______503020(.DIN1 (_________32131), .DIN2 (__9_____29818),
       .Q (_________32258));
  nor2s1 _______503021(.DIN1 (_________31878), .DIN2 (_________32110),
       .Q (_________32257));
  nnd2s1 ______503022(.DIN1 (_________32123), .DIN2 (_________32135),
       .Q (_________32256));
  nnd2s1 _______503023(.DIN1 (______9__32107), .DIN2 (____09__28480),
       .Q (_________32255));
  nor2s1 ______503024(.DIN1 (______0__32253), .DIN2 (______9__32252),
       .Q (_________32254));
  nor2s1 _______503025(.DIN1 (________29519), .DIN2 (_________32111),
       .Q (_________32251));
  nor2s1 _______503026(.DIN1 (________29531), .DIN2 (______0__32118),
       .Q (_________32250));
  nor2s1 ______503027(.DIN1 (__99____30531), .DIN2 (_________32132), .Q
       (_________32249));
  nor2s1 _______503028(.DIN1 (___0_____30962), .DIN2 (_________32106),
       .Q (_________32248));
  or2s1 _______503029(.DIN1 (_________32246), .DIN2 (_________32125),
       .Q (_________32247));
  nor2s1 _______503030(.DIN1 (_____0___34102), .DIN2 (_________32115),
       .Q (_________32245));
  nnd2s1 _______503031(.DIN1 (_________32120), .DIN2 (______9__32330),
       .Q (_________32244));
  nnd2s1 ______503032(.DIN1 (_________32109), .DIN2 (__9_____30332), .Q
       (______0__32243));
  nor2s1 _______503033(.DIN1 (___0____25136), .DIN2 (_____9___32180),
       .Q (______9__32242));
  nor2s1 _______503034(.DIN1 (_________32241), .DIN2 (_________32133),
       .Q (____9____32398));
  nnd2s1 _______503035(.DIN1 (_________32066), .DIN2 (_________32239),
       .Q (_________32240));
  nnd2s1 _____9_503036(.DIN1 (_____9___32081), .DIN2 (______9__32753),
       .Q (_________32238));
  nor2s1 _____9_503037(.DIN1 (_________32100), .DIN2 (___0_00__31023),
       .Q (_________32237));
  nnd2s1 _______503038(.DIN1 (_________32235), .DIN2 (________27457),
       .Q (_________32236));
  nnd2s1 _______503039(.DIN1 (_____0___32095), .DIN2 (___0_____31049),
       .Q (______0__32234));
  nnd2s1 _____9_503040(.DIN1 (_________32048), .DIN2 (________29029),
       .Q (______9__32233));
  nnd2s1 ______503041(.DIN1 (_________32235), .DIN2 (_____9__28940), .Q
       (_________32232));
  nnd2s1 _______503042(.DIN1 (_____0___32092), .DIN2 (____9____32424),
       .Q (_________32231));
  or2s1 _____9_503043(.DIN1 (________28986), .DIN2 (______0__32060), .Q
       (_________32230));
  nor2s1 _______503044(.DIN1 (___0_____31190), .DIN2 (_____9___32083),
       .Q (_________32229));
  nnd2s1 ______503045(.DIN1 (_________40942), .DIN2 (________29079), .Q
       (_________32228));
  nnd2s1 _______503046(.DIN1 (_____0___32090), .DIN2 (___9____29566),
       .Q (_________32227));
  nnd2s1 _______503047(.DIN1 (_____9___32087), .DIN2 (_____0__29204),
       .Q (_________32226));
  hi1s1 _______503048(.DIN (______0__32224), .Q (_________32225));
  nor2s1 _______503049(.DIN1 (______0__31970), .DIN2 (______0__40944),
       .Q (______9__32223));
  nnd2s1 _______503050(.DIN1 (_____9___32088), .DIN2 (__9_____29976),
       .Q (_________32222));
  nnd2s1 _______503051(.DIN1 (_________32064), .DIN2 (__9__9__30215),
       .Q (_________32221));
  nnd2s1 _______503052(.DIN1 (______9__32069), .DIN2 (_________32004),
       .Q (_________32220));
  or2s1 ______503053(.DIN1 (_________32218), .DIN2 (_____9___32085), .Q
       (_________32219));
  nor2s1 _______503054(.DIN1 (___0_0___30746), .DIN2 (_____9___32086),
       .Q (_________32217));
  nor2s1 _______503055(.DIN1 (__990___30459), .DIN2 (_________32063),
       .Q (_________32216));
  or2s1 _______503056(.DIN1 (______0__32214), .DIN2 (_____9___32084),
       .Q (_________32215));
  hi1s1 _____9_503057(.DIN (____90___32382), .Q (____90___32384));
  nor2s1 _______503058(.DIN1 (____0____32541), .DIN2 (_____0___32093),
       .Q (_____9___32375));
  hi1s1 _______503059(.DIN (______9__32213), .Q (_________32358));
  xor2s1 _______503060(.DIN1 (________28893), .DIN2 (_________32161),
       .Q (_________33080));
  nor2s1 _____9_503061(.DIN1 (_________32142), .DIN2 (______9__32079),
       .Q (_________32212));
  nor2s1 _____0_503062(.DIN1 (____0___29017), .DIN2 (_________32103),
       .Q (_________32211));
  and2s1 _____0_503063(.DIN1 (_________32051), .DIN2 (__9_____30305),
       .Q (_________32210));
  nnd2s1 _____0_503064(.DIN1 (_____0___32091), .DIN2 (____0____31577),
       .Q (_________32209));
  nnd2s1 ____0__503065(.DIN1 (_________32037), .DIN2 (________25544),
       .Q (_________32208));
  nnd2s1 _______503066(.DIN1 (______0__32070), .DIN2 (__9__0__30130),
       .Q (_________32207));
  nnd2s1 _______503067(.DIN1 (_________32072), .DIN2 (______0__32205),
       .Q (_________32206));
  nor2s1 _______503068(.DIN1 (_____9__28368), .DIN2 (_________32052),
       .Q (______9__32204));
  nor2s1 _______503069(.DIN1 (___0_____31086), .DIN2 (_________32047),
       .Q (_________32203));
  nnd2s1 _______503070(.DIN1 (_____99__32089), .DIN2 (__9_____30241),
       .Q (_________32202));
  nnd2s1 ______503071(.DIN1 (______9__32059), .DIN2 (___9____26906), .Q
       (_________32201));
  nor2s1 _______503072(.DIN1 (___00____30610), .DIN2 (_________32045),
       .Q (_________32200));
  nor2s1 _______503073(.DIN1 (____0____32541), .DIN2 (_________32068),
       .Q (_________32199));
  nor2s1 _______503074(.DIN1 (____9____33386), .DIN2 (_________32054),
       .Q (_________32198));
  and2s1 _______503075(.DIN1 (_________32057), .DIN2 (______0__32196),
       .Q (_________32197));
  nor2s1 _______503076(.DIN1 (__9_0___29728), .DIN2 (_________32044),
       .Q (_____09__32195));
  nor2s1 _______503077(.DIN1 (__99_9__30527), .DIN2 (______9__32049),
       .Q (_____0___32194));
  nor2s1 ______503078(.DIN1 (________28909), .DIN2 (_________32061), .Q
       (_____0___32193));
  nor2s1 _______503079(.DIN1 (____0____31547), .DIN2 (_________32046),
       .Q (_____0___32192));
  nor2s1 _______503080(.DIN1 (_________31843), .DIN2 (_____9___32082),
       .Q (_____0___32191));
  nor2s1 ______503081(.DIN1 (____0____32539), .DIN2 (______0__32050),
       .Q (_____0___32190));
  nnd2s1 _______503082(.DIN1 (_________32043), .DIN2 (______9__31765),
       .Q (_____0___32189));
  and2s1 _______503083(.DIN1 (_________32041), .DIN2 (__90____29647),
       .Q (_____0___32188));
  nnd2s1 _____9_503084(.DIN1 (______9__32039), .DIN2 (________28338),
       .Q (_____0___32187));
  or2s1 ____9__503085(.DIN1 (________29291), .DIN2 (______0__32040), .Q
       (_____00__32186));
  nor2s1 ____9__503086(.DIN1 (_________31667), .DIN2 (_________32038),
       .Q (_____99__32185));
  or2s1 ______503087(.DIN1 (_____9___32184), .DIN2 (_________32077), .Q
       (_________32334));
  nnd2s1 _______503088(.DIN1 (_________32034), .DIN2 (___99____39861),
       .Q (_____9___32183));
  xor2s1 ______503089(.DIN1 (______9__31930), .DIN2 (______0__35853),
       .Q (_____9___32182));
  or2s1 _______503090(.DIN1 (_________32241), .DIN2 (_____90__31980),
       .Q (_____9___32181));
  nor2s1 _______503091(.DIN1 (_________31870), .DIN2 (_____9___31981),
       .Q (_____9___32180));
  xor2s1 _______503092(.DIN1 (_________31927), .DIN2 (___9_____39301),
       .Q (_____9___32179));
  nor2s1 _______503093(.DIN1 (_________32613), .DIN2 (_____90__32176),
       .Q (_____9___32178));
  nor2s1 ______503094(.DIN1 (_____90__32176), .DIN2 (______9__32175),
       .Q (_____9___32177));
  nor2s1 _______503095(.DIN1 (___0_____31227), .DIN2 (_________31975),
       .Q (_________32174));
  nor2s1 _______503096(.DIN1 (__9_____30128), .DIN2 (_____0___31993),
       .Q (_________32173));
  or2s1 _______503097(.DIN1 (_________33580), .DIN2 (______0__32020),
       .Q (_________32172));
  xor2s1 _____0_503098(.DIN1 (_________31914), .DIN2 (___009___39979),
       .Q (_________32171));
  nnd2s1 ______503099(.DIN1 (_________32035), .DIN2 (____00___31507),
       .Q (_________32170));
  xor2s1 _______503100(.DIN1
       (____________________________________________21834), .DIN2
       (_____9___34281), .Q (_________32169));
  nnd2s1 ______503101(.DIN1 (_________32006), .DIN2 (______9__31660),
       .Q (_________32168));
  nnd2s1 ______503102(.DIN1 (_________32007), .DIN2 (___90___28649), .Q
       (_________32167));
  nor2s1 _______503103(.DIN1 (___00____30615), .DIN2 (_________32005),
       .Q (______0__32166));
  nnd2s1 _______503104(.DIN1 (______0__32137), .DIN2 (____0___27393),
       .Q (______9__32165));
  nnd2s1 ______503105(.DIN1 (_________32003), .DIN2 (________28402), .Q
       (_________32164));
  nnd2s1 _______503106(.DIN1 (_________32158), .DIN2 (_________31648),
       .Q (_________32163));
  nnd2s1 _______503107(.DIN1 (_________32161), .DIN2 (________28892),
       .Q (_________32162));
  or2s1 ______503108(.DIN1 (_________32159), .DIN2 (_________32158), .Q
       (_________32160));
  and2s1 ______503109(.DIN1 (______0__32000), .DIN2 (__9_90__30169), .Q
       (_________32157));
  nor2s1 _____9_503110(.DIN1 (___0_____31262), .DIN2 (_________32008),
       .Q (______0__32156));
  nnd2s1 _____9_503111(.DIN1 (_____0___31997), .DIN2 (________25544),
       .Q (______9__32155));
  nnd2s1 _____9_503112(.DIN1 (_____0___31996), .DIN2 (________26422),
       .Q (_________32154));
  nnd2s1 _____0_503113(.DIN1 (_____0___31995), .DIN2 (____0____31566),
       .Q (_________32153));
  nnd2s1 _____0_503114(.DIN1 (_____0___31992), .DIN2 (_________31973),
       .Q (_________32152));
  nor2s1 _______503115(.DIN1 (___09____31480), .DIN2 (_____00__31990),
       .Q (_________32151));
  nor2s1 _______503116(.DIN1 (______0__41140), .DIN2 (_________32023),
       .Q (_________32150));
  nnd2s1 _______503117(.DIN1 (_________32028), .DIN2 (_________32022),
       .Q (_________32149));
  nor2s1 _______503118(.DIN1 (_________31809), .DIN2 (______9__32029),
       .Q (_________32148));
  nor2s1 _______503119(.DIN1 (__9_____30106), .DIN2 (_____0___31998),
       .Q (______0__32147));
  nnd2s1 _______503120(.DIN1 (_________32027), .DIN2 (_____0___32287),
       .Q (_________32314));
  xor2s1 _______503121(.DIN1 (_________31926), .DIN2 (____0_0__38064),
       .Q (______9__32213));
  nnd2s1 _______503122(.DIN1 (_________32017), .DIN2 (_________31642),
       .Q (_____0___32285));
  and2s1 _______503123(.DIN1 (______9__32146), .DIN2
       (____________________________________________21789), .Q
       (_________32315));
  nor2s1 _______503124(.DIN1
       (____________________________________________21789), .DIN2
       (______9__32146), .Q (______0__32224));
  xor2s1 _______503125(.DIN1 (_________31915), .DIN2 (_________32145),
       .Q (____90___32382));
  nnd2s1 _______503126(.DIN1 (_________31978), .DIN2 (_____9___31694),
       .Q (_________32144));
  nor2s1 _______503127(.DIN1 (_________32142), .DIN2 (_________31976),
       .Q (_________32143));
  nnd2s1 _______503128(.DIN1 (______9__31979), .DIN2 (_________32140),
       .Q (_________32141));
  nor2s1 _______503129(.DIN1 (________28500), .DIN2 (_____9___31982),
       .Q (_________32139));
  nor2s1 _______503130(.DIN1 (_____9___32376), .DIN2 (______0__32137),
       .Q (_________32138));
  nor2s1 _______503131(.DIN1 (___09____31467), .DIN2 (_________32021),
       .Q (______9__32136));
  nnd2s1 ______503132(.DIN1 (_________32036), .DIN2 (____9_9__32410),
       .Q (_________32135));
  nnd2s1 ____0__503133(.DIN1 (______0__31940), .DIN2 (___0_____31297),
       .Q (_________32134));
  or2s1 ____00_503134(.DIN1 (_________32142), .DIN2 (_________31943),
       .Q (_________32133));
  nor2s1 ____00_503135(.DIN1 (_________33897), .DIN2 (_________31948),
       .Q (_________32132));
  nor2s1 _____9_503136(.DIN1 (_________32130), .DIN2 (______9__31949),
       .Q (_________32131));
  or2s1 _____503137(.DIN1 (___09____31451), .DIN2 (_________31951), .Q
       (_________32129));
  nor2s1 ____90_503138(.DIN1 (_____9___32376), .DIN2 (______0__31960),
       .Q (_________32128));
  nor2s1 ____90_503139(.DIN1 (__9__9__30419), .DIN2 (______9__31969),
       .Q (______0__32127));
  nnd2s1 ____90_503140(.DIN1 (_________31974), .DIN2 (_____9___31891),
       .Q (______9__32126));
  nnd2s1 ____9__503141(.DIN1 (_________31971), .DIN2 (_________41238),
       .Q (_________32125));
  or2s1 ____9__503142(.DIN1 (__9_____29790), .DIN2 (_________31946), .Q
       (_________32124));
  nnd2s1 ____9__503143(.DIN1 (_________31963), .DIN2 (____0____32543),
       .Q (_________32123));
  nor2s1 ____9__503144(.DIN1 (_________41168), .DIN2 (_________31965),
       .Q (_________32122));
  nor2s1 ____9_503145(.DIN1 (___0_____31132), .DIN2 (_________31968),
       .Q (_________32121));
  nor2s1 ____9__503146(.DIN1 (____0____31584), .DIN2 (_________31972),
       .Q (_________32120));
  and2s1 ____9__503147(.DIN1 (_________31962), .DIN2 (____0____31579),
       .Q (_________32119));
  or2s1 ____9__503148(.DIN1 (______9__32117), .DIN2 (_________31967),
       .Q (______0__32118));
  nnd2s1 ____00_503149(.DIN1 (_________31941), .DIN2 (_________32266),
       .Q (_________32116));
  nnd2s1 ____9_503150(.DIN1 (______9__31959), .DIN2 (_________32114),
       .Q (_________32115));
  nnd2s1 ____9_503151(.DIN1 (_________31961), .DIN2 (_________32140),
       .Q (_________32113));
  nor2s1 ____9_503152(.DIN1 (____9____33386), .DIN2 (_________31956),
       .Q (_________32112));
  nnd2s1 ____9__503153(.DIN1 (_________31954), .DIN2 (___9____29592),
       .Q (_________32111));
  nor2s1 ____9__503154(.DIN1 (___99___25116), .DIN2 (_________31957),
       .Q (_________32110));
  and2s1 ____9__503155(.DIN1 (_________31952), .DIN2 (______0__32108),
       .Q (_________32109));
  nor2s1 ____9__503156(.DIN1 (__9__9__30262), .DIN2 (_________31964),
       .Q (______9__32107));
  or2s1 ____503157(.DIN1 (_________32105), .DIN2 (_________31945), .Q
       (_________32106));
  or2s1 ____9__503158(.DIN1 (_________32142), .DIN2 (_________31966),
       .Q (_________32267));
  nnd2s1 _______503159(.DIN1 (_____9___31988), .DIN2 (_________32104),
       .Q (_____9___32281));
  nor2s1 ____0__503160(.DIN1 (_________32142), .DIN2 (_________31947),
       .Q (______9__32252));
  nnd2s1 _______503161(.DIN1 (_____9___31987), .DIN2 (____9_9__32410),
       .Q (_____9___32275));
  nor2s1 _______503162(.DIN1 (____0_9__31532), .DIN2 (_____9___31984),
       .Q (_____9___36007));
  xor2s1 _______503163(.DIN1 (_________31883), .DIN2
       (______________22067), .Q (_____0___32286));
  nnd2s1 ____9__503164(.DIN1 (______0__31875), .DIN2 (___009___30639),
       .Q (_________32103));
  xor2s1 _______503165(.DIN1 (___0_____40548), .DIN2 (_________32031),
       .Q (_________32102));
  xor2s1 _______503166(.DIN1 (___0009__30554), .DIN2 (_________32026),
       .Q (_________32101));
  xor2s1 _______503167(.DIN1 (_________31819), .DIN2 (___0_0___30647),
       .Q (_________32100));
  xor2s1 _______503168(.DIN1 (_________32016), .DIN2 (_____9___35917),
       .Q (_________32099));
  nor2s1 _______503169(.DIN1
       (____________________________________________21761), .DIN2
       (_____9___34281), .Q (______0__32098));
  nnd2s1 _______503170(.DIN1 (_____9___34281), .DIN2
       (____________________________________________21761), .Q
       (_____09__32097));
  nor2s1 _______503171(.DIN1
       (____________________________________________21834), .DIN2
       (_____9___34281), .Q (_____0___32096));
  nnd2s1 _____9_503172(.DIN1 (_________31923), .DIN2 (_________32159),
       .Q (_____0___32095));
  and2s1 _______503173(.DIN1 (_____9___34281), .DIN2
       (____________________________________________21834), .Q
       (_____0___32094));
  nnd2s1 _______503174(.DIN1 (_________31922), .DIN2 (_________33000),
       .Q (_____0___32093));
  nnd2s1 ______503175(.DIN1 (_________31918), .DIN2 (_________32296),
       .Q (_____0___32092));
  nor2s1 ____9__503176(.DIN1 (___0_0___30649), .DIN2 (_________31872),
       .Q (_____0___32091));
  nor2s1 ______503177(.DIN1 (________28087), .DIN2 (______0__31865), .Q
       (_____0___32090));
  nor2s1 _____9_503178(.DIN1 (_________32071), .DIN2 (_________31908),
       .Q (_____99__32089));
  nor2s1 ____503179(.DIN1 (_________33742), .DIN2 (_________31907), .Q
       (_____9___32088));
  nor2s1 ____90_503180(.DIN1 (___090___31408), .DIN2 (______9__31874),
       .Q (_____9___32087));
  nnd2s1 ____90_503181(.DIN1 (_________31904), .DIN2 (___0_____31151),
       .Q (_____9___32086));
  or2s1 ____90_503182(.DIN1 (___0____28762), .DIN2 (_________31905), .Q
       (_____9___32085));
  or2s1 ____503183(.DIN1 (___9____27793), .DIN2 (_____0___31901), .Q
       (_____9___32084));
  nnd2s1 ____9_503184(.DIN1 (_________31863), .DIN2 (____9___28195), .Q
       (_____9___32083));
  nnd2s1 ____9_503185(.DIN1 (_____0___31897), .DIN2 (____0___28020), .Q
       (_____9___32082));
  nnd2s1 ____9_503186(.DIN1 (_____90__31885), .DIN2 (_____90__32080),
       .Q (_____9___32081));
  nnd2s1 ____9__503187(.DIN1 (_________31932), .DIN2 (_________32078),
       .Q (______9__32079));
  or2s1 ____9__503188(.DIN1 (___0_____30866), .DIN2 (_________31853),
       .Q (_________32077));
  nor2s1 ______503189(.DIN1 (_________32075), .DIN2 (_________32074),
       .Q (_________32076));
  and2s1 _______503190(.DIN1 (_________32073), .DIN2
       (____________________________________________21804), .Q
       (_________32318));
  nor2s1 ______503191(.DIN1
       (____________________________________________21804), .DIN2
       (_________32073), .Q (____9_0__32460));
  nor2s1 ______503192(.DIN1 (_________31924), .DIN2 (_________31919),
       .Q (_________32235));
  nor2s1 ____9__503193(.DIN1 (_________32071), .DIN2 (_____00__31894),
       .Q (_________32072));
  nor2s1 ____9__503194(.DIN1 (____0___28380), .DIN2 (_________31861),
       .Q (______0__32070));
  nor2s1 ____9__503195(.DIN1 (________28582), .DIN2 (_________31929),
       .Q (______9__32069));
  nor2s1 ____9__503196(.DIN1 (___00____30605), .DIN2 (_____0___31896),
       .Q (_________32068));
  nnd2s1 ____9__503197(.DIN1 (_____9___31889), .DIN2 (____9_9__32410),
       .Q (_________32067));
  nor2s1 ____9__503198(.DIN1 (_________32065), .DIN2 (_________31909),
       .Q (_________32066));
  nnd2s1 ____9__503199(.DIN1 (_________31880), .DIN2 (____9____32424),
       .Q (_________32064));
  nor2s1 ____9__503200(.DIN1 (___0____25136), .DIN2 (_____09__31902),
       .Q (_________32063));
  nnd2s1 ____9__503201(.DIN1 (_________31867), .DIN2 (___9____26906),
       .Q (_________32062));
  nnd2s1 ____9__503202(.DIN1 (_________31876), .DIN2 (__9_____29775),
       .Q (_________32061));
  nor2s1 ____9__503203(.DIN1 (___0____25136), .DIN2 (_________31871),
       .Q (______0__32060));
  nor2s1 ____9_503204(.DIN1 (_________32058), .DIN2 (_________31862),
       .Q (______9__32059));
  nor2s1 ____9__503205(.DIN1 (_________32056), .DIN2 (_________31869),
       .Q (_________32057));
  nnd2s1 ____9__503206(.DIN1 (_____9___31893), .DIN2 (____9_9__32410),
       .Q (_________32055));
  nor2s1 ____9__503207(.DIN1 (_________32130), .DIN2 (_________31858),
       .Q (_________32054));
  nor2s1 ____9__503208(.DIN1 (____9____33386), .DIN2 (_________40946),
       .Q (_________32053));
  nnd2s1 ____9__503209(.DIN1 (_____9___31887), .DIN2 (________29033),
       .Q (_________32052));
  nor2s1 ____9_503210(.DIN1 (__9_90__29887), .DIN2 (_________31859), .Q
       (_________32051));
  nor2s1 ____9_503211(.DIN1 (_____0___41315), .DIN2 (_____9___31892),
       .Q (______0__32050));
  nnd2s1 ____9__503212(.DIN1 (______9__31920), .DIN2 (___0_____30900),
       .Q (______9__32049));
  nor2s1 ____99_503213(.DIN1 (________27266), .DIN2 (_________31877),
       .Q (_________32048));
  nnd2s1 ____99_503214(.DIN1 (______0__31911), .DIN2 (_____0__29296),
       .Q (_________32047));
  nnd2s1 ____99_503215(.DIN1 (______9__31864), .DIN2 (____00___31511),
       .Q (_________32046));
  nnd2s1 ____00_503216(.DIN1 (_________31860), .DIN2 (________29299),
       .Q (_________32045));
  nnd2s1 ____00_503217(.DIN1 (______0__31931), .DIN2 (_____9__28580),
       .Q (_________32044));
  nor2s1 ____503218(.DIN1 (_________32042), .DIN2 (_____9___31890), .Q
       (_________32043));
  nor2s1 ____0__503219(.DIN1 (___99___29635), .DIN2 (_____0___31899),
       .Q (_________32041));
  nor2s1 ____0__503220(.DIN1 (___0900), .DIN2 (_________31857), .Q
       (______0__32040));
  nor2s1 ____09_503221(.DIN1 (________27199), .DIN2 (______9__31854),
       .Q (______9__32039));
  nnd2s1 _______503222(.DIN1 (_________31934), .DIN2 (________29181),
       .Q (_________32038));
  nnd2s1 _______503223(.DIN1 (_________31936), .DIN2 (_________31749),
       .Q (_________32037));
  nnd2s1 _______503224(.DIN1 (_____0___31801), .DIN2 (_____09__31708),
       .Q (_________32036));
  nor2s1 ____9__503225(.DIN1 (____00___31505), .DIN2 (_____0___31799),
       .Q (_________32035));
  xor2s1 _____0_503226(.DIN1 (_________31729), .DIN2 (_________38385),
       .Q (_________32034));
  nor2s1 _______503227(.DIN1 (_________32032), .DIN2 (_________32031),
       .Q (_________32033));
  and2s1 ______503228(.DIN1 (_________32031), .DIN2 (_________32032),
       .Q (______0__32030));
  nnd2s1 ____9_503229(.DIN1 (_____99__31794), .DIN2 (_____0__29175), .Q
       (______9__32029));
  nor2s1 ____9__503230(.DIN1 (_________31673), .DIN2 (_________31826),
       .Q (_________32028));
  nnd2s1 _______503231(.DIN1 (_________32026), .DIN2 (_________32024),
       .Q (_________32027));
  nor2s1 _______503232(.DIN1 (_________32024), .DIN2 (_________32026),
       .Q (_________32025));
  nnd2s1 ____9__503233(.DIN1 (_________31830), .DIN2 (_________32022),
       .Q (_________32023));
  nnd2s1 ____9__503234(.DIN1 (_____09__31804), .DIN2 (___0_____30943),
       .Q (_________32021));
  nnd2s1 _______503235(.DIN1 (_________31829), .DIN2 (______9__32019),
       .Q (______0__32020));
  or2s1 _______503236(.DIN1 (_____9___32376), .DIN2 (_________31828),
       .Q (_________32018));
  or2s1 _____503237(.DIN1 (______0__31641), .DIN2 (_________32016), .Q
       (_________32017));
  nnd2s1 _______503238(.DIN1 (_________32012), .DIN2 (______0__34524),
       .Q (_________32015));
  xor2s1 _______503239(.DIN1 (___90____39055), .DIN2 (_________36578),
       .Q (_________32014));
  nor2s1 _______503240(.DIN1 (___0_9___31399), .DIN2 (_________32012),
       .Q (_________32013));
  nor2s1 _______503241(.DIN1 (_________33973), .DIN2 (_________32016),
       .Q (_________32011));
  and2s1 _______503242(.DIN1 (_________32016), .DIN2 (_________33973),
       .Q (______0__32010));
  nor2s1 _______503243(.DIN1 (_________32159), .DIN2 (______0__31805),
       .Q (______9__32009));
  nnd2s1 _______503244(.DIN1 (_____9___31788), .DIN2 (_____9__28246),
       .Q (_________32008));
  nor2s1 _______503245(.DIN1 (___90___28652), .DIN2 (______9__31814),
       .Q (_________32007));
  nor2s1 _____9_503246(.DIN1 (__9_____30318), .DIN2 (_________31777),
       .Q (_________32006));
  nnd2s1 _____9_503247(.DIN1 (_____00__31795), .DIN2 (_________32004),
       .Q (_________32005));
  nor2s1 _____9_503248(.DIN1 (___0____27887), .DIN2 (_________31810),
       .Q (_________32003));
  nor2s1 ____90_503249(.DIN1 (_________32001), .DIN2 (_____0___31797),
       .Q (_________32002));
  nor2s1 ____9__503250(.DIN1 (_____09__31999), .DIN2 (_________31816),
       .Q (______0__32000));
  nnd2s1 ____9__503251(.DIN1 (_____9___31787), .DIN2 (___0_____30753),
       .Q (_____0___31998));
  nnd2s1 ____9__503252(.DIN1 (_________31818), .DIN2 (_________31731),
       .Q (_____0___31997));
  nor2s1 ____9__503253(.DIN1 (____0___27576), .DIN2 (_________31812),
       .Q (_____0___31996));
  nor2s1 ____9__503254(.DIN1 (_____0___31994), .DIN2 (_________31832),
       .Q (_____0___31995));
  nnd2s1 ____9__503255(.DIN1 (_________31852), .DIN2 (__9__9__30290),
       .Q (_____0___31993));
  nor2s1 ____9_503256(.DIN1 (_____0___31991), .DIN2 (_____0___31800),
       .Q (_____0___31992));
  nnd2s1 ____9__503257(.DIN1 (_____0___31798), .DIN2 (___0_____30997),
       .Q (_____00__31990));
  and2s1 ______503258(.DIN1 (_____99__31989), .DIN2 (________28845), .Q
       (______9__32175));
  hi1s1 _____9_503259(.DIN (_________32073), .Q (______9__32146));
  nor2s1 ____9__503260(.DIN1 (___009__25134), .DIN2 (_________31806),
       .Q (_________32158));
  nnd2s1 ____9_503261(.DIN1 (_________31808), .DIN2 (_________31882),
       .Q (_________32161));
  nor2s1 _____9_503262(.DIN1 (___0__0__31033), .DIN2 (______0__31835),
       .Q (_____0___36733));
  nor2s1 ______503263(.DIN1 (________27603), .DIN2 (_____99__31989), .Q
       (_____90__32176));
  dffacs1 _______________________503264(.CLRB (reset), .CLK (clk), .DIN
       (_________31807), .QN (_____________________21705));
  nor2s1 ____9__503265(.DIN1 (_____0___33821), .DIN2 (_____9___31786),
       .Q (_____9___31988));
  and2s1 ____9__503266(.DIN1 (_____0___31796), .DIN2 (_____90__32080),
       .Q (_____9___31987));
  or2s1 ____9__503267(.DIN1 (_____9___32376), .DIN2 (_____9___31985),
       .Q (_____9___31986));
  nnd2s1 ____9_503268(.DIN1 (_________31772), .DIN2 (_________31771),
       .Q (_____9___31984));
  nor2s1 ____99_503269(.DIN1 (___09___27028), .DIN2 (_____90__31785),
       .Q (_____9___31983));
  nnd2s1 ____99_503270(.DIN1 (______0__31776), .DIN2 (____9____32417),
       .Q (_____9___31982));
  nnd2s1 ____503271(.DIN1 (_________31779), .DIN2 (_____9___31697), .Q
       (_____9___31981));
  nnd2s1 ____503272(.DIN1 (_________31770), .DIN2 (_________32078), .Q
       (_____90__31980));
  nor2s1 ____00_503273(.DIN1 (_________31942), .DIN2 (_________31769),
       .Q (______9__31979));
  nor2s1 ____00_503274(.DIN1 (_________32071), .DIN2 (_________31780),
       .Q (_________31978));
  nnd2s1 ____0_503275(.DIN1 (_________31773), .DIN2 (____0____32543),
       .Q (_________31977));
  or2s1 ____0__503276(.DIN1 (______9__32852), .DIN2 (_________31768),
       .Q (_________31976));
  nor2s1 ____9__503277(.DIN1 (_____90__32273), .DIN2 (_________31784),
       .Q (_________31975));
  and2s1 ____0__503278(.DIN1 (______0__31766), .DIN2 (_________31973),
       .Q (_________31974));
  nnd2s1 ____0_503279(.DIN1 (_________31761), .DIN2 (__9__0__29814), .Q
       (_________31972));
  nor2s1 ____0__503280(.DIN1 (______0__31970), .DIN2 (_________31760),
       .Q (_________31971));
  nnd2s1 ____0__503281(.DIN1 (_________31767), .DIN2 (___0__9__30671),
       .Q (______9__31969));
  nnd2s1 ____0__503282(.DIN1 (_________31764), .DIN2 (___0__0__31168),
       .Q (_________31968));
  nnd2s1 ____0__503283(.DIN1 (_________31759), .DIN2 (________28261),
       .Q (_________31967));
  nnd2s1 ____0_503284(.DIN1 (_________31758), .DIN2 (_________32078),
       .Q (_________31966));
  nnd2s1 ____0__503285(.DIN1 (_________31757), .DIN2 (________28386),
       .Q (_________31965));
  nnd2s1 ____0__503286(.DIN1 (______0__31756), .DIN2 (___0_____31204),
       .Q (_________31964));
  or2s1 ____0_503287(.DIN1 (_________32042), .DIN2 (______9__31755), .Q
       (_________31963));
  nor2s1 ____503288(.DIN1 (_____0__28863), .DIN2 (_________31833), .Q
       (_________31962));
  nor2s1 _____0_503289(.DIN1 (___09_9__31446), .DIN2 (_________31839),
       .Q (_________31961));
  nor2s1 _____0_503290(.DIN1 (_________31827), .DIN2 (_________31763),
       .Q (______0__31960));
  nor2s1 _____503291(.DIN1 (_________31958), .DIN2 (_________31840), .Q
       (______9__31959));
  nor2s1 _______503292(.DIN1 (___0_____30656), .DIN2 (_________31842),
       .Q (_________31957));
  nor2s1 _______503293(.DIN1 (_________31955), .DIN2 (_________31754),
       .Q (_________31956));
  and2s1 ______503294(.DIN1 (______9__31844), .DIN2 (_________31953),
       .Q (_________31954));
  nor2s1 _______503295(.DIN1 (________28936), .DIN2 (_________31837),
       .Q (_________31952));
  or2s1 _______503296(.DIN1 (______0__31950), .DIN2 (_____9___31790),
       .Q (_________31951));
  nnd2s1 _______503297(.DIN1 (_________31847), .DIN2 (___0_____31237),
       .Q (______9__31949));
  nor2s1 ______503298(.DIN1 (_________33742), .DIN2 (______0__31845),
       .Q (_________31948));
  nnd2s1 _______503299(.DIN1 (_________31838), .DIN2 (_________31868),
       .Q (_________31947));
  nnd2s1 _______503300(.DIN1 (_________31849), .DIN2 (__9_0_), .Q
       (_________31946));
  nnd2s1 ______503301(.DIN1 (_________31850), .DIN2 (_________31944),
       .Q (_________31945));
  or2s1 _______503302(.DIN1 (_________31942), .DIN2 (_________31841),
       .Q (_________31943));
  nnd2s1 _______503303(.DIN1 (_________31851), .DIN2 (______0__32196),
       .Q (_________31941));
  nor2s1 _____9_503304(.DIN1 (___0_____31277), .DIN2 (_________31753),
       .Q (______0__31940));
  nor2s1 ____0__503305(.DIN1 (___9____27788), .DIN2 (_________31782),
       .Q (______0__32137));
  dffacs1 _______________________503306(.CLRB (reset), .CLK (clk), .DIN
       (_________31774), .QN (_____________________21708));
  nor2s1 ____0__503307(.DIN1 (_________31938), .DIN2 (_________31913),
       .Q (______9__31939));
  nnd2s1 ______503308(.DIN1 (_________31674), .DIN2 (________26299), .Q
       (_________31937));
  and2s1 _______503309(.DIN1 (______0__31671), .DIN2 (_________31935),
       .Q (_________31936));
  and2s1 _______503310(.DIN1 (_________31669), .DIN2 (_________31933),
       .Q (_________31934));
  nor2s1 ____0__503311(.DIN1 (___0_____31268), .DIN2 (_____9___31692),
       .Q (_________31932));
  nor2s1 ____0__503312(.DIN1 (___09____31457), .DIN2 (_____9___31691),
       .Q (______0__31931));
  xnr2s1 _______503313(.DIN1
       (__________________________________________________________________21986),
       .DIN2 (______9__31834), .Q (______9__31930));
  nnd2s1 ____0__503314(.DIN1 (______0__31737), .DIN2 (___90___27744),
       .Q (_________31929));
  nor2s1 _______503315(.DIN1 (________26545), .DIN2 (____0_9__32507),
       .Q (_________31928));
  nor2s1 _______503316(.DIN1 (_________36578), .DIN2 (_________31925),
       .Q (_________31927));
  and2s1 _______503317(.DIN1 (_________31925), .DIN2 (_________36578),
       .Q (_________31926));
  nor2s1 _____9_503318(.DIN1 (_________32918), .DIN2 (_________31713),
       .Q (_________31924));
  nnd2s1 ____9__503319(.DIN1 (_________31723), .DIN2 (____0___27396),
       .Q (_________31923));
  and2s1 ____9_503320(.DIN1 (_________31722), .DIN2 (______0__31921),
       .Q (_________31922));
  nor2s1 ____0__503321(.DIN1 (__990___30455), .DIN2 (_________31730),
       .Q (______9__31920));
  nor2s1 ____9__503322(.DIN1
       (______________________________________________________________________________________0__22096),
       .DIN2 (_________31719), .Q (_________31919));
  nor2s1 ____99_503323(.DIN1 (___0_____31282), .DIN2 (_________31714),
       .Q (_________31918));
  nor2s1 ____99_503324(.DIN1 (___09_9__31475), .DIN2 (______9__31717),
       .Q (_________31917));
  nor2s1 _______503325(.DIN1 (______9__31670), .DIN2 (___09____31491),
       .Q (_________31916));
  nnd2s1 ____0__503326(.DIN1 (_________31712), .DIN2 (_________31628),
       .Q (_________31915));
  nnd2s1 ____0_503327(.DIN1 (_________31913), .DIN2 (_________32145),
       .Q (_________31914));
  xnr2s1 ____0_503328(.DIN1 (______0__35711), .DIN2 (____9____36110),
       .Q (_________31912));
  and2s1 ____0__503329(.DIN1 (_____9___31693), .DIN2 (______9__31910),
       .Q (______0__31911));
  nnd2s1 ____0__503330(.DIN1 (_____0___31704), .DIN2 (___0_____30968),
       .Q (_________31909));
  or2s1 ____0__503331(.DIN1 (_________32042), .DIN2 (______9__31679),
       .Q (_________31908));
  or2s1 ____0__503332(.DIN1 (_________31906), .DIN2 (_____0___31703),
       .Q (_________31907));
  nnd2s1 ____0__503333(.DIN1 (_____0___31700), .DIN2 (_____0___31702),
       .Q (_________31905));
  nor2s1 ____0__503334(.DIN1 (______0__31903), .DIN2 (_____0___31701),
       .Q (_________31904));
  nor2s1 ____0_503335(.DIN1 (_________32058), .DIN2 (_____99__31698),
       .Q (_____09__31902));
  nnd2s1 ____0__503336(.DIN1 (_____9___31696), .DIN2 (____99__28107),
       .Q (_____0___31901));
  and2s1 _____9_503337(.DIN1 (_____0___31900), .DIN2
       (____________________________________________21805), .Q
       (_________32075));
  nor2s1 _____9_503338(.DIN1
       (____________________________________________21805), .DIN2
       (_____0___31900), .Q (_________32074));
  xor2s1 _______503339(.DIN1 (___0__9__40638), .DIN2 (_____9___33157),
       .Q (_________32073));
  hi1s1 ____9__503340(.DIN (____9____34309), .Q (_____9___34281));
  nor2s1 _______503341(.DIN1 (___0900), .DIN2 (______0__31855), .Q
       (_____0___31899));
  nor2s1 ____0__503342(.DIN1 (______0__32253), .DIN2 (_____90__31689),
       .Q (_____0___31898));
  nor2s1 ____0__503343(.DIN1 (__9_____30385), .DIN2 (_________31685),
       .Q (_____0___31897));
  nnd2s1 ____0_503344(.DIN1 (_________31750), .DIN2 (_____0___31895),
       .Q (_____0___31896));
  or2s1 ____0__503345(.DIN1 (_____0___41315), .DIN2 (______0__31709),
       .Q (_____00__31894));
  nnd2s1 ____0__503346(.DIN1 (_________31683), .DIN2 (____09___31595),
       .Q (_____9___31893));
  nnd2s1 ____0__503347(.DIN1 (_________31682), .DIN2 (_____9___31891),
       .Q (_____9___31892));
  nnd2s1 ____0__503348(.DIN1 (_________31681), .DIN2 (___0_____31175),
       .Q (_____9___31890));
  or2s1 ____09_503349(.DIN1 (______0__41140), .DIN2 (_____9___31695),
       .Q (_____9___31889));
  nnd2s1 ____09_503350(.DIN1 (_________31735), .DIN2 (inData[31]), .Q
       (_____9___31888));
  nor2s1 ____09_503351(.DIN1 (_____9___31886), .DIN2 (_____0___31706),
       .Q (_____9___31887));
  nor2s1 ____09_503352(.DIN1 (______9__31884), .DIN2 (_________31751),
       .Q (_____90__31885));
  and2s1 ____503353(.DIN1 (______0__31728), .DIN2 (_________31882), .Q
       (_________31883));
  nnd2s1 _______503354(.DIN1 (_________31677), .DIN2 (________29248),
       .Q (_________31881));
  nnd2s1 _______503355(.DIN1 (______9__31736), .DIN2 (_________31879),
       .Q (_________31880));
  nor2s1 _______503356(.DIN1 (____0____32539), .DIN2 (_________31676),
       .Q (_________31878));
  nnd2s1 _______503357(.DIN1 (_________31742), .DIN2 (___99___26953),
       .Q (_________31877));
  nor2s1 ______503358(.DIN1 (_____9___33155), .DIN2 (_________31726),
       .Q (_________31876));
  nor2s1 ______503359(.DIN1 (_____0__28220), .DIN2 (_________31744), .Q
       (______0__31875));
  nnd2s1 _______503360(.DIN1 (_____00__31699), .DIN2 (_________31873),
       .Q (______9__31874));
  nnd2s1 _______503361(.DIN1 (_________31684), .DIN2 (___0_00__30740),
       .Q (_________31872));
  nor2s1 _______503362(.DIN1 (_________31870), .DIN2 (______9__31746),
       .Q (_________31871));
  nnd2s1 _______503363(.DIN1 (_________31733), .DIN2 (_________31868),
       .Q (_________31869));
  or2s1 _______503364(.DIN1 (_________31866), .DIN2 (_________31745),
       .Q (_________31867));
  nnd2s1 _______503365(.DIN1 (_________31748), .DIN2 (___0_____30700),
       .Q (______0__31865));
  nor2s1 ______503366(.DIN1 (_________32658), .DIN2 (_________31743),
       .Q (______9__31864));
  nor2s1 _______503367(.DIN1 (__9_____30231), .DIN2 (_________31741),
       .Q (_________31863));
  nnd2s1 ______503368(.DIN1 (_________31739), .DIN2 (_____9__27609), .Q
       (_________31862));
  nnd2s1 _______503369(.DIN1 (_________31740), .DIN2 (__9__9__30056),
       .Q (_________31861));
  nor2s1 ______503370(.DIN1 (___0_9___30731), .DIN2 (_________31752),
       .Q (_________31860));
  nor2s1 _______503371(.DIN1 (____0____32541), .DIN2 (_________31732),
       .Q (_________31859));
  or2s1 _______503372(.DIN1 (_________32056), .DIN2 (_________31686),
       .Q (_________31858));
  nor2s1 ______503373(.DIN1 (________29210), .DIN2 (_________31675), .Q
       (_________31857));
  nnd2s1 _______503374(.DIN1 (______0__31855), .DIN2 (___9____28704),
       .Q (_________31856));
  nnd2s1 _______503375(.DIN1 (_________31672), .DIN2 (__9__0__30206),
       .Q (______9__31854));
  nnd2s1 ____0_503376(.DIN1 (______0__31747), .DIN2 (________28870), .Q
       (_________31853));
  nor2s1 ____0__503377(.DIN1 (___0_____31342), .DIN2 (_____0___31611),
       .Q (_________31852));
  nor2s1 _______503378(.DIN1 (______9__31884), .DIN2 (____0____31561),
       .Q (_________31851));
  and2s1 _______503379(.DIN1 (____0____31585), .DIN2 (_________31873),
       .Q (_________31850));
  nor2s1 _______503380(.DIN1 (________28969), .DIN2 (____0____31564),
       .Q (_________31849));
  nnd2s1 _______503381(.DIN1 (____0____31570), .DIN2 (_________32266),
       .Q (_________31848));
  nor2s1 _______503382(.DIN1 (_________31846), .DIN2 (____0____31567),
       .Q (_________31847));
  or2s1 ______503383(.DIN1 (_________32311), .DIN2 (____0_9__31562), .Q
       (______0__31845));
  nor2s1 _______503384(.DIN1 (_________31843), .DIN2 (____0____31568),
       .Q (______9__31844));
  nnd2s1 _______503385(.DIN1 (____0____31578), .DIN2 (___0_____30654),
       .Q (_________31842));
  nnd2s1 _______503386(.DIN1 (____0_9__31572), .DIN2 (__99____30516),
       .Q (_________31841));
  or2s1 _______503387(.DIN1 (_________33106), .DIN2 (____0____31590),
       .Q (_________31840));
  nnd2s1 _______503388(.DIN1 (____0____31565), .DIN2 (___09____31487),
       .Q (_________31839));
  nor2s1 _______503389(.DIN1 (__99____30485), .DIN2 (____0____31555),
       .Q (_________31838));
  or2s1 _____0_503390(.DIN1 (_________31836), .DIN2 (____0____31557),
       .Q (_________31837));
  and2s1 _______503391(.DIN1 (______9__31834), .DIN2 (___0_0___31030),
       .Q (______0__31835));
  nnd2s1 _____9_503392(.DIN1 (____0____31576), .DIN2 (___0_09__30651),
       .Q (_________31833));
  nnd2s1 ____0__503393(.DIN1 (______0__31613), .DIN2 (_________31831),
       .Q (_________31832));
  nor2s1 ____0__503394(.DIN1 (__9_00__30272), .DIN2 (____09___31601),
       .Q (_________31830));
  nor2s1 _____503395(.DIN1 (________28937), .DIN2 (_________31634), .Q
       (_________31829));
  nor2s1 ____90_503396(.DIN1 (_________31827), .DIN2 (______0__31633),
       .Q (_________31828));
  nnd2s1 ____0_503397(.DIN1 (_____0___31610), .DIN2 (______0__31825),
       .Q (_________31826));
  xor2s1 ____9__503398(.DIN1 (____0____31551), .DIN2 (______9__34088),
       .Q (______9__31824));
  xor2s1 ____99_503399(.DIN1 (____0____31529), .DIN2 (_________38860),
       .Q (_________31823));
  nnd2s1 ____0__503400(.DIN1 (_________31711), .DIN2 (_________31821),
       .Q (_________31822));
  xor2s1 ____0__503401(.DIN1 (_________37687), .DIN2
       (______________________________________________21902), .Q
       (_________31820));
  xnr2s1 ____0__503402(.DIN1
       (__________________________________________________________________21990),
       .DIN2 (______________________________________________21902), .Q
       (_________31819));
  nor2s1 ____0_503403(.DIN1 (_________31817), .DIN2 (____09___31599),
       .Q (_________31818));
  nnd2s1 ____0__503404(.DIN1 (_____9___31791), .DIN2 (______0__31815),
       .Q (_________31816));
  nnd2s1 ____0_503405(.DIN1 (_________31656), .DIN2 (___0____28822), .Q
       (______9__31814));
  nor2s1 ____0_503406(.DIN1 (_________32159), .DIN2 (_________31687),
       .Q (_________31813));
  nnd2s1 ____0__503407(.DIN1 (______0__31623), .DIN2 (_________31811),
       .Q (_________31812));
  nor2s1 ____0__503408(.DIN1 (_________31809), .DIN2 (_________31629),
       .Q (_________31810));
  or2s1 ____0__503409(.DIN1 (______________22067), .DIN2
       (______9__31727), .Q (_________31808));
  nnd2s1 ____0__503410(.DIN1 (_________31619), .DIN2 (_________34163),
       .Q (_________31807));
  nnd2s1 ____0__503411(.DIN1 (_________31662), .DIN2 (___0_9__28814),
       .Q (_________31806));
  nor2s1 ____0__503412(.DIN1 (_____0___33821), .DIN2 (_________31652),
       .Q (______0__31805));
  nor2s1 ____0__503413(.DIN1 (_____0___31803), .DIN2 (_________31621),
       .Q (_____09__31804));
  nnd2s1 ____0__503414(.DIN1 (_________31734), .DIN2 (___0____26094),
       .Q (_____0___31802));
  nnd2s1 ____9_503415(.DIN1 (_________31631), .DIN2 (_________33000),
       .Q (_________32012));
  hi1s1 _______503416(.DIN (_____0___31900), .Q (_________32031));
  xor2s1 ____0__503417(.DIN1 (___0_____40642), .DIN2 (______0__31718),
       .Q (____9____34309));
  nor2s1 ______503418(.DIN1 (_____9__28137), .DIN2 (_________31637), .Q
       (_________32026));
  nor2s1 _______503419(.DIN1 (_________31666), .DIN2 (_________31925),
       .Q (_____99__31989));
  xor2s1 ____0__503420(.DIN1 (____0____31525), .DIN2 (___9_____39384),
       .Q (_________32016));
  and2s1 _______503421(.DIN1 (____09___31596), .DIN2 (_________31678),
       .Q (_____0___31801));
  nnd2s1 ____0__503422(.DIN1 (_____0___31606), .DIN2 (_____0___31609),
       .Q (_____0___31800));
  nnd2s1 ____0__503423(.DIN1 (____099__31602), .DIN2 (___0_____31362),
       .Q (_____0___31799));
  nor2s1 ____0__503424(.DIN1 (_____0___31991), .DIN2 (_____0___31607),
       .Q (_____0___31798));
  nor2s1 ____0_503425(.DIN1 (__9_____30339), .DIN2 (_________31638), .Q
       (_____0___31797));
  nor2s1 _____0_503426(.DIN1 (_____9__26275), .DIN2 (_________31653),
       .Q (_____0___31796));
  nor2s1 _____0_503427(.DIN1 (___0_____30697), .DIN2 (_________31618),
       .Q (_____00__31795));
  nor2s1 ______503428(.DIN1 (___0_____31073), .DIN2 (_________31654),
       .Q (_____99__31794));
  nor2s1 _______503429(.DIN1 (___0__9__30890), .DIN2 (_____0___31605),
       .Q (_____9___31793));
  nor2s1 _______503430(.DIN1 (_________32159), .DIN2 (_____9___31791),
       .Q (_____9___31792));
  or2s1 _____0_503431(.DIN1 (_____9___31789), .DIN2 (____0____31558),
       .Q (_____9___31790));
  nor2s1 _______503432(.DIN1 (__9_0___30179), .DIN2 (_________31644),
       .Q (_____9___31788));
  nnd2s1 _______503433(.DIN1 (_____00__31603), .DIN2 (________25544),
       .Q (_____9___31787));
  nnd2s1 _______503434(.DIN1 (______9__31650), .DIN2 (_________32114),
       .Q (_____9___31786));
  or2s1 _______503435(.DIN1 (______0__41150), .DIN2 (_________31649),
       .Q (_____90__31785));
  nor2s1 ______503436(.DIN1 (_________31783), .DIN2 (_________31614),
       .Q (_________31784));
  nnd2s1 _______503437(.DIN1 (_________31664), .DIN2 (_________31781),
       .Q (_________31782));
  nnd2s1 _______503438(.DIN1 (____09___31600), .DIN2 (__9_0___29899),
       .Q (_________31780));
  and2s1 _______503439(.DIN1 (_________31659), .DIN2 (_________31778),
       .Q (_________31779));
  nnd2s1 _______503440(.DIN1 (____090__31593), .DIN2 (____99__28199),
       .Q (_________31777));
  nor2s1 _______503441(.DIN1 (__999___30543), .DIN2 (_________31658),
       .Q (______0__31776));
  nor2s1 _______503442(.DIN1 (____0____32539), .DIN2 (______0__31651),
       .Q (______9__31775));
  nnd2s1 _______503443(.DIN1 (______0__31661), .DIN2 (_________34163),
       .Q (_________31774));
  or2s1 _______503444(.DIN1 (______0__41140), .DIN2 (_________31615),
       .Q (_________31773));
  nnd2s1 ______503445(.DIN1 (____9____36110), .DIN2 (_____9___38610),
       .Q (_________31772));
  nnd2s1 _______503446(.DIN1 (____0____31571), .DIN2 (____0_9__31552),
       .Q (_________31771));
  nor2s1 _______503447(.DIN1 (_________31783), .DIN2 (_________31663),
       .Q (_________31770));
  or2s1 _______503448(.DIN1 (______9__32852), .DIN2 (_________31636),
       .Q (_________31769));
  nnd2s1 ____0__503449(.DIN1 (_____0___31608), .DIN2 (___0_____31040),
       .Q (_________31768));
  nor2s1 _______503450(.DIN1 (___00_9__30621), .DIN2 (____09___31594),
       .Q (_________31767));
  and2s1 _____9_503451(.DIN1 (____0____31575), .DIN2 (______9__31765),
       .Q (______0__31766));
  nor2s1 _____9_503452(.DIN1 (________27040), .DIN2 (____0____31580),
       .Q (_________31764));
  or2s1 _____0_503453(.DIN1 (_________31762), .DIN2 (____0_9__31592),
       .Q (_________31763));
  and2s1 _______503454(.DIN1 (____0____31588), .DIN2 (___9____28693),
       .Q (_________31761));
  nnd2s1 _______503455(.DIN1 (____0____31587), .DIN2 (______0__31815),
       .Q (_________31760));
  nor2s1 _______503456(.DIN1 (________29217), .DIN2 (____0_0__31573),
       .Q (_________31759));
  nor2s1 ______503457(.DIN1 (_____9___33059), .DIN2 (____0____31586),
       .Q (_________31758));
  nor2s1 ______503458(.DIN1 (________28060), .DIN2 (____0_0__31563), .Q
       (_________31757));
  and2s1 ______503459(.DIN1 (____0____31569), .DIN2 (___00____30556),
       .Q (______0__31756));
  or2s1 _______503460(.DIN1 (___0_____31381), .DIN2 (____0_9__31582),
       .Q (______9__31755));
  nnd2s1 _____0_503461(.DIN1 (____0_0__31583), .DIN2 (___0_____31084),
       .Q (_________31754));
  nnd2s1 _______503462(.DIN1 (____09___31597), .DIN2 (__9_9___29801),
       .Q (_________31753));
  and2s1 _______503463(.DIN1 (_________31645), .DIN2 (______0__31921),
       .Q (_____9___31985));
  dffacs1 ________________________________________________503464(.CLRB
       (reset), .CLK (clk), .DIN (_________31635), .Q
       (_______________________________________________________________9__21995));
  nor2s1 _______503465(.DIN1 (___0____25136), .DIN2 (____00___31510),
       .Q (_________31752));
  nnd2s1 _____503466(.DIN1 (___0999__31502), .DIN2 (____9_9__32410), .Q
       (_________31751));
  and2s1 _____9_503467(.DIN1 (___09____31482), .DIN2 (_________31749),
       .Q (_________31750));
  nor2s1 _____9_503468(.DIN1 (________29230), .DIN2 (___09_0__31486),
       .Q (_________31748));
  nor2s1 ______503469(.DIN1 (_________31958), .DIN2 (____0____31528),
       .Q (______0__31747));
  nnd2s1 _______503470(.DIN1 (___09____31490), .DIN2 (___0_____31266),
       .Q (______9__31746));
  nnd2s1 _____503471(.DIN1 (___09____31488), .DIN2 (_____90__32080), .Q
       (_________31745));
  nor2s1 _______503472(.DIN1 (____0____32541), .DIN2 (___09____31489),
       .Q (_________31744));
  nnd2s1 _______503473(.DIN1 (___09____31474), .DIN2 (___0_____30917),
       .Q (_________31743));
  nor2s1 _______503474(.DIN1 (________26649), .DIN2 (____009__31512),
       .Q (_________31742));
  nnd2s1 ______503475(.DIN1 (___0_0___31121), .DIN2 (___09____31473),
       .Q (_________31741));
  nor2s1 _______503476(.DIN1 (_________41128), .DIN2 (_________41361),
       .Q (_________31740));
  and2s1 _______503477(.DIN1 (___099___31500), .DIN2 (_________31738),
       .Q (_________31739));
  nnd2s1 _______503478(.DIN1 (___09_0__31476), .DIN2 (________25545),
       .Q (______0__31737));
  nor2s1 _______503479(.DIN1 (_________32058), .DIN2 (___099___31498),
       .Q (______9__31736));
  hi1s1 ______503480(.DIN (_________31734), .Q (_________31735));
  nor2s1 _____503481(.DIN1 (_________31846), .DIN2 (___099___31495), .Q
       (_________31733));
  and2s1 _______503482(.DIN1 (___09____31479), .DIN2 (_________31731),
       .Q (_________31732));
  nor2s1 _____0_503483(.DIN1 (___0____25136), .DIN2 (___099___31497),
       .Q (_________31730));
  xor2s1 _______503484(.DIN1 (___09____31454), .DIN2 (___0_____31247),
       .Q (_________31729));
  hi1s1 ______503485(.DIN (______9__31727), .Q (______0__31728));
  nnd2s1 _______503486(.DIN1 (___09____31470), .DIN2 (_________31725),
       .Q (_________31726));
  nnd2s1 ____0_503487(.DIN1 (____0____31537), .DIN2 (_________41196),
       .Q (_________31724));
  and2s1 ____0__503488(.DIN1 (____0____31536), .DIN2 (________26629),
       .Q (_________31723));
  and2s1 ____09_503489(.DIN1 (____0____31548), .DIN2 (_________33692),
       .Q (_________31722));
  nnd2s1 ____09_503490(.DIN1 (_________31624), .DIN2 (_________31720),
       .Q (_________31721));
  nor2s1 _______503491(.DIN1 (___99___26044), .DIN2 (______0__31718),
       .Q (_________31719));
  and2s1 _______503492(.DIN1 (_________31716), .DIN2 (_________31715),
       .Q (______9__31717));
  nnd2s1 _______503493(.DIN1 (____0_0__31543), .DIN2 (__99____30513),
       .Q (_________31714));
  nor2s1 _______503494(.DIN1 (________25275), .DIN2 (______0__31718),
       .Q (_________31713));
  nor2s1 _______503495(.DIN1 (____0____31541), .DIN2 (____0____31544),
       .Q (_________31712));
  hi1s1 _____0_503496(.DIN (_________31711), .Q (_________31913));
  xor2s1 _______503497(.DIN1 (____9___28468), .DIN2 (_________40949),
       .Q (_____0___31900));
  or2s1 ____0__503498(.DIN1 (___9_____39582), .DIN2 (_________31710),
       .Q (____0_9__32507));
  nor2s1 ______503499(.DIN1 (____0_0__31533), .DIN2 (___09____31441),
       .Q (_________36578));
  nnd2s1 _______503500(.DIN1 (___09____31481), .DIN2 (_____09__31708),
       .Q (______0__31709));
  nnd2s1 _______503501(.DIN1 (____0____31521), .DIN2 (________27711),
       .Q (_____0___31707));
  nnd2s1 _____9_503502(.DIN1 (____0____31549), .DIN2 (________29338),
       .Q (_____0___31706));
  and2s1 _____9_503503(.DIN1 (___09____31492), .DIN2 (__9_____30104),
       .Q (_____0___31705));
  nor2s1 _____9_503504(.DIN1 (___09____31429), .DIN2 (____0____31518),
       .Q (_____0___31704));
  or2s1 _____0_503505(.DIN1 (____0____31591), .DIN2 (____0____31516),
       .Q (_____0___31703));
  nor2s1 _____0_503506(.DIN1 (___0_____30815), .DIN2 (___09____31471),
       .Q (_____0___31702));
  nnd2s1 ______503507(.DIN1 (____0____31515), .DIN2 (________28583), .Q
       (_____0___31701));
  nor2s1 _______503508(.DIN1 (__9__0__29936), .DIN2 (___09____31477),
       .Q (_____0___31700));
  nor2s1 _______503509(.DIN1 (__9__0__29956), .DIN2 (___09____31483),
       .Q (_____00__31699));
  nnd2s1 _______503510(.DIN1 (____0____31514), .DIN2 (_____9___31697),
       .Q (_____99__31698));
  nor2s1 _______503511(.DIN1 (________28343), .DIN2 (____0_0__31513),
       .Q (_____9___31696));
  nnd2s1 ______503512(.DIN1 (____0____31546), .DIN2 (_____9___31694),
       .Q (_____9___31695));
  and2s1 _______503513(.DIN1 (___09_9__31485), .DIN2 (____0___29371),
       .Q (_____9___31693));
  nnd2s1 _______503514(.DIN1 (____0____31524), .DIN2 (____0____31554),
       .Q (_____9___31692));
  or2s1 _______503515(.DIN1 (_____9___31690), .DIN2 (____0____31526),
       .Q (_____9___31691));
  and2s1 _______503516(.DIN1 (____0_9__31522), .DIN2 (______9__31688),
       .Q (_____90__31689));
  nnd2s1 _______503517(.DIN1 (____00___31504), .DIN2 (___0_0___31119),
       .Q (_________31686));
  or2s1 _______503518(.DIN1 (__9_9___29799), .DIN2 (____0____31539), .Q
       (_________31685));
  nor2s1 _______503519(.DIN1 (___0_____31191), .DIN2 (____0____31540),
       .Q (_________31684));
  and2s1 ______503520(.DIN1 (___09____31484), .DIN2 (___090___31415),
       .Q (_________31683));
  and2s1 _______503521(.DIN1 (____00___31508), .DIN2 (___0_____30903),
       .Q (_________31682));
  and2s1 _______503522(.DIN1 (___09_9__31493), .DIN2 (___0_____30979),
       .Q (_________31681));
  nor2s1 _______503523(.DIN1 (___0_9___31018), .DIN2 (____0____31520),
       .Q (______0__31680));
  nnd2s1 ______503524(.DIN1 (____00___31506), .DIN2 (_________31678),
       .Q (______9__31679));
  nor2s1 ______503525(.DIN1 (________29346), .DIN2 (___099___31501), .Q
       (_________31677));
  and2s1 _____9_503526(.DIN1 (___09____31468), .DIN2 (_____0___41313),
       .Q (_________31676));
  nnd2s1 _______503527(.DIN1 (___09_0__31466), .DIN2 (___00____30562),
       .Q (_________31675));
  or2s1 _______503528(.DIN1 (_________31673), .DIN2 (___09____31463),
       .Q (_________31674));
  nor2s1 _______503529(.DIN1 (________28975), .DIN2 (___09____31459),
       .Q (_________31672));
  nor2s1 _____503530(.DIN1 (___09___27915), .DIN2 (___09____31462), .Q
       (______0__31671));
  nor2s1 _______503531(.DIN1 (___0__9__30890), .DIN2 (___09____31460),
       .Q (______9__31670));
  nor2s1 _______503532(.DIN1 (_________31668), .DIN2 (___09____31464),
       .Q (_________31669));
  nor2s1 _______503533(.DIN1 (_________31667), .DIN2 (___09____31458),
       .Q (______0__31855));
  xor2s1 ____00_503534(.DIN1 (___0_____31332), .DIN2 (_________41264),
       .Q (_________31666));
  nor2s1 _____9_503535(.DIN1 (___99___25116), .DIN2 (___090___31411),
       .Q (_________31665));
  nor2s1 _____9_503536(.DIN1 (___0_90__31108), .DIN2 (___0_____31393),
       .Q (_________31664));
  or2s1 _______503537(.DIN1 (_________32056), .DIN2 (___0_____31386),
       .Q (_________31663));
  and2s1 _____9_503538(.DIN1 (___0_9___31402), .DIN2 (_____90__33327),
       .Q (_________31662));
  and2s1 _______503539(.DIN1 (___09____31433), .DIN2 (______9__31660),
       .Q (______0__31661));
  and2s1 _______503540(.DIN1 (___09_9__31436), .DIN2 (_________31738),
       .Q (_________31659));
  nnd2s1 _______503541(.DIN1 (___09____31423), .DIN2 (___0__9__30661),
       .Q (_________31658));
  xor2s1 _______503542(.DIN1 (___0_____31248), .DIN2 (_____9___34189),
       .Q (_________31657));
  and2s1 _______503543(.DIN1 (___09____31439), .DIN2 (_________31655),
       .Q (_________31656));
  nnd2s1 _______503544(.DIN1 (___0__9__31397), .DIN2 (________28281),
       .Q (_________31654));
  nnd2s1 ______503545(.DIN1 (___09____31425), .DIN2 (______9__33575),
       .Q (_________31653));
  nnd2s1 _____503546(.DIN1 (___09_0__31427), .DIN2 (_________33016), .Q
       (_________31652));
  nor2s1 _____0_503547(.DIN1 (___9____27800), .DIN2 (___0_____31395),
       .Q (______0__31651));
  and2s1 ______503548(.DIN1 (___0_____31384), .DIN2 (_____0___33721),
       .Q (______9__31650));
  nnd2s1 _____0_503549(.DIN1 (_________31646), .DIN2 (_________31648),
       .Q (_________31649));
  nor2s1 _____0_503550(.DIN1 (_________32159), .DIN2 (_________31646),
       .Q (_________31647));
  nor2s1 ______503551(.DIN1 (_________31762), .DIN2 (___0_____31392),
       .Q (_________31645));
  nnd2s1 _______503552(.DIN1 (___0__0__31388), .DIN2 (________27495),
       .Q (_________31644));
  nnd2s1 _______503553(.DIN1 (___099___31499), .DIN2 (______9__32753),
       .Q (_________31643));
  nnd2s1 ____9__503554(.DIN1 (_________31639), .DIN2 (______9__31640),
       .Q (_________31642));
  nor2s1 ____9__503555(.DIN1 (______9__31640), .DIN2 (_________31639),
       .Q (______0__31641));
  nnd2s1 _____0_503556(.DIN1 (___09____31430), .DIN2 (________27179),
       .Q (_________31638));
  nor2s1 ____9__503557(.DIN1 (_____0__28138), .DIN2 (_________40949),
       .Q (_________31637));
  or2s1 _______503558(.DIN1 (_________31783), .DIN2 (___09_0__31447),
       .Q (_________31636));
  or2s1 _____0_503559(.DIN1 (________25794), .DIN2 (___0_____31389), .Q
       (_________31635));
  nnd2s1 ____0_503560(.DIN1 (___09____31445), .DIN2 (___0_____31162),
       .Q (_________31634));
  nnd2s1 ____0__503561(.DIN1 (___09____31442), .DIN2 (______9__31632),
       .Q (______0__31633));
  nor2s1 ____0__503562(.DIN1 (_________33742), .DIN2 (___09____31444),
       .Q (_________31631));
  hi1s1 _____0_503563(.DIN (_________31710), .Q (_________31630));
  nor2s1 _____503564(.DIN1 (____0___28479), .DIN2 (___09____31421), .Q
       (_________31629));
  xor2s1 _______503565(.DIN1 (___0_0___31313), .DIN2 (_________38533),
       .Q (_________31628));
  xor2s1 _______503566(.DIN1 (___9_0__26873), .DIN2 (_________34034),
       .Q (_________31627));
  or2s1 _____503567(.DIN1 (_________32001), .DIN2 (___09____31432), .Q
       (_________31626));
  hi1s1 _______503568(.DIN (_________31624), .Q (_________31625));
  and2s1 _______503569(.DIN1 (___09____31448), .DIN2 (_________31935),
       .Q (______0__31623));
  nor2s1 _______503570(.DIN1 (____9___26773), .DIN2 (___09____31440),
       .Q (______9__31622));
  nnd2s1 ______503571(.DIN1 (___0_____31382), .DIN2 (___0__9__31260),
       .Q (_________31621));
  nnd2s1 _____503572(.DIN1 (___09____31452), .DIN2 (_________31715), .Q
       (_________31620));
  and2s1 _____9_503573(.DIN1 (___0_99__31407), .DIN2 (___99___29636),
       .Q (_________31619));
  nnd2s1 _____9_503574(.DIN1 (___09____31434), .DIN2 (___0_9__27902),
       .Q (_________31618));
  nnd2s1 _______503575(.DIN1 (_________31616), .DIN2 (______9__32360),
       .Q (_________31882));
  hi1s1 _____0_503576(.DIN (_________31617), .Q (______0__32843));
  nor2s1 _______503577(.DIN1 (_________34207), .DIN2 (___09_0__31437),
       .Q (_________31687));
  nnd2s1 ____9__503578(.DIN1 (___09____31450), .DIN2 (___09____31453),
       .Q (______9__31834));
  nnd2s1 _______503579(.DIN1 (___09_0__31456), .DIN2 (______0__35853),
       .Q (_________31711));
  nor2s1 _______503580(.DIN1 (______9__32360), .DIN2 (_________31616),
       .Q (______9__31727));
  xor2s1 ____0__503581(.DIN1 (___0_____31331), .DIN2 (_________37864),
       .Q (_________31925));
  dffacs1 _______________________________________________503582(.CLRB
       (reset), .CLK (clk), .DIN (___09____31431), .QN
       (_____________________________________________21928));
  or2s1 _____9_503583(.DIN1 (_____0___41315), .DIN2 (___0_90__31398),
       .Q (_________31615));
  nnd2s1 _______503584(.DIN1 (___0_____31390), .DIN2 (___0__0__30787),
       .Q (_________31614));
  and2s1 _______503585(.DIN1 (___09____31422), .DIN2 (_____09__31612),
       .Q (______0__31613));
  nor2s1 _______503586(.DIN1 (____0____32541), .DIN2 (___09____31420),
       .Q (_____0___31611));
  and2s1 _______503587(.DIN1 (___0__9__31387), .DIN2 (_____0___31609),
       .Q (_____0___31610));
  nor2s1 _______503588(.DIN1 (___0__0__30872), .DIN2 (___09____31419),
       .Q (_____0___31608));
  nnd2s1 ______503589(.DIN1 (___09____31418), .DIN2 (___0_____31173),
       .Q (_____0___31607));
  nor2s1 _______503590(.DIN1 (___00____30589), .DIN2 (___09_0__31417),
       .Q (_____0___31606));
  nor2s1 _______503591(.DIN1 (_____0___31604), .DIN2 (___0909__31416),
       .Q (_____0___31605));
  nnd2s1 _______503592(.DIN1 (___090___31414), .DIN2 (_____9__29542),
       .Q (_____00__31603));
  nor2s1 _______503593(.DIN1 (_________41156), .DIN2 (___090___31412),
       .Q (____099__31602));
  nnd2s1 _______503594(.DIN1 (___0_9___31406), .DIN2 (_____9___31891),
       .Q (____09___31601));
  and2s1 _______503595(.DIN1 (___090___31409), .DIN2 (______0__31825),
       .Q (____09___31600));
  nnd2s1 _______503596(.DIN1 (___09____31424), .DIN2 (____09___31598),
       .Q (____09___31599));
  nor2s1 ______503597(.DIN1 (____0___28206), .DIN2 (___09_9__31455), .Q
       (____09___31597));
  and2s1 _____0_503598(.DIN1 (___0_9___31404), .DIN2 (____09___31595),
       .Q (____09___31596));
  nnd2s1 ______503599(.DIN1 (___0__9__31377), .DIN2 (_____9___32868),
       .Q (____09___31594));
  nor2s1 _____503600(.DIN1 (__9_____30026), .DIN2 (___09____31435), .Q
       (____090__31593));
  or2s1 _______503601(.DIN1 (____0____31591), .DIN2 (___0__0__31378),
       .Q (____0_9__31592));
  or2s1 _______503602(.DIN1 (____0____31589), .DIN2 (___0_____31355),
       .Q (____0____31590));
  nor2s1 _______503603(.DIN1 (__9_____30378), .DIN2 (___0_____31344),
       .Q (____0____31588));
  nor2s1 _____9_503604(.DIN1 (____0____31559), .DIN2 (___0_____31375),
       .Q (____0____31587));
  nnd2s1 _____9_503605(.DIN1 (___0_____31351), .DIN2 (__9_____30285),
       .Q (____0____31586));
  nor2s1 _____0_503606(.DIN1 (____0____31584), .DIN2 (___0_____31372),
       .Q (____0____31585));
  nor2s1 _____0_503607(.DIN1 (____000__31503), .DIN2 (___0_____31371),
       .Q (____0_0__31583));
  nnd2s1 ______503608(.DIN1 (___0_____31364), .DIN2 (____0____31581),
       .Q (____0_9__31582));
  nnd2s1 _______503609(.DIN1 (___0_____31354), .DIN2 (____0____31579),
       .Q (____0____31580));
  and2s1 _______503610(.DIN1 (___0_____31363), .DIN2 (____0____31577),
       .Q (____0____31578));
  nor2s1 _______503611(.DIN1 (__9_____30430), .DIN2 (___0_____31352),
       .Q (____0____31576));
  nor2s1 ______503612(.DIN1 (________29183), .DIN2 (___0__0__31358), .Q
       (____0____31575));
  nor2s1 _______503613(.DIN1 (___0_____30673), .DIN2 (___0_____31374),
       .Q (____0____31574));
  nnd2s1 _______503614(.DIN1 (___0__0__31348), .DIN2 (______0__32108),
       .Q (____0_0__31573));
  nor2s1 ______503615(.DIN1 (________25932), .DIN2 (___0__9__31357), .Q
       (____0_9__31572));
  nor2s1 _______503616(.DIN1 (_____9___38610), .DIN2 (______9__35888),
       .Q (____0____31571));
  nnd2s1 ______503617(.DIN1 (___0_____31356), .DIN2 (____9_9__32410),
       .Q (____0____31570));
  nor2s1 ______503618(.DIN1 (___0__9__31050), .DIN2 (___0_____31365),
       .Q (____0____31569));
  nnd2s1 _______503619(.DIN1 (___0_____31350), .DIN2 (_____9__28350),
       .Q (____0____31568));
  nnd2s1 _______503620(.DIN1 (___0__9__31367), .DIN2 (____0____31566),
       .Q (____0____31567));
  nor2s1 _______503621(.DIN1 (____00___33437), .DIN2 (___0_____31370),
       .Q (____0____31565));
  nnd2s1 _______503622(.DIN1 (___0_____31359), .DIN2 (___0__0__31339),
       .Q (____0____31564));
  nnd2s1 _______503623(.DIN1 (___0_____31373), .DIN2 (___00____30568),
       .Q (____0_0__31563));
  nnd2s1 _______503624(.DIN1 (___0_____31379), .DIN2 (_________33692),
       .Q (____0_9__31562));
  or2s1 _______503625(.DIN1 (_________32130), .DIN2 (___0_____31346),
       .Q (____0____31561));
  nor2s1 _____503626(.DIN1 (____0____31559), .DIN2 (___0_____31369), .Q
       (____0____31560));
  nnd2s1 _____9_503627(.DIN1 (___0_____31353), .DIN2 (___0_____31391),
       .Q (____0____31558));
  nnd2s1 _____9_503628(.DIN1 (___0_____31360), .DIN2 (____0____31556),
       .Q (____0____31557));
  nnd2s1 _____9_503629(.DIN1 (___0_____31380), .DIN2 (____0____31554),
       .Q (____0____31555));
  nnd2s1 _____0_503630(.DIN1 (___0_____31361), .DIN2 (________29541),
       .Q (____0_0__31553));
  nor2s1 _______503631(.DIN1 (____0_0__32518), .DIN2 (___0_____31396),
       .Q (_____9___31791));
  nor2s1 ______503632(.DIN1 (_________34207), .DIN2 (___090___31410),
       .Q (_________31734));
  nor2s1 _______503633(.DIN1 (____0_9__31552), .DIN2 (______9__35888),
       .Q (____9____36110));
  nor2s1 _______503634(.DIN1 (____0____31530), .DIN2 (_________31821),
       .Q (____0____31551));
  nnd2s1 _______503635(.DIN1 (___0_09__31319), .DIN2 (_________32266),
       .Q (____0____31550));
  nor2s1 _______503636(.DIN1 (__9_____30167), .DIN2 (______0__40953),
       .Q (____0____31549));
  nor2s1 _____0_503637(.DIN1 (____0____31547), .DIN2 (___0_____31325),
       .Q (____0____31548));
  nor2s1 _____503638(.DIN1 (____0____31545), .DIN2 (___0_____31298), .Q
       (____0____31546));
  and2s1 ______503639(.DIN1 (___0_0___31315), .DIN2 (______0__35853),
       .Q (____0____31544));
  nor2s1 _____0_503640(.DIN1 (____0_9__31542), .DIN2 (___0_____31328),
       .Q (____0_0__31543));
  nor2s1 ______503641(.DIN1 (____0_9__31552), .DIN2 (___0_0___31316),
       .Q (____0____31541));
  or2s1 _____0_503642(.DIN1 (___0_0___30743), .DIN2 (___0_____31264),
       .Q (____0____31540));
  nnd2s1 _____0_503643(.DIN1 (___0_____31288), .DIN2 (________27549),
       .Q (____0____31539));
  or2s1 _______503644(.DIN1
       (____________________________________________21833), .DIN2
       (_________34034), .Q (____0____31538));
  and2s1 _____0_503645(.DIN1 (___0_____31327), .DIN2 (________29452),
       .Q (____0____31537));
  nor2s1 _______503646(.DIN1 (_________33170), .DIN2 (___0_____31326),
       .Q (____0____31536));
  nnd2s1 _______503647(.DIN1 (_________34034), .DIN2
       (____________________________________________21833), .Q
       (____0____31535));
  nor2s1 _____0_503648(.DIN1 (___0990__31494), .DIN2 (___0_____31322),
       .Q (____0____31534));
  nor2s1 _______503649(.DIN1 (___0_0___31311), .DIN2 (___0_0___31318),
       .Q (____0_0__31533));
  nor2s1 _______503650(.DIN1 (___0909__40655), .DIN2 (_________31821),
       .Q (____0_9__31532));
  nor2s1 _______503651(.DIN1 (_________32145), .DIN2 (____0____31530),
       .Q (____0____31531));
  nnd2s1 _______503652(.DIN1 (____0____31530), .DIN2 (_________31938),
       .Q (____0____31529));
  nnd2s1 _____9_503653(.DIN1 (___0_00__31310), .DIN2 (____0____31527),
       .Q (____0____31528));
  nnd2s1 _____9_503654(.DIN1 (___0_____31285), .DIN2 (__9090), .Q
       (____0____31526));
  xor2s1 _______503655(.DIN1 (___0_____31136), .DIN2
       (______________22066), .Q (____0____31525));
  nor2s1 _____9_503656(.DIN1 (____0_0__31523), .DIN2 (___0_90__31300),
       .Q (____0____31524));
  and2s1 _______503657(.DIN1 (___0_____31321), .DIN2 (___0_____31366),
       .Q (____0_9__31522));
  nor2s1 ______503658(.DIN1 (___999__29637), .DIN2 (___0_9___31307), .Q
       (____0____31521));
  and2s1 _______503659(.DIN1 (____0____31519), .DIN2 (_________31715),
       .Q (____0____31520));
  nnd2s1 _______503660(.DIN1 (___0_9___31305), .DIN2 (____0____31517),
       .Q (____0____31518));
  nnd2s1 _______503661(.DIN1 (___0_9___31303), .DIN2 (_________32239),
       .Q (____0____31516));
  nor2s1 _______503662(.DIN1 (___09_9__31465), .DIN2 (___0_9___31308),
       .Q (____0____31515));
  nor2s1 _______503663(.DIN1 (___0_____30764), .DIN2 (___0_9___31306),
       .Q (____0____31514));
  nnd2s1 _______503664(.DIN1 (___0_9___31302), .DIN2 (___00____30575),
       .Q (____0_0__31513));
  nnd2s1 _____9_503665(.DIN1 (___0_99__31309), .DIN2 (__90_9), .Q
       (____009__31512));
  xor2s1 _______503666(.DIN1 (___0_9___31210), .DIN2 (_________38463),
       .Q (_________31617));
  nnd2s1 _______503667(.DIN1 (_________34034), .DIN2 (___0_0___40564),
       .Q (_________31624));
  nnd2s1 _______503668(.DIN1 (___0__0__31320), .DIN2 (____00___31511),
       .Q (_________31716));
  or2s1 _______503669(.DIN1 (___0_0___40564), .DIN2 (_________34034),
       .Q (_________31720));
  hi1s1 ____9__503670(.DIN (____9____33371), .Q (____9____33400));
  xor2s1 _______503671(.DIN1 (___0_9___31212), .DIN2 (___9_0___39077),
       .Q (_________31710));
  xor2s1 _______503672(.DIN1 (___0_____31171), .DIN2 (___9_____39784),
       .Q (______0__31718));
  dffacs1 ________________________________________________503673(.CLRB
       (reset), .CLK (clk), .DIN (___0__9__31329), .Q
       (______________________________________________21902));
  nor2s1 _______503674(.DIN1 (____00___31509), .DIN2 (___0_____31267),
       .Q (____00___31510));
  and2s1 ______503675(.DIN1 (___0_____31291), .DIN2 (____00___31507),
       .Q (____00___31508));
  nor2s1 _______503676(.DIN1 (____00___31505), .DIN2 (___0__9__31289),
       .Q (____00___31506));
  nor2s1 _______503677(.DIN1 (____000__31503), .DIN2 (___0_____31323),
       .Q (____00___31504));
  nor2s1 _______503678(.DIN1 (_________31866), .DIN2 (___0_____31287),
       .Q (___0999__31502));
  nnd2s1 _______503679(.DIN1 (___0_____31257), .DIN2 (_____0___32577),
       .Q (___099___31501));
  nor2s1 _______503680(.DIN1 (___0____27897), .DIN2 (___0_____31286),
       .Q (___099___31500));
  nnd2s1 _______503681(.DIN1 (___0_____31263), .DIN2 (__9_____30162),
       .Q (___099___31498));
  nor2s1 _______503682(.DIN1 (___099___31496), .DIN2 (_________40951),
       .Q (___099___31497));
  or2s1 _______503683(.DIN1 (___0990__31494), .DIN2 (___0__0__31281),
       .Q (___099___31495));
  nor2s1 _______503684(.DIN1 (___0_____30956), .DIN2 (___0_____31278),
       .Q (___09_9__31493));
  nor2s1 _______503685(.DIN1 (_________32344), .DIN2 (___0__0__31271),
       .Q (___09____31492));
  nor2s1 _______503686(.DIN1 (___99___25116), .DIN2 (___0_____31276),
       .Q (___09____31491));
  nor2s1 _______503687(.DIN1 (__909___29719), .DIN2 (___0_____31273),
       .Q (___09____31490));
  nor2s1 ______503688(.DIN1 (____00__29009), .DIN2 (___0__9__31270), .Q
       (___09____31489));
  and2s1 ______503689(.DIN1 (___0_____31269), .DIN2 (___09____31487),
       .Q (___09____31488));
  nor2s1 _______503690(.DIN1 (_________31809), .DIN2 (___0_____31275),
       .Q (___09_0__31486));
  nnd2s1 _______503691(.DIN1 (___0_____31272), .DIN2 (________25544),
       .Q (___09_9__31485));
  nor2s1 ______503692(.DIN1 (__9_____29835), .DIN2 (___0_____31292), .Q
       (___09____31484));
  nnd2s1 _______503693(.DIN1 (___0__0__31251), .DIN2 (____9___29188),
       .Q (___09____31483));
  nor2s1 ______503694(.DIN1 (_________41285), .DIN2 (___0_____31279),
       .Q (___09____31482));
  nor2s1 _____9_503695(.DIN1 (___09____31480), .DIN2 (___0__0__31261),
       .Q (___09____31481));
  nor2s1 _____9_503696(.DIN1 (___09____31478), .DIN2 (___0_____31265),
       .Q (___09____31479));
  nnd2s1 _____503697(.DIN1 (___0_____31283), .DIN2 (____0___29286), .Q
       (___09____31477));
  nnd2s1 _____0_503698(.DIN1 (___0_____31259), .DIN2 (____9___26491),
       .Q (___09_0__31476));
  nor2s1 _____0_503699(.DIN1 (_________32001), .DIN2 (___0_____31255),
       .Q (___09_9__31475));
  and2s1 _____0_503700(.DIN1 (___0_9___31304), .DIN2 (______9__31632),
       .Q (___09____31474));
  and2s1 _____0_503701(.DIN1 (___0_____31256), .DIN2 (___09____31472),
       .Q (___09____31473));
  nor2s1 _______503702(.DIN1 (___0_____31336), .DIN2 (___0_____31254),
       .Q (___09____31471));
  and2s1 _______503703(.DIN1 (___0_____31284), .DIN2 (___09____31469),
       .Q (___09____31470));
  nor2s1 _______503704(.DIN1 (___09____31467), .DIN2 (___0__9__31250),
       .Q (___09____31468));
  nor2s1 _______503705(.DIN1 (___09_9__31465), .DIN2 (___0_____31245),
       .Q (___09_0__31466));
  nnd2s1 _______503706(.DIN1 (___0_____31249), .DIN2 (___9____28696),
       .Q (___09____31464));
  or2s1 _______503707(.DIN1 (__9_____29881), .DIN2 (___0_____31294), .Q
       (___09____31463));
  nnd2s1 _______503708(.DIN1 (___0_____31341), .DIN2 (___09____31461),
       .Q (___09____31462));
  nor2s1 _______503709(.DIN1 (___00____30608), .DIN2 (___0_____31343),
       .Q (___09____31460));
  nnd2s1 _______503710(.DIN1 (___0_____31338), .DIN2 (___9____29575),
       .Q (___09____31459));
  nnd2s1 ______503711(.DIN1 (___0_____31246), .DIN2 (__9_____30163), .Q
       (___09____31458));
  nor2s1 _______503712(.DIN1 (___0900), .DIN2 (___0_____31152), .Q
       (___09____31457));
  xor2s1 _____0_503713(.DIN1 (___0_0___31314), .DIN2 (_____9___36360),
       .Q (___09_0__31456));
  nnd2s1 ______503714(.DIN1 (___0_____31224), .DIN2 (______0__41032),
       .Q (___09_9__31455));
  nnd2s1 ____09_503715(.DIN1 (___09____31449), .DIN2 (___09____31453),
       .Q (___09____31454));
  or2s1 ______503716(.DIN1 (___09____31451), .DIN2 (___0_____31142), .Q
       (___09____31452));
  nnd2s1 ______503717(.DIN1 (___09____31449), .DIN2 (________29487), .Q
       (___09____31450));
  nor2s1 ______503718(.DIN1 (________27681), .DIN2 (___0__9__31157), .Q
       (___09____31448));
  or2s1 _______503719(.DIN1 (___09_9__31446), .DIN2 (___0_____31144),
       .Q (___09_0__31447));
  nor2s1 _______503720(.DIN1 (___0_____30821), .DIN2 (___0_9___31213),
       .Q (___09____31445));
  nnd2s1 ______503721(.DIN1 (___0_0___31217), .DIN2 (___09____31443),
       .Q (___09____31444));
  nor2s1 _______503722(.DIN1 (____0____31547), .DIN2 (___0_99__31215),
       .Q (___09____31442));
  nor2s1 ______503723(.DIN1 (___0_0___31317), .DIN2 (___0_____31296),
       .Q (___09____31441));
  or2s1 ______503724(.DIN1 (_____0__28591), .DIN2 (___0__9__31177), .Q
       (___09____31440));
  and2s1 _______503725(.DIN1 (___0_____31159), .DIN2 (___09____31438),
       .Q (___09____31439));
  or2s1 _______503726(.DIN1 (_____0___34102), .DIN2 (___0_9___31207),
       .Q (___09_0__31437));
  nor2s1 _______503727(.DIN1 (__9__0__30394), .DIN2 (___0_____31145),
       .Q (___09_9__31436));
  nnd2s1 _______503728(.DIN1 (___0_____31146), .DIN2 (___0_____30864),
       .Q (___09____31435));
  nor2s1 _______503729(.DIN1 (________28231), .DIN2 (___0_____31201),
       .Q (___09____31434));
  nor2s1 _______503730(.DIN1 (___0_9__28795), .DIN2 (___0_____31155),
       .Q (___09____31433));
  nor2s1 _______503731(.DIN1 (_________32311), .DIN2 (___0_9___31209),
       .Q (___09____31432));
  nnd2s1 _______503732(.DIN1 (___0_____31203), .DIN2 (________25846),
       .Q (___09____31431));
  nor2s1 ______503733(.DIN1 (___09____31429), .DIN2 (___0__9__31196),
       .Q (___09____31430));
  or2s1 ______503734(.DIN1 (__9_____30105), .DIN2 (___0_____31161), .Q
       (___09____31428));
  and2s1 _______503735(.DIN1 (___0_____31193), .DIN2 (___09_9__31426),
       .Q (___09_0__31427));
  nor2s1 _____503736(.DIN1 (________26632), .DIN2 (___0_____31189), .Q
       (___09____31425));
  nor2s1 _____9_503737(.DIN1 (____0____32521), .DIN2 (___0__0__31188),
       .Q (___09____31424));
  nor2s1 _____9_503738(.DIN1 (___9____28667), .DIN2 (___0_0___31219),
       .Q (___09____31423));
  and2s1 _____503739(.DIN1 (___0_____31184), .DIN2 (___0__9__30851), .Q
       (___09____31422));
  nnd2s1 _____503740(.DIN1 (___0_____31199), .DIN2 (________28230), .Q
       (___09____31421));
  nor2s1 _____0_503741(.DIN1 (__9_00__29993), .DIN2 (___0_____31183),
       .Q (___09____31420));
  nnd2s1 _____0_503742(.DIN1 (___0_____31181), .DIN2 (__90____29649),
       .Q (___09____31419));
  and2s1 _____0_503743(.DIN1 (___0_____31150), .DIN2 (__9_____30189),
       .Q (___09____31418));
  nnd2s1 _______503744(.DIN1 (___0_____31179), .DIN2 (__9_9___30451),
       .Q (___09_0__31417));
  nnd2s1 _______503745(.DIN1 (___0__0__31178), .DIN2 (___090___31415),
       .Q (___0909__31416));
  nor2s1 _______503746(.DIN1 (___090___31413), .DIN2 (___0__0__31158),
       .Q (___090___31414));
  nnd2s1 _______503747(.DIN1 (___0_____31192), .DIN2 (___0_____30870),
       .Q (___090___31412));
  nor2s1 _______503748(.DIN1 (_________31673), .DIN2 (___0_____31172),
       .Q (___090___31411));
  nnd2s1 _______503749(.DIN1 (___0__9__31187), .DIN2 (____9____33362),
       .Q (___090___31410));
  and2s1 _______503750(.DIN1 (___0_____31169), .DIN2 (____09___31595),
       .Q (___090___31409));
  nor2s1 ______503751(.DIN1 (___0900), .DIN2 (___0_____31166), .Q
       (___090___31408));
  nor2s1 _______503752(.DIN1 (__99____30496), .DIN2 (___0_90__31206),
       .Q (___0_99__31407));
  nor2s1 _______503753(.DIN1 (___0_9___31405), .DIN2 (___0_____31133),
       .Q (___0_9___31406));
  nnd2s1 _______503754(.DIN1 (___0_09__31221), .DIN2 (___0_____30893),
       .Q (_________31639));
  xor2s1 _______503755(.DIN1 (_____0___36368), .DIN2 (______9__35584),
       .Q (_____0___36370));
  nnd2s1 _______503756(.DIN1 (___0_____31200), .DIN2 (___0_____31134),
       .Q (_________31616));
  xor2s1 ____0__503757(.DIN1 (___0_____31039), .DIN2 (_________33321),
       .Q (____9____33371));
  hi1s1 _______503758(.DIN (_________31821), .Q (______9__35888));
  and2s1 _____0_503759(.DIN1 (___0_____31225), .DIN2 (___0_9___31403),
       .Q (___0_9___31404));
  nor2s1 _______503760(.DIN1 (___0_9___31401), .DIN2 (___0_____31195),
       .Q (___0_9___31402));
  and2s1 _______503761(.DIN1 (___0_9___31399), .DIN2 (_________31715),
       .Q (___0_9___31400));
  nnd2s1 _______503762(.DIN1 (___0_____31176), .DIN2 (_____0___41313),
       .Q (___0_90__31398));
  nor2s1 _______503763(.DIN1 (_____9__29174), .DIN2 (___0_____31170),
       .Q (___0__9__31397));
  nnd2s1 ______503764(.DIN1 (___0__0__31148), .DIN2 (____9_0__32391),
       .Q (___0_____31396));
  nnd2s1 _______503765(.DIN1 (___0_____31174), .DIN2 (___0_____31394),
       .Q (___0_____31395));
  or2s1 _______503766(.DIN1 (_________31906), .DIN2 (___0_____31202),
       .Q (___0_____31393));
  nnd2s1 _____9_503767(.DIN1 (___0_____31163), .DIN2 (___0_____31391),
       .Q (___0_____31392));
  and2s1 _____9_503768(.DIN1 (___0_____31141), .DIN2 (____0____31554),
       .Q (___0_____31390));
  nor2s1 _____9_503769(.DIN1 (___0__0__31197), .DIN2 (________26249),
       .Q (___0_____31389));
  nor2s1 _____503770(.DIN1 (___00_0__30612), .DIN2 (___0_____31143), .Q
       (___0__0__31388));
  nor2s1 _____0_503771(.DIN1 (__9_____30260), .DIN2 (___0__9__31205),
       .Q (___0__9__31387));
  nnd2s1 _____0_503772(.DIN1 (___0_____31149), .DIN2 (___0_____31385),
       .Q (___0_____31386));
  and2s1 _______503773(.DIN1 (___0_____31165), .DIN2 (____9____33353),
       .Q (___0_____31384));
  nor2s1 _______503774(.DIN1 (________29307), .DIN2 (___0_9___31208),
       .Q (___0_____31383));
  nor2s1 _______503775(.DIN1 (___0_____31381), .DIN2 (___0_____31139),
       .Q (___0_____31382));
  nor2s1 _____0_503776(.DIN1 (___0_____31140), .DIN2 (___0_9___31114),
       .Q (___0_____31380));
  nor2s1 _______503777(.DIN1 (_________31906), .DIN2 (___0_____31131),
       .Q (___0_____31379));
  nnd2s1 _______503778(.DIN1 (___0__9__31231), .DIN2 (__9_9___29986),
       .Q (___0__0__31378));
  and2s1 ______503779(.DIN1 (___0__0__31128), .DIN2 (___0_____31376),
       .Q (___0__9__31377));
  nnd2s1 ______503780(.DIN1 (___0__0__31368), .DIN2 (___0__0__30662),
       .Q (___0_____31375));
  nnd2s1 _______503781(.DIN1 (___0_99__31117), .DIN2 (________29242),
       .Q (___0_____31374));
  nor2s1 _______503782(.DIN1 (__9_____29914), .DIN2 (___0_9___31115),
       .Q (___0_____31373));
  or2s1 _____9_503783(.DIN1 (__9_____29781), .DIN2 (___0_9___31113), .Q
       (___0_____31372));
  nnd2s1 _____9_503784(.DIN1 (___0_9___31112), .DIN2 (__9_____29911),
       .Q (___0_____31371));
  nnd2s1 _____9_503785(.DIN1 (___0_9___31110), .DIN2 (______9__33575),
       .Q (___0_____31370));
  nnd2s1 _____9_503786(.DIN1 (___0__0__31368), .DIN2 (_________40965),
       .Q (___0_____31369));
  and2s1 _____503787(.DIN1 (___0_0___31122), .DIN2 (___0_____31366), .Q
       (___0__9__31367));
  nnd2s1 _____0_503788(.DIN1 (___0_9___31109), .DIN2 (____09__28022),
       .Q (___0_____31365));
  nor2s1 _____0_503789(.DIN1 (_________41126), .DIN2 (___0_00__31118),
       .Q (___0_____31364));
  and2s1 _____503790(.DIN1 (___0_____31185), .DIN2 (___0_____31362), .Q
       (___0_____31363));
  nor2s1 _______503791(.DIN1 (________29239), .DIN2 (___0_0___31218),
       .Q (___0_____31361));
  nor2s1 _______503792(.DIN1 (__9_0___30373), .DIN2 (___0_____31349),
       .Q (___0_____31360));
  nnd2s1 _______503793(.DIN1 (___0__9__31240), .DIN2 (__9_____29735),
       .Q (___0_____31359));
  nnd2s1 _______503794(.DIN1 (___0_0___31126), .DIN2 (________26735),
       .Q (___0__0__31358));
  nnd2s1 _______503795(.DIN1 (___0_0___31120), .DIN2 (__9__9__30319),
       .Q (___0__9__31357));
  nor2s1 _______503796(.DIN1 (_________32130), .DIN2 (___0_____31235),
       .Q (___0_____31356));
  nnd2s1 _______503797(.DIN1 (___0_____31243), .DIN2 (_________32811),
       .Q (___0_____31355));
  nor2s1 _______503798(.DIN1 (__9__9__30337), .DIN2 (___0_____31233),
       .Q (___0_____31354));
  nor2s1 _______503799(.DIN1 (___0_0___31031), .DIN2 (___0_____31130),
       .Q (___0_____31353));
  nnd2s1 _______503800(.DIN1 (___0_____31234), .DIN2 (__9_99__29895),
       .Q (___0_____31352));
  nor2s1 ______503801(.DIN1 (________27181), .DIN2 (___0_____31226), .Q
       (___0_____31351));
  nor2s1 ______503802(.DIN1 (__9__9__29925), .DIN2 (___0_____31349), .Q
       (___0_____31350));
  nor2s1 _______503803(.DIN1 (___0__9__31347), .DIN2 (___0_____31228),
       .Q (___0__0__31348));
  or2s1 _____9_503804(.DIN1 (___0_____31345), .DIN2 (___0_____31238),
       .Q (___0_____31346));
  nor2s1 _____0_503805(.DIN1 (___0900), .DIN2 (___0_____31236), .Q
       (___0_____31344));
  nnd2s1 ______503806(.DIN1 (___0__9__31137), .DIN2 (______0__32196),
       .Q (___099___31499));
  and2s1 ______503807(.DIN1 (___0__0__31138), .DIN2 (_________32114),
       .Q (_________31646));
  nnd2s1 ______503808(.DIN1 (___0__0__31051), .DIN2 (______0__41032),
       .Q (___0_____31343));
  nnd2s1 _______503809(.DIN1 (___0_____31056), .DIN2 (__99_0__30489),
       .Q (___0_____31342));
  nor2s1 _______503810(.DIN1 (__9_____30312), .DIN2 (___0_____31055),
       .Q (___0_____31341));
  nnd2s1 _______503811(.DIN1 (___0_____31054), .DIN2 (inData[12]), .Q
       (___0_____31340));
  nnd2s1 _______503812(.DIN1 (___0_____31048), .DIN2 (________26723),
       .Q (___0__0__31339));
  nor2s1 ______503813(.DIN1 (________27183), .DIN2 (___0_____31044), .Q
       (___0_____31338));
  nor2s1 ____90_503814(.DIN1 (___0_____31336), .DIN2 (___0_9___31020),
       .Q (___0_____31337));
  xor2s1 _______503815(.DIN1 (______0__36056), .DIN2 (_________36928),
       .Q (___0_____31335));
  xor2s1 _______503816(.DIN1 (___0_____30885), .DIN2 (_________22046),
       .Q (___0_____31334));
  or2s1 _______503817(.DIN1 (_____9__26546), .DIN2 (_________32806), .Q
       (___0_____31333));
  and2s1 _______503818(.DIN1 (_____0___36368), .DIN2 (___0__0__31330),
       .Q (___0_____31332));
  nor2s1 ______503819(.DIN1 (___0__0__31330), .DIN2 (_____0___36368),
       .Q (___0_____31331));
  nnd2s1 ______503820(.DIN1 (___0_0___31024), .DIN2 (________25845), .Q
       (___0__9__31329));
  or2s1 _______503821(.DIN1 (_________32602), .DIN2 (___0_0___31029),
       .Q (___0_____31328));
  nor2s1 _______503822(.DIN1 (________29450), .DIN2 (___0_0___31025),
       .Q (___0_____31327));
  nnd2s1 ______503823(.DIN1 (___0_0___31028), .DIN2 (_____0__25938), .Q
       (___0_____31326));
  or2s1 _______503824(.DIN1 (___0_____31324), .DIN2 (___0_09__31032),
       .Q (___0_____31325));
  nnd2s1 _____9_503825(.DIN1 (___0_____31036), .DIN2 (________28066),
       .Q (___0_____31323));
  nnd2s1 _____9_503826(.DIN1 (___0_0___31027), .DIN2 (____9___28290),
       .Q (___0_____31322));
  nor2s1 _____503827(.DIN1 (_____0__28502), .DIN2 (___0_0___31026), .Q
       (___0_____31321));
  nor2s1 _______503828(.DIN1 (_________31827), .DIN2 (___0_9___31021),
       .Q (___0__0__31320));
  or2s1 ______503829(.DIN1 (_________32241), .DIN2 (_________40957), .Q
       (___0_09__31319));
  nor2s1 _____0_503830(.DIN1 (___0_0___31312), .DIN2 (___0_0___31317),
       .Q (___0_0___31318));
  nnd2s1 ______503831(.DIN1 (___0_99__31022), .DIN2 (_____09__35744),
       .Q (___0_0___31316));
  nor2s1 _______503832(.DIN1 (_____09__35744), .DIN2 (___0_0___31314),
       .Q (___0_0___31315));
  nnd2s1 _______503833(.DIN1 (___0_0___31312), .DIN2 (___0_0___31311),
       .Q (___0_0___31313));
  nor2s1 _______503834(.DIN1 (_________33551), .DIN2 (___0_____31001),
       .Q (___0_00__31310));
  and2s1 _______503835(.DIN1 (_________40959), .DIN2 (________27583),
       .Q (___0_99__31309));
  nnd2s1 _______503836(.DIN1 (___0_9___31014), .DIN2 (___0__9__30984),
       .Q (___0_9___31308));
  nnd2s1 ______503837(.DIN1 (___0_____31091), .DIN2 (__9_____29748), .Q
       (___0_9___31307));
  nnd2s1 ______503838(.DIN1 (___0_____31009), .DIN2 (________27180), .Q
       (___0_9___31306));
  nor2s1 ______503839(.DIN1 (___0_____31129), .DIN2 (___0_____31068),
       .Q (___0_9___31305));
  nor2s1 _______503840(.DIN1 (________25753), .DIN2 (___0_____31097),
       .Q (___0_9___31304));
  nor2s1 _______503841(.DIN1 (_________32903), .DIN2 (___0_____31083),
       .Q (___0_9___31303));
  and2s1 ______503842(.DIN1 (___0_9___31019), .DIN2 (___0_9___31301),
       .Q (___0_9___31302));
  nnd2s1 _______503843(.DIN1 (___0__9__31089), .DIN2 (___0__9__31299),
       .Q (___0_90__31300));
  nnd2s1 _______503844(.DIN1 (___0__0__31099), .DIN2 (___0_____31297),
       .Q (___0_____31298));
  hi1s1 _______503845(.DIN (___0_____31296), .Q (____0____31530));
  xor2s1 _______503846(.DIN1 (_________32145), .DIN2 (_________41264),
       .Q (_________31821));
  hi1s1 _______503847(.DIN (___0_____31295), .Q (_________34034));
  nnd2s1 _______503848(.DIN1 (___0_____31057), .DIN2 (___0_99__30832),
       .Q (___0_____31294));
  nnd2s1 _____0_503849(.DIN1 (___0_____31043), .DIN2 (__9_0___30277),
       .Q (___0_____31293));
  nnd2s1 _______503850(.DIN1 (___0_____31106), .DIN2 (________28528),
       .Q (___0_____31292));
  and2s1 _______503851(.DIN1 (___0_____31105), .DIN2 (___0__0__31290),
       .Q (___0_____31291));
  nnd2s1 _______503852(.DIN1 (___0_____31103), .DIN2 (___00____30606),
       .Q (___0__9__31289));
  nor2s1 _____503853(.DIN1 (________28631), .DIN2 (___0__0__31042), .Q
       (___0_____31288));
  nnd2s1 _______503854(.DIN1 (___0_____31002), .DIN2 (___0_____31385),
       .Q (___0_____31287));
  nnd2s1 _______503855(.DIN1 (___0_____31004), .DIN2 (___09____31469),
       .Q (___0_____31286));
  nor2s1 ______503856(.DIN1 (________28964), .DIN2 (___0_____31000), .Q
       (___0_____31285));
  nor2s1 _______503857(.DIN1 (_________41158), .DIN2 (___0_____31005),
       .Q (___0_____31284));
  nor2s1 _______503858(.DIN1 (________29081), .DIN2 (___0_____31082),
       .Q (___0_____31283));
  nnd2s1 _______503859(.DIN1 (___0_____31081), .DIN2 (___0__9__31280),
       .Q (___0__0__31281));
  nnd2s1 ______503860(.DIN1 (___0__9__31098), .DIN2 (__99____30533), .Q
       (___0_____31279));
  or2s1 _______503861(.DIN1 (___0_____31277), .DIN2 (___0_____31104),
       .Q (___0_____31278));
  nor2s1 _______503862(.DIN1 (__9_____30432), .DIN2 (___0_____31007),
       .Q (___0_____31276));
  nor2s1 ______503863(.DIN1 (___0_____31274), .DIN2 (___0_____31095),
       .Q (___0_____31275));
  nnd2s1 _______503864(.DIN1 (___0__9__31107), .DIN2 (___0_____30810),
       .Q (___0_____31273));
  nnd2s1 _______503865(.DIN1 (___0_____31074), .DIN2 (_________31731),
       .Q (___0_____31272));
  nnd2s1 _______503866(.DIN1 (___0_____31093), .DIN2 (________29121),
       .Q (___0__0__31271));
  nnd2s1 _______503867(.DIN1 (___0__0__31090), .DIN2 (___9____27766),
       .Q (___0__9__31270));
  nor2s1 _______503868(.DIN1 (___0_____31268), .DIN2 (___0_____31085),
       .Q (___0_____31269));
  nnd2s1 _______503869(.DIN1 (___0_____31069), .DIN2 (___0_____31266),
       .Q (___0_____31267));
  nnd2s1 _____9_503870(.DIN1 (___0_____31079), .DIN2 (___009___30634),
       .Q (___0_____31265));
  nnd2s1 _____9_503871(.DIN1 (_________40955), .DIN2 (_____0__29227),
       .Q (___0_____31264));
  nor2s1 _____9_503872(.DIN1 (___0_____31262), .DIN2 (___0__9__31070),
       .Q (___0_____31263));
  nnd2s1 _____9_503873(.DIN1 (___0_____31077), .DIN2 (___0__9__31260),
       .Q (___0__0__31261));
  and2s1 _____503874(.DIN1 (___0__0__31071), .DIN2 (___0_____31258), .Q
       (___0_____31259));
  nor2s1 _____503875(.DIN1 (____99__28923), .DIN2 (___0_____31087), .Q
       (___0_____31257));
  nor2s1 _____0_503876(.DIN1 (_________33002), .DIN2 (___0_____31101),
       .Q (___0_____31256));
  and2s1 _____0_503877(.DIN1 (___0_9___31016), .DIN2 (___0_9___31214),
       .Q (___0_____31255));
  nor2s1 _____0_503878(.DIN1 (_________32058), .DIN2 (___0_____31072),
       .Q (___0_____31254));
  nnd2s1 _____0_503879(.DIN1 (___0_____31067), .DIN2 (_________32266),
       .Q (___0_____31253));
  nor2s1 _____0_503880(.DIN1 (____9____33386), .DIN2 (___0__9__31041),
       .Q (___0_____31252));
  nor2s1 ______503881(.DIN1 (___0__9__30908), .DIN2 (___0_90__31013),
       .Q (___0__0__31251));
  or2s1 _______503882(.DIN1 (___09____31480), .DIN2 (___0_____31065),
       .Q (___0__9__31250));
  and2s1 ______503883(.DIN1 (___0_____31058), .DIN2 (_____9__25937), .Q
       (___0_____31249));
  nor2s1 _______503884(.DIN1 (___0_____31247), .DIN2 (___0_____31102),
       .Q (___0_____31248));
  nor2s1 _______503885(.DIN1 (__9_0___30000), .DIN2 (___0_____31062),
       .Q (___0_____31246));
  nnd2s1 _______503886(.DIN1 (___0_____31059), .DIN2 (____9___29190),
       .Q (___0_____31245));
  nnd2s1 _______503887(.DIN1 (___0_9___31017), .DIN2 (_________31781),
       .Q (____0____31519));
  nor2s1 _______503888(.DIN1 (____0____32539), .DIN2 (___0_____30992),
       .Q (___0_____31244));
  nor2s1 ______503889(.DIN1 (___0_____31242), .DIN2 (___0_____30897),
       .Q (___0_____31243));
  nor2s1 _______503890(.DIN1 (__9__0__30150), .DIN2 (___0_____30942),
       .Q (___0__0__31241));
  nnd2s1 _______503891(.DIN1 (___0_0___30932), .DIN2 (___9____26916),
       .Q (___0__9__31240));
  nor2s1 _______503892(.DIN1 (___0_____30950), .DIN2 (__999___30541),
       .Q (___0_____31239));
  nnd2s1 _______503893(.DIN1 (___0_9___30924), .DIN2 (___0_____31237),
       .Q (___0_____31238));
  nor2s1 _______503894(.DIN1 (__9_0___29726), .DIN2 (___0__0__30935),
       .Q (___0_____31236));
  or2s1 _______503895(.DIN1 (___0_____31268), .DIN2 (___0_0___30928),
       .Q (___0_____31235));
  and2s1 _______503896(.DIN1 (___0_____30906), .DIN2 (___0_____31006),
       .Q (___0_____31234));
  or2s1 ____90_503897(.DIN1 (_________41156), .DIN2 (___0_____30936),
       .Q (___0_____31233));
  nnd2s1 ____90_503898(.DIN1 (___0_____30904), .DIN2 (____9_9__32410),
       .Q (___0__0__31232));
  nor2s1 ____90_503899(.DIN1 (________28223), .DIN2 (___0__9__30918),
       .Q (___0__9__31231));
  nor2s1 ____90_503900(.DIN1 (___0_____31229), .DIN2 (___0_____30995),
       .Q (___0_____31230));
  nnd2s1 ____9__503901(.DIN1 (___0__0__30994), .DIN2 (________29511),
       .Q (___0_____31228));
  nor2s1 ____9__503902(.DIN1 (____9____33386), .DIN2 (___0_____30907),
       .Q (___0_____31227));
  or2s1 ____9_503903(.DIN1 (____000__31503), .DIN2 (___0__0__30909), .Q
       (___0_____31226));
  nor2s1 ____0__503904(.DIN1 (___0_____31223), .DIN2 (___0_____30895),
       .Q (___0_____31225));
  nor2s1 ____0__503905(.DIN1 (___0_____31223), .DIN2 (___0_____30896),
       .Q (___0_____31224));
  dffacs1 _______________503906(.CLRB (reset), .CLK (clk), .DIN
       (_________31938), .Q (outData[5]));
  nnd2s1 _______503907(.DIN1 (___0_____30848), .DIN2 (_________32266),
       .Q (___0__0__31222));
  or2s1 _______503908(.DIN1 (_________32024), .DIN2 (___0_____30892),
       .Q (___0_09__31221));
  nnd2s1 _______503909(.DIN1 (___0_____31153), .DIN2 (___00___26956),
       .Q (___0_0___31219));
  nor2s1 _______503910(.DIN1 (___0_____30961), .DIN2 (___0_9___31116),
       .Q (___0_0___31218));
  and2s1 _______503911(.DIN1 (___0__0__30881), .DIN2 (___0_00__31216),
       .Q (___0_0___31217));
  nnd2s1 _______503912(.DIN1 (___0_____30883), .DIN2 (___0_9___31214),
       .Q (___0_99__31215));
  nnd2s1 _______503913(.DIN1 (___0_____30877), .DIN2 (___0_____30912),
       .Q (___0_9___31213));
  nor2s1 _______503914(.DIN1 (___0_____30716), .DIN2 (___0_9___31211),
       .Q (___0_9___31212));
  or2s1 _______503915(.DIN1 (___0_____30878), .DIN2 (______0__36056),
       .Q (___0_9___31210));
  nnd2s1 _______503916(.DIN1 (___0_____30969), .DIN2 (___0_____31096),
       .Q (___0_9___31209));
  nnd2s1 _______503917(.DIN1 (___0_____30868), .DIN2 (___0____28817),
       .Q (___0_9___31208));
  nnd2s1 _______503918(.DIN1 (___0_____30867), .DIN2 (___09_9__31426),
       .Q (___0_9___31207));
  nnd2s1 _______503919(.DIN1 (___0_____30865), .DIN2 (____99__29552),
       .Q (___0_90__31206));
  nnd2s1 _______503920(.DIN1 (___0__9__30871), .DIN2 (___0_____31204),
       .Q (___0__9__31205));
  nnd2s1 _______503921(.DIN1 (___0_____30859), .DIN2 (inData[18]), .Q
       (___0_____31203));
  nnd2s1 _______503922(.DIN1 (___0__0__30862), .DIN2 (___0_____30888),
       .Q (___0_____31202));
  nor2s1 ______503923(.DIN1 (_________31809), .DIN2 (___0__9__30861),
       .Q (___0_____31201));
  nnd2s1 _______503924(.DIN1 (___0_____31135), .DIN2
       (______________22066), .Q (___0_____31200));
  nor2s1 _______503925(.DIN1 (___0_____31198), .DIN2 (___0_____30860),
       .Q (___0_____31199));
  nor2s1 _______503926(.DIN1 (__99____30501), .DIN2 (___0_____30857),
       .Q (___0__0__31197));
  or2s1 _______503927(.DIN1 (_____9___31789), .DIN2 (___0_____30876),
       .Q (___0__9__31196));
  or2s1 _______503928(.DIN1 (___0_____31194), .DIN2 (___0_____30987),
       .Q (___0_____31195));
  nor2s1 _______503929(.DIN1 (____9____34365), .DIN2 (___0__9__30974),
       .Q (___0_____31193));
  nor2s1 ______503930(.DIN1 (___0_____31191), .DIN2 (___0_____30988),
       .Q (___0_____31192));
  nor2s1 _______503931(.DIN1 (___0____25136), .DIN2 (___0_____30855),
       .Q (___0_____31190));
  or2s1 _______503932(.DIN1 (________28310), .DIN2 (___0__0__30852), .Q
       (___0_____31189));
  nnd2s1 _______503933(.DIN1 (___0_____30850), .DIN2 (__9__0__29966),
       .Q (___0__0__31188));
  nor2s1 ______503934(.DIN1 (____0____33496), .DIN2 (___0_____30879),
       .Q (___0__9__31187));
  xor2s1 _______503935(.DIN1 (___0_9___30831), .DIN2 (______9__37429),
       .Q (___0_____31295));
  xor2s1 _______503936(.DIN1 (___0_____30718), .DIN2 (___9__9__39731),
       .Q (___09____31449));
  nor2s1 ____9__503937(.DIN1 (___0_____31186), .DIN2 (___0_____30916),
       .Q (___0__0__31368));
  nnd2s1 ____9__503938(.DIN1 (___0__9__30993), .DIN2 (________28982),
       .Q (___0_____31349));
  nnd2s1 ______503939(.DIN1 (___0_____30999), .DIN2 (___0_0___31311),
       .Q (___0_____31296));
  dffacs1 ________________0_503940(.CLRB (reset), .CLK (clk), .DIN
       (___0_____30946), .QN
       (______________________________________________________________________________________0));
  dffacs1 ________________9_(.CLRB (reset), .CLK (clk), .DIN
       (___0_____30947), .QN (___________9___22071));
  and2s1 _______503941(.DIN1 (___0_0___30931), .DIN2 (___0_____31204),
       .Q (___0_____31185));
  nor2s1 ______503942(.DIN1 (_____0__26804), .DIN2 (___0_____30843), .Q
       (___0_____31184));
  nnd2s1 _____9_503943(.DIN1 (___0_____30874), .DIN2 (___0_____31182),
       .Q (___0_____31183));
  nor2s1 _____9_503944(.DIN1 (____9___29544), .DIN2 (___0_____30875),
       .Q (___0_____31181));
  nnd2s1 _____0_503945(.DIN1 (___0_____30998), .DIN2 (________26299),
       .Q (___0_____31180));
  nor2s1 _____0_503946(.DIN1 (___0_____30981), .DIN2 (___00_0__30603),
       .Q (___0_____31179));
  nor2s1 ______503947(.DIN1 (___00____30587), .DIN2 (___0_9___30920),
       .Q (___0__0__31178));
  nnd2s1 _______503948(.DIN1 (___0_____30869), .DIN2 (__9_____30250),
       .Q (___0__9__31177));
  and2s1 _______503949(.DIN1 (___0_____30989), .DIN2 (___0_____31175),
       .Q (___0_____31176));
  and2s1 _______503950(.DIN1 (___0_____30996), .DIN2 (___0_____31173),
       .Q (___0_____31174));
  or2s1 ______503951(.DIN1 (___0_0___31125), .DIN2 (___0_____30957), .Q
       (___0_____31172));
  nor2s1 _______503952(.DIN1 (____9___28466), .DIN2 (___0__0__30955),
       .Q (___0_____31171));
  nnd2s1 _______503953(.DIN1 (___0__9__30964), .DIN2 (________28189),
       .Q (___0_____31170));
  and2s1 _______503954(.DIN1 (___0_____30980), .DIN2 (___0__0__31168),
       .Q (___0_____31169));
  nor2s1 ______503955(.DIN1 (__999_), .DIN2 (___0_____30973), .Q
       (___0__9__31167));
  nor2s1 _______503956(.DIN1 (________26303), .DIN2 (___0__0__30985),
       .Q (___0_____31166));
  and2s1 _______503957(.DIN1 (___0_____30847), .DIN2 (___0_____31164),
       .Q (___0_____31165));
  and2s1 ______503958(.DIN1 (___0_____30963), .DIN2 (___0_____31162),
       .Q (___0_____31163));
  nnd2s1 _______503959(.DIN1 (___0_____30972), .DIN2 (__9_90__29985),
       .Q (___0_____31161));
  nnd2s1 _______503960(.DIN1 (___0_____30983), .DIN2 (____9_9__32410),
       .Q (___0_____31160));
  nor2s1 _______503961(.DIN1 (________27962), .DIN2 (___0_____30982),
       .Q (___0_____31159));
  nnd2s1 _______503962(.DIN1 (___0_____30960), .DIN2 (__9_99__29992),
       .Q (___0__0__31158));
  nnd2s1 _______503963(.DIN1 (___0_____30849), .DIN2 (___0_____31156),
       .Q (___0__9__31157));
  nnd2s1 ______503964(.DIN1 (___0_____30976), .DIN2 (___0__0__30711),
       .Q (___0_____31155));
  or2s1 _______503965(.DIN1 (_________32159), .DIN2 (___0_____31153),
       .Q (___0_____31154));
  and2s1 _______503966(.DIN1 (___0_____30959), .DIN2 (___0_____31151),
       .Q (___0_____31152));
  nor2s1 _______503967(.DIN1 (___9____29573), .DIN2 (___0_____30845),
       .Q (___0_____31150));
  nor2s1 _______503968(.DIN1 (_____9___33059), .DIN2 (___0_____30990),
       .Q (___0_____31149));
  nor2s1 _______503969(.DIN1 (___0__9__31147), .DIN2 (___0_____30978),
       .Q (___0__0__31148));
  nnd2s1 _______503970(.DIN1 (___0__0__30965), .DIN2 (__9_____30255),
       .Q (___0_____31146));
  nnd2s1 _____503971(.DIN1 (___0_____30966), .DIN2 (___0__0__31003), .Q
       (___0_____31145));
  or2s1 _____9_503972(.DIN1 (___0_____31345), .DIN2 (___0__9__30954),
       .Q (___0_____31144));
  nnd2s1 _____9_503973(.DIN1 (___0_____30853), .DIN2 (___0_____30805),
       .Q (___0_____31143));
  nnd2s1 _____9_503974(.DIN1 (___0_____30953), .DIN2 (___0_00__31216),
       .Q (___0_____31142));
  nor2s1 _____0_503975(.DIN1 (___0_____31140), .DIN2 (___0_____30846),
       .Q (___0_____31141));
  or2s1 _____503976(.DIN1 (___0_____31277), .DIN2 (___0__0__30975), .Q
       (___0_____31139));
  nor2s1 _______503977(.DIN1 (________26293), .DIN2 (___0_____30858),
       .Q (___0__0__31138));
  nor2s1 _______503978(.DIN1 (_________31955), .DIN2 (___0_____30873),
       .Q (___0__9__31137));
  nnd2s1 _______503979(.DIN1 (___0_____31135), .DIN2 (___0_____31134),
       .Q (___0_____31136));
  or2s1 _______503980(.DIN1 (___0_____31132), .DIN2 (___0_____30863),
       .Q (___0_____31133));
  or2s1 _______503981(.DIN1 (____0____31591), .DIN2 (___0__0__30945),
       .Q (___0_____31131));
  or2s1 _______503982(.DIN1 (___0_____31129), .DIN2 (___0_____30913),
       .Q (___0_____31130));
  nor2s1 _______503983(.DIN1 (___0_09__31127), .DIN2 (___0_____30940),
       .Q (___0__0__31128));
  nor2s1 ______503984(.DIN1 (___0_0___31125), .DIN2 (___0__9__30944),
       .Q (___0_0___31126));
  nor2s1 ______503985(.DIN1 (__99_9__30537), .DIN2 (___0_____30938), .Q
       (___0_0___31124));
  nnd2s1 _______503986(.DIN1 (___0_____30914), .DIN2 (__9_____29787),
       .Q (___0_0___31123));
  and2s1 _______503987(.DIN1 (___0_9___30922), .DIN2 (___0_____30789),
       .Q (___0_0___31122));
  nnd2s1 ______503988(.DIN1 (___0_09__30934), .DIN2 (___0_0___30748),
       .Q (___0_0___31121));
  and2s1 ______503989(.DIN1 (___0_0___30929), .DIN2 (___0_0___31119),
       .Q (___0_0___31120));
  nnd2s1 _______503990(.DIN1 (___0_____30952), .DIN2 (___0_____31175),
       .Q (___0_00__31118));
  and2s1 _______503991(.DIN1 (___0_9___31116), .DIN2 (__9_____30321),
       .Q (___0_99__31117));
  nnd2s1 _____9_503992(.DIN1 (___0_____31046), .DIN2 (_________40961),
       .Q (___0_9___31115));
  nnd2s1 _____9_503993(.DIN1 (___0_00__30927), .DIN2 (___0_0___31119),
       .Q (___0_9___31114));
  nnd2s1 _____503994(.DIN1 (___0_9___30925), .DIN2 (___9_0__29593), .Q
       (___0_9___31113));
  nor2s1 _____0_503995(.DIN1 (___0_9___31111), .DIN2 (___0_____30902),
       .Q (___0_9___31112));
  nor2s1 _____0_503996(.DIN1 (_________32931), .DIN2 (___0_9___30923),
       .Q (___0_9___31110));
  nor2s1 _____0_503997(.DIN1 (_____0__27270), .DIN2 (___0_____30951),
       .Q (___0_9___31109));
  or2s1 ______503998(.DIN1 (___0_90__31108), .DIN2 (___0_____30889), .Q
       (___0_9___31399));
  nor2s1 _____503999(.DIN1 (__9_0___29995), .DIN2 (___0_____30802), .Q
       (___0__9__31107));
  nor2s1 _______504000(.DIN1 (____0___28207), .DIN2 (___0_____30794),
       .Q (___0_____31106));
  and2s1 _______504001(.DIN1 (___0_0___30839), .DIN2 (_____0___31609),
       .Q (___0_____31105));
  nnd2s1 _______504002(.DIN1 (___0_____30818), .DIN2 (___0_____30894),
       .Q (___0_____31104));
  nor2s1 _______504003(.DIN1 (___0_____31223), .DIN2 (___0_9___30829),
       .Q (___0_____31103));
  hi1s1 _______504004(.DIN (_________32145), .Q (___0_____31102));
  or2s1 _______504005(.DIN1 (___0_____31100), .DIN2 (___0__0__30804),
       .Q (___0_____31101));
  nor2s1 _______504006(.DIN1 (_____0___31803), .DIN2 (___0_00__30833),
       .Q (___0__0__31099));
  nor2s1 _______504007(.DIN1 (__9_____29908), .DIN2 (___0_____30775),
       .Q (___0__9__31098));
  nnd2s1 _______504008(.DIN1 (___0__0__30814), .DIN2 (___0_____31096),
       .Q (___0_____31097));
  nnd2s1 _______504009(.DIN1 (___0_9___30825), .DIN2 (___0_____31094),
       .Q (___0_____31095));
  nor2s1 ______504010(.DIN1 (___0_____31092), .DIN2 (___0__0__30769),
       .Q (___0_____31093));
  nor2s1 _______504011(.DIN1 (__9_9___30360), .DIN2 (___0_9___30828),
       .Q (___0_____31091));
  nor2s1 ______504012(.DIN1 (________29142), .DIN2 (___0_9___30738), .Q
       (___0__0__31090));
  nor2s1 ______504013(.DIN1 (___0_____31088), .DIN2 (___0__9__30795),
       .Q (___0__9__31089));
  nnd2s1 _______504014(.DIN1 (___0_____30784), .DIN2 (__9__9), .Q
       (___0_____31087));
  nor2s1 _______504015(.DIN1 (________27149), .DIN2 (___0_____30774),
       .Q (___0_____31086));
  nnd2s1 _______504016(.DIN1 (___0_____30772), .DIN2 (___0_____31084),
       .Q (___0_____31085));
  nnd2s1 _______504017(.DIN1 (___0__9__30822), .DIN2 (_________32260),
       .Q (___0_____31083));
  nor2s1 _____9_504018(.DIN1 (___0____25136), .DIN2 (___0_____30779),
       .Q (___0_____31082));
  nor2s1 _____9_504019(.DIN1 (___0__0__31080), .DIN2 (___0__9__30777),
       .Q (___0_____31081));
  and2s1 _____9_504020(.DIN1 (___0__0__30759), .DIN2 (___0_____31078),
       .Q (___0_____31079));
  nor2s1 ______504021(.DIN1 (__9_9___29991), .DIN2 (___0_____30785), .Q
       (___0_____31077));
  nnd2s1 ____90_504022(.DIN1 (___0_____30755), .DIN2 (________28186),
       .Q (___0_____31076));
  nnd2s1 ____504023(.DIN1 (___0_____30762), .DIN2 (____0____32543), .Q
       (___0_____31075));
  nor2s1 ____9_504024(.DIN1 (___0_____31073), .DIN2 (___0__9__30768),
       .Q (___0_____31074));
  or2s1 ____9__504025(.DIN1 (___099___31496), .DIN2 (___0_____30761),
       .Q (___0_____31072));
  nor2s1 ____9__504026(.DIN1 (________28392), .DIN2 (___0_____30799),
       .Q (___0__0__31071));
  nnd2s1 ____9__504027(.DIN1 (___0_____30765), .DIN2 (___0____27853),
       .Q (___0__9__31070));
  nor2s1 ____9__504028(.DIN1 (___9____27783), .DIN2 (___0_____30766),
       .Q (___0_____31069));
  nnd2s1 ____9__504029(.DIN1 (___0_90__30823), .DIN2 (___9____27782),
       .Q (___0_____31068));
  or2s1 ____9__504030(.DIN1 (_________31955), .DIN2 (___0_____30756),
       .Q (___0_____31067));
  nnd2s1 ____9__504031(.DIN1 (___0__9__30758), .DIN2 (________24879),
       .Q (___0_____31066));
  nnd2s1 ____9__504032(.DIN1 (_________40969), .DIN2 (____00___31507),
       .Q (___0_____31065));
  nnd2s1 ____9__504033(.DIN1 (___0_____30782), .DIN2 (___0_____30770),
       .Q (___0_____31064));
  nor2s1 ____9__504034(.DIN1 (_________36852), .DIN2 (___0_____31053),
       .Q (___0_____31063));
  or2s1 ____99_504035(.DIN1 (___0__0__31061), .DIN2 (___0_____30751),
       .Q (___0_____31062));
  nor2s1 ____504036(.DIN1 (__9__9__29877), .DIN2 (___0__0__30750), .Q
       (___0__9__31060));
  nor2s1 ____00_504037(.DIN1 (__9__0__29916), .DIN2 (___0_9___30732),
       .Q (___0_____31059));
  nor2s1 ____0__504038(.DIN1 (________25573), .DIN2 (___0_0___30745),
       .Q (___0_____31058));
  and2s1 ____0__504039(.DIN1 (___0_0___30742), .DIN2 (_________41178),
       .Q (___0_____31057));
  nor2s1 _____0_504040(.DIN1 (__9_____29865), .DIN2 (___0_9___30733),
       .Q (___0_____31056));
  nnd2s1 ______504041(.DIN1 (___0_99__30739), .DIN2 (________28955), .Q
       (___0_____31055));
  nor2s1 _______504042(.DIN1 (________22562), .DIN2 (___0_____31053),
       .Q (___0_____31054));
  nnd2s1 _______504043(.DIN1 (___0_____30776), .DIN2 (____9_9__32410),
       .Q (___0_____31052));
  nor2s1 _______504044(.DIN1 (___0__9__31050), .DIN2 (___0_0___30744),
       .Q (___0__0__31051));
  nnd2s1 _______504045(.DIN1 (___0_9___30736), .DIN2 (inData[31]), .Q
       (___0_____31049));
  nnd2s1 _______504046(.DIN1 (___0_0___30747), .DIN2 (____9___28922),
       .Q (___0_____31048));
  or2s1 _____9_504047(.DIN1 (__9_____30417), .DIN2 (___0_____31046), .Q
       (___0_____31047));
  nnd2s1 _____9_504048(.DIN1 (___0_0___30741), .DIN2 (____9_9__32410),
       .Q (___0_____31045));
  nnd2s1 _____0_504049(.DIN1 (___0_9___30735), .DIN2 (_____0__27103),
       .Q (___0_____31044));
  nor2s1 ______504050(.DIN1 (__9_____29940), .DIN2 (___0_____30754), .Q
       (___0_____31043));
  nnd2s1 _____0_504051(.DIN1 (___0__9__30786), .DIN2 (________28597),
       .Q (___0__0__31042));
  dffacs1 _______________504052(.CLRB (reset), .CLK (clk), .DIN
       (______0__35853), .Q (outData[4]));
  and2s1 _____0_504053(.DIN1 (___0_____30788), .DIN2 (___0_____31040),
       .Q (___0__9__31041));
  xnr2s1 _______504054(.DIN1 (____9____37036), .DIN2 (__99____30519),
       .Q (___0_____31039));
  xor2s1 _______504055(.DIN1 (____0_9__31552), .DIN2 (_____9___38610),
       .Q (___0_____31037));
  and2s1 _____0_504056(.DIN1 (_________40967), .DIN2 (___0_____31035),
       .Q (___0_____31036));
  nor2s1 _____504057(.DIN1 (__9__9__30309), .DIN2 (___0_0___30834), .Q
       (___0_____31034));
  nor2s1 _______504058(.DIN1
       (__________________________________________________________________21986),
       .DIN2 (______0__35853), .Q (___0__0__31033));
  or2s1 ______504059(.DIN1 (___0_0___31031), .DIN2 (___0__9__30720), .Q
       (___0_09__31032));
  nnd2s1 _______504060(.DIN1 (______0__35853), .DIN2
       (__________________________________________________________________21986),
       .Q (___0_0___31030));
  nnd2s1 _______504061(.DIN1 (___0_90__30730), .DIN2 (__90____29657),
       .Q (___0_0___31029));
  nor2s1 _______504062(.DIN1 (___0__9__31147), .DIN2 (___0_____30713),
       .Q (___0_0___31028));
  nor2s1 _____9_504063(.DIN1 (__9_____30441), .DIN2 (___0_____30790),
       .Q (___0_0___31027));
  nnd2s1 _____9_504064(.DIN1 (___0_____30780), .DIN2 (_____0__29407),
       .Q (___0_0___31026));
  nnd2s1 _______504065(.DIN1 (___0_____30714), .DIN2 (__99____30522),
       .Q (___0_0___31025));
  or2s1 _______504066(.DIN1 (___0_0___30835), .DIN2 (___0_00__31023),
       .Q (___0_0___31024));
  nnd2s1 _______504067(.DIN1 (______0__35853), .DIN2 (________28849),
       .Q (___0_99__31022));
  nnd2s1 _______504068(.DIN1 (___0_____30712), .DIN2 (_________31781),
       .Q (___0_9___31021));
  nor2s1 _______504069(.DIN1 (___099___31496), .DIN2 (___0_9___30737),
       .Q (___0_9___31020));
  nor2s1 _______504070(.DIN1 (___0_____30809), .DIN2 (___0_09__30749),
       .Q (___0_9___31019));
  nor2s1 _______504071(.DIN1 (_________32001), .DIN2 (___0_9___30827),
       .Q (___0_9___31018));
  and2s1 _______504072(.DIN1 (___0_9___30826), .DIN2 (______9__31632),
       .Q (___0_9___31017));
  nor2s1 ______504073(.DIN1 (___0_9___31015), .DIN2 (___0_9___30824),
       .Q (___0_9___31016));
  nor2s1 _______504074(.DIN1 (___9____27809), .DIN2 (___0_____30819),
       .Q (___0_9___31014));
  nnd2s1 _______504075(.DIN1 (___0_____30820), .DIN2 (___0_9__28785),
       .Q (___0_90__31013));
  nor2s1 _______504076(.DIN1 (__9_____30062), .DIN2 (___0_____30817),
       .Q (___0__9__31012));
  or2s1 _______504077(.DIN1 (___0_____31010), .DIN2 (___0_____30773),
       .Q (___0_____31011));
  nor2s1 _______504078(.DIN1 (___0_____30760), .DIN2 (___0_____30811),
       .Q (___0_____31009));
  or2s1 _______504079(.DIN1 (___9____29625), .DIN2 (___0_9___30830), .Q
       (___0_____31008));
  nnd2s1 _______504080(.DIN1 (______0__40963), .DIN2 (___0_____31006),
       .Q (___0_____31007));
  nnd2s1 _______504081(.DIN1 (___0_____30808), .DIN2 (___9____26925),
       .Q (___0_____31005));
  and2s1 _______504082(.DIN1 (___0_____30806), .DIN2 (___0__0__31003),
       .Q (___0_____31004));
  and2s1 _______504083(.DIN1 (___0_____30797), .DIN2 (_________31831),
       .Q (___0_____31002));
  nnd2s1 _____504084(.DIN1 (___0_____30791), .DIN2 (________26523), .Q
       (___0_____31001));
  nnd2s1 _____9_504085(.DIN1 (___0_____30792), .DIN2 (_________31944),
       .Q (___0_____31000));
  hi1s1 _______504086(.DIN (___0_____30999), .Q (___0_0___31312));
  hi1s1 ______504087(.DIN (___0_0___31317), .Q (___0_0___31314));
  and2s1 _______504088(.DIN1 (___0__0__31330), .DIN2 (__9_90__30357),
       .Q (_________32806));
  dffacs1 ________________________________________________504089(.CLRB
       (reset), .CLK (clk), .DIN (___0_____30715), .Q
       (______________________________________________21931));
  xor2s1 ______504090(.DIN1 (_____0__29165), .DIN2 (____0_9__31552), .Q
       (_____0___36368));
  dffacs1 ________________________________________________504091(.CLRB
       (reset), .CLK (clk), .DIN (___0__9__30710), .Q
       (_______________________________________________________________9));
  dffacs1 __________________504092(.CLRB (reset), .CLK (clk), .DIN
       (___0_0___30838), .QN (___0_____40411));
  nnd2s1 _______504093(.DIN1 (___0_0___30650), .DIN2 (___0_____30997),
       .Q (___0_____30998));
  and2s1 _______504094(.DIN1 (___0_____30703), .DIN2 (___0_90__30919),
       .Q (___0_____30996));
  nnd2s1 ____09_504095(.DIN1 (__99____30529), .DIN2 (_____9__29362), .Q
       (___0_____30995));
  nor2s1 ____504096(.DIN1 (__9_0___29904), .DIN2 (___000___30552), .Q
       (___0__0__30994));
  nor2s1 ____0__504097(.DIN1 (________28866), .DIN2 (___00____30569),
       .Q (___0__9__30993));
  nor2s1 ____0__504098(.DIN1 (___0_____31132), .DIN2 (__99____30532),
       .Q (___0_____30992));
  nnd2s1 ______504099(.DIN1 (___00____30594), .DIN2 (__9_____30416), .Q
       (___0_____30991));
  nnd2s1 _______504100(.DIN1 (___009___30636), .DIN2 (_____0__29417),
       .Q (___0_____30990));
  nor2s1 _______504101(.DIN1 (___0____27878), .DIN2 (______0__40973),
       .Q (___0_____30989));
  nnd2s1 _______504102(.DIN1 (___0_____30653), .DIN2 (_________41178),
       .Q (___0_____30988));
  or2s1 _______504103(.DIN1 (___0_____30986), .DIN2 (___00_9__30631),
       .Q (___0_____30987));
  nnd2s1 ______504104(.DIN1 (___009___30638), .DIN2 (___0__9__30984),
       .Q (___0__0__30985));
  nnd2s1 _______504105(.DIN1 (___00____30609), .DIN2 (______0__32205),
       .Q (___0_____30983));
  nnd2s1 _______504106(.DIN1 (___00____30599), .DIN2 (________26603),
       .Q (___0_____30982));
  nnd2s1 _______504107(.DIN1 (___0_____30658), .DIN2 (________27605),
       .Q (___0_____30981));
  and2s1 ______504108(.DIN1 (___00____30600), .DIN2 (___0_____30979),
       .Q (___0_____30980));
  or2s1 _______504109(.DIN1 (___0_____30977), .DIN2 (___0__9__30681),
       .Q (___0_____30978));
  nor2s1 _______504110(.DIN1 (__9_____30103), .DIN2 (___00____30617),
       .Q (___0_____30976));
  nnd2s1 _______504111(.DIN1 (___00____30616), .DIN2 (____0____31577),
       .Q (___0__0__30975));
  nnd2s1 ______504112(.DIN1 (___00____30626), .DIN2 (____0____31527),
       .Q (___0__9__30974));
  nnd2s1 _______504113(.DIN1 (___00____30623), .DIN2 (________28957),
       .Q (___0_____30973));
  or2s1 _______504114(.DIN1 (__9_____30401), .DIN2 (___0_____30971), .Q
       (___0_____30972));
  nnd2s1 _______504115(.DIN1 (___0_____30680), .DIN2 (__9990), .Q
       (___0_____30970));
  and2s1 _______504116(.DIN1 (___00____30598), .DIN2 (___0_____30968),
       .Q (___0_____30969));
  nor2s1 _______504117(.DIN1 (_________32001), .DIN2 (___0_____30685),
       .Q (___0_____30967));
  nor2s1 _____504118(.DIN1 (__9__9__29743), .DIN2 (___00____30613), .Q
       (___0_____30966));
  nnd2s1 _____9_504119(.DIN1 (___0_____30694), .DIN2 (____9____32424),
       .Q (___0__0__30965));
  nor2s1 _____9_504120(.DIN1 (________29359), .DIN2 (___0_0___30648),
       .Q (___0__9__30964));
  nor2s1 _____9_504121(.DIN1 (____9___26402), .DIN2 (___00_0__30622),
       .Q (___0_____30963));
  nor2s1 ____504122(.DIN1 (___0_____30961), .DIN2 (___00____30558), .Q
       (___0_____30962));
  nor2s1 ____90_504123(.DIN1 (___0__9__31347), .DIN2 (___00_9__30611),
       .Q (___0_____30960));
  and2s1 ____9__504124(.DIN1 (___00_9__30602), .DIN2 (___0_____30958),
       .Q (___0_____30959));
  or2s1 ____9__504125(.DIN1 (___0_____30956), .DIN2 (___00____30607),
       .Q (___0_____30957));
  nnd2s1 ____9_504126(.DIN1 (___00____30597), .DIN2 (___990__26041), .Q
       (___0__0__30955));
  nnd2s1 ____9__504127(.DIN1 (___00____30601), .DIN2 (___0_____31237),
       .Q (___0__9__30954));
  nor2s1 ____9__504128(.DIN1 (____0___25769), .DIN2 (_________40971),
       .Q (___0_____30953));
  nor2s1 ____0__504129(.DIN1 (_____0___31991), .DIN2 (___00____30590),
       .Q (___0_____30952));
  nnd2s1 ____0__504130(.DIN1 (___00____30604), .DIN2 (________27156),
       .Q (___0_____30951));
  nnd2s1 ____9__504131(.DIN1 (__9_9___30080), .DIN2 (___00____30591),
       .Q (___0_____30950));
  nnd2s1 ____9__504132(.DIN1 (___0_____30708), .DIN2 (___0_____30948),
       .Q (___0_____30949));
  nnd2s1 ____9__504133(.DIN1 (_________40975), .DIN2 (__9_90), .Q
       (___0_____30947));
  or2s1 ____9__504134(.DIN1 (___00____30586), .DIN2 (__99____30476), .Q
       (___0_____30946));
  nnd2s1 ____9__504135(.DIN1 (___00_0__30584), .DIN2 (______9__32019),
       .Q (___0__0__30945));
  nnd2s1 ____9__504136(.DIN1 (___00____30581), .DIN2 (___0_____30943),
       .Q (___0__9__30944));
  nnd2s1 ____9__504137(.DIN1 (__99____30523), .DIN2 (________29451), .Q
       (___0_____30942));
  nnd2s1 ____9__504138(.DIN1 (___00____30579), .DIN2 (________26299),
       .Q (___0_____30941));
  or2s1 ____9__504139(.DIN1 (___0_____30939), .DIN2 (__99____30526), .Q
       (___0_____30940));
  and2s1 ____99_504140(.DIN1 (___0_____30937), .DIN2 (________29537),
       .Q (___0_____30938));
  nnd2s1 ____504141(.DIN1 (___00____30557), .DIN2 (___0_____30844), .Q
       (___0_____30936));
  or2s1 ____00_504142(.DIN1 (___09_9__31465), .DIN2 (___00_0__30574),
       .Q (___0__0__30935));
  nnd2s1 ____00_504143(.DIN1 (___00_9__30573), .DIN2 (_________31725),
       .Q (___0_09__30934));
  nnd2s1 ____0__504144(.DIN1 (___00____30571), .DIN2 (__9_9___30079),
       .Q (___0_0___30933));
  and2s1 ____0__504145(.DIN1 (___00____30567), .DIN2 (___0_____30958),
       .Q (___0_0___30932));
  nor2s1 ____0__504146(.DIN1 (_________41156), .DIN2 (___00____30572),
       .Q (___0_0___30931));
  and2s1 ____0_504147(.DIN1 (___00____30588), .DIN2 (________26299), .Q
       (___0_0___30930));
  and2s1 ____0__504148(.DIN1 (___00____30566), .DIN2 (___0_99__30926),
       .Q (___0_0___30929));
  nnd2s1 ____0_504149(.DIN1 (___00_0__30565), .DIN2 (___99___27826), .Q
       (___0_0___30928));
  and2s1 ____0__504150(.DIN1 (__99____30530), .DIN2 (___0_99__30926),
       .Q (___0_00__30927));
  nnd2s1 ____0__504151(.DIN1 (___00____30563), .DIN2 (________26723),
       .Q (___0_9___30925));
  and2s1 ____0_504152(.DIN1 (___00____30561), .DIN2 (_________31868),
       .Q (___0_9___30924));
  nnd2s1 ____0_504153(.DIN1 (___00____30560), .DIN2 (_________41321),
       .Q (___0_9___30923));
  nor2s1 ____0__504154(.DIN1 (____0___27488), .DIN2 (___00____30577),
       .Q (___0_9___30922));
  nnd2s1 ____9__504155(.DIN1 (___0_0___30646), .DIN2 (_________32611),
       .Q (___0_____31135));
  nor2s1 ____9__504156(.DIN1 (________27161), .DIN2 (___00____30629),
       .Q (___0_____31153));
  nnd2s1 _______504157(.DIN1 (___00____30595), .DIN2 (____0____32532),
       .Q (_________32818));
  nnd2s1 _______504158(.DIN1 (___0_____30687), .DIN2 (_______22172), .Q
       (_________35696));
  hi1s1 _______504159(.DIN (___0_9___30921), .Q (_________31938));
  nb1s1 _______504160(.DIN (___0_9___30921), .Q (_________32145));
  nnd2s1 _______504161(.DIN1 (___0_____30655), .DIN2 (___0_90__30919),
       .Q (___0_9___30920));
  nnd2s1 _____0_504162(.DIN1 (___00____30582), .DIN2 (___0_____30917),
       .Q (___0__9__30918));
  or2s1 _______504163(.DIN1 (_________33986), .DIN2 (___0000__30545),
       .Q (___0_____30916));
  nor2s1 _______504164(.DIN1 (___0____27837), .DIN2 (__999___30540), .Q
       (___0_____30915));
  nor2s1 _______504165(.DIN1 (________28958), .DIN2 (__999___30538), .Q
       (___0_____30914));
  nnd2s1 ______504166(.DIN1 (__99_0__30528), .DIN2 (___0_____30912), .Q
       (___0_____30913));
  nnd2s1 _______504167(.DIN1 (____9____37998), .DIN2 (__99____30535),
       .Q (___0_____30911));
  nnd2s1 _______504168(.DIN1 (__999___30542), .DIN2 (________29266), .Q
       (___0_____30910));
  nnd2s1 _______504169(.DIN1 (___000___30550), .DIN2 (___0_0__26092),
       .Q (___0__0__30909));
  nnd2s1 ______504170(.DIN1 (___000___30548), .DIN2 (____9___28638), .Q
       (___0__9__30908));
  nor2s1 ______504171(.DIN1 (_________31866), .DIN2 (___000___30546),
       .Q (___0_____30907));
  nor2s1 ______504172(.DIN1 (___0_00__30642), .DIN2 (___00____30585),
       .Q (___0_____30906));
  and2s1 ______504173(.DIN1 (___00____30580), .DIN2 (_____0___32676),
       .Q (___0_____30905));
  nnd2s1 _______504174(.DIN1 (___00____30559), .DIN2 (___0_____30903),
       .Q (___0_____30904));
  nnd2s1 _______504175(.DIN1 (__99____30524), .DIN2 (___0__9__31280),
       .Q (___0_____30902));
  nor2s1 _______504176(.DIN1 (________27153), .DIN2 (__99____30534), .Q
       (___0_____30901));
  nor2s1 _______504177(.DIN1 (__9_____30028), .DIN2 (__99____30521), .Q
       (___0_____30900));
  nor2s1 _____9_504178(.DIN1 (______0__32253), .DIN2 (___0__9__30898),
       .Q (___0__0__30899));
  nnd2s1 _____0_504179(.DIN1 (__999___30544), .DIN2 (______0__41180),
       .Q (___0_____30897));
  nnd2s1 _______504180(.DIN1 (__99_9__30517), .DIN2 (________27339), .Q
       (___0_____30896));
  nnd2s1 _______504181(.DIN1 (__99_0__30518), .DIN2 (___0_____30894),
       .Q (___0_____30895));
  dffacs1 _______________504182(.CLRB (reset), .CLK (clk), .DIN
       (____0_9__31552), .Q (outData[3]));
  or2s1 _______504183(.DIN1 (____________), .DIN2 (_________40977), .Q
       (___0_____30893));
  and2s1 _______504184(.DIN1 (_________40977), .DIN2 (____________), .Q
       (___0_____30892));
  nor2s1 _______504185(.DIN1 (___0__9__30890), .DIN2 (___0_____30657),
       .Q (___0__0__30891));
  nnd2s1 _______504186(.DIN1 (___00____30618), .DIN2 (___0_____30888),
       .Q (___0_____30889));
  xor2s1 _______504187(.DIN1 (________28120), .DIN2 (___0_____30886),
       .Q (___0_____30887));
  xor2s1 _______504188(.DIN1 (___0_____30886), .DIN2 (_________38573),
       .Q (___0_____30885));
  xor2s1 _______504189(.DIN1 (________27673), .DIN2 (___0_____30886),
       .Q (___0_____30884));
  nor2s1 _______504190(.DIN1 (___0_____30882), .DIN2 (___00_0__30555),
       .Q (___0_____30883));
  and2s1 _______504191(.DIN1 (___0_____30706), .DIN2 (___0__9__30880),
       .Q (___0__0__30881));
  or2s1 _____504192(.DIN1 (_________33551), .DIN2 (___0099__30641), .Q
       (___0_____30879));
  nor2s1 _______504193(.DIN1 (________27603), .DIN2 (___0_0___31311),
       .Q (___0_____30878));
  nor2s1 ______504194(.DIN1 (__9_0___30274), .DIN2 (___0_____30704), .Q
       (___0_____30877));
  or2s1 _____0_504195(.DIN1 (____0____31591), .DIN2 (___0__0__30672),
       .Q (___0_____30876));
  nnd2s1 _____9_504196(.DIN1 (___00_0__30593), .DIN2 (__9_____30314),
       .Q (___0_____30875));
  nor2s1 _____9_504197(.DIN1 (____0___29011), .DIN2 (___009___30635),
       .Q (___0_____30874));
  or2s1 ______504198(.DIN1 (___0__0__30872), .DIN2 (___0_____30660), .Q
       (___0_____30873));
  and2s1 ______504199(.DIN1 (___0_0___30643), .DIN2 (___0_____30870),
       .Q (___0__9__30871));
  nor2s1 _______504200(.DIN1 (____9___28103), .DIN2 (___00____30614),
       .Q (___0_____30869));
  nor2s1 _______504201(.DIN1 (________29515), .DIN2 (___0__0__30701),
       .Q (___0_____30868));
  nor2s1 _______504202(.DIN1 (___0_____30866), .DIN2 (___009___30633),
       .Q (___0_____30867));
  and2s1 _______504203(.DIN1 (___0_____30698), .DIN2 (__9_____30345),
       .Q (___0_____30865));
  nnd2s1 _______504204(.DIN1 (___0_____30696), .DIN2 (________25545),
       .Q (___0_____30864));
  or2s1 _______504205(.DIN1 (________27504), .DIN2 (___0_____30702), .Q
       (___0_____30863));
  and2s1 _______504206(.DIN1 (___0_____30693), .DIN2 (__9_____29968),
       .Q (___0__0__30862));
  nor2s1 _______504207(.DIN1 (________29173), .DIN2 (___0__0__30692),
       .Q (___0__9__30861));
  nnd2s1 _______504208(.DIN1 (___00____30628), .DIN2 (____9___29463),
       .Q (___0_____30860));
  nor2s1 ______504209(.DIN1 (___0_____30699), .DIN2 (________26787), .Q
       (___0_____30859));
  nnd2s1 ______504210(.DIN1 (___009___30640), .DIN2 (________29441), .Q
       (___0_____30858));
  nnd2s1 _______504211(.DIN1 (___0__9__30691), .DIN2 (___0____26120),
       .Q (___0_____30857));
  nor2s1 _______504212(.DIN1 (___0__9__30890), .DIN2 (___0_____30659),
       .Q (___0_____30856));
  nor2s1 ______504213(.DIN1 (__9_____29742), .DIN2 (___0__0__30682), .Q
       (___0_____30855));
  and2s1 _______504214(.DIN1 (___00____30620), .DIN2 (___909__28654),
       .Q (___0_____30854));
  nor2s1 _______504215(.DIN1 (___0_____30801), .DIN2 (___0_____30678),
       .Q (___0_____30853));
  nnd2s1 _______504216(.DIN1 (___00____30624), .DIN2 (___0__9__30851),
       .Q (___0__0__30852));
  nor2s1 _______504217(.DIN1 (________29053), .DIN2 (___0_____30677),
       .Q (___0_____30850));
  nor2s1 _______504218(.DIN1 (___9_0__26940), .DIN2 (___0_____30670),
       .Q (___0_____30849));
  nnd2s1 _______504219(.DIN1 (___0_____30668), .DIN2 (________25926),
       .Q (___0_____30848));
  and2s1 _______504220(.DIN1 (___0_____30664), .DIN2 (_________32720),
       .Q (___0_____30847));
  nnd2s1 _______504221(.DIN1 (___0_____30667), .DIN2 (_____09__31612),
       .Q (___0_____30846));
  nnd2s1 ______504222(.DIN1 (___0__0__30652), .DIN2 (___0_____30844),
       .Q (___0_____30845));
  nnd2s1 _____9_504223(.DIN1 (___0_____30666), .DIN2 (____9___28642),
       .Q (___0_____30843));
  nor2s1 _____0_504224(.DIN1 (_________31667), .DIN2 (___000___30547),
       .Q (___0_9___31116));
  nnd2s1 ______504225(.DIN1 (___0_0___30840), .DIN2 (___0_09__30841),
       .Q (___0_____31038));
  nnd2s1 _______504226(.DIN1 (____0_9__31552), .DIN2 (________29483),
       .Q (___0_____30999));
  hi1s1 ______504227(.DIN (___0__0__30842), .Q (___0_9___31211));
  nor2s1 _______504228(.DIN1 (___0_09__30841), .DIN2 (___0_0___30840),
       .Q (___0_0___31220));
  nor2s1 _______504229(.DIN1 (________28848), .DIN2 (____0_9__31552),
       .Q (___0_0___31317));
  and2s1 _______504230(.DIN1 (___0_0___31311), .DIN2 (________27603),
       .Q (______0__36056));
  and2s1 ____504231(.DIN1 (__9_9___30452), .DIN2 (____0____31581), .Q
       (___0_0___30839));
  nnd2s1 _______504232(.DIN1 (____0____37147), .DIN2 (__9_____30406),
       .Q (___0_0___30838));
  nnd2s1 ____9__504233(.DIN1 (__99____30483), .DIN2 (________29322), .Q
       (___0_0___30837));
  or2s1 ____9_504234(.DIN1 (___0_9___40270), .DIN2 (__99_0__30509), .Q
       (___0_0___30836));
  xor2s1 ____9_504235(.DIN1
       (________________________________________________________________),
       .DIN2
       (__________________________________________________________________21990),
       .Q (___0_0___30835));
  nor2s1 _______504236(.DIN1 (_________32159), .DIN2 (___0_____30803),
       .Q (___0_0___30834));
  nnd2s1 ______504237(.DIN1 (__99_9__30478), .DIN2 (___0_99__30832), .Q
       (___0_00__30833));
  xor2s1 ____9__504238(.DIN1 (___00____30596), .DIN2 (____9___28467),
       .Q (___0_9___30831));
  nnd2s1 _______504239(.DIN1 (__9_____30408), .DIN2 (__90____29671), .Q
       (___0_9___30830));
  nnd2s1 ____9__504240(.DIN1 (__9__0__30403), .DIN2 (___0_____30793),
       .Q (___0_9___30829));
  nnd2s1 ____9__504241(.DIN1 (__99____30475), .DIN2 (________28133), .Q
       (___0_9___30828));
  nor2s1 ____9__504242(.DIN1 (__9__0__29946), .DIN2 (__99____30474), .Q
       (___0_9___30827));
  and2s1 ____9__504243(.DIN1 (__9__0__30420), .DIN2 (___09____31443),
       .Q (___0_9___30826));
  nor2s1 ____9_504244(.DIN1 (__9_____30400), .DIN2 (__99____30472), .Q
       (___0_9___30825));
  or2s1 ____9__504245(.DIN1 (__99____30525), .DIN2 (__99____30471), .Q
       (___0_9___30824));
  nor2s1 ____9__504246(.DIN1 (____00__25586), .DIN2 (__9_____30397), .Q
       (___0_90__30823));
  nor2s1 ____9__504247(.DIN1 (___0_____30821), .DIN2 (__99____30464),
       .Q (___0__9__30822));
  nnd2s1 ____9__504248(.DIN1 (__99____30462), .DIN2 (___0_____30783),
       .Q (___0_____30820));
  nnd2s1 ____504249(.DIN1 (__990___30460), .DIN2 (__99__), .Q
       (___0_____30819));
  and2s1 ____99_504250(.DIN1 (__9909), .DIN2 (___0_____30844), .Q
       (___0_____30818));
  and2s1 ____99_504251(.DIN1 (___0_____30816), .DIN2 (_____9__27471),
       .Q (___0_____30817));
  nnd2s1 ____99_504252(.DIN1 (__9_____30424), .DIN2 (________27980), .Q
       (___0_____30815));
  nor2s1 ____99_504253(.DIN1 (___0__9__30813), .DIN2 (__99_9), .Q
       (___0__0__30814));
  nnd2s1 ____99_504254(.DIN1 (__990___30458), .DIN2 (___0_9__27864), .Q
       (___0_____30812));
  nnd2s1 ____99_504255(.DIN1 (__99_0), .DIN2 (___0_____30810), .Q
       (___0_____30811));
  nnd2s1 ____00_504256(.DIN1 (__990___30457), .DIN2 (__9_____29876), .Q
       (___0_____30809));
  and2s1 ____00_504257(.DIN1 (__9_____30412), .DIN2 (___0_____30807),
       .Q (___0_____30808));
  and2s1 ____00_504258(.DIN1 (__9_9___30453), .DIN2 (___0_____30805),
       .Q (___0_____30806));
  nnd2s1 _______504259(.DIN1 (__9_____30383), .DIN2 (___0____27861), .Q
       (___0__0__30804));
  or2s1 ____0__504260(.DIN1 (___0_____30801), .DIN2 (__9_9___30450), .Q
       (___0_____30802));
  nor2s1 ____0__504261(.DIN1 (__9_0___30184), .DIN2 (__9_9___30448), .Q
       (___0_____30800));
  or2s1 ____0__504262(.DIN1 (___0_____30798), .DIN2 (__99____30470), .Q
       (___0_____30799));
  and2s1 ____0__504263(.DIN1 (__9_90__30445), .DIN2 (___0__0__30796),
       .Q (___0_____30797));
  nnd2s1 ____0_504264(.DIN1 (__9__0__30411), .DIN2 (__9_____30306), .Q
       (___0__9__30795));
  nnd2s1 ____0__504265(.DIN1 (__9_____30431), .DIN2 (___0_____30793),
       .Q (___0_____30794));
  and2s1 ____0__504266(.DIN1 (__9_____30387), .DIN2 (__9_____30316), .Q
       (___0_____30792));
  nor2s1 ____0_504267(.DIN1 (________26449), .DIN2 (__9__9__30384), .Q
       (___0_____30791));
  nnd2s1 ____0__504268(.DIN1 (__9_____30443), .DIN2 (___0_____30789),
       .Q (___0_____30790));
  and2s1 ____0__504269(.DIN1 (__9_____30435), .DIN2 (___0__0__30787),
       .Q (___0_____30788));
  nor2s1 ____0__504270(.DIN1 (__9_____30399), .DIN2 (_____9___41008),
       .Q (___0__9__30786));
  nnd2s1 ____0__504271(.DIN1 (__9_____30433), .DIN2 (___0_90__30919),
       .Q (___0_____30785));
  nnd2s1 _______504272(.DIN1 (__9_99__30454), .DIN2 (___0_____30783),
       .Q (___0_____30784));
  nor2s1 ____0__504273(.DIN1 (___0_0__28776), .DIN2 (__9_____30440), .Q
       (___0_____30782));
  nor2s1 ____09_504274(.DIN1 (____9___27475), .DIN2 (__990_), .Q
       (___0_____30781));
  nor2s1 ____09_504275(.DIN1 (__9_____30115), .DIN2 (__9_____30389), .Q
       (___0_____30780));
  nor2s1 ____09_504276(.DIN1 (_____9___33155), .DIN2 (__9_____30413),
       .Q (___0_____30779));
  nnd2s1 ____504277(.DIN1 (__9__9__30410), .DIN2 (___0____28782), .Q
       (___0__0__30778));
  nnd2s1 _______504278(.DIN1 (__99____30466), .DIN2 (__9__0__30234), .Q
       (___0__9__30777));
  nnd2s1 ____9__504279(.DIN1 (___0_0___30645), .DIN2
       (______________22065), .Q (___0_____31134));
  xor2s1 ____9_504280(.DIN1 (___0_____30686), .DIN2 (__9_____29972), .Q
       (___0_9___30921));
  nnd2s1 ____9__504281(.DIN1 (__99____30494), .DIN2 (_________34154),
       .Q (____0____31559));
  dffacs1 _______________________________________504282(.CLRB (reset),
       .CLK (clk), .DIN (__99____30510), .QN (______________22105));
  nnd2s1 ____0__504283(.DIN1 (__9_____30442), .DIN2 (____9___25578), .Q
       (_________36643));
  hi1s1 _______504284(.DIN (___0_0___31311), .Q (______0__35853));
  nnd2s1 _______504285(.DIN1 (__9_____30376), .DIN2 (__9_____30035), .Q
       (___0_____30776));
  nnd2s1 _______504286(.DIN1 (__99____30512), .DIN2 (___900__29553), .Q
       (___0_____30775));
  nor2s1 _______504287(.DIN1 (_________41291), .DIN2 (__9_____30391),
       .Q (___0_____30774));
  nnd2s1 _______504288(.DIN1 (__9_____30404), .DIN2 (________28272), .Q
       (___0_____30773));
  and2s1 _______504289(.DIN1 (__9_____30388), .DIN2 (___0_____30771),
       .Q (___0_____30772));
  nor2s1 _______504290(.DIN1 (__9_9___29800), .DIN2 (__9__9__30402), .Q
       (___0_____30770));
  nor2s1 _______504291(.DIN1 (____0___29372), .DIN2 (_________40981),
       .Q (___0__0__30769));
  nnd2s1 _______504292(.DIN1 (__9_9___30447), .DIN2 (______0__32108),
       .Q (___0__9__30768));
  nnd2s1 ______504293(.DIN1 (__9_____30395), .DIN2 (____0___29010), .Q
       (___0_____30767));
  nnd2s1 _______504294(.DIN1 (__9_____30392), .DIN2 (____9___27294), .Q
       (___0_____30766));
  nor2s1 _______504295(.DIN1 (___0_____30764), .DIN2 (__9_____30390),
       .Q (___0_____30765));
  nnd2s1 _______504296(.DIN1 (__9_____30386), .DIN2 (________29298), .Q
       (___0_____30763));
  or2s1 _______504297(.DIN1 (___09____31480), .DIN2 (__9_____30439), .Q
       (___0_____30762));
  or2s1 ______504298(.DIN1 (___0_____30760), .DIN2 (__9_____30405), .Q
       (___0_____30761));
  nor2s1 _______504299(.DIN1 (________28277), .DIN2 (__99____30481), .Q
       (___0__0__30759));
  nnd2s1 _______504300(.DIN1 (__99____30511), .DIN2 (____00___31511),
       .Q (___0__9__30758));
  nor2s1 _____504301(.DIN1 (_____90__32273), .DIN2 (__9_____30425), .Q
       (___0_____30757));
  nnd2s1 _____9_504302(.DIN1 (__9_____30381), .DIN2 (__99____30465), .Q
       (___0_____30756));
  nnd2s1 _____9_504303(.DIN1 (__9_____30382), .DIN2 (_____9__27471), .Q
       (___0_____30755));
  nor2s1 _____504304(.DIN1 (________27149), .DIN2 (__9_____30427), .Q
       (___0_____30754));
  and2s1 _______504305(.DIN1 (__99_9__30498), .DIN2 (___0_____30752),
       .Q (___0_____30753));
  nnd2s1 _______504306(.DIN1 (___0_9___30734), .DIN2 (________29501),
       .Q (___0_____30751));
  and2s1 _______504307(.DIN1 (___0_09__30749), .DIN2 (___0_0___30748),
       .Q (___0__0__30750));
  nor2s1 _____9_504308(.DIN1 (___0_0___30746), .DIN2 (__9_____30377),
       .Q (___0_0___30747));
  nnd2s1 _____0_504309(.DIN1 (__9_____30379), .DIN2 (________28030), .Q
       (___0_0___30745));
  or2s1 _______504310(.DIN1 (___0_0___30743), .DIN2 (__9_0___30367), .Q
       (___0_0___30744));
  nor2s1 _____9_504311(.DIN1 (__9_____30071), .DIN2 (__9_0___30371), .Q
       (___0_0___30742));
  nnd2s1 _______504312(.DIN1 (__9__0__30375), .DIN2 (___0_00__30740),
       .Q (___0_0___30741));
  and2s1 _______504313(.DIN1 (__9_09__30374), .DIN2 (_________31953),
       .Q (___0_99__30739));
  nnd2s1 _______504314(.DIN1 (__9_____30422), .DIN2 (________28543), .Q
       (___0_9___30738));
  nnd2s1 ______504315(.DIN1 (__9__0__30429), .DIN2 (___0_____30679), .Q
       (___0_9___30737));
  or2s1 _______504316(.DIN1 (___0_____30866), .DIN2 (__9_0___30368), .Q
       (___0_9___30736));
  and2s1 _______504317(.DIN1 (___0_9___30734), .DIN2 (________28211),
       .Q (___0_9___30735));
  or2s1 _____9_504318(.DIN1 (_________32854), .DIN2 (__9_0___30370), .Q
       (___0_9___30733));
  nnd2s1 _____504319(.DIN1 (__9_0___30372), .DIN2 (___9____29574), .Q
       (___0_9___30732));
  nor2s1 _______504320(.DIN1 (__9_____29827), .DIN2 (__9_0___30369), .Q
       (___0_9___30731));
  nor2s1 _______504321(.DIN1 (________28535), .DIN2 (__99____30495), .Q
       (___0_90__30730));
  nnd2s1 _______504322(.DIN1 (___0_____30886), .DIN2 (___0_____30727),
       .Q (___0__9__30729));
  nor2s1 _______504323(.DIN1 (___0_____30727), .DIN2 (___0_____30886),
       .Q (___0_____30728));
  nor2s1 _______504324(.DIN1
       (__________________________________________), .DIN2
       (__9__9__30437), .Q (___0_____30726));
  nnd2s1 _______504325(.DIN1 (__9__9__30437), .DIN2
       (__________________________________________), .Q
       (___0_____30725));
  and2s1 _______504326(.DIN1 (___0_____30886), .DIN2 (_________22046),
       .Q (___0_____30724));
  nor2s1 _______504327(.DIN1 (_________22046), .DIN2 (___0_____30886),
       .Q (___0_____30723));
  nor2s1 _____0_504328(.DIN1
       (____________________________________________21818), .DIN2
       (__9__9__30437), .Q (___0_____30722));
  nnd2s1 _____0_504329(.DIN1 (__9__9__30437), .DIN2
       (____________________________________________21818), .Q
       (___0__0__30721));
  nnd2s1 _______504330(.DIN1 (__99____30493), .DIN2 (___0_____30719),
       .Q (___0__9__30720));
  nor2s1 _______504331(.DIN1
       (_________________________________________0___21895), .DIN2
       (___0_____30717), .Q (___0_____30718));
  nor2s1 _______504332(.DIN1 (___0_____30709), .DIN2 (___0_____30717),
       .Q (___0_____30716));
  nnd2s1 _______504333(.DIN1 (__99____30502), .DIN2 (___09___26138), .Q
       (___0_____30715));
  nor2s1 _______504334(.DIN1 (________29300), .DIN2 (__99____30503), .Q
       (___0_____30714));
  or2s1 _______504335(.DIN1 (______0__32892), .DIN2 (__99_9__30488), .Q
       (___0_____30713));
  nor2s1 ______504336(.DIN1 (________26840), .DIN2 (__99____30507), .Q
       (___0_____30712));
  nor2s1 _______504337(.DIN1 (___0_0__28805), .DIN2 (__99____30505), .Q
       (___0__0__30711));
  or2s1 _______504338(.DIN1 (__99____30504), .DIN2 (________27674), .Q
       (___0__9__30710));
  nnd2s1 _______504339(.DIN1 (___0_____30717), .DIN2
       (_________________________________________0___21895), .Q
       (___09____31453));
  nnd2s1 _______504340(.DIN1 (___0_____30717), .DIN2 (___0_____30709),
       .Q (___0__0__30842));
  hi1s1 _____0_504341(.DIN (___0_____30708), .Q (___0_____31053));
  nor2s1 _______504342(.DIN1 (_________31809), .DIN2 (__9_____30434),
       .Q (___0_____31046));
  xor2s1 _______504343(.DIN1 (__9_____30353), .DIN2 (___0_____40308),
       .Q (___0__0__31330));
  nor2s1 _______504344(.DIN1 (____9____33386), .DIN2 (__9_____30245),
       .Q (___0_____30707));
  nor2s1 _____9_504345(.DIN1 (________26424), .DIN2 (__9_____30355), .Q
       (___0_____30706));
  xor2s1 ____9__504346(.DIN1 (_________22045), .DIN2 (__9_____30118),
       .Q (___0_____30705));
  nnd2s1 ______504347(.DIN1 (__9_9___30359), .DIN2 (_____0__25379), .Q
       (___0_____30704));
  nor2s1 ____9__504348(.DIN1 (__9_____30198), .DIN2 (__9__0__30338), .Q
       (___0_____30703));
  nnd2s1 ____9_504349(.DIN1 (__9_____30283), .DIN2 (___0_____31175), .Q
       (___0_____30702));
  nnd2s1 ____9__504350(.DIN1 (__9__0__30347), .DIN2 (__9_____29863), .Q
       (___0__0__30701));
  nor2s1 ____9__504351(.DIN1 (__9_____30346), .DIN2 (________29076), .Q
       (___0_____30700));
  nor2s1 ____9__504352(.DIN1 (__900___29642), .DIN2 (___0_____30690),
       .Q (___0_____30699));
  nor2s1 ____9__504353(.DIN1 (___0_____30697), .DIN2 (__9_____30284),
       .Q (___0_____30698));
  or2s1 ____9__504354(.DIN1 (___0_____30695), .DIN2 (__9_____30343), .Q
       (___0_____30696));
  nor2s1 ____9_504355(.DIN1 (___9____29571), .DIN2 (__9_____30342), .Q
       (___0_____30694));
  nor2s1 ____9_504356(.DIN1 (__99____30492), .DIN2 (__9_____30341), .Q
       (___0_____30693));
  nnd2s1 ____9__504357(.DIN1 (__9_9___30266), .DIN2 (________28596), .Q
       (___0__0__30692));
  nor2s1 ____9_504358(.DIN1 (________22440), .DIN2 (___0_____30690), .Q
       (___0__9__30691));
  nor2s1 ____9_504359(.DIN1 (__9_0___30279), .DIN2 (___0_____30688), .Q
       (___0_____30689));
  or2s1 ____9__504360(.DIN1 (_______22244), .DIN2 (___0_____30686), .Q
       (___0_____30687));
  and2s1 ____9__504361(.DIN1 (__9_____30344), .DIN2 (___0_____30684),
       .Q (___0_____30685));
  nor2s1 ____9__504362(.DIN1 (_________32001), .DIN2 (__9_____30336),
       .Q (___0_____30683));
  nnd2s1 ____00_504363(.DIN1 (______0__40983), .DIN2 (__9_____30058),
       .Q (___0__0__30682));
  nnd2s1 ____00_504364(.DIN1 (__9_____30331), .DIN2 (________28084), .Q
       (___0__9__30681));
  nnd2s1 ____0__504365(.DIN1 (__9_____30327), .DIN2 (___0_____30679),
       .Q (___0_____30680));
  or2s1 ____0__504366(.DIN1 (____0___28201), .DIN2 (__9_____30326), .Q
       (___0_____30678));
  nnd2s1 ____0__504367(.DIN1 (__9_____30287), .DIN2 (___0_____30676),
       .Q (___0_____30677));
  nor2s1 ____0_504368(.DIN1 (____9____32439), .DIN2 (__9__0__30282), .Q
       (___0_____30675));
  nnd2s1 ____0__504369(.DIN1 (___0_____30673), .DIN2 (___0_____30783),
       .Q (___0_____30674));
  nnd2s1 ____0__504370(.DIN1 (__9_____30301), .DIN2 (___0__9__30671),
       .Q (___0__0__30672));
  or2s1 ____0__504371(.DIN1 (___0_____30669), .DIN2 (__9_____30323), .Q
       (___0_____30670));
  nor2s1 ____0_504372(.DIN1 (___09_9__31446), .DIN2 (__9__0__30320), .Q
       (___0_____30668));
  nor2s1 ____0__504373(.DIN1 (__9_____30098), .DIN2 (__9_____30317), .Q
       (___0_____30667));
  nor2s1 ____0__504374(.DIN1 (________27951), .DIN2 (__9_____30428), .Q
       (___0_____30666));
  nnd2s1 ____0__504375(.DIN1 (__9_____30315), .DIN2 (___9____26906), .Q
       (___0_____30665));
  nor2s1 ____0__504376(.DIN1 (___00____30630), .DIN2 (__9_9___30363),
       .Q (___0_____30664));
  nor2s1 ____0__504377(.DIN1 (___00___27833), .DIN2 (__9__0__30310), .Q
       (___0_____30663));
  and2s1 ____0__504378(.DIN1 (__9_0___30278), .DIN2 (___0__9__30661),
       .Q (___0__0__30662));
  or2s1 ____0__504379(.DIN1 (_____0___31994), .DIN2 (__9_____30307), .Q
       (___0_____30660));
  nor2s1 ____0__504380(.DIN1 (________26734), .DIN2 (__9_____30289), .Q
       (___0_____30659));
  nor2s1 ____0_504381(.DIN1 (________27982), .DIN2 (__9_____30304), .Q
       (___0_____30658));
  nor2s1 ____0_504382(.DIN1 (___0_____30656), .DIN2 (__9_____30302), .Q
       (___0_____30657));
  and2s1 ____0__504383(.DIN1 (__9_90__30263), .DIN2 (___0_____30654),
       .Q (___0_____30655));
  nor2s1 ____0__504384(.DIN1 (__9_____30303), .DIN2 (_________40985),
       .Q (___0_____30653));
  and2s1 ____0__504385(.DIN1 (__9__9__30329), .DIN2 (___0_09__30651),
       .Q (___0__0__30652));
  nor2s1 ____0__504386(.DIN1 (___0_0___30649), .DIN2 (__9_____30299),
       .Q (___0_0___30650));
  nnd2s1 _______504387(.DIN1 (__9_9___30265), .DIN2 (_________31811),
       .Q (___0_0___30648));
  nnd2s1 ____0_504388(.DIN1
       (________________________________________________________________),
       .DIN2 (__________________________________________9_), .Q
       (___0_0___30647));
  hi1s1 ____0__504389(.DIN (___0_0___30645), .Q (___0_0___30646));
  nnd2s1 ____0__504390(.DIN1 (__9_____29872), .DIN2 (__9_____30352), .Q
       (___0_0___30644));
  nor2s1 ____0__504391(.DIN1 (___0_00__30642), .DIN2 (__9_____30351),
       .Q (___0_0___30643));
  or2s1 ____0__504392(.DIN1 (_________33217), .DIN2 (__9_____30257), .Q
       (___0099__30641));
  and2s1 ____0_504393(.DIN1 (__9_____30240), .DIN2 (___0_____31164), .Q
       (___009___30640));
  nnd2s1 ____0_504394(.DIN1 (__9_____30308), .DIN2 (__9_9___30270), .Q
       (___009___30639));
  nor2s1 ____0__504395(.DIN1 (___9____25999), .DIN2 (__9_____30334), .Q
       (___009___30638));
  nnd2s1 ____0__504396(.DIN1 (__9_____30286), .DIN2 (_________32266),
       .Q (___009___30637));
  nor2s1 ____0_504397(.DIN1 (__9_____30039), .DIN2 (__9__0__30244), .Q
       (___009___30636));
  nnd2s1 ____09_504398(.DIN1 (__9_____30313), .DIN2 (___009___30634),
       .Q (___009___30635));
  nnd2s1 ____09_504399(.DIN1 (__9_____30297), .DIN2 (___0090__30632),
       .Q (___009___30633));
  or2s1 ____09_504400(.DIN1 (___00____30630), .DIN2 (__9_0___30280), .Q
       (___00_9__30631));
  nnd2s1 _____504401(.DIN1 (__9_____30324), .DIN2 (____9_0__32391), .Q
       (___00____30629));
  and2s1 _____0_504402(.DIN1 (__9_9___30268), .DIN2 (___00____30627),
       .Q (___00____30628));
  nor2s1 _____0_504403(.DIN1 (___00____30625), .DIN2 (__9_0___30276),
       .Q (___00____30626));
  nor2s1 _____0_504404(.DIN1 (________26278), .DIN2 (__9_____30296), .Q
       (___00____30624));
  nor2s1 _____0_504405(.DIN1 (________28456), .DIN2 (__9_9___30269), .Q
       (___00____30623));
  or2s1 _______504406(.DIN1 (___00_9__30621), .DIN2 (__9_0___30275), .Q
       (___00_0__30622));
  nnd2s1 _______504407(.DIN1 (__9_____30328), .DIN2 (___0_0___30748),
       .Q (___00____30620));
  nor2s1 ______504408(.DIN1 (___0__9__30890), .DIN2 (__9_0___30273), .Q
       (___00____30619));
  and2s1 _______504409(.DIN1 (__9_____30258), .DIN2 (___0_____31096),
       .Q (___00____30618));
  nnd2s1 _______504410(.DIN1 (__9_____30256), .DIN2 (________29302), .Q
       (___00____30617));
  nor2s1 ______504411(.DIN1 (__9_____29870), .DIN2 (_________40990), .Q
       (___00____30616));
  nor2s1 _______504412(.DIN1 (__9_____29862), .DIN2 (__9_____30294), .Q
       (___00____30615));
  nnd2s1 _______504413(.DIN1 (_________41363), .DIN2 (_____0__29117),
       .Q (___00____30614));
  or2s1 _______504414(.DIN1 (___00_0__30612), .DIN2 (__9__0__30330), .Q
       (___00____30613));
  nnd2s1 ______504415(.DIN1 (_________40988), .DIN2 (___0_____31156),
       .Q (___00_9__30611));
  nor2s1 ______504416(.DIN1 (___0_____31336), .DIN2 (__9_____30249), .Q
       (___00____30610));
  nor2s1 _______504417(.DIN1 (___00____30608), .DIN2 (__9_____30261),
       .Q (___00____30609));
  nnd2s1 _______504418(.DIN1 (__9_____30298), .DIN2 (___00____30606),
       .Q (___00____30607));
  nor2s1 ____0_504419(.DIN1 (___00____30605), .DIN2 (__9_____30333), .Q
       (___0_____30971));
  xor2s1 ____9__504420(.DIN1 (__9__9__30119), .DIN2 (_________38860),
       .Q (___0_0___31311));
  hi1s1 _______504421(.DIN (___0_____30717), .Q (____0_9__31552));
  nor2s1 _______504422(.DIN1 (________27983), .DIN2 (___00_0__30603),
       .Q (___00____30604));
  nor2s1 ______504423(.DIN1 (________29170), .DIN2 (__9_____30246), .Q
       (___00_9__30602));
  and2s1 _______504424(.DIN1 (__9__0__30254), .DIN2 (___0_____31366),
       .Q (___00____30601));
  nor2s1 _______504425(.DIN1 (________28153), .DIN2 (__9_9___30264), .Q
       (___00____30600));
  nor2s1 _______504426(.DIN1 (___0_0__26112), .DIN2 (__9_____30350), .Q
       (___00____30599));
  nor2s1 ______504427(.DIN1 (________28587), .DIN2 (__9_____30340), .Q
       (___00____30598));
  or2s1 _____9_504428(.DIN1 (____90), .DIN2 (___00____30596), .Q
       (___00____30597));
  nnd2s1 _____9_504429(.DIN1 (__9_____30242), .DIN2 (____9_9__32410),
       .Q (___00____30595));
  nor2s1 _____9_504430(.DIN1 (__9__9__30129), .DIN2 (__9_____30426), .Q
       (___00____30594));
  nor2s1 _____0_504431(.DIN1 (__9__9__30010), .DIN2 (__9_____30311), .Q
       (___00_0__30593));
  xor2s1 _____0_504432(.DIN1 (___0_____40640), .DIN2 (___00____39929),
       .Q (___00_9__30592));
  nnd2s1 _____504433(.DIN1 (___00____30570), .DIN2 (__9_9___30174), .Q
       (___00____30591));
  or2s1 ______504434(.DIN1 (___00____30589), .DIN2 (__9_____30190), .Q
       (___00____30590));
  or2s1 _______504435(.DIN1 (___00____30587), .DIN2 (__9_____30210), .Q
       (___00____30588));
  nor2s1 ______504436(.DIN1 (___9_0__27752), .DIN2 (_________36870), .Q
       (___00____30586));
  or2s1 _______504437(.DIN1 (____9___29003), .DIN2 (___00_0__30603), .Q
       (___00____30585));
  and2s1 _______504438(.DIN1 (__9_____30203), .DIN2 (____9____33393),
       .Q (___00_0__30584));
  nnd2s1 _______504439(.DIN1 (__9_____30221), .DIN2 (__9_____30349), .Q
       (___00_9__30583));
  and2s1 _______504440(.DIN1 (__9_____30219), .DIN2 (___0_____31391),
       .Q (___00____30582));
  and2s1 _______504441(.DIN1 (__9_____30199), .DIN2 (___0_____30654),
       .Q (___00____30581));
  nor2s1 _______504442(.DIN1 (___9_9__29619), .DIN2 (__9_9___30172), .Q
       (___00____30580));
  nnd2s1 _______504443(.DIN1 (__9_____30187), .DIN2 (_________32022),
       .Q (___00____30579));
  nor2s1 _______504444(.DIN1 (__90____29695), .DIN2 (__9_____30214), .Q
       (___00____30578));
  nnd2s1 _______504445(.DIN1 (__9_____30223), .DIN2 (___0__0__30796),
       .Q (___00____30577));
  nor2s1 _______504446(.DIN1 (__999___30539), .DIN2 (___00____30575),
       .Q (___00____30576));
  or2s1 ______504447(.DIN1 (________26392), .DIN2 (__9_____30211), .Q
       (___00_0__30574));
  nor2s1 ______504448(.DIN1 (________27724), .DIN2 (__9_0___30181), .Q
       (___00_9__30573));
  nnd2s1 _______504449(.DIN1 (__9_0___30183), .DIN2 (___0_____30793),
       .Q (___00____30572));
  nor2s1 _____9_504450(.DIN1 (__9_____30007), .DIN2 (___00____30570),
       .Q (___00____30571));
  nnd2s1 _____9_504451(.DIN1 (___00____30568), .DIN2 (__99____30480),
       .Q (___00____30569));
  and2s1 _____504452(.DIN1 (__9_____30209), .DIN2 (________28533), .Q
       (___00____30567));
  nor2s1 _____0_504453(.DIN1 (__9__9__30444), .DIN2 (__9__9__30205), .Q
       (___00____30566));
  and2s1 ______504454(.DIN1 (__9_____30201), .DIN2 (________26358), .Q
       (___00_0__30565));
  nnd2s1 _______504455(.DIN1 (___9____29596), .DIN2 (__9_____30164), .Q
       (___00_9__30564));
  nnd2s1 ______504456(.DIN1 (__9_____30194), .DIN2 (___00____30562), .Q
       (___00____30563));
  and2s1 _______504457(.DIN1 (__9_____30193), .DIN2 (________26240), .Q
       (___00____30561));
  and2s1 _______504458(.DIN1 (__9_____30192), .DIN2 (_____09__31612),
       .Q (___00____30560));
  nor2s1 _______504459(.DIN1 (__9__0__30120), .DIN2 (__9_____30200), .Q
       (___00____30559));
  nor2s1 _______504460(.DIN1 (________28046), .DIN2 (__9_____30293), .Q
       (___00____30558));
  and2s1 _______504461(.DIN1 (__9_____30188), .DIN2 (___00____30556),
       .Q (___00____30557));
  nnd2s1 _______504462(.DIN1 (__9_9___30361), .DIN2 (___0_9__26081), .Q
       (___00_0__30555));
  xnr2s1 ______504463(.DIN1 (_________35084), .DIN2 (_________32024),
       .Q (___0009__30554));
  or2s1 _______504464(.DIN1 (_________32105), .DIN2 (__9_99__30176), .Q
       (___000___30553));
  nnd2s1 _____9_504465(.DIN1 (__9__0__30186), .DIN2 (_________41064),
       .Q (___000___30552));
  nnd2s1 _____0_504466(.DIN1 (__9_____30227), .DIN2 (_________36556),
       .Q (___000___30551));
  nor2s1 _____0_504467(.DIN1 (________27192), .DIN2 (__9_____30224), .Q
       (___000___30550));
  nor2s1 _____504468(.DIN1 (___0__9__40412), .DIN2 (_________35966), .Q
       (___000___30549));
  nor2s1 _______504469(.DIN1 (________29329), .DIN2 (__9_9___30173), .Q
       (___000___30548));
  nnd2s1 ______504470(.DIN1 (__9_9___30171), .DIN2 (___00____30562), .Q
       (___000___30547));
  nnd2s1 _______504471(.DIN1 (__9_____30235), .DIN2 (__9__0__29760), .Q
       (___000___30546));
  or2s1 _______504472(.DIN1 (_________33549), .DIN2 (__9_____30202), .Q
       (___0000__30545));
  nor2s1 ______504473(.DIN1 (___099), .DIN2 (_________35966), .Q
       (__9999));
  nor2s1 _______504474(.DIN1 (__999___30543), .DIN2 (__9_9___30170), .Q
       (__999___30544));
  nor2s1 _______504475(.DIN1 (________27278), .DIN2 (__9__9__30168), .Q
       (__999___30542));
  nnd2s1 _______504476(.DIN1 (__9_____30230), .DIN2 (________27527), .Q
       (__999___30541));
  nor2s1 _______504477(.DIN1 (__999___30539), .DIN2 (__9_____30217), .Q
       (__999___30540));
  and2s1 _______504478(.DIN1 (__999_), .DIN2 (__9990), .Q
       (__999___30538));
  nor2s1 _______504479(.DIN1 (__9_____29827), .DIN2 (__99____30536), .Q
       (__99_9__30537));
  nnd2s1 _______504480(.DIN1 (__9__0__30226), .DIN2 (inData[22]), .Q
       (__99____30535));
  and2s1 ______504481(.DIN1 (__9_0___30178), .DIN2 (__99____30533), .Q
       (__99____30534));
  nnd2s1 _______504482(.DIN1 (__9_09__30185), .DIN2 (__9__9__30300), .Q
       (__99____30532));
  nor2s1 _______504483(.DIN1 (_________32001), .DIN2 (______0__40992),
       .Q (__99____30531));
  nor2s1 _______504484(.DIN1 (__9_____30380), .DIN2 (__9_____30197), .Q
       (__99____30530));
  nnd2s1 _______504485(.DIN1 (_________40994), .DIN2 (________27151),
       .Q (__99____30529));
  nor2s1 _______504486(.DIN1 (_________32748), .DIN2 (__9_____30220),
       .Q (__99_0__30528));
  nnd2s1 _______504487(.DIN1 (__9_____30165), .DIN2 (___00___27832), .Q
       (__99_9__30527));
  or2s1 _______504488(.DIN1 (__99____30525), .DIN2 (_________40996), .Q
       (__99____30526));
  nor2s1 _______504489(.DIN1 (__9_____30222), .DIN2 (__9__9__30233), .Q
       (__99____30524));
  or2s1 _____0_504490(.DIN1 (___0____28820), .DIN2 (__99____30522), .Q
       (__99____30523));
  nnd2s1 ______504491(.DIN1 (________29522), .DIN2 (__9_____30236), .Q
       (__99____30521));
  nnd2s1 _______504492(.DIN1 (__9_____30207), .DIN2 (___0_____30783),
       .Q (__99____30520));
  nnd2s1 _______504493(.DIN1 (__99____30515), .DIN2 (__9__0__30159), .Q
       (__99____30519));
  nor2s1 _______504494(.DIN1 (__990___30461), .DIN2 (__9_____30238), .Q
       (__99_0__30518));
  nor2s1 _______504495(.DIN1 (________26764), .DIN2 (__9_____30237), .Q
       (__99_9__30517));
  and2s1 _______504496(.DIN1 (__9__9__30195), .DIN2 (__99____30516), .Q
       (___0__9__30898));
  nnd2s1 _______504497(.DIN1 (__99____30515), .DIN2 (__9_____30160), .Q
       (___0_0___30840));
  nor2s1 _______504498(.DIN1 (__99____30514), .DIN2 (_________36870),
       .Q (___0_____30708));
  nnd2s1 _______504499(.DIN1 (__9_0___30180), .DIN2 (__99____30513), .Q
       (___0_____30937));
  nor2s1 _______504500(.DIN1 (____9___27560), .DIN2 (__9_____30232), .Q
       (__99____30512));
  nor2s1 ______504501(.DIN1 (________27939), .DIN2 (__9_____30069), .Q
       (__99____30511));
  nnd2s1 ____9__504502(.DIN1 (__9_____30154), .DIN2 (________25514), .Q
       (__99____30510));
  nor2s1 ____9__504503(.DIN1 (__99_9__30508), .DIN2 (__9_____30152), .Q
       (__99_0__30509));
  nnd2s1 ____9__504504(.DIN1 (__9_____30136), .DIN2 (__99____30506), .Q
       (__99____30507));
  or2s1 ____9__504505(.DIN1 (________28097), .DIN2 (__9_____30151), .Q
       (__99____30505));
  nnd2s1 ____9__504506(.DIN1 (___090__26132), .DIN2 (__9_____30125), .Q
       (__99____30504));
  nnd2s1 ____9__504507(.DIN1 (__9_____30132), .DIN2 (___0____28797), .Q
       (__99____30503));
  or2s1 ____9__504508(.DIN1 (__99____30501), .DIN2 (__9_____30148), .Q
       (__99____30502));
  nnd2s1 ____0__504509(.DIN1 (________29022), .DIN2 (__9_____30144), .Q
       (__99____30500));
  nnd2s1 ____0__504510(.DIN1 (__9__0__30140), .DIN2 (___0_____30752),
       .Q (__99_0__30499));
  nor2s1 ____0__504511(.DIN1 (_________33143), .DIN2 (__9_____30138),
       .Q (__99_9__30498));
  nor2s1 ____0__504512(.DIN1 (____0___29102), .DIN2 (__9_____30146), .Q
       (__99____30497));
  nor2s1 ____09_504513(.DIN1 (_________31809), .DIN2 (__9__9__30139),
       .Q (__99____30496));
  nnd2s1 _____504514(.DIN1 (__9_____30131), .DIN2 (___9____27778), .Q
       (__99____30495));
  and2s1 _______504515(.DIN1 (__9_____30134), .DIN2 (____9_0__32391),
       .Q (__99____30494));
  nor2s1 _______504516(.DIN1 (__99____30492), .DIN2 (__9_____30141), .Q
       (__99____30493));
  and2s1 _______504517(.DIN1 (__9_____30123), .DIN2 (__99____30490), .Q
       (__99____30491));
  nnd2s1 _______504518(.DIN1 (__9_____30143), .DIN2 (__9_9___30270), .Q
       (__99_0__30489));
  or2s1 _______504519(.DIN1 (__99____30487), .DIN2 (__9_____30133), .Q
       (__99_9__30488));
  nor2s1 _______504520(.DIN1 (__99____30485), .DIN2 (__9_____30122), .Q
       (__99____30486));
  nor2s1 _______504521(.DIN1 (____0___28296), .DIN2 (__9_____30127), .Q
       (__99____30484));
  or2s1 _______504522(.DIN1 (__9__9__29935), .DIN2 (__99____30482), .Q
       (__99____30483));
  nnd2s1 _______504523(.DIN1 (__9_____30044), .DIN2 (__99____30480), .Q
       (__99____30481));
  nor2s1 _______504524(.DIN1 (inData[15]), .DIN2 (_________36288), .Q
       (__99_0__30479));
  nor2s1 _______504525(.DIN1 (__9__9__29751), .DIN2 (__9_____30121), .Q
       (__99_9__30478));
  nor2s1 _______504526(.DIN1 (inData[16]), .DIN2 (_________36288), .Q
       (__99____30477));
  nor2s1 ______504527(.DIN1 (inData[20]), .DIN2 (____9_9__36114), .Q
       (__99____30476));
  nor2s1 _______504528(.DIN1 (________28250), .DIN2 (__9_____30050), .Q
       (__99____30475));
  nnd2s1 _______504529(.DIN1 (__9__9__30110), .DIN2 (__99____30473), .Q
       (__99____30474));
  nnd2s1 _______504530(.DIN1 (__9_____30043), .DIN2 (___0____28811), .Q
       (__99____30472));
  nnd2s1 ______504531(.DIN1 (__9_____30396), .DIN2 (_________41146), .Q
       (__99____30471));
  nnd2s1 _______504532(.DIN1 (__9__0__30102), .DIN2 (__99_0__30469), .Q
       (__99____30470));
  nnd2s1 _______504533(.DIN1 (__9__9__30101), .DIN2 (__99____30468), .Q
       (__99_9));
  nnd2s1 _______504534(.DIN1 (__9_____30100), .DIN2 (________27965), .Q
       (__99____30467));
  and2s1 _______504535(.DIN1 (__9_____30099), .DIN2 (__99____30465), .Q
       (__99____30466));
  or2s1 _______504536(.DIN1 (__99____30463), .DIN2 (__9_____30017), .Q
       (__99____30464));
  nnd2s1 ______504537(.DIN1 (__9_____30009), .DIN2 (__99__), .Q
       (__99____30462));
  nor2s1 _______504538(.DIN1 (___9____29608), .DIN2 (__9_0___30088), .Q
       (__99_0));
  nor2s1 ______504539(.DIN1 (__990___30461), .DIN2 (__9_____30072), .Q
       (__9909));
  nor2s1 ______504540(.DIN1 (__9_____30054), .DIN2 (__9_____30094), .Q
       (__990___30460));
  and2s1 _______504541(.DIN1 (__9_0___30090), .DIN2 (__9990), .Q
       (__990___30459));
  nnd2s1 _______504542(.DIN1 (__9_0___30089), .DIN2 (__9_____30019), .Q
       (__990___30458));
  and2s1 _______504543(.DIN1 (__90____29712), .DIN2 (__9_____30407), .Q
       (__990___30457));
  nnd2s1 _______504544(.DIN1 (__9_0___30084), .DIN2 (__9_____30423), .Q
       (__990___30456));
  nnd2s1 _______504545(.DIN1 (__9_00__30083), .DIN2 (________28622), .Q
       (__990___30455));
  nnd2s1 _______504546(.DIN1 (__9_99__30082), .DIN2 (__9900), .Q
       (__990_));
  nnd2s1 _______504547(.DIN1 (__9_9___30081), .DIN2 (________28495), .Q
       (__9_99__30454));
  nor2s1 ______504548(.DIN1 (_____0__28148), .DIN2 (__9_____30161), .Q
       (__9_9___30453));
  and2s1 _____504549(.DIN1 (__9__0__30064), .DIN2 (__9_9___30451), .Q
       (__9_9___30452));
  or2s1 _____9_504550(.DIN1 (__9_9___30449), .DIN2 (__9_0___30087), .Q
       (__9_9___30450));
  nor2s1 _____9_504551(.DIN1 (__999___30539), .DIN2 (__9_9___30077), .Q
       (__9_9___30448));
  nor2s1 _____0_504552(.DIN1 (________28879), .DIN2 (_________41000),
       .Q (__9_9___30447));
  nor2s1 _____0_504553(.DIN1 (________28855), .DIN2 (__9_____30021), .Q
       (__9_9___30446));
  nor2s1 _____504554(.DIN1 (__9__9__30444), .DIN2 (__9_____30040), .Q
       (__9_90__30445));
  nor2s1 _______504555(.DIN1 (____0___26503), .DIN2 (__9_____30116), .Q
       (__9_____30443));
  and2s1 _______504556(.DIN1 (_________36288), .DIN2 (________27408),
       .Q (__9_____30442));
  and2s1 _______504557(.DIN1 (_____9___41008), .DIN2 (__9_9___30270),
       .Q (__9_____30440));
  or2s1 _______504558(.DIN1 (__9__0__30438), .DIN2 (_____9___41004), .Q
       (__9_____30439));
  nnd2s1 _____0_504559(.DIN1 (__9_____30124), .DIN2 (__90____29655), .Q
       (___0_0___30645));
  xor2s1 ____9__504560(.DIN1 (__9_____29973), .DIN2 (___9_0___39624),
       .Q (___0_____30717));
  hi1s1 _______504561(.DIN (__9__9__30437), .Q (___0_____30886));
  and2s1 _______504562(.DIN1 (___0____28801), .DIN2 (__9__0__30048), .Q
       (__9_____30436));
  and2s1 _______504563(.DIN1 (__9_____30097), .DIN2 (___0__9__30851),
       .Q (__9_____30435));
  nnd2s1 ______504564(.DIN1 (__9_____30060), .DIN2 (_____0__28530), .Q
       (__9_____30434));
  nor2s1 _______504565(.DIN1 (__9_____30432), .DIN2 (__9_____30066), .Q
       (__9_____30433));
  nor2s1 _______504566(.DIN1 (__9_____30430), .DIN2 (__9_____30065), .Q
       (__9_____30431));
  nor2s1 _______504567(.DIN1 (___9____29622), .DIN2 (__9_____30059), .Q
       (__9__0__30429));
  hi1s1 _______504568(.DIN (__9_____30426), .Q (__9_____30427));
  nor2s1 _______504569(.DIN1 (___0__0__30872), .DIN2 (__9_____30157),
       .Q (__9_____30425));
  nnd2s1 _______504570(.DIN1 (__9_____30042), .DIN2 (__9_____30423), .Q
       (__9_____30424));
  nor2s1 ______504571(.DIN1 (___9____27803), .DIN2 (__9_____30041), .Q
       (__9_____30422));
  nor2s1 ______504572(.DIN1 (inData[14]), .DIN2 (_________36288), .Q
       (__9_____30421));
  nor2s1 _______504573(.DIN1 (__9__9__30419), .DIN2 (__9_____30107), .Q
       (__9__0__30420));
  nor2s1 _______504574(.DIN1 (__9_____30417), .DIN2 (__9_____30416), .Q
       (__9_____30418));
  nnd2s1 _____504575(.DIN1 (__9_____30012), .DIN2 (_____9__29126), .Q
       (__9_____30415));
  nor2s1 _____9_504576(.DIN1 (________29245), .DIN2 (__9_____30008), .Q
       (__9_____30414));
  nnd2s1 _____9_504577(.DIN1 (__9__0__30038), .DIN2 (__9_0___29729), .Q
       (__9_____30413));
  nor2s1 _____0_504578(.DIN1 (_________41128), .DIN2 (__9__9__30393),
       .Q (__9_____30412));
  nor2s1 _____0_504579(.DIN1 (__9_____30204), .DIN2 (__9_____30045), .Q
       (__9__0__30411));
  nnd2s1 ______504580(.DIN1 (__9_9___30078), .DIN2 (___0_____30783), .Q
       (__9__9__30410));
  nnd2s1 _______504581(.DIN1 (__9__9__30020), .DIN2 (________28954), .Q
       (__9_____30409));
  or2s1 _______504582(.DIN1 (__9_____29827), .DIN2 (__9_____30407), .Q
       (__9_____30408));
  nor2s1 _______504583(.DIN1 (__9_0___29809), .DIN2 (__9_____30032), .Q
       (__9_____30406));
  nnd2s1 _______504584(.DIN1 (__9_0___30091), .DIN2 (__9900), .Q
       (__9_____30405));
  nnd2s1 _______504585(.DIN1 (__9_____30025), .DIN2 (________27151), .Q
       (__9_____30404));
  nor2s1 ______504586(.DIN1 (__9_0___30182), .DIN2 (__9_____30037), .Q
       (__9__0__30403));
  nor2s1 _______504587(.DIN1 (__9_____30401), .DIN2 (__9_____30398), .Q
       (__9__9__30402));
  nnd2s1 _______504588(.DIN1 (__9_____30398), .DIN2 (________29297), .Q
       (__9_____30399));
  nnd2s1 _______504589(.DIN1 (__9_____30396), .DIN2 (________28169), .Q
       (__9_____30397));
  nor2s1 ______504590(.DIN1 (__9__0__30394), .DIN2 (__9__9__30393), .Q
       (__9_____30395));
  nor2s1 _______504591(.DIN1 (__9_____29773), .DIN2 (__9_____30033), .Q
       (__9_____30392));
  nnd2s1 _______504592(.DIN1 (__9_____30034), .DIN2 (________28122), .Q
       (__9_____30391));
  nnd2s1 _______504593(.DIN1 (__9_____30013), .DIN2 (___09____31469),
       .Q (__9_____30390));
  nnd2s1 _______504594(.DIN1 (__9_90__30074), .DIN2 (___0____27011), .Q
       (__9_____30389));
  nor2s1 ______504595(.DIN1 (________27582), .DIN2 (__9__0__30011), .Q
       (__9_____30388));
  nnd2s1 _____9_504596(.DIN1 (__9_____30014), .DIN2 (___0_____30783),
       .Q (__9_____30387));
  nnd2s1 _____504597(.DIN1 (__9_____30385), .DIN2 (_____9__27471), .Q
       (__9_____30386));
  or2s1 _____0_504598(.DIN1 (___0_____31242), .DIN2 (__9_9___30075), .Q
       (__9__9__30384));
  nor2s1 _____0_504599(.DIN1 (__90____29664), .DIN2 (__9_____30006), .Q
       (__9_____30383));
  or2s1 _____0_504600(.DIN1 (___0__9__31347), .DIN2 (__9_____30015), .Q
       (__9_____30382));
  nor2s1 _______504601(.DIN1 (__9_____30380), .DIN2 (__9_9___30076), .Q
       (__9_____30381));
  nor2s1 _______504602(.DIN1 (___0_9__26966), .DIN2 (__9_00__30366), .Q
       (__9_____30379));
  nor2s1 ______504603(.DIN1 (___0_____30961), .DIN2 (__9_0___30001), .Q
       (__9_____30378));
  or2s1 _______504604(.DIN1 (____0___27925), .DIN2 (__9_____30004), .Q
       (__9_____30377));
  nor2s1 _____0_504605(.DIN1 (_____9___41006), .DIN2 (_____0__29387),
       .Q (__9_____30376));
  nor2s1 _______504606(.DIN1 (___0_____30956), .DIN2 (__9_____30052),
       .Q (__9__0__30375));
  nor2s1 _______504607(.DIN1 (__9_0___30373), .DIN2 (__9_____30005), .Q
       (__9_09__30374));
  nor2s1 ______504608(.DIN1 (__9_____30208), .DIN2 (__9_____30055), .Q
       (__9_0___30372));
  or2s1 _______504609(.DIN1 (____9___27651), .DIN2 (_____9___41006), .Q
       (__9_0___30371));
  nnd2s1 _______504610(.DIN1 (____9___29189), .DIN2 (__9_____30057), .Q
       (__9_0___30370));
  nor2s1 _______504611(.DIN1 (________29149), .DIN2 (__9_0___29999), .Q
       (__9_0___30369));
  nnd2s1 _______504612(.DIN1 (__9_09__30002), .DIN2 (_________34243),
       .Q (__9_0___30368));
  or2s1 _______504613(.DIN1 (___0_00__30642), .DIN2 (__9_____30061), .Q
       (__9_0___30367));
  nor2s1 ______504614(.DIN1 (___0900), .DIN2 (__9_____30023), .Q
       (___0_____30803));
  nnd2s1 ______504615(.DIN1 (__9_09__30092), .DIN2 (__9__0__29878), .Q
       (___0_____30816));
  nor2s1 ____9__504616(.DIN1 (____9___29547), .DIN2 (__9_00__30366), .Q
       (___0_9___30734));
  nnd2s1 ____9__504617(.DIN1 (_____90__41002), .DIN2 (___0____27892),
       .Q (___0_09__30749));
  dffacs1 ____________________________________9_504618(.CLRB (reset),
       .CLK (clk), .DIN (__9_____30156), .Q (_________9_));
  dffacs1 _______________________________________504619(.CLRB (reset),
       .CLK (clk), .DIN (__9_____30155), .Q (______________22103));
  dffacs1 _________________________________________0_____504620(.CLRB
       (reset), .CLK (clk), .DIN (__9_____30113), .QN (___0_0___40566));
  dffacs1 _______________________________________504621(.CLRB (reset),
       .CLK (clk), .DIN (__9_____30153), .Q (______________22106));
  dffacs1 _________________________________________0_____504622(.CLRB
       (reset), .CLK (clk), .DIN (__9_____30018), .Q (___0_____40572));
  dffacs1 __________________504623(.CLRB (reset), .CLK (clk), .DIN
       (__9__0__30111), .QN (_______________22072));
  nnd2s1 _______504624(.DIN1 (__9_9___30364), .DIN2 (________23121), .Q
       (__9_9___30365));
  or2s1 _______504625(.DIN1 (__9_9___30362), .DIN2 (__9_0___29902), .Q
       (__9_9___30363));
  nor2s1 ____9__504626(.DIN1 (__9_9___30360), .DIN2 (__9_9___29987), .Q
       (__9_9___30361));
  nor2s1 ____9__504627(.DIN1 (_____0__26428), .DIN2 (__9_____29982), .Q
       (__9_9___30359));
  nor2s1 _____0_504628(.DIN1 (________29521), .DIN2 (__9_____29978), .Q
       (__9_9___30358));
  or2s1 _______504629(.DIN1 (______9__32949), .DIN2 (_________36082),
       .Q (__9_90__30357));
  nnd2s1 ______504630(.DIN1 (__9_____29983), .DIN2 (________27152), .Q
       (__9__9__30356));
  or2s1 _______504631(.DIN1 (___0_09__31127), .DIN2 (__9_____29977), .Q
       (__9_____30355));
  and2s1 _______504632(.DIN1 (__9_____29980), .DIN2 (_________33137),
       .Q (__9_____30354));
  and2s1 _____0_504633(.DIN1 (_________36082), .DIN2 (______9__32949),
       .Q (__9_____30353));
  nor2s1 _______504634(.DIN1 (________28630), .DIN2 (__9_____29930), .Q
       (__9_____30352));
  nnd2s1 _______504635(.DIN1 (__9_____29928), .DIN2 (________28242), .Q
       (__9_____30351));
  nnd2s1 _______504636(.DIN1 (__9_____29962), .DIN2 (__9_____30349), .Q
       (__9_____30350));
  nor2s1 _______504637(.DIN1 (__9_____29858), .DIN2 (__9_____29864), .Q
       (__9_____30348));
  nor2s1 _______504638(.DIN1 (__9_____29857), .DIN2 (__9_____29961), .Q
       (__9__0__30347));
  nnd2s1 _______504639(.DIN1 (__9_____29958), .DIN2 (__90____29666), .Q
       (__9_____30346));
  nor2s1 _______504640(.DIN1 (__9_____29875), .DIN2 (____00__29466), .Q
       (__9_____30345));
  nor2s1 _______504641(.DIN1 (___0_____30821), .DIN2 (__9_____29943),
       .Q (__9_____30344));
  nnd2s1 ______504642(.DIN1 (__9_____29954), .DIN2 (___0____27016), .Q
       (__9_____30343));
  nnd2s1 _______504643(.DIN1 (__9_9___29988), .DIN2 (________29112), .Q
       (__9_____30342));
  nnd2s1 _______504644(.DIN1 (__9_____29929), .DIN2 (________26151), .Q
       (__9_____30341));
  or2s1 ______504645(.DIN1 (__9_____30339), .DIN2 (__9_____29947), .Q
       (__9_____30340));
  or2s1 _______504646(.DIN1 (__9__9__30337), .DIN2 (__9_9___29890), .Q
       (__9__0__30338));
  nor2s1 _______504647(.DIN1 (__9_____30335), .DIN2 (_____0___41014),
       .Q (__9_____30336));
  nnd2s1 _______504648(.DIN1 (__9__9__29955), .DIN2 (________28029), .Q
       (__9_____30334));
  nnd2s1 _______504649(.DIN1 (__9_____29939), .DIN2 (__9_____30332), .Q
       (__9_____30333));
  and2s1 _______504650(.DIN1 (__9_____29933), .DIN2 (_________33934),
       .Q (__9_____30331));
  nnd2s1 _______504651(.DIN1 (__9_____29931), .DIN2 (_____0__29213), .Q
       (__9__0__30330));
  and2s1 _____9_504652(.DIN1 (__9_____29853), .DIN2 (_________41178),
       .Q (__9__9__30329));
  nnd2s1 _____9_504653(.DIN1 (__9_____29927), .DIN2 (__9900), .Q
       (__9_____30328));
  nor2s1 _____9_504654(.DIN1 (_____9___41301), .DIN2 (__9_____29874),
       .Q (__9_____30327));
  nnd2s1 _____504655(.DIN1 (__9_____29934), .DIN2 (__9_____30325), .Q
       (__9_____30326));
  nor2s1 _____0_504656(.DIN1 (________26733), .DIN2 (__9_____29922), .Q
       (__9_____30324));
  nnd2s1 _____0_504657(.DIN1 (__9_____29920), .DIN2 (__9_____30322), .Q
       (__9_____30323));
  nor2s1 _____0_504658(.DIN1 (________29238), .DIN2 (__9_____29919), .Q
       (__9_____30321));
  nnd2s1 ______504659(.DIN1 (__9_____29918), .DIN2 (__9__9__30319), .Q
       (__9__0__30320));
  nnd2s1 _______504660(.DIN1 (__9__9__29840), .DIN2 (____99__29096), .Q
       (__9_____30318));
  nnd2s1 _______504661(.DIN1 (________28504), .DIN2 (__9_____30295), .Q
       (__9_____30317));
  nor2s1 _______504662(.DIN1 (_____9__28946), .DIN2 (__9_____29836), .Q
       (__9_____30316));
  nnd2s1 _______504663(.DIN1 (__9_____29912), .DIN2 (__9_____30314), .Q
       (__9_____30315));
  nor2s1 _______504664(.DIN1 (__9_____30312), .DIN2 (__9_____29910), .Q
       (__9_____30313));
  nnd2s1 _______504665(.DIN1 (________29408), .DIN2 (__9_____30117), .Q
       (__9_____30311));
  nor2s1 _______504666(.DIN1 (__9__0__30291), .DIN2 (__9_____29909), .Q
       (__9__0__30310));
  nor2s1 _______504667(.DIN1 (inData[31]), .DIN2 (____0____33493), .Q
       (__9__9__30309));
  nnd2s1 _______504668(.DIN1 (__9_09__29905), .DIN2 (__9_____29845), .Q
       (__9_____30308));
  nnd2s1 ______504669(.DIN1 (__9_____29963), .DIN2 (__9_____30306), .Q
       (__9_____30307));
  nnd2s1 _______504670(.DIN1 (__9_____29967), .DIN2 (_____9__27471), .Q
       (__9_____30305));
  or2s1 _______504671(.DIN1 (__9_____30303), .DIN2 (__9_0___29898), .Q
       (__9_____30304));
  nnd2s1 _______504672(.DIN1 (__9_00__29896), .DIN2 (__9_9___30451), .Q
       (__9_____30302));
  nor2s1 _______504673(.DIN1 (____0___29202), .DIN2 (__9_____29942), .Q
       (__9_____30301));
  nnd2s1 _______504674(.DIN1 (__9_9___29891), .DIN2 (________29389), .Q
       (__9_____30299));
  nor2s1 _______504675(.DIN1 (___9____29580), .DIN2 (__9_0___29903), .Q
       (__9_____30298));
  nor2s1 _______504676(.DIN1 (___00____30625), .DIN2 (__9__0__29850),
       .Q (__9_____30297));
  nnd2s1 _______504677(.DIN1 (__9_____30295), .DIN2 (________28267), .Q
       (__9_____30296));
  nor2s1 _______504678(.DIN1 (_____9__25947), .DIN2 (__9_____29838), .Q
       (__9_____30294));
  nnd2s1 _______504679(.DIN1 (__9_____29907), .DIN2 (________28523), .Q
       (__9_____30293));
  nor2s1 _______504680(.DIN1 (__9__0__30291), .DIN2 (__9_____29880), .Q
       (__9_____30292));
  nor2s1 _______504681(.DIN1 (____90__28005), .DIN2 (_____00__41012),
       .Q (__9__9__30290));
  nnd2s1 _______504682(.DIN1 (__9_____29825), .DIN2 (______0__41032),
       .Q (__9_____30289));
  nor2s1 _______504683(.DIN1 (__9_____30401), .DIN2 (__9_____29879), .Q
       (__9_____30288));
  nor2s1 _______504684(.DIN1 (_____0__29037), .DIN2 (__9_____29924), .Q
       (__9_____30287));
  nnd2s1 _____9_504685(.DIN1 (__9__0__29906), .DIN2 (__9_____30285), .Q
       (__9_____30286));
  nnd2s1 _____9_504686(.DIN1 (__9_____29951), .DIN2 (________29357), .Q
       (__9_____30284));
  and2s1 _____9_504687(.DIN1 (__9_____29826), .DIN2 (___0_____30943),
       .Q (__9_____30283));
  nnd2s1 _____9_504688(.DIN1 (__9_____29822), .DIN2 (__9_09__30281), .Q
       (__9__0__30282));
  nnd2s1 _____504689(.DIN1 (__9_____29842), .DIN2 (________29439), .Q
       (__9_0___30280));
  nor2s1 _____504690(.DIN1 (________22485), .DIN2 (__9_____29869), .Q
       (__9_0___30279));
  nor2s1 _____0_504691(.DIN1 (____9___28007), .DIN2 (__9_____29861), .Q
       (__9_0___30278));
  nor2s1 _____0_504692(.DIN1 (________29514), .DIN2 (__9_____29848), .Q
       (__9_0___30277));
  or2s1 _______504693(.DIN1 (___0_____30977), .DIN2 (__9_____29837), .Q
       (__9_0___30276));
  or2s1 _______504694(.DIN1 (__9_0___30274), .DIN2 (__9_____29969), .Q
       (__9_0___30275));
  nor2s1 _______504695(.DIN1 (__9_00__30272), .DIN2 (__9_0___29900), .Q
       (__9_0___30273));
  nnd2s1 _______504696(.DIN1 (__9_____29854), .DIN2 (__9_9___30270), .Q
       (__9_99__30271));
  nnd2s1 _______504697(.DIN1 (__9_____29937), .DIN2 (____90__28285), .Q
       (__9_9___30269));
  and2s1 ______504698(.DIN1 (__9__0__29868), .DIN2 (__9_9___30267), .Q
       (__9_9___30268));
  nor2s1 _______504699(.DIN1 (________27243), .DIN2 (__9__9__29867), .Q
       (__9_9___30266));
  nor2s1 _______504700(.DIN1 (_________31836), .DIN2 (__9_____29846),
       .Q (__9_9___30265));
  nnd2s1 ______504701(.DIN1 (__9_____29829), .DIN2 (__9__9__30063), .Q
       (__9_9___30264));
  nor2s1 _______504702(.DIN1 (__9__9__30262), .DIN2 (__9_____29871), .Q
       (__9_90__30263));
  or2s1 _______504703(.DIN1 (__9_____30260), .DIN2 (__9_9___29894), .Q
       (__9_____30261));
  nnd2s1 _______504704(.DIN1 (__9_____30259), .DIN2 (__9_____29856), .Q
       (_________32834));
  nnd2s1 _______504705(.DIN1 (__9__9__29965), .DIN2 (________29399), .Q
       (___0_____30690));
  nor2s1 _______504706(.DIN1 (________22724), .DIN2 (__9_____29960), .Q
       (___0_____30686));
  xor2s1 ____9__504707(.DIN1 (__90____29715), .DIN2 (__9_____29851), .Q
       (__9__9__30437));
  xor2s1 ____9_504708(.DIN1 (__90____29714), .DIN2 (___9_____39312), .Q
       (__99____30515));
  dffacs1 ________________________________________________504709(.CLRB
       (reset), .CLK (clk), .DIN (__9_____29950), .QN
       (________________________________________________________________));
  nor2s1 _______504710(.DIN1 (__9_0___30274), .DIN2 (__9_____29923), .Q
       (__9_____30258));
  nnd2s1 _______504711(.DIN1 (__9_____29913), .DIN2 (______9__34050),
       .Q (__9_____30257));
  nnd2s1 ______504712(.DIN1 (__9_____29948), .DIN2 (__9_____30255), .Q
       (__9_____30256));
  and2s1 _______504713(.DIN1 (__9_____30295), .DIN2 (_________41148),
       .Q (__9__0__30254));
  nor2s1 ______504714(.DIN1 (________29289), .DIN2 (__9_____29828), .Q
       (__9__9__30253));
  nnd2s1 _______504715(.DIN1 (__9_____29816), .DIN2 (_____0__28581), .Q
       (__9_____30252));
  or2s1 _______504716(.DIN1 (___09___28829), .DIN2 (__9_____30250), .Q
       (__9_____30251));
  nor2s1 _____504717(.DIN1 (_________31870), .DIN2 (__9_0___29810), .Q
       (__9_____30249));
  nor2s1 _____9_504718(.DIN1 (_____0__27552), .DIN2 (__9__9__29823), .Q
       (__9_____30248));
  nnd2s1 _____9_504719(.DIN1 (__9_____29820), .DIN2 (__9_0___29808), .Q
       (__9_____30247));
  nnd2s1 _____9_504720(.DIN1 (__9_____29917), .DIN2 (___0____26989), .Q
       (__9_____30246));
  nor2s1 _____9_504721(.DIN1 (_________31942), .DIN2 (__9_____29819),
       .Q (__9_____30245));
  nnd2s1 _____9_504722(.DIN1 (__9_____29821), .DIN2 (___9____25975), .Q
       (__9__0__30244));
  nnd2s1 _____0_504723(.DIN1 (__9_09__29813), .DIN2 (________28633), .Q
       (__9__9__30243));
  nnd2s1 _____504724(.DIN1 (__9_____29882), .DIN2 (__9_____30241), .Q
       (__9_____30242));
  and2s1 _______504725(.DIN1 (__9_____29944), .DIN2 (__9_____30239), .Q
       (__9_____30240));
  nnd2s1 ______504726(.DIN1 (__9_0___29806), .DIN2 (________29379), .Q
       (__9_____30238));
  nnd2s1 ______504727(.DIN1 (__9_0___29807), .DIN2 (__9_____29843), .Q
       (__9_____30237));
  nor2s1 ____90_504728(.DIN1 (___900__28646), .DIN2 (__9_9___29803), .Q
       (__9_____30236));
  and2s1 _____9_504729(.DIN1 (__9_____29741), .DIN2 (__9__0__30234), .Q
       (__9_____30235));
  nnd2s1 _____504730(.DIN1 (__9_____29746), .DIN2 (________28152), .Q
       (__9__9__30233));
  nor2s1 ______504731(.DIN1 (__9_____29827), .DIN2 (__9_____29753), .Q
       (__9_____30231));
  or2s1 _______504732(.DIN1 (__999___30539), .DIN2 (__9_____30229), .Q
       (__9_____30230));
  nnd2s1 _______504733(.DIN1 (____9_0__37080), .DIN2 (inData[13]), .Q
       (__9_____30228));
  nor2s1 ______504734(.DIN1 (___09___22360), .DIN2 (_________36618), .Q
       (__9_____30227));
  nor2s1 _______504735(.DIN1 (__9__9__30225), .DIN2 (__9_9_), .Q
       (__9__0__30226));
  nnd2s1 _______504736(.DIN1 (__9_____29738), .DIN2 (________27611), .Q
       (__9_____30224));
  nor2s1 _______504737(.DIN1 (__9_____30222), .DIN2 (__9__9__29759), .Q
       (__9_____30223));
  nor2s1 _____9_504738(.DIN1 (_________41066), .DIN2 (__9_____29794),
       .Q (__9_____30221));
  or2s1 _____9_504739(.DIN1 (___0_9___31015), .DIN2 (__9_____29793), .Q
       (__9_____30220));
  and2s1 _____9_504740(.DIN1 (__9_____29791), .DIN2 (___0_____30888),
       .Q (__9_____30219));
  nnd2s1 _____0_504741(.DIN1 (__9_____29765), .DIN2 (_____9__27471), .Q
       (__9_____30218));
  and2s1 _______504742(.DIN1 (__9__9__29788), .DIN2 (__9__0__30216), .Q
       (__9_____30217));
  nnd2s1 _______504743(.DIN1 (__9_____29785), .DIN2 (___0_0___30748),
       .Q (__9__9__30215));
  nor2s1 ______504744(.DIN1 (__999___30539), .DIN2 (__9_____29833), .Q
       (__9_____30214));
  nnd2s1 _______504745(.DIN1 (__9_____29782), .DIN2 (________29084), .Q
       (__9_____30213));
  nor2s1 _______504746(.DIN1 (________23522), .DIN2 (____9_0__37080),
       .Q (__9_____30212));
  nnd2s1 _______504747(.DIN1 (__9099), .DIN2 (__9_____29771), .Q
       (__9_____30211));
  or2s1 _______504748(.DIN1 (___0_____30956), .DIN2 (__9_____29768), .Q
       (__9_____30210));
  nor2s1 ______504749(.DIN1 (__9_____30208), .DIN2 (__9_____29772), .Q
       (__9_____30209));
  nnd2s1 _______504750(.DIN1 (__9__0__29770), .DIN2 (__9__0__30206), .Q
       (__9_____30207));
  or2s1 _______504751(.DIN1 (__9_____30204), .DIN2 (__9__9__29769), .Q
       (__9__9__30205));
  nor2s1 _______504752(.DIN1 (___0_____31324), .DIN2 (__9_____29795),
       .Q (__9_____30203));
  or2s1 _______504753(.DIN1 (___0_____31194), .DIN2 (__9_____29747), .Q
       (__9_____30202));
  and2s1 _______504754(.DIN1 (__9_____29749), .DIN2 (_________41321),
       .Q (__9_____30201));
  or2s1 _______504755(.DIN1 (__9_0___29897), .DIN2 (__9_____29736), .Q
       (__9_____30200));
  nor2s1 _______504756(.DIN1 (__9_____30198), .DIN2 (_________41026),
       .Q (__9_____30199));
  nnd2s1 ______504757(.DIN1 (__9_____29734), .DIN2 (__9__0__30196), .Q
       (__9_____30197));
  nor2s1 _______504758(.DIN1 (________29233), .DIN2 (__9_____29763), .Q
       (__9__9__30195));
  nor2s1 _______504759(.DIN1 (__9_____29777), .DIN2 (__9_____29762), .Q
       (__9_____30194));
  nor2s1 _______504760(.DIN1 (___0990__31494), .DIN2 (__9_____29761),
       .Q (__9_____30193));
  and2s1 ______504761(.DIN1 (__9_____29730), .DIN2 (___0__0__30796), .Q
       (__9_____30192));
  nor2s1 _____504762(.DIN1 (___0_____40486), .DIN2 (____9_0__37080), .Q
       (__9_____30191));
  nnd2s1 _____0_504763(.DIN1 (__9_____30189), .DIN2 (__9_____29755), .Q
       (__9_____30190));
  nor2s1 _____0_504764(.DIN1 (____0___27924), .DIN2 (_____0___41018),
       .Q (__9_____30188));
  and2s1 _______504765(.DIN1 (_____0___41020), .DIN2 (___0_____30654),
       .Q (__9_____30187));
  nor2s1 ______504766(.DIN1 (____9___29093), .DIN2 (__9_____29732), .Q
       (__9__0__30186));
  nor2s1 _______504767(.DIN1 (_____9__28570), .DIN2 (__9_9___29802), .Q
       (__9_09__30185));
  nor2s1 _______504768(.DIN1 (__9_____29827), .DIN2 (_________41028),
       .Q (__9_0___30184));
  nor2s1 _______504769(.DIN1 (__9_0___30182), .DIN2 (__9__0__29752), .Q
       (__9_0___30183));
  nnd2s1 _______504770(.DIN1 (__9_00__29804), .DIN2 (________29428), .Q
       (__9_0___30181));
  nor2s1 _______504771(.DIN1 (__9_0___30179), .DIN2 (__9_09), .Q
       (__9_0___30180));
  and2s1 ______504772(.DIN1 (______0__41022), .DIN2 (__9_00__30177), .Q
       (__9_0___30178));
  nnd2s1 _______504773(.DIN1 (__9__0), .DIN2 (_____9__28914), .Q
       (__9_99__30176));
  nnd2s1 _______504774(.DIN1 (__9_____29776), .DIN2 (__9_9___30174), .Q
       (__9_9___30175));
  nor2s1 _______504775(.DIN1 (________29051), .DIN2 (__9_____29778), .Q
       (__9_9___30173));
  nor2s1 _______504776(.DIN1 (___0_____30961), .DIN2 (__9_____29786),
       .Q (__9_9___30172));
  nor2s1 _____9_504777(.DIN1 (________29249), .DIN2 (__9_0___29725), .Q
       (__9_9___30171));
  nnd2s1 _____0_504778(.DIN1 (__9__0__29780), .DIN2 (__9_90__30169), .Q
       (__9_9___30170));
  and2s1 _____0_504779(.DIN1 (__9_____30167), .DIN2 (__9990), .Q
       (__9__9__30168));
  nor2s1 ______504780(.DIN1 (____9___23879), .DIN2 (____9_0__37080), .Q
       (__9_____30166));
  nnd2s1 ______504781(.DIN1 (_____0___41016), .DIN2 (__9_____30423), .Q
       (__9_____30165));
  nnd2s1 _______504782(.DIN1 (__9_0___29727), .DIN2 (________29323), .Q
       (__9_____30164));
  nnd2s1 _______504783(.DIN1 (__9_____29839), .DIN2 (__9_____30163), .Q
       (___0_____30673));
  nnd2s1 _______504784(.DIN1 (_____9___41010), .DIN2 (______9__33575),
       .Q (__9_____30428));
  nor2s1 _______504785(.DIN1 (________29110), .DIN2 (__9__9__29796), .Q
       (___00____30568));
  nor2s1 _______504786(.DIN1 (__9__0__30394), .DIN2 (_________41024),
       .Q (___00____30575));
  nnd2s1 ______504787(.DIN1 (__9_____29774), .DIN2 (__9_____30162), .Q
       (___00____30570));
  nnd2s1 _______504788(.DIN1 (__9_____29767), .DIN2 (__9_____30332), .Q
       (__9_____30426));
  nor2s1 ____9__504789(.DIN1 (___9____27774), .DIN2 (_________41030),
       .Q (__99____30522));
  or2s1 ____9__504790(.DIN1 (___0_____30760), .DIN2 (__9__0__29744), .Q
       (__999_));
  nnd2s1 _______504791(.DIN1 (__9_____29852), .DIN2 (____0___28839), .Q
       (___00____30596));
  nnd2s1 ____9__504792(.DIN1 (__9_____29784), .DIN2 (________27537), .Q
       (___0_____31100));
  nor2s1 ____9_504793(.DIN1 (__90____29692), .DIN2 (__909___29723), .Q
       (__99____30536));
  nnd2s1 _______504794(.DIN1 (__9_____30189), .DIN2 (___0_____31394),
       .Q (___00_0__30603));
  nor2s1 _______504795(.DIN1 (_____0___34102), .DIN2 (__9__9__29831),
       .Q (____0____32524));
  or2s1 _______504796(.DIN1 (__9_9___29989), .DIN2 (____9_0__37080), .Q
       (____0____37173));
  hi1s1 ______504797(.DIN (_________36288), .Q (_________35966));
  hi1s1 _______504798(.DIN (____9_9__36114), .Q (_________36870));
  nnd2s1 ______504799(.DIN1 (__9_____30325), .DIN2 (________29528), .Q
       (__9_____30161));
  nnd2s1 ____0__504800(.DIN1 (__9__0__30159), .DIN2 (_________33321),
       .Q (__9_____30160));
  or2s1 _____504801(.DIN1 (__90____29716), .DIN2 (_________35186), .Q
       (__9__9__30158));
  nnd2s1 _______504802(.DIN1 (___9____29594), .DIN2 (__9_____29737), .Q
       (__9_____30157));
  nnd2s1 _______504803(.DIN1 (__90____29711), .DIN2 (________23776), .Q
       (__9_____30156));
  or2s1 _______504804(.DIN1 (________23817), .DIN2 (__90_0__29660), .Q
       (__9_____30155));
  nnd2s1 _______504805(.DIN1 (__90____29710), .DIN2 (inData[0]), .Q
       (__9_____30154));
  nnd2s1 ______504806(.DIN1 (__90_0__29709), .DIN2 (____00__25678), .Q
       (__9_____30153));
  nnd2s1 ______504807(.DIN1 (____99__27741), .DIN2 (__90____29682), .Q
       (__9_____30152));
  nor2s1 _______504808(.DIN1 (_________31809), .DIN2 (__90____29706),
       .Q (__9_____30151));
  nnd2s1 ______504809(.DIN1 (__90____29656), .DIN2 (________29453), .Q
       (__9__0__30150));
  nnd2s1 _______504810(.DIN1 (_________38377), .DIN2 (__90____29700),
       .Q (__9__9__30149));
  nnd2s1 _______504811(.DIN1 (_________38377), .DIN2 (__90____29703),
       .Q (__9_____30148));
  nor2s1 _______504812(.DIN1 (________29144), .DIN2 (__90_9__29669), .Q
       (__9_____30147));
  nor2s1 _______504813(.DIN1 (__9_____29827), .DIN2 (__90____29693), .Q
       (__9_____30146));
  nnd2s1 _______504814(.DIN1 (__90____29702), .DIN2 (____0____37165),
       .Q (__9_____30145));
  nor2s1 _______504815(.DIN1 (____0___27656), .DIN2 (__90____29676), .Q
       (__9_____30144));
  or2s1 ______504816(.DIN1 (__9_____30142), .DIN2 (__90____29687), .Q
       (__9_____30143));
  nnd2s1 ______504817(.DIN1 (__90____29691), .DIN2 (__9_____29792), .Q
       (__9_____30141));
  nor2s1 _______504818(.DIN1 (____9___28193), .DIN2 (__90____29677), .Q
       (__9__0__30140));
  nor2s1 _______504819(.DIN1 (___9_9__27776), .DIN2 (__90_0__29689), .Q
       (__9__9__30139));
  nnd2s1 _______504820(.DIN1 (__90____29686), .DIN2 (__9_09__30281), .Q
       (__9_____30138));
  nnd2s1 _____0_504821(.DIN1 (__90____29683), .DIN2 (________28949), .Q
       (__9_____30137));
  nor2s1 _______504822(.DIN1 (___00_9__30621), .DIN2 (__90____29707),
       .Q (__9_____30136));
  nnd2s1 ______504823(.DIN1 (__90____29713), .DIN2 (____0____37165), .Q
       (__9_____30135));
  and2s1 _______504824(.DIN1 (__90_9__29679), .DIN2 (______0__33736),
       .Q (__9_____30134));
  or2s1 _______504825(.DIN1 (_________33549), .DIN2 (__90____29673), .Q
       (__9_____30133));
  nor2s1 _______504826(.DIN1 (____0___29471), .DIN2 (__90____29674), .Q
       (__9_____30132));
  and2s1 _______504827(.DIN1 (__90____29681), .DIN2 (__9__0__30130), .Q
       (__9_____30131));
  nnd2s1 ______504828(.DIN1 (____90__29543), .DIN2 (__9_____30126), .Q
       (__9__9__30129));
  nnd2s1 _______504829(.DIN1 (__90____29662), .DIN2 (___0____27869), .Q
       (__9_____30128));
  nor2s1 _____9_504830(.DIN1 (__9_____30126), .DIN2 (__9__0__30291), .Q
       (__9_____30127));
  nnd2s1 _____0_504831(.DIN1 (____0___26234), .DIN2 (__90_0__29680), .Q
       (__9_____30125));
  or2s1 _____0_504832(.DIN1 (_________36858), .DIN2 (__90____29704), .Q
       (__9_____30124));
  nor2s1 _______504833(.DIN1 (________28243), .DIN2 (__90____29668), .Q
       (__9_____30123));
  or2s1 _______504834(.DIN1 (_____9___33059), .DIN2 (__90____29667), .Q
       (__9_____30122));
  or2s1 _______504835(.DIN1 (__9__0__30120), .DIN2 (____9___29550), .Q
       (__9_____30121));
  xor2s1 ______504836(.DIN1 (________22726), .DIN2 (__9_____29959), .Q
       (__9__9__30119));
  xor2s1 _______504837(.DIN1 (____9___29005), .DIN2 (_________37884),
       .Q (__9_____30118));
  or2s1 _______504838(.DIN1 (__9_____30115), .DIN2 (___9____29595), .Q
       (__9_____30116));
  nnd2s1 _______504839(.DIN1 (__9_____30031), .DIN2 (___0_____40509),
       .Q (__9_____30114));
  nnd2s1 ______504840(.DIN1 (___99___29631), .DIN2 (_________38262), .Q
       (__9_____30113));
  nnd2s1 _______504841(.DIN1 (_________41034), .DIN2 (inData[26]), .Q
       (__9_____30112));
  nnd2s1 _______504842(.DIN1 (__900___29643), .DIN2 (_____0__25389), .Q
       (__9__0__30111));
  nor2s1 ______504843(.DIN1 (__9_____30109), .DIN2 (__900___29639), .Q
       (__9__9__30110));
  nor2s1 _______504844(.DIN1 (________29516), .DIN2 (___0____28791), .Q
       (__9_____30108));
  or2s1 _______504845(.DIN1 (___0_____31129), .DIN2 (__900___29638), .Q
       (__9_____30107));
  nnd2s1 _______504846(.DIN1 (________29479), .DIN2 (___9____29587), .Q
       (__9_____30106));
  nnd2s1 _______504847(.DIN1 (____99__28645), .DIN2 (___9____29624), .Q
       (__9_____30105));
  nnd2s1 _______504848(.DIN1 (__90____29665), .DIN2 (___99___29634), .Q
       (__9_____30104));
  nnd2s1 _______504849(.DIN1 (___99___29632), .DIN2 (________29070), .Q
       (__9_____30103));
  and2s1 _______504850(.DIN1 (___9_0__29570), .DIN2 (________28308), .Q
       (__9__0__30102));
  and2s1 _______504851(.DIN1 (___99___29630), .DIN2 (___0_____30719),
       .Q (__9__9__30101));
  nnd2s1 _____504852(.DIN1 (__9_____29957), .DIN2 (_________41066), .Q
       (__9_____30100));
  nor2s1 _____9_504853(.DIN1 (__9_____30098), .DIN2 (__90_0__29650), .Q
       (__9_____30099));
  and2s1 _____504854(.DIN1 (___990__29628), .DIN2 (__9_____30096), .Q
       (__9_____30097));
  nnd2s1 _____0_504855(.DIN1 (___9_0__29620), .DIN2 (________29180), .Q
       (__9_____30095));
  or2s1 _____0_504856(.DIN1 (__9__0__30093), .DIN2 (___9____29617), .Q
       (__9_____30094));
  nor2s1 _______504857(.DIN1 (____99__28013), .DIN2 (___9____29618), .Q
       (__9_09__30092));
  nor2s1 _______504858(.DIN1 (________29319), .DIN2 (___9____29623), .Q
       (__9_0___30091));
  nnd2s1 _______504859(.DIN1 (__900___29640), .DIN2 (__9_____29873), .Q
       (__9_0___30090));
  nnd2s1 _______504860(.DIN1 (__9_0___30085), .DIN2 (___90___26868), .Q
       (__9_0___30089));
  nnd2s1 _______504861(.DIN1 (___9____29616), .DIN2 (________29140), .Q
       (__9_0___30088));
  or2s1 _______504862(.DIN1 (_________32602), .DIN2 (___9____29567), .Q
       (__9_0___30087));
  nnd2s1 ______504863(.DIN1 (__9_0___30085), .DIN2 (___9____29612), .Q
       (__9_0___30086));
  nnd2s1 _______504864(.DIN1 (___9_0__29611), .DIN2 (____9___27477), .Q
       (__9_0___30084));
  nnd2s1 _______504865(.DIN1 (___9_9__29610), .DIN2 (__9990), .Q
       (__9_00__30083));
  nor2s1 _______504866(.DIN1 (________28441), .DIN2 (___9____29609), .Q
       (__9_99__30082));
  and2s1 ______504867(.DIN1 (___9____29607), .DIN2 (________28519), .Q
       (__9_9___30081));
  or2s1 _______504868(.DIN1 (___0_____31336), .DIN2 (__9_9___30079), .Q
       (__9_9___30080));
  nnd2s1 _______504869(.DIN1 (___9____29605), .DIN2 (________28507), .Q
       (__9_9___30078));
  nor2s1 _______504870(.DIN1 (___9____26914), .DIN2 (___9____29604), .Q
       (__9_9___30077));
  or2s1 _______504871(.DIN1 (__9__9__30444), .DIN2 (__90____29654), .Q
       (__9_9___30076));
  or2s1 _______504872(.DIN1 (___0_____31194), .DIN2 (___9____29598), .Q
       (__9_9___30075));
  nor2s1 ______504873(.DIN1 (________29540), .DIN2 (__9__9__30073), .Q
       (__9_90__30074));
  nor2s1 _______504874(.DIN1 (_________31870), .DIN2 (__90____29658),
       .Q (__99____30482));
  xor2s1 _____0_504875(.DIN1 (________29480), .DIN2 (________29123), .Q
       (_________32024));
  dffacs1 _____________________________________________9_504876(.CLRB
       (reset), .CLK (clk), .DIN (__90_9__29698), .Q
       (_________________________________________________________________22000));
  or2s1 _____9_504877(.DIN1 (__9_____30071), .DIN2 (___9____29579), .Q
       (__9_____30072));
  nor2s1 _____9_504878(.DIN1 (________28317), .DIN2 (___9_9__29569), .Q
       (__9_____30070));
  nnd2s1 _____9_504879(.DIN1 (__9_____30049), .DIN2 (__9_0___29994), .Q
       (__9_____30069));
  nor2s1 _____9_504880(.DIN1 (________29205), .DIN2 (____9___29549), .Q
       (__9_____30068));
  nnd2s1 _____9_504881(.DIN1 (___9____29589), .DIN2 (____9___28919), .Q
       (__9_____30067));
  nnd2s1 _______504882(.DIN1 (___9____29583), .DIN2 (___0_99__30832),
       .Q (__9_____30066));
  nnd2s1 _______504883(.DIN1 (___9____29582), .DIN2 (__9_9___29893), .Q
       (__9_____30065));
  and2s1 _______504884(.DIN1 (___9____29581), .DIN2 (__9__9__30063), .Q
       (__9__0__30064));
  nor2s1 ______504885(.DIN1 (____0___28295), .DIN2 (______0__41062), .Q
       (__9_____30062));
  nnd2s1 _______504886(.DIN1 (__9_____30051), .DIN2 (_________41138),
       .Q (__9_____30061));
  nor2s1 _______504887(.DIN1 (__9_____29750), .DIN2 (___9_0__29576), .Q
       (__9_____30060));
  nnd2s1 _____0_504888(.DIN1 (_____9__29509), .DIN2 (__9_____30058), .Q
       (__9_____30059));
  nnd2s1 _______504889(.DIN1 (________27152), .DIN2 (________29512), .Q
       (__9_____30057));
  or2s1 _______504890(.DIN1 (__9_____30054), .DIN2 (_____9__29502), .Q
       (__9_____30055));
  nnd2s1 _______504891(.DIN1 (________29506), .DIN2 (___9_9__28688), .Q
       (__9_____30053));
  nnd2s1 _______504892(.DIN1 (__9_____30051), .DIN2 (____0___29098), .Q
       (__9_____30052));
  nnd2s1 _______504893(.DIN1 (__9_____30049), .DIN2 (_________41154),
       .Q (__9_____30050));
  nnd2s1 ______504894(.DIN1 (__9_____30255), .DIN2 (___9____29572), .Q
       (__9__0__30048));
  and2s1 _______504895(.DIN1 (__9_____30046), .DIN2 (___90___29557), .Q
       (__9__9__30047));
  nnd2s1 ______504896(.DIN1 (__90____29652), .DIN2 (___0____26093), .Q
       (__9_____30045));
  and2s1 _______504897(.DIN1 (_________41038), .DIN2 (__9_9___29990),
       .Q (__9_____30044));
  nor2s1 ______504898(.DIN1 (___0_____30798), .DIN2 (___9____29562), .Q
       (__9_____30043));
  nnd2s1 _______504899(.DIN1 (_________41044), .DIN2 (________28154),
       .Q (__9_____30042));
  nnd2s1 _______504900(.DIN1 (________29520), .DIN2 (_____0__27620), .Q
       (__9_____30041));
  or2s1 _______504901(.DIN1 (__9_____30039), .DIN2 (____9___29545), .Q
       (__9_____30040));
  nor2s1 _______504902(.DIN1 (___9_9__27767), .DIN2 (_____0__29527), .Q
       (__9__0__30038));
  nnd2s1 _____0_504903(.DIN1 (______0__41052), .DIN2 (____9___29002),
       .Q (__9_____30037));
  nnd2s1 _____0_504904(.DIN1 (___9_9__29585), .DIN2 (__9_____30035), .Q
       (__9_____30036));
  nor2s1 _______504905(.DIN1 (___099__27921), .DIN2 (________29539), .Q
       (__9_____30034));
  nnd2s1 _______504906(.DIN1 (___9____29565), .DIN2 (________28952), .Q
       (__9_____30033));
  nor2s1 _______504907(.DIN1 (inData[22]), .DIN2 (__9_____30031), .Q
       (__9_____30032));
  nnd2s1 _______504908(.DIN1 (________29538), .DIN2 (___90___28647), .Q
       (__9_____30030));
  and2s1 ______504909(.DIN1 (________29530), .DIN2 (__9_____30423), .Q
       (__9__9__30029));
  nor2s1 _______504910(.DIN1 (___0_____31336), .DIN2 (_________41036),
       .Q (__9_____30028));
  nnd2s1 _______504911(.DIN1 (_________41054), .DIN2 (___0_0___30748),
       .Q (__9_____30027));
  nor2s1 _______504912(.DIN1 (____0___29104), .DIN2 (___9____29599), .Q
       (__9_____30026));
  nnd2s1 _______504913(.DIN1 (_________41046), .DIN2 (__9_____30024),
       .Q (__9_____30025));
  nnd2s1 _______504914(.DIN1 (___90___29560), .DIN2 (__9_____29921), .Q
       (__9_____30023));
  nnd2s1 _______504915(.DIN1 (________29532), .DIN2 (___0_0___30748),
       .Q (__9_____30022));
  nor2s1 _______504916(.DIN1 (________27153), .DIN2 (________29517), .Q
       (__9_____30021));
  nnd2s1 _______504917(.DIN1 (__9_____30019), .DIN2 (________29524), .Q
       (__9__9__30020));
  nnd2s1 _______504918(.DIN1 (___90___29554), .DIN2 (_____0___37283),
       .Q (__9_____30018));
  or2s1 _______504919(.DIN1 (__9_____30016), .DIN2 (___9____29626), .Q
       (__9_____30017));
  nnd2s1 _______504920(.DIN1 (______0__41042), .DIN2 (___0____27858),
       .Q (__9_____30015));
  nnd2s1 _______504921(.DIN1 (________29536), .DIN2 (__9_____30163), .Q
       (__9_____30014));
  nor2s1 _______504922(.DIN1 (____0_9__31542), .DIN2 (_____9__29526),
       .Q (__9_____30013));
  nnd2s1 _____9_504923(.DIN1 (________29518), .DIN2 (__9_9___30270), .Q
       (__9_____30012));
  or2s1 _____9_504924(.DIN1 (__9__9__30010), .DIN2 (_________41050), .Q
       (__9__0__30011));
  nor2s1 _____9_504925(.DIN1 (___9____29606), .DIN2 (________29535), .Q
       (__9_____30009));
  and2s1 ____90_504926(.DIN1 (__9_____30007), .DIN2 (________27151), .Q
       (__9_____30008));
  nor2s1 ____90_504927(.DIN1 (__9_____29783), .DIN2 (___90___29555), .Q
       (__9_____30006));
  nnd2s1 _______504928(.DIN1 (_____0__29510), .DIN2 (___9____28722), .Q
       (__9_____30005));
  nnd2s1 ____0_504929(.DIN1 (___9____29577), .DIN2 (__9__0__30003), .Q
       (__9_____30004));
  nor2s1 ____0_504930(.DIN1 (___0____28754), .DIN2 (_________41060), .Q
       (__9_09__30002));
  nor2s1 ____0_504931(.DIN1 (__9_0___30000), .DIN2 (_________41058), .Q
       (__9_0___30001));
  nnd2s1 ____0__504932(.DIN1 (_________41056), .DIN2 (________28484),
       .Q (__9_0___29999));
  nnd2s1 ____9__504933(.DIN1 (__9_0___29997), .DIN2 (____09___35375),
       .Q (__9_0___29998));
  xor2s1 ____9__504934(.DIN1 (______9__35773), .DIN2 (___9_____39397),
       .Q (__9_0___29996));
  and2s1 _______504935(.DIN1 (___99___29633), .DIN2 (____0____32499),
       .Q (______0__32940));
  nnd2s1 ____9__504936(.DIN1 (____9_9__34346), .DIN2 (___9____29564),
       .Q (_________34013));
  or2s1 ____9__504937(.DIN1 (__9_0___29995), .DIN2 (___9_0__29586), .Q
       (__9__9__30393));
  and2s1 ____9__504938(.DIN1 (__9_0___29994), .DIN2 (_____0__27251), .Q
       (__9_____30396));
  nor2s1 ____9__504939(.DIN1 (__9_00__29993), .DIN2 (_________41048),
       .Q (__9_____30398));
  nnd2s1 ____504940(.DIN1 (_________41040), .DIN2 (__9_99__29992), .Q
       (__9_____30385));
  nor2s1 _______504941(.DIN1 (_________33175), .DIN2 (________29504),
       .Q (_________32797));
  nnd2s1 _____0_504942(.DIN1 (________29507), .DIN2 (___0_____31151),
       .Q (__9_00__30366));
  nnd2s1 ______504943(.DIN1 (__9_9___29990), .DIN2 (_________41064), .Q
       (__9_____30232));
  nor2s1 ______504944(.DIN1 (___0_____31073), .DIN2 (__90____29646), .Q
       (__9_____30416));
  nnd2s1 ______504945(.DIN1 (__909_), .DIN2 (__9_9___29989), .Q
       (______9__35498));
  and2s1 _______504946(.DIN1 (___9____29621), .DIN2 (___09____31472),
       .Q (____99___32478));
  and2s1 _______504947(.DIN1 (___9____29613), .DIN2 (__9_____30024), .Q
       (__9_____30407));
  nor2s1 _______504948(.DIN1 (__9_____29827), .DIN2 (_____0__29503), .Q
       (_________32598));
  dffacs1 _______________________________________________504949(.CLRB
       (reset), .CLK (clk), .DIN (__90____29678), .Q
       (_________________________________________________________________22001));
  dffacs1 _________________________________________0____504950(.CLRB
       (reset), .CLK (clk), .DIN (___909__29561), .QN (___0_____40579));
  nnd2s1 _______504951(.DIN1 (__900___29644), .DIN2 (____0___29012), .Q
       (____9_9__36114));
  nnd2s1 ____9__504952(.DIN1 (__9_____30031), .DIN2 (________27259), .Q
       (____0____37147));
  nnd2s1 ______504953(.DIN1 (__90_0), .DIN2 (________28454), .Q
       (_________36288));
  nor2s1 _______504954(.DIN1 (___09___27917), .DIN2 (____00__29369), .Q
       (__9_9___29988));
  nnd2s1 _______504955(.DIN1 (_____0__29486), .DIN2 (__9_9___29986), .Q
       (__9_9___29987));
  nnd2s1 _______504956(.DIN1 (__9__9__29984), .DIN2 (__90____29661), .Q
       (__9_90__29985));
  nnd2s1 _____0_504957(.DIN1 (________29492), .DIN2 (___9_0__27768), .Q
       (__9_____29983));
  nnd2s1 ______504958(.DIN1 (________29493), .DIN2 (__9_____29981), .Q
       (__9_____29982));
  nor2s1 _______504959(.DIN1 (________29481), .DIN2 (__9_____29979), .Q
       (__9_____29980));
  nor2s1 _____0_504960(.DIN1 (___0_0__27855), .DIN2 (_____9__29485), .Q
       (__9_____29978));
  nnd2s1 _____0_504961(.DIN1 (________29491), .DIN2 (__9_____29976), .Q
       (__9_____29977));
  xor2s1 ______504962(.DIN1
       (____________________________________________21831), .DIN2
       (______0__33640), .Q (__9__0__29975));
  xnr2s1 _______504963(.DIN1 (___0_9___40553), .DIN2 (_____9___38611),
       .Q (__9__9__29974));
  xor2s1 ______504964(.DIN1 (____9___29095), .DIN2
       (_____________22099), .Q (__9_____29973));
  xor2s1 _______504965(.DIN1 (____9___22449), .DIN2 (_____9___38611),
       .Q (__9_____29972));
  nnd2s1 _______504966(.DIN1 (____0___29473), .DIN2 (__9_____29968), .Q
       (__9_____29969));
  nnd2s1 _______504967(.DIN1 (____0___29375), .DIN2 (__9__0__29966), .Q
       (__9_____29967));
  nnd2s1 _______504968(.DIN1 (________29430), .DIN2
       (______________________________________________21930), .Q
       (__9__9__29965));
  nnd2s1 _______504969(.DIN1 (_________37414), .DIN2 (inData[23]), .Q
       (__9_____29964));
  nor2s1 _______504970(.DIN1 (___0____27849), .DIN2 (________29337), .Q
       (__9_____29963));
  and2s1 _______504971(.DIN1 (____0___29472), .DIN2 (________28407), .Q
       (__9_____29962));
  nnd2s1 _______504972(.DIN1 (____0___29470), .DIN2 (________28634), .Q
       (__9_____29961));
  nor2s1 _______504973(.DIN1 (________22725), .DIN2 (__9_____29959), .Q
       (__9_____29960));
  nnd2s1 _______504974(.DIN1 (__9_____29957), .DIN2 (__90____29648), .Q
       (__9_____29958));
  nor2s1 ______504975(.DIN1 (___0_____30961), .DIN2 (_____9__29445), .Q
       (__9__0__29956));
  nor2s1 _______504976(.DIN1 (___9____26010), .DIN2 (____9___29457), .Q
       (__9__9__29955));
  nor2s1 _______504977(.DIN1 (________28094), .DIN2 (____9___29464), .Q
       (__9_____29954));
  nor2s1 _______504978(.DIN1 (______9__22017), .DIN2 (___0_____40583),
       .Q (__9_____29953));
  nnd2s1 _______504979(.DIN1 (___0_____40583), .DIN2 (______9__22017),
       .Q (__9_____29952));
  nor2s1 ______504980(.DIN1 (________28336), .DIN2 (____99__29465), .Q
       (__9_____29951));
  nnd2s1 _______504981(.DIN1 (_____0__29446), .DIN2 (__9_____29949), .Q
       (__9_____29950));
  nnd2s1 _______504982(.DIN1 (____9___29460), .DIN2 (__9_____29866), .Q
       (__9_____29948));
  or2s1 _____9_504983(.DIN1 (__9__0__29946), .DIN2 (________29454), .Q
       (__9_____29947));
  nor2s1 _____9_504984(.DIN1 (________29301), .DIN2 (___0____28798), .Q
       (__9__9__29945));
  nor2s1 _____9_504985(.DIN1 (__9_____29932), .DIN2 (________29449), .Q
       (__9_____29944));
  nnd2s1 _____0_504986(.DIN1 (________29394), .DIN2 (__9_____29941), .Q
       (__9_____29943));
  nnd2s1 _____0_504987(.DIN1 (________29404), .DIN2 (__9_____29941), .Q
       (__9_____29942));
  nnd2s1 _____0_504988(.DIN1 (________29382), .DIN2 (___0____27839), .Q
       (__9_____29940));
  nor2s1 _____0_504989(.DIN1 (__9_____29766), .DIN2 (________29443), .Q
       (__9_____29939));
  nnd2s1 _____504990(.DIN1 (____09__29475), .DIN2 (inData[6]), .Q
       (__9_____29938));
  nor2s1 ______504991(.DIN1 (________29039), .DIN2 (__9__0__29926), .Q
       (__9_____29937));
  nor2s1 _______504992(.DIN1 (__9__9__29935), .DIN2 (________29444), .Q
       (__9__0__29936));
  nor2s1 _______504993(.DIN1 (________28283), .DIN2 (________29427), .Q
       (__9_____29934));
  nor2s1 _______504994(.DIN1 (__9_____29932), .DIN2 (_____9__29435), .Q
       (__9_____29933));
  and2s1 _______504995(.DIN1 (________29434), .DIN2 (________29533), .Q
       (__9_____29931));
  nor2s1 ______504996(.DIN1 (________29432), .DIN2 (________27172), .Q
       (__9_____29930));
  nor2s1 _______504997(.DIN1 (___0_0__26999), .DIN2 (_____9__29344), .Q
       (__9_____29929));
  nor2s1 _______504998(.DIN1 (___9____29584), .DIN2 (________29414), .Q
       (__9_____29928));
  nor2s1 _______504999(.DIN1 (___0_9__28765), .DIN2 (__9__0__29926), .Q
       (__9_____29927));
  nnd2s1 _______505000(.DIN1 (________29494), .DIN2 (________29350), .Q
       (__9__9__29925));
  nnd2s1 _______505001(.DIN1 (_____0__29426), .DIN2 (___09____31461),
       .Q (__9_____29924));
  nnd2s1 _______505002(.DIN1 (________29343), .DIN2 (________26520), .Q
       (__9_____29923));
  nnd2s1 _______505003(.DIN1 (________29422), .DIN2 (__9_____29921), .Q
       (__9_____29922));
  and2s1 _______505004(.DIN1 (________29421), .DIN2 (__99____30480), .Q
       (__9_____29920));
  nnd2s1 ______505005(.DIN1 (________29419), .DIN2 (___0____28784), .Q
       (__9_____29919));
  nor2s1 ______505006(.DIN1 (__9_____30380), .DIN2 (________29418), .Q
       (__9_____29918));
  nor2s1 _______505007(.DIN1 (__9__0__29916), .DIN2 (_____9__29416), .Q
       (__9_____29917));
  and2s1 _______505008(.DIN1 (__9_____29914), .DIN2 (_____9__27471), .Q
       (__9__9__29915));
  nor2s1 _______505009(.DIN1 (___9____27798), .DIN2 (________29440), .Q
       (__9_____29913));
  and2s1 ______505010(.DIN1 (________29413), .DIN2 (__9_____29911), .Q
       (__9_____29912));
  nnd2s1 _______505011(.DIN1 (________29412), .DIN2 (________27287), .Q
       (__9_____29910));
  nor2s1 ______505012(.DIN1 (__9_____29908), .DIN2 (________29496), .Q
       (__9_____29909));
  nor2s1 _______505013(.DIN1 (________28337), .DIN2 (________29403), .Q
       (__9_____29907));
  nor2s1 _______505014(.DIN1 (___0____28758), .DIN2 (________29401), .Q
       (__9__0__29906));
  nor2s1 _______505015(.DIN1 (__9_0___29904), .DIN2 (________29400), .Q
       (__9_09__29905));
  nnd2s1 _____505016(.DIN1 (_____0__29353), .DIN2 (___9____27791), .Q
       (__9_0___29903));
  nnd2s1 _____9_505017(.DIN1 (________29388), .DIN2 (___0____28788), .Q
       (__9_0___29902));
  nor2s1 _____505018(.DIN1 (_______22226), .DIN2 (____9____37049), .Q
       (__9_0___29901));
  nnd2s1 _____0_505019(.DIN1 (________29383), .DIN2 (__9_0___29899), .Q
       (__9_0___29900));
  or2s1 _____0_505020(.DIN1 (__9_0___29897), .DIN2 (_____9__29352), .Q
       (__9_0___29898));
  and2s1 _____0_505021(.DIN1 (________29380), .DIN2 (__9_99__29895), .Q
       (__9_00__29896));
  nnd2s1 _____0_505022(.DIN1 (__9_9___29893), .DIN2 (____09__29377), .Q
       (__9_9___29894));
  and2s1 _______505023(.DIN1 (_____0__29378), .DIN2 (________26190), .Q
       (__9_9___29891));
  or2s1 _______505024(.DIN1 (__9__9__30262), .DIN2 (_____9__29396), .Q
       (__9_9___29890));
  nor2s1 _______505025(.DIN1 (________29340), .DIN2 (__9_9___29888), .Q
       (__9_9___29889));
  nor2s1 ______505026(.DIN1 (________27153), .DIN2 (________29398), .Q
       (__9_90__29887));
  nor2s1 _______505027(.DIN1 (_________37321), .DIN2 (_________37414),
       .Q (__9__9__29886));
  nor2s1 _______505028(.DIN1 (________22418), .DIN2 (_________37414),
       .Q (__9_____29885));
  or2s1 _______505029(.DIN1 (__9_____29883), .DIN2 (____9___29459), .Q
       (__9_____29884));
  nor2s1 _______505030(.DIN1 (__9_____29881), .DIN2 (______0__41082),
       .Q (__9_____29882));
  nor2s1 _______505031(.DIN1 (___9____27772), .DIN2 (________29360), .Q
       (__9_____29880));
  and2s1 _______505032(.DIN1 (_____0__29397), .DIN2 (__9__0__29878), .Q
       (__9_____29879));
  nor2s1 _______505033(.DIN1 (__90____29663), .DIN2 (__9_____29876), .Q
       (__9__9__29877));
  nor2s1 _______505034(.DIN1 (________29433), .DIN2 (________29119), .Q
       (__9_____29875));
  nnd2s1 ______505035(.DIN1 (________29429), .DIN2 (__9_____29873), .Q
       (__9_____29874));
  nor2s1 _______505036(.DIN1 (____0___29105), .DIN2 (____0___29468), .Q
       (__9_____29872));
  or2s1 _______505037(.DIN1 (__9_____29870), .DIN2 (____99__29368), .Q
       (__9_____29871));
  xnr2s1 _______505038(.DIN1 (________28985), .DIN2
       (_____________________________________________21927), .Q
       (__9_____29869));
  nor2s1 ______505039(.DIN1 (__909___29720), .DIN2 (____90__29456), .Q
       (__9__0__29868));
  nnd2s1 _______505040(.DIN1 (________29355), .DIN2 (__9_____29866), .Q
       (__9__9__29867));
  nor2s1 _______505041(.DIN1 (________29411), .DIN2 (__9_____30417), .Q
       (__9_____29865));
  nor2s1 _______505042(.DIN1 (__9_____29863), .DIN2 (__9_____29862), .Q
       (__9_____29864));
  or2s1 ______505043(.DIN1 (__9_____29860), .DIN2 (_________41070), .Q
       (__9_____29861));
  and2s1 _______505044(.DIN1 (__9_____29857), .DIN2 (__9_____29957), .Q
       (__9_____29858));
  nnd2s1 _______505045(.DIN1 (__9_9___30270), .DIN2 (__9_____29855), .Q
       (__9_____29856));
  nnd2s1 _____9_505046(.DIN1 (________29356), .DIN2 (__9_00__30177), .Q
       (__9_____29854));
  nor2s1 _____9_505047(.DIN1 (__9_____29754), .DIN2 (_____0__29476), .Q
       (__9_____29853));
  or2s1 _____9_505048(.DIN1 (__9_____29851), .DIN2 (________28421), .Q
       (__9_____29852));
  nnd2s1 _____0_505049(.DIN1 (____0___29469), .DIN2 (__9__9__29849), .Q
       (__9__0__29850));
  and2s1 _____0_505050(.DIN1 (__9_____29847), .DIN2 (__9_9___30270), .Q
       (__9_____29848));
  nnd2s1 ______505051(.DIN1 (________29333), .DIN2 (__9_____29845), .Q
       (__9_____29846));
  nnd2s1 _______505052(.DIN1 (_____0__29335), .DIN2 (__9_____29843), .Q
       (__9_____29844));
  nor2s1 _______505053(.DIN1 (__9__0__29841), .DIN2 (________29306), .Q
       (__9_____29842));
  nor2s1 _______505054(.DIN1 (____9___28640), .DIN2 (_____9__29304), .Q
       (__9__9__29840));
  nor2s1 _______505055(.DIN1 (________29225), .DIN2 (________29310), .Q
       (__9_____29839));
  nnd2s1 _______505056(.DIN1 (____9___29462), .DIN2 (________26622), .Q
       (__9_____29838));
  nnd2s1 _______505057(.DIN1 (________29442), .DIN2 (____999__33432),
       .Q (__9_____29837));
  nor2s1 _______505058(.DIN1 (___0_____30961), .DIN2 (________29488),
       .Q (__9_____29836));
  nnd2s1 _______505059(.DIN1 (____9___29363), .DIN2 (__9_____29834), .Q
       (_________32364));
  nor2s1 _______505060(.DIN1 (________27934), .DIN2 (________29448), .Q
       (_________32639));
  nor2s1 _______505061(.DIN1 (___0____27881), .DIN2 (________29347), .Q
       (_________32004));
  nor2s1 _______505062(.DIN1 (___0_9___31111), .DIN2 (________29410),
       .Q (__9_____30117));
  nor2s1 _______505063(.DIN1 (_____9___32184), .DIN2 (________29423),
       .Q (____0____33493));
  nor2s1 _______505064(.DIN1 (____90__28462), .DIN2 (________29484), .Q
       (_________36082));
  and2s1 ____505065(.DIN1 (__9__0__29832), .DIN2 (________27494), .Q
       (__9_____29833));
  nnd2s1 ______505066(.DIN1 (________29437), .DIN2 (_________32114), .Q
       (__9__9__29831));
  nor2s1 _______505067(.DIN1 (________29327), .DIN2 (___0_0__27855), .Q
       (__9_____29830));
  and2s1 ______505068(.DIN1 (__9_9___29893), .DIN2 (_________41134), .Q
       (__9_____29829));
  nor2s1 ______505069(.DIN1 (__9_____29827), .DIN2 (________29318), .Q
       (__9_____29828));
  nor2s1 _______505070(.DIN1 (___0_____30656), .DIN2 (_____9__29406),
       .Q (__9_____29826));
  nor2s1 _______505071(.DIN1 (__9__0__29824), .DIN2 (________29390), .Q
       (__9_____29825));
  nor2s1 _______505072(.DIN1 (__9_____29827), .DIN2 (________29317), .Q
       (__9__9__29823));
  nor2s1 _______505073(.DIN1 (___0____27862), .DIN2 (________29294), .Q
       (__9_____29822));
  nor2s1 _______505074(.DIN1 (___009__27835), .DIN2 (____0___29474), .Q
       (__9_____29821));
  nnd2s1 _______505075(.DIN1 (_________41068), .DIN2 (__9_9___30270),
       .Q (__9_____29820));
  nnd2s1 _______505076(.DIN1 (_____0__29325), .DIN2 (__9_____29818), .Q
       (__9_____29819));
  nnd2s1 _______505077(.DIN1 (________29308), .DIN2 (_____0__29315), .Q
       (__9_____29817));
  nnd2s1 _____9_505078(.DIN1 (________29303), .DIN2 (___0_0___30748),
       .Q (__9_____29816));
  or2s1 _____9_505079(.DIN1 (___0_____40156), .DIN2 (________29438), .Q
       (__9_____29815));
  nnd2s1 _____9_505080(.DIN1 (__90_9__29717), .DIN2 (____0___29376), .Q
       (__9__0__29814));
  nnd2s1 _____9_505081(.DIN1 (________29332), .DIN2 (________29361), .Q
       (__9_09__29813));
  nor2s1 ____505082(.DIN1 (_____9__28190), .DIN2 (________29328), .Q
       (__9_0___29812));
  and2s1 ____90_505083(.DIN1 (_________38743), .DIN2 (___0_____40583),
       .Q (__9_0___29811));
  nnd2s1 ____90_505084(.DIN1 (________29320), .DIN2 (__9_____29873), .Q
       (__9_0___29810));
  nor2s1 ____90_505085(.DIN1 (_____0__23319), .DIN2 (____9____37049),
       .Q (__9_0___29809));
  nnd2s1 ____90_505086(.DIN1 (_____9__27471), .DIN2 (________29312), .Q
       (__9_0___29808));
  nor2s1 _______505087(.DIN1 (___9_0__28698), .DIN2 (__9_0___29805), .Q
       (__9_0___29807));
  nor2s1 ______505088(.DIN1 (__9_0___29805), .DIN2 (_____9__29386), .Q
       (__9_0___29806));
  nor2s1 _______505089(.DIN1 (___9____27770), .DIN2 (____9___29187), .Q
       (__9_00__29804));
  xor2s1 ____9_505090(.DIN1 (________28883), .DIN2 (___0_00__40461), .Q
       (__9_99));
  nor2s1 _______505091(.DIN1 (__9_____29827), .DIN2 (________29179), .Q
       (__9_9___29803));
  nnd2s1 _______505092(.DIN1 (__9_9___29801), .DIN2 (_____9__29184), .Q
       (__9_9___29802));
  and2s1 _______505093(.DIN1 (__9_9___29799), .DIN2 (__9_____30019), .Q
       (__9_9___29800));
  nnd2s1 ____9__505094(.DIN1 (_________34225), .DIN2 (___0_____40620),
       .Q (__9_9___29798));
  nnd2s1 ____9__505095(.DIN1 (_________34225), .DIN2 (_________22032),
       .Q (__9_9___29797));
  nnd2s1 ____9__505096(.DIN1 (____9___29274), .DIN2 (_____0__28276), .Q
       (__9_9_));
  nnd2s1 ____9_505097(.DIN1 (__9_____29739), .DIN2 (inData[19]), .Q
       (__9_90));
  or2s1 ____9__505098(.DIN1 (_________41285), .DIN2 (__9_____29731), .Q
       (__9__9__29796));
  or2s1 ____9__505099(.DIN1 (__99____30463), .DIN2 (____09__29203), .Q
       (__9_____29795));
  nnd2s1 ____99_505100(.DIN1 (_________41080), .DIN2 (________29447),
       .Q (__9_____29794));
  nnd2s1 ____00_505101(.DIN1 (_____0__29219), .DIN2 (__9_____29792), .Q
       (__9_____29793));
  nor2s1 ____00_505102(.DIN1 (___00_9__30621), .DIN2 (________29265),
       .Q (__9_____29791));
  nnd2s1 ____00_505103(.DIN1 (________29267), .DIN2 (___9____28685), .Q
       (__9_____29790));
  nor2s1 ____0_505104(.DIN1 (________29182), .DIN2 (________29047), .Q
       (__9__0__29789));
  nor2s1 ____0__505105(.DIN1 (__9_0___30179), .DIN2 (________29258), .Q
       (__9__9__29788));
  nor2s1 ____0__505106(.DIN1 (________28527), .DIN2 (________29260), .Q
       (__9_____29787));
  nor2s1 ____0__505107(.DIN1 (__9_0___29724), .DIN2 (________29257), .Q
       (__9_____29786));
  nnd2s1 ____0_505108(.DIN1 (________29255), .DIN2 (___9____26932), .Q
       (__9_____29785));
  or2s1 ____0__505109(.DIN1 (__9_____29783), .DIN2 (_________41074), .Q
       (__9_____29784));
  nnd2s1 ____0__505110(.DIN1 (____9___29275), .DIN2 (________28460), .Q
       (__9_____29782));
  nnd2s1 ____0__505111(.DIN1 (____0___28925), .DIN2 (____0___29196), .Q
       (__9_____29781));
  and2s1 ____0__505112(.DIN1 (________29254), .DIN2 (__9__9__29779), .Q
       (__9__0__29780));
  nor2s1 ____0__505113(.DIN1 (__9_____29777), .DIN2 (________29226), .Q
       (__9_____29778));
  nnd2s1 ____0__505114(.DIN1 (_____9__29252), .DIN2 (__9_____29775), .Q
       (__9_____29776));
  nor2s1 ____0__505115(.DIN1 (__9_____29773), .DIN2 (________29247), .Q
       (__9_____29774));
  nnd2s1 ____0__505116(.DIN1 (_____9__29244), .DIN2 (__9_____29771), .Q
       (__9_____29772));
  nor2s1 ____0__505117(.DIN1 (________28934), .DIN2 (______0__41072),
       .Q (__9__0__29770));
  or2s1 ____0__505118(.DIN1 (________26656), .DIN2 (________29240), .Q
       (__9__9__29769));
  nnd2s1 ____0__505119(.DIN1 (_____9__29271), .DIN2 (___9____27763), .Q
       (__9_____29768));
  nor2s1 _______505120(.DIN1 (__9_____29766), .DIN2 (________29381), .Q
       (__9_____29767));
  or2s1 ____09_505121(.DIN1 (___0_____30669), .DIN2 (____00__29279), .Q
       (__9_____29765));
  nnd2s1 ____09_505122(.DIN1 (__9_____29756), .DIN2 (_______22277), .Q
       (__9_____29764));
  or2s1 _______505123(.DIN1 (__90____29653), .DIN2 (____0___29199), .Q
       (__9_____29763));
  nnd2s1 _______505124(.DIN1 (________29211), .DIN2 (__9_____30163), .Q
       (__9_____29762));
  nnd2s1 _______505125(.DIN1 (________29232), .DIN2 (__9__0__29760), .Q
       (__9_____29761));
  nnd2s1 _______505126(.DIN1 (________29228), .DIN2 (__9_____29758), .Q
       (__9__9__29759));
  nnd2s1 _______505127(.DIN1 (__9_____29756), .DIN2 (___0___22170), .Q
       (__9_____29757));
  nor2s1 _______505128(.DIN1 (________28614), .DIN2 (__9__0__30438), .Q
       (__9_____29755));
  nor2s1 _______505129(.DIN1 (____00___31509), .DIN2 (____90__29185),
       .Q (__9_____29753));
  or2s1 _______505130(.DIN1 (__9__9__29751), .DIN2 (________29206), .Q
       (__9__0__29752));
  and2s1 _____0_505131(.DIN1 (_____9__29234), .DIN2 (___0__9__30851),
       .Q (__9_____29749));
  nnd2s1 _______505132(.DIN1 (________29263), .DIN2 (______0__41180),
       .Q (__9_____29747));
  nor2s1 ______505133(.DIN1 (__9_____29745), .DIN2 (___09____40683), .Q
       (__9_____29746));
  or2s1 _______505134(.DIN1 (__9__9__29743), .DIN2 (________29214), .Q
       (__9__0__29744));
  nor2s1 _______505135(.DIN1 (___9____27754), .DIN2 (________29224), .Q
       (__9_____29741));
  nnd2s1 _______505136(.DIN1 (__9_____29739), .DIN2 (____9____38963),
       .Q (__9_____29740));
  and2s1 _______505137(.DIN1 (________29237), .DIN2 (__9_____29737), .Q
       (__9_____29738));
  nnd2s1 _______505138(.DIN1 (____9___29186), .DIN2 (_____0__27157), .Q
       (__9_____29736));
  nor2s1 _______505139(.DIN1 (____0___29197), .DIN2 (___0____28777), .Q
       (__9__0));
  nnd2s1 _______505140(.DIN1 (________29207), .DIN2 (__9_____29735), .Q
       (__9__9));
  nor2s1 _______505141(.DIN1 (________29236), .DIN2 (_________41076),
       .Q (__9_____29734));
  nor2s1 ______505142(.DIN1 (_____0__23826), .DIN2 (_________34225), .Q
       (__9_____29733));
  or2s1 ______505143(.DIN1 (____09__28843), .DIN2 (__9_____29731), .Q
       (__9_____29732));
  nor2s1 _______505144(.DIN1 (__9_____30039), .DIN2 (________29330), .Q
       (__9_____29730));
  nnd2s1 _______505145(.DIN1 (____0___29195), .DIN2 (___0_0___30748),
       .Q (__9___));
  nnd2s1 _____9_505146(.DIN1 (____9___29192), .DIN2 (__9_0___29729), .Q
       (__9_09));
  nnd2s1 _____505147(.DIN1 (________28908), .DIN2 (____9___29191), .Q
       (__9_0___29728));
  or2s1 _____0_505148(.DIN1 (__9_0___29726), .DIN2 (________29250), .Q
       (__9_0___29727));
  or2s1 _____505149(.DIN1 (__9_0___29724), .DIN2 (________29212), .Q
       (__9_0___29725));
  nor2s1 _______505150(.DIN1 (________29209), .DIN2 (________28594), .Q
       (__9_0_));
  nnd2s1 _______505151(.DIN1 (________29215), .DIN2 (_____9__28965), .Q
       (__9_00));
  nor2s1 _______505152(.DIN1 (________29049), .DIN2 (____0___29282), .Q
       (__9099));
  nnd2s1 _______505153(.DIN1 (____99__29193), .DIN2 (________28895), .Q
       (__909___29723));
  nnd2s1 _______505154(.DIN1 (_____0__28627), .DIN2 (____0___29284), .Q
       (__909___29722));
  nor2s1 ____9_505155(.DIN1 (__909___29721), .DIN2 (________29351), .Q
       (__9__9__30300));
  nnd2s1 ______505156(.DIN1 (___0____28771), .DIN2 (____0___29281), .Q
       (____0____31584));
  nnd2s1 _______505157(.DIN1 (__9_____30259), .DIN2 (________28992), .Q
       (_____0___32775));
  nor2s1 ____9__505158(.DIN1 (__909___29720), .DIN2 (_____0__29345), .Q
       (__9_____30250));
  nor2s1 _____9_505159(.DIN1 (__909___29719), .DIN2 (________29270), .Q
       (__9_____30229));
  and2s1 _____0_505160(.DIN1 (_____0__29288), .DIN2 (_________33128),
       .Q (____0____32512));
  nor2s1 _____0_505161(.DIN1 (________28935), .DIN2 (__909___29718), .Q
       (_________32325));
  or2s1 _______505162(.DIN1 (___0_____30760), .DIN2 (_____9__29261), .Q
       (__9_____30167));
  nor2s1 ____9_505163(.DIN1 (___9____29600), .DIN2 (_________37414), .Q
       (__9_9___30364));
  nor2s1 ____9__505164(.DIN1 (__99____30485), .DIN2 (________29424), .Q
       (__9_____30295));
  nnd2s1 _______505165(.DIN1 (__9_____29756), .DIN2 (___09___28825), .Q
       (_________37322));
  nor2s1 _______505166(.DIN1 (_____0___41315), .DIN2 (___0_____31132),
       .Q (__9_____30189));
  nor2s1 ____9__505167(.DIN1 (_________37317), .DIN2 (________29478),
       .Q (_________37576));
  or2s1 ______505168(.DIN1 (__9_____29739), .DIN2 (_________36713), .Q
       (_________36618));
  dffacs1 _________________________________________0_____505169(.CLRB
       (reset), .CLK (clk), .DIN (____9___29461), .Q (___0_____40574));
  hi1s1 ____9__505170(.DIN (__909_), .Q (____9_0__37080));
  nnd2s1 ____09_505171(.DIN1 (__90_9__29717), .DIN2 (________29021), .Q
       (__9090));
  nor2s1 _______505172(.DIN1 (________26530), .DIN2 (________29163), .Q
       (__90____29716));
  xor2s1 _______505173(.DIN1 (____0___28840), .DIN2 (_____0___36285),
       .Q (__90____29715));
  nor2s1 _______505174(.DIN1 (_________41365), .DIN2 (___9_9__29601),
       .Q (__90____29714));
  nor2s1 _______505175(.DIN1
       (_____________________________________________21857), .DIN2
       (__90____29701), .Q (__90____29713));
  nor2s1 _______505176(.DIN1 (________29040), .DIN2 (__90_0__29670), .Q
       (__90____29712));
  nnd2s1 ______505177(.DIN1 (________28995), .DIN2 (inData[22]), .Q
       (__90____29711));
  nor2s1 _______505178(.DIN1 (________29133), .DIN2 (__90_9__29708), .Q
       (__90____29710));
  or2s1 _______505179(.DIN1 (____9___29004), .DIN2 (__90_9__29708), .Q
       (__90_0__29709));
  or2s1 ______505180(.DIN1 (__9_0___30274), .DIN2 (________29159), .Q
       (__90____29707));
  nor2s1 ______505181(.DIN1 (___0____26115), .DIN2 (_____0__29155), .Q
       (__90____29706));
  nor2s1 _______505182(.DIN1 (________28329), .DIN2 (________29120), .Q
       (__90____29705));
  nor2s1 ______505183(.DIN1 (_____0__22869), .DIN2 (________29154), .Q
       (__90____29704));
  nor2s1 _____9_505184(.DIN1 (________29132), .DIN2 (__90_0__29699), .Q
       (__90____29703));
  nor2s1 _____505185(.DIN1 (___0_0___40466), .DIN2 (__90____29701), .Q
       (__90____29702));
  nor2s1 _____0_505186(.DIN1 (________29131), .DIN2 (__90_0__29699), .Q
       (__90____29700));
  nnd2s1 _______505187(.DIN1 (________29147), .DIN2 (___9_____39494),
       .Q (__90_9__29698));
  nnd2s1 _______505188(.DIN1 (_____9___34279), .DIN2 (_________22045),
       .Q (__90____29697));
  nor2s1 ______505189(.DIN1 (_________22045), .DIN2 (_____9___34279),
       .Q (__90____29696));
  and2s1 _______505190(.DIN1 (_____9__29145), .DIN2 (__9_9___30174), .Q
       (__90____29695));
  nnd2s1 _______505191(.DIN1 (___0_____40386), .DIN2 (________23118),
       .Q (__90____29694));
  nor2s1 _______505192(.DIN1 (__90____29692), .DIN2 (________29141), .Q
       (__90____29693));
  nor2s1 _______505193(.DIN1 (______0__41270), .DIN2 (________29125),
       .Q (__90____29691));
  nnd2s1 _______505194(.DIN1 (______0__33640), .DIN2
       (____________________________________________21831), .Q
       (__90____29690));
  nnd2s1 _______505195(.DIN1 (________29160), .DIN2 (__90_9__29688), .Q
       (__90_0__29689));
  nnd2s1 _______505196(.DIN1 (________29134), .DIN2 (____0___28109), .Q
       (__90____29687));
  nor2s1 _____505197(.DIN1 (________29151), .DIN2 (_____0__28981), .Q
       (__90____29686));
  nor2s1 ______505198(.DIN1
       (____________________________________________21831), .DIN2
       (______0__33640), .Q (__90____29685));
  nor2s1 _______505199(.DIN1 (___99___27825), .DIN2 (________28993), .Q
       (__90____29683));
  xor2s1 _______505200(.DIN1 (___9____28683), .DIN2
       (______________22105), .Q (__90____29682));
  nor2s1 _______505201(.DIN1 (________29269), .DIN2 (____9___29364), .Q
       (__90____29681));
  xor2s1 _______505202(.DIN1
       (__________________________________________________________________21983),
       .DIN2 (______________________________________________21904), .Q
       (__90_0__29680));
  nor2s1 _____505203(.DIN1 (____9____34365), .DIN2 (________29130), .Q
       (__90_9__29679));
  nnd2s1 _____9_505204(.DIN1 (________29148), .DIN2 (___9_____39494),
       .Q (__90____29678));
  nor2s1 _____9_505205(.DIN1 (___0_0__27855), .DIN2 (________29143), .Q
       (__90____29677));
  nor2s1 _____9_505206(.DIN1 (__90____29675), .DIN2 (__9__0__30291), .Q
       (__90____29676));
  nnd2s1 _____0_505207(.DIN1 (________29122), .DIN2 (_____9__28167), .Q
       (__90____29674));
  nnd2s1 _____0_505208(.DIN1 (________29139), .DIN2 (__90____29672), .Q
       (__90____29673));
  nnd2s1 _______505209(.DIN1 (__90_0__29670), .DIN2 (__9_____30423), .Q
       (__90____29671));
  nor2s1 ______505210(.DIN1 (__9_____29827), .DIN2 (________29150), .Q
       (__90_9__29669));
  nor2s1 ______505211(.DIN1 (________29111), .DIN2 (__9_____30401), .Q
       (__90____29668));
  nnd2s1 _______505212(.DIN1 (_____0__29127), .DIN2 (________29231), .Q
       (__90____29667));
  nnd2s1 _______505213(.DIN1 (__90____29665), .DIN2 (________29113), .Q
       (__90____29666));
  nor2s1 _______505214(.DIN1 (__90____29663), .DIN2 (_____9__29116), .Q
       (__90____29664));
  nnd2s1 _______505215(.DIN1 (__90____29661), .DIN2 (________29114), .Q
       (__90____29662));
  nor2s1 _______505216(.DIN1 (________29129), .DIN2 (________28994), .Q
       (__90_0__29660));
  nnd2s1 ______505217(.DIN1 (________29118), .DIN2 (________28593), .Q
       (__90_9__29659));
  nnd2s1 ______505218(.DIN1 (____9___29365), .DIN2 (__90____29657), .Q
       (__90____29658));
  nnd2s1 _____505219(.DIN1 (_________33030), .DIN2 (_____9__29314), .Q
       (__90____29656));
  nnd2s1 ____90_505220(.DIN1 (________29124), .DIN2 (_________36858),
       .Q (__90____29655));
  or2s1 ____09_505221(.DIN1 (__90____29651), .DIN2 (__90____29653), .Q
       (__90____29654));
  nor2s1 ____09_505222(.DIN1 (_________41132), .DIN2 (__90____29651),
       .Q (__90____29652));
  nnd2s1 ____0_505223(.DIN1 (__90_9), .DIN2 (__90____29649), .Q
       (__90_0__29650));
  nor2s1 ____0__505224(.DIN1 (________29063), .DIN2 (________28976), .Q
       (__90____29647));
  nnd2s1 ____9__505225(.DIN1 (____0___28929), .DIN2 (________29176), .Q
       (__90____29646));
  or2s1 ____9__505226(.DIN1 (inData[17]), .DIN2 (______0__36766), .Q
       (__90____29645));
  nnd2s1 ____9__505227(.DIN1 (_________37317), .DIN2 (inData[25]), .Q
       (__90__));
  nor2s1 ____9__505228(.DIN1 (________28859), .DIN2 (________28903), .Q
       (__90_0));
  nor2s1 ____9_505229(.DIN1 (________27058), .DIN2 (_____9__29082), .Q
       (__900___29644));
  nnd2s1 ____9__505230(.DIN1 (_________37223), .DIN2 (inData[21]), .Q
       (__900___29643));
  nor2s1 ____9__505231(.DIN1
       (______________________________________________21930), .DIN2
       (__900___29641), .Q (__900___29642));
  nor2s1 ____9__505232(.DIN1 (________27522), .DIN2 (______0__41092),
       .Q (__900___29640));
  nnd2s1 ____9__505233(.DIN1 (____9___29277), .DIN2 (_________41144),
       .Q (__900___29639));
  or2s1 ____9_505234(.DIN1 (__900_), .DIN2 (________29080), .Q
       (__900___29638));
  nnd2s1 ____9__505235(.DIN1 (__90____29665), .DIN2 (_________41084),
       .Q (___99___29636));
  nnd2s1 ____9__505236(.DIN1 (________29061), .DIN2 (___9____28694), .Q
       (___99___29635));
  nnd2s1 ____9__505237(.DIN1 (________29073), .DIN2 (___90___28653), .Q
       (___99___29634));
  and2s1 ____9__505238(.DIN1 (________29042), .DIN2 (___0____27848), .Q
       (___99___29633));
  nnd2s1 ____505239(.DIN1 (________29067), .DIN2 (____9___29551), .Q
       (___99___29632));
  and2s1 ____99_505240(.DIN1 (________29071), .DIN2 (________24056), .Q
       (___99___29631));
  and2s1 ____99_505241(.DIN1 (________28933), .DIN2 (___99___29629), .Q
       (___99___29630));
  and2s1 ____00_505242(.DIN1 (___9_9__29627), .DIN2 (________29420), .Q
       (___990__29628));
  nnd2s1 ____00_505243(.DIN1 (_________41146), .DIN2 (_____0__29065),
       .Q (___9____29626));
  nnd2s1 ____0_505244(.DIN1 (________27529), .DIN2 (________28945), .Q
       (___9____29625));
  nnd2s1 ____0__505245(.DIN1 (__9_9___30270), .DIN2 (_________41098),
       .Q (___9____29624));
  or2s1 ____0__505246(.DIN1 (_________41158), .DIN2 (___9____29622), .Q
       (___9____29623));
  and2s1 ____0__505247(.DIN1 (________28411), .DIN2 (________29059), .Q
       (___9____29621));
  nnd2s1 ____0__505248(.DIN1 (_____0__29055), .DIN2 (___0_____30783),
       .Q (___9_0__29620));
  nnd2s1 ____0__505249(.DIN1 (________28967), .DIN2 (___9____28665), .Q
       (___9_9__29619));
  nnd2s1 ____0__505250(.DIN1 (____99__29278), .DIN2 (________27954), .Q
       (___9____29618));
  nnd2s1 ____0__505251(.DIN1 (________29050), .DIN2 (____9___28917), .Q
       (___9____29617));
  nor2s1 ____0_505252(.DIN1 (___9____29615), .DIN2 (________29044), .Q
       (___9____29616));
  or2s1 ____0__505253(.DIN1 (___0_9___40354), .DIN2 (________29085), .Q
       (___9____29614));
  and2s1 ____0_505254(.DIN1 (_____0__28941), .DIN2 (___9_0__27805), .Q
       (___9____29613));
  nor2s1 ____0__505255(.DIN1 (___9____27780), .DIN2 (_________41098),
       .Q (___9____29612));
  nor2s1 ____0__505256(.DIN1 (____0___28377), .DIN2 (________29038), .Q
       (___9_0__29611));
  nnd2s1 ____0__505257(.DIN1 (_________41086), .DIN2 (___0____28748),
       .Q (___9_9__29610));
  or2s1 ____0_505258(.DIN1 (___9____29608), .DIN2 (_____9__29036), .Q
       (___9____29609));
  nor2s1 ____0__505259(.DIN1 (___9____29606), .DIN2 (________29035), .Q
       (___9____29607));
  and2s1 ____0__505260(.DIN1 (____9___28918), .DIN2 (________28887), .Q
       (___9____29605));
  nnd2s1 ____0__505261(.DIN1 (________29032), .DIN2 (________29171), .Q
       (___9____29604));
  or2s1 ____0__505262(.DIN1 (___9_0__29602), .DIN2 (____9___29001), .Q
       (___9____29603));
  nnd2s1 _______505263(.DIN1 (___9_9__29601), .DIN2 (_________41365),
       .Q (__9__0__30159));
  nor2s1 ____9__505264(.DIN1 (____0____32521), .DIN2 (________29109),
       .Q (__9_____30126));
  hi1s1 ____9__505265(.DIN (____9____37049), .Q (__9_____30031));
  or2s1 ____9__505266(.DIN1 (_________37317), .DIN2 (________29477), .Q
       (_________37405));
  nnd2s1 ____9_505267(.DIN1 (_________41090), .DIN2 (___9____29600), .Q
       (_________37504));
  nnd2s1 ____9_505268(.DIN1 (__90____29701), .DIN2 (____0____37165), .Q
       (_____9___36996));
  nor2s1 _____0_505269(.DIN1 (________29354), .DIN2 (_____0__29075), .Q
       (___9____29599));
  nnd2s1 _____0_505270(.DIN1 (____00__28924), .DIN2 (___9____29597), .Q
       (___9____29598));
  nnd2s1 _____0_505271(.DIN1 (________29077), .DIN2 (___0_____30783),
       .Q (___9____29596));
  or2s1 _____0_505272(.DIN1 (________26637), .DIN2 (____09__29018), .Q
       (___9____29595));
  and2s1 _______505273(.DIN1 (____0___29016), .DIN2 (_____0__27419), .Q
       (___9____29594));
  nnd2s1 _______505274(.DIN1 (__90_9__29717), .DIN2 (_____9__29091), .Q
       (___9_0__29593));
  nor2s1 _______505275(.DIN1 (________28977), .DIN2 (__9__0__30291), .Q
       (___9____29591));
  nnd2s1 ______505276(.DIN1 (_____9__27471), .DIN2 (____9___29094), .Q
       (___9____29589));
  or2s1 _______505277(.DIN1 (____0___29200), .DIN2 (_____9__29054), .Q
       (___9____29588));
  nnd2s1 _______505278(.DIN1 (__9_9___30270), .DIN2 (________29060), .Q
       (___9____29587));
  or2s1 _______505279(.DIN1 (___9____29608), .DIN2 (________28997), .Q
       (___9_0__29586));
  nor2s1 _______505280(.DIN1 (___9____29584), .DIN2 (_____9__29135), .Q
       (___9_9__29585));
  and2s1 _______505281(.DIN1 (_____0__29136), .DIN2 (___0_09__30651),
       .Q (___9____29583));
  and2s1 _______505282(.DIN1 (_________41096), .DIN2 (________28483),
       .Q (___9____29582));
  nor2s1 ______505283(.DIN1 (___9____29580), .DIN2 (________29137), .Q
       (___9____29581));
  or2s1 ______505284(.DIN1 (___9____29578), .DIN2 (________29167), .Q
       (___9____29579));
  nor2s1 ____9__505285(.DIN1 (________27079), .DIN2 (________28983), .Q
       (___9____29577));
  nnd2s1 ____9__505286(.DIN1 (_____0__28990), .DIN2 (_____0__29495), .Q
       (___9_0__29576));
  and2s1 _____9_505287(.DIN1 (________28984), .DIN2 (___9____29574), .Q
       (___9____29575));
  or2s1 _____505288(.DIN1 (___9____29571), .DIN2 (____0___29099), .Q
       (___9____29572));
  nor2s1 _____0_505289(.DIN1 (_____0__27706), .DIN2 (_________32982),
       .Q (___9_0__29570));
  nnd2s1 _______505290(.DIN1 (___099__28833), .DIN2 (________28944), .Q
       (___9_9__29569));
  nnd2s1 _______505291(.DIN1 (____0___28928), .DIN2 (____90__28637), .Q
       (___9____29568));
  nnd2s1 _______505292(.DIN1 (________29034), .DIN2 (________27538), .Q
       (___9____29567));
  nor2s1 _______505293(.DIN1 (________27974), .DIN2 (_____9__29064), .Q
       (___9____29566));
  nor2s1 _______505294(.DIN1 (_____9___34186), .DIN2 (________28970),
       .Q (___9____29565));
  nnd2s1 ______505295(.DIN1 (_________34136), .DIN2 (__99____30501), .Q
       (___9____29564));
  nnd2s1 _______505296(.DIN1 (________28913), .DIN2 (inData[12]), .Q
       (___9____29563));
  nnd2s1 _______505297(.DIN1 (_________41088), .DIN2 (________28074),
       .Q (___9____29562));
  nnd2s1 _______505298(.DIN1 (________28948), .DIN2 (_________37722),
       .Q (___909__29561));
  nor2s1 _______505299(.DIN1 (___9_0__26920), .DIN2 (___90___29559), .Q
       (___90___29560));
  nnd2s1 _______505300(.DIN1 (________27152), .DIN2 (_____9__28956), .Q
       (___90___29558));
  nnd2s1 _______505301(.DIN1 (_____0__28973), .DIN2 (inData[10]), .Q
       (___90___29557));
  nor2s1 _______505302(.DIN1 (________22575), .DIN2 (_________37317),
       .Q (___90___29556));
  and2s1 ______505303(.DIN1 (________28953), .DIN2 (__99____30513), .Q
       (___90___29555));
  nor2s1 ______505304(.DIN1 (________27053), .DIN2 (____00__29097), .Q
       (___90___29554));
  nnd2s1 ______505305(.DIN1 (____9___29551), .DIN2 (________29069), .Q
       (____99__29552));
  nnd2s1 _____505306(.DIN1 (____9___29548), .DIN2 (___09____40684), .Q
       (____9___29550));
  nnd2s1 _____9_505307(.DIN1 (____9___29548), .DIN2 (___9____28719), .Q
       (____9___29549));
  nnd2s1 _____9_505308(.DIN1 (________28971), .DIN2 (________29208), .Q
       (____9___29547));
  nor2s1 _____9_505309(.DIN1 (_________37320), .DIN2 (_________37317),
       .Q (____9___29546));
  or2s1 _____9_505310(.DIN1 (____9___29544), .DIN2 (________29024), .Q
       (____9___29545));
  and2s1 _____505311(.DIN1 (________29513), .DIN2 (_____9__29542), .Q
       (____90__29543));
  nor2s1 _____0_505312(.DIN1 (________28902), .DIN2 (________28943), .Q
       (________29541));
  or2s1 _____505313(.DIN1 (____0___27658), .DIN2 (________29019), .Q
       (________29540));
  or2s1 _______505314(.DIN1 (_________31836), .DIN2 (________28962), .Q
       (________29539));
  nnd2s1 ______505315(.DIN1 (________28901), .DIN2 (________29537), .Q
       (________29538));
  nor2s1 _______505316(.DIN1 (___09_9__31465), .DIN2 (____9___28921),
       .Q (________29536));
  or2s1 _______505317(.DIN1 (_____0__29534), .DIN2 (________29062), .Q
       (________29535));
  or2s1 _______505318(.DIN1 (____0___29013), .DIN2 (___9____29622), .Q
       (________29532));
  or2s1 _______505319(.DIN1 (________29529), .DIN2 (_________41094), .Q
       (________29530));
  nor2s1 _______505320(.DIN1 (_____9___31886), .DIN2 (________29041),
       .Q (________29528));
  nnd2s1 _______505321(.DIN1 (________28899), .DIN2 (________28987), .Q
       (_____0__29527));
  nnd2s1 _______505322(.DIN1 (____9___28916), .DIN2 (________29525), .Q
       (_____9__29526));
  nnd2s1 _______505323(.DIN1 (________28904), .DIN2 (________29523), .Q
       (________29524));
  nnd2s1 _______505324(.DIN1 (________28910), .DIN2 (____0___29285), .Q
       (________29522));
  nor2s1 _______505325(.DIN1 (__9_____30417), .DIN2 (________28951), .Q
       (________29521));
  nor2s1 _______505326(.DIN1 (________29519), .DIN2 (________28907), .Q
       (________29520));
  or2s1 _______505327(.DIN1 (_________31817), .DIN2 (_____0__28932), .Q
       (________29518));
  nor2s1 ______505328(.DIN1 (____9____32449), .DIN2 (_____0__28906), .Q
       (________29517));
  and2s1 _______505329(.DIN1 (________29515), .DIN2 (________28592), .Q
       (________29516));
  nor2s1 _______505330(.DIN1 (________29513), .DIN2 (__9_____30401), .Q
       (________29514));
  nnd2s1 _______505331(.DIN1 (_____9__28880), .DIN2 (________29511), .Q
       (________29512));
  nor2s1 ______505332(.DIN1 (________28878), .DIN2 (________29505), .Q
       (_____0__29510));
  nor2s1 _______505333(.DIN1 (________29508), .DIN2 (________28988), .Q
       (_____9__29509));
  nor2s1 _____9_505334(.DIN1 (________27554), .DIN2 (________28884), .Q
       (________29507));
  nnd2s1 _______505335(.DIN1 (________29505), .DIN2 (__9_____30019), .Q
       (________29506));
  or2s1 _______505336(.DIN1 (____9____32439), .DIN2 (________28978), .Q
       (________29504));
  nor2s1 _______505337(.DIN1 (___0_____31262), .DIN2 (________28885),
       .Q (_____0__29503));
  nnd2s1 _______505338(.DIN1 (________28888), .DIN2 (________29501), .Q
       (_____9__29502));
  nor2s1 _______505339(.DIN1 (____0____31547), .DIN2 (________29216),
       .Q (__9_____30049));
  nor2s1 ____0__505340(.DIN1 (________26714), .DIN2 (________29499), .Q
       (__9_____30051));
  nnd2s1 _______505341(.DIN1 (________29089), .DIN2 (________29498), .Q
       (__9_____30007));
  nor2s1 ______505342(.DIN1 (_____0__28947), .DIN2 (________28584), .Q
       (____9____32413));
  and2s1 _____505343(.DIN1 (________28938), .DIN2 (___0_____30917), .Q
       (__9_0___29994));
  xor2s1 _____9_505344(.DIN1 (________29497), .DIN2 (_________38203),
       .Q (__9_0___29997));
  nnd2s1 _______505345(.DIN1 (________29020), .DIN2 (________27421), .Q
       (__909_));
  nor2s1 _______505346(.DIN1 (___00___28744), .DIN2 (_____9__29045), .Q
       (__9_0___30085));
  nor2s1 _______505347(.DIN1 (___099___31496), .DIN2 (____0___29014),
       .Q (__9_9___30079));
  nor2s1 _______505348(.DIN1 (___0__9__30890), .DIN2 (________29177),
       .Q (_____9___32771));
  nnd2s1 ______505349(.DIN1 (_________34136), .DIN2 (______0__41260),
       .Q (____9_9__34346));
  nnd2s1 ______505350(.DIN1 (___0_____30870), .DIN2 (___0__0__31290),
       .Q (_____0___31991));
  dffacs1 _______________________________________505351(.CLRB (reset),
       .CLK (clk), .DIN (________29161), .Q (______________22104));
  nnd2s1 ______505352(.DIN1 (________28599), .DIN2 (________27726), .Q
       (________29496));
  nor2s1 _______505353(.DIN1 (_____9__26437), .DIN2 (________29490), .Q
       (________29493));
  nor2s1 ______505354(.DIN1 (________29326), .DIN2 (________28856), .Q
       (________29492));
  nor2s1 _____9_505355(.DIN1 (_____9__27731), .DIN2 (________29490), .Q
       (________29491));
  and2s1 _____9_505356(.DIN1 (_____9__28853), .DIN2 (__90____29661), .Q
       (________29489));
  nor2s1 _______505357(.DIN1 (_________31667), .DIN2 (________28619),
       .Q (________29488));
  hi1s1 _______505358(.DIN (___0_____31247), .Q (________29487));
  nor2s1 _______505359(.DIN1 (________27520), .DIN2 (________29490), .Q
       (_____0__29486));
  nor2s1 _______505360(.DIN1 (________28131), .DIN2 (_____0__28854), .Q
       (_____9__29485));
  nor2s1 ______505361(.DIN1 (___0_____30709), .DIN2 (________28847), .Q
       (________29484));
  nor2s1 _____505362(.DIN1 (________28846), .DIN2 (____99__29008), .Q
       (________29483));
  nnd2s1 _______505363(.DIN1 (__90____29661), .DIN2 (____0___28842), .Q
       (________29482));
  nnd2s1 _______505364(.DIN1 (____0___28841), .DIN2 (________28494), .Q
       (________29481));
  xor2s1 ____9__505365(.DIN1 (________29153), .DIN2 (_________35084),
       .Q (________29480));
  nnd2s1 _______505366(.DIN1 (_____9__27471), .DIN2 (________28601), .Q
       (________29479));
  hi1s1 ____9__505367(.DIN (________29477), .Q (________29478));
  or2s1 ____9__505368(.DIN1 (___9____29580), .DIN2 (___9____28725), .Q
       (_____0__29476));
  nor2s1 ____9_505369(.DIN1 (___0_____40419), .DIN2 (___0_____40166),
       .Q (____09__29475));
  nnd2s1 ____9__505370(.DIN1 (___00___28743), .DIN2 (____0___29015), .Q
       (____0___29474));
  nor2s1 ____9__505371(.DIN1 (___9____27789), .DIN2 (___9____28656), .Q
       (____0___29473));
  nor2s1 ____9__505372(.DIN1 (___0_9__28824), .DIN2 (____0___29471), .Q
       (____0___29472));
  nor2s1 ____9__505373(.DIN1 (___0____28816), .DIN2 (________29313), .Q
       (____0___29470));
  nor2s1 ____9__505374(.DIN1 (____0____31589), .DIN2 (___0_0__28815),
       .Q (____0___29469));
  and2s1 ____9__505375(.DIN1 (____0___29467), .DIN2 (__9_____30255), .Q
       (____0___29468));
  nor2s1 ____9__505376(.DIN1 (___0____28813), .DIN2 (__9_____29862), .Q
       (____00__29466));
  nor2s1 ____9_505377(.DIN1 (___0____28812), .DIN2 (________27172), .Q
       (____99__29465));
  nnd2s1 ____9__505378(.DIN1 (___0____28808), .DIN2 (____9___29463), .Q
       (____9___29464));
  nor2s1 ____9__505379(.DIN1 (________26561), .DIN2 (___0____28807), .Q
       (____9___29462));
  nnd2s1 ____9_505380(.DIN1 (___0____28803), .DIN2 (_____90__35555), .Q
       (____9___29461));
  nor2s1 ____99_505381(.DIN1 (________29072), .DIN2 (___0____28802), .Q
       (____9___29460));
  or2s1 ____99_505382(.DIN1 (____9___29458), .DIN2 (___09___28832), .Q
       (____9___29459));
  nnd2s1 ____99_505383(.DIN1 (___9____28711), .DIN2 (_________31933),
       .Q (____9___29457));
  nnd2s1 ____99_505384(.DIN1 (___9____28690), .DIN2 (_____9__29455), .Q
       (____90__29456));
  nnd2s1 ____505385(.DIN1 (___0____28799), .DIN2 (___0____26123), .Q
       (________29454));
  or2s1 ____505386(.DIN1 (________29452), .DIN2 (__9_____29862), .Q
       (________29453));
  nnd2s1 ____00_505387(.DIN1 (__90____29665), .DIN2 (________29450), .Q
       (________29451));
  nnd2s1 ____00_505388(.DIN1 (___0____28789), .DIN2 (_____9___33329),
       .Q (________29449));
  nor2s1 ____505389(.DIN1 (________29447), .DIN2 (__9_____29862), .Q
       (________29448));
  and2s1 ____0__505390(.DIN1 (_____0__28618), .DIN2 (___0____26130), .Q
       (_____0__29446));
  nor2s1 ____0__505391(.DIN1 (_________32001), .DIN2 (___0_0__28786),
       .Q (_____9__29445));
  nor2s1 ____0__505392(.DIN1 (___0____27860), .DIN2 (___0____28749), .Q
       (________29444));
  nnd2s1 ____0__505393(.DIN1 (___0____28769), .DIN2 (__9_99__29992), .Q
       (________29443));
  and2s1 ____0__505394(.DIN1 (___0____28780), .DIN2 (________29441), .Q
       (________29442));
  nnd2s1 ____0__505395(.DIN1 (___0____28747), .DIN2 (________29439), .Q
       (________29440));
  nor2s1 ____0__505396(.DIN1 (__99_9__30508), .DIN2 (____0___28835), .Q
       (________29438));
  nor2s1 ____0_505397(.DIN1 (___0_____30977), .DIN2 (___0____28774), .Q
       (________29437));
  nor2s1 ____0__505398(.DIN1 (__9_____29783), .DIN2 (___0____28772), .Q
       (_____0__29436));
  or2s1 ____0__505399(.DIN1 (___0_____30986), .DIN2 (___0____28770), .Q
       (_____9__29435));
  nor2s1 ____0__505400(.DIN1 (_____9__27344), .DIN2 (_____90__41100),
       .Q (________29434));
  nor2s1 ____0__505401(.DIN1 (___0_____30695), .DIN2 (_____9___41106),
       .Q (________29433));
  nor2s1 ____0__505402(.DIN1 (________29431), .DIN2 (____9___29092), .Q
       (________29432));
  nor2s1 ____0__505403(.DIN1
       (_________________________________________9___21929), .DIN2
       (_____________________________________________21928), .Q
       (________29430));
  and2s1 ____0__505404(.DIN1 (___0____28768), .DIN2 (________29428), .Q
       (________29429));
  nnd2s1 ____0__505405(.DIN1 (___0_0__28766), .DIN2 (___0____27847), .Q
       (________29427));
  and2s1 ____0__505406(.DIN1 (___0____28764), .DIN2 (_____9__29425), .Q
       (_____0__29426));
  or2s1 ____0_505407(.DIN1 (___0_9___31111), .DIN2 (___0____28759), .Q
       (________29424));
  or2s1 ____0_505408(.DIN1 (_________33106), .DIN2 (___0_9__28755), .Q
       (________29423));
  nor2s1 ____0__505409(.DIN1 (___0__9__31147), .DIN2 (___0____28751),
       .Q (________29422));
  and2s1 ____0__505410(.DIN1 (___0____28752), .DIN2 (________26732), .Q
       (________29421));
  and2s1 ____09_505411(.DIN1 (___9____28669), .DIN2 (________28942), .Q
       (________29419));
  nnd2s1 ____09_505412(.DIN1 (___0_0__28746), .DIN2 (_____0__29417), .Q
       (________29418));
  or2s1 ____09_505413(.DIN1 (________29415), .DIN2 (___0____28767), .Q
       (_____9__29416));
  nnd2s1 ____505414(.DIN1 (___9____28706), .DIN2 (________29166), .Q
       (________29414));
  and2s1 _____0_505415(.DIN1 (___09___28828), .DIN2 (___99___28730), .Q
       (________29413));
  nor2s1 _____0_505416(.DIN1 (___0____28763), .DIN2 (___00___28742), .Q
       (________29412));
  nor2s1 _____0_505417(.DIN1 (____9____32449), .DIN2 (___00___28739),
       .Q (________29411));
  or2s1 _____0_505418(.DIN1 (________29409), .DIN2 (___00___28738), .Q
       (________29410));
  and2s1 _____0_505419(.DIN1 (___000__28736), .DIN2 (_____0__29407), .Q
       (________29408));
  nnd2s1 _____505420(.DIN1 (___9_0__28708), .DIN2 (________29405), .Q
       (_____9__29406));
  nor2s1 ____00_505421(.DIN1 (____0___27214), .DIN2 (___0____28810), .Q
       (________29404));
  nnd2s1 _______505422(.DIN1 (___99___28733), .DIN2 (___9____27769), .Q
       (________29403));
  nor2s1 _______505423(.DIN1 (_____9___41102), .DIN2 (__9_____30401),
       .Q (________29402));
  or2s1 _______505424(.DIN1 (__9__9__30073), .DIN2 (_____9___41104), .Q
       (________29401));
  nnd2s1 _______505425(.DIN1 (___99___28729), .DIN2 (___9____29592), .Q
       (________29400));
  nnd2s1 ______505426(.DIN1
       (_____________________________________________21928), .DIN2
       (_________________________________________9___21929), .Q
       (________29399));
  nor2s1 _______505427(.DIN1 (__9_____29750), .DIN2 (_____0___41112),
       .Q (________29398));
  nor2s1 ______505428(.DIN1 (___0_____30669), .DIN2 (___9____28723), .Q
       (_____0__29397));
  nnd2s1 _______505429(.DIN1 (_____0__28571), .DIN2 (________29395), .Q
       (_____9__29396));
  and2s1 _______505430(.DIN1 (___0____28800), .DIN2 (________29393), .Q
       (________29394));
  nor2s1 _______505431(.DIN1 (________28263), .DIN2 (___9____28721), .Q
       (________29392));
  nor2s1 _______505432(.DIN1 (________26441), .DIN2 (___9____28720), .Q
       (________29391));
  nnd2s1 _______505433(.DIN1 (________28980), .DIN2 (________29389), .Q
       (________29390));
  and2s1 _______505434(.DIN1 (___9____28713), .DIN2 (_________33020),
       .Q (________29388));
  or2s1 _______505435(.DIN1 (_____9__29386), .DIN2 (___0_0__28756), .Q
       (_____0__29387));
  or2s1 _______505436(.DIN1 (________29384), .DIN2 (___9_9__28707), .Q
       (________29385));
  nor2s1 _______505437(.DIN1 (___0_0___31125), .DIN2 (___0____28787),
       .Q (________29383));
  nnd2s1 _______505438(.DIN1 (___9_0__28718), .DIN2 (_____9__29295), .Q
       (________29382));
  nnd2s1 _______505439(.DIN1 (___9_9__28717), .DIN2 (_________31935),
       .Q (________29381));
  and2s1 ______505440(.DIN1 (___9____28699), .DIN2 (________29379), .Q
       (________29380));
  and2s1 _______505441(.DIN1 (____09__29377), .DIN2 (___9____27796), .Q
       (_____0__29378));
  nnd2s1 _______505442(.DIN1 (___0_9__28775), .DIN2 (____90__29272), .Q
       (____0___29376));
  nor2s1 ______505443(.DIN1 (____0___29374), .DIN2 (___9____28700), .Q
       (____0___29375));
  nor2s1 _____0_505444(.DIN1 (___9____28677), .DIN2 (____0___29372), .Q
       (____0___29373));
  nnd2s1 _____0_505445(.DIN1 (________28621), .DIN2 (__9_____30019), .Q
       (____0___29371));
  nor2s1 _____9_505446(.DIN1 (________28632), .DIN2 (___0____27856), .Q
       (____0___29370));
  nnd2s1 _____9_505447(.DIN1 (_____9__28607), .DIN2 (___0____27889), .Q
       (____00__29369));
  nnd2s1 _______505448(.DIN1 (___9____28714), .DIN2 (____9___29367), .Q
       (____99__29368));
  nor2s1 _______505449(.DIN1 (________28273), .DIN2 (________28623), .Q
       (____9___29366));
  nor2s1 _______505450(.DIN1 (________28574), .DIN2 (____9___28643), .Q
       (____9___29363));
  nnd2s1 _____9_505451(.DIN1 (________29361), .DIN2 (___0____28778), .Q
       (_____9__29362));
  or2s1 _____0_505452(.DIN1 (________29359), .DIN2 (_____9__28598), .Q
       (________29360));
  nnd2s1 _____0_505453(.DIN1 (__9_9___30270), .DIN2 (________29349), .Q
       (________29358));
  nor2s1 _____505454(.DIN1 (________27998), .DIN2 (___0____28821), .Q
       (________29357));
  and2s1 ______505455(.DIN1 (___0____28750), .DIN2 (________29523), .Q
       (________29356));
  nor2s1 _______505456(.DIN1 (________29354), .DIN2 (___9_0__28681), .Q
       (________29355));
  nor2s1 _______505457(.DIN1 (________27333), .DIN2 (_____9__29334), .Q
       (_____0__29353));
  or2s1 _______505458(.DIN1 (________28486), .DIN2 (_________41126), .Q
       (_____9__29352));
  nnd2s1 _______505459(.DIN1 (____0___28836), .DIN2 (_____0___41313),
       .Q (________29351));
  nor2s1 _______505460(.DIN1 (________28125), .DIN2 (________29349), .Q
       (________29350));
  nor2s1 _______505461(.DIN1 (___0____28818), .DIN2 (___0_9__28804), .Q
       (________29348));
  nor2s1 _______505462(.DIN1 (___9____28658), .DIN2 (________27172), .Q
       (________29347));
  nnd2s1 _______505463(.DIN1 (________28577), .DIN2 (___9____28666), .Q
       (________29346));
  nnd2s1 _______505464(.DIN1 (___9____28659), .DIN2 (________27989), .Q
       (_____0__29345));
  nnd2s1 ______505465(.DIN1 (________29342), .DIN2 (________27614), .Q
       (_____9__29344));
  and2s1 ______505466(.DIN1 (________29342), .DIN2 (________29341), .Q
       (________29343));
  nor2s1 _______505467(.DIN1 (_____00__34847), .DIN2 (___9_9__28672),
       .Q (________29340));
  and2s1 _______505468(.DIN1 (____0___28383), .DIN2 (________29338), .Q
       (________29339));
  or2s1 _______505469(.DIN1 (________29336), .DIN2 (_____0___41116), .Q
       (________29337));
  nor2s1 _______505470(.DIN1 (___9____28710), .DIN2 (_____9__29334), .Q
       (_____0__29335));
  nor2s1 _______505471(.DIN1 (________28609), .DIN2 (________27985), .Q
       (________29333));
  nnd2s1 _______505472(.DIN1 (________28606), .DIN2 (________27545), .Q
       (________29332));
  nnd2s1 _______505473(.DIN1 (________28858), .DIN2 (________27694), .Q
       (__90____29648));
  nnd2s1 _______505474(.DIN1 (_____0__28844), .DIN2 (_____0__28481), .Q
       (__9__9__29984));
  xor2s1 ____9__505475(.DIN1 (______________22109), .DIN2
       (___0_____40585), .Q (__90____29684));
  nnd2s1 _______505476(.DIN1 (___009__28745), .DIN2 (________29331), .Q
       (__9_____29855));
  nor2s1 _______505477(.DIN1 (___0____26114), .DIN2 (___0____28823), .Q
       (__9_____29863));
  nor2s1 ______505478(.DIN1 (_________22038), .DIN2 (___00___28740), .Q
       (__9_____29970));
  or2s1 ______505479(.DIN1 (________28961), .DIN2 (___0____28794), .Q
       (__9_____29914));
  nor2s1 _______505480(.DIN1 (___09___28830), .DIN2 (________27594), .Q
       (_________32738));
  nnd2s1 _______505481(.DIN1 (____0____35363), .DIN2 (______0__35537),
       .Q (____9____35254));
  nnd2s1 _______505482(.DIN1 (____0___28837), .DIN2 (____9___29006), .Q
       (___0_____40376));
  dffacs1 ____________________________________9_505483(.CLRB (reset),
       .CLK (clk), .DIN (___0____28809), .Q (___0_____40583));
  hi1s1 _____9_505484(.DIN (_________41090), .Q (_________37414));
  nor2s1 _______505485(.DIN1 (________28860), .DIN2 (___09___28826), .Q
       (____9____37049));
  nnd2s1 _______505486(.DIN1 (________28517), .DIN2 (__9_____29758), .Q
       (________29330));
  nor2s1 _______505487(.DIN1 (________28624), .DIN2 (________28968), .Q
       (________29329));
  nor2s1 ______505488(.DIN1 (________28603), .DIN2 (________27149), .Q
       (________29328));
  nor2s1 ______505489(.DIN1 (________29326), .DIN2 (___9____28687), .Q
       (________29327));
  nor2s1 _______505490(.DIN1 (_________41152), .DIN2 (___9_9__28680),
       .Q (_____0__29325));
  nnd2s1 ______505491(.DIN1 (________29323), .DIN2 (________28595), .Q
       (_____9__29324));
  nnd2s1 _______505492(.DIN1 (________29321), .DIN2 (__9_____30423), .Q
       (________29322));
  nor2s1 _______505493(.DIN1 (________29319), .DIN2 (___9____28701), .Q
       (________29320));
  and2s1 ______505494(.DIN1 (________28576), .DIN2 (__9_____30162), .Q
       (________29318));
  and2s1 _______505495(.DIN1 (________28611), .DIN2 (__9_____30162), .Q
       (________29317));
  or2s1 _______505496(.DIN1 (___0____22331), .DIN2 (___0_____40166), .Q
       (________29316));
  nnd2s1 _______505497(.DIN1 (_____9__29314), .DIN2 (________29313), .Q
       (_____0__29315));
  nnd2s1 ______505498(.DIN1 (________28575), .DIN2 (________29311), .Q
       (________29312));
  nnd2s1 ______505499(.DIN1 (___9____28697), .DIN2 (________29309), .Q
       (________29310));
  nnd2s1 _______505500(.DIN1 (________29307), .DIN2 (__90____29665), .Q
       (________29308));
  or2s1 _______505501(.DIN1 (_____0__29305), .DIN2 (_____9__28590), .Q
       (________29306));
  nor2s1 _______505502(.DIN1 (_____00__41110), .DIN2 (________27172),
       .Q (_____9__29304));
  or2s1 _______505503(.DIN1 (___0_____30760), .DIN2 (________28586), .Q
       (________29303));
  nnd2s1 ______505504(.DIN1 (_____0___41118), .DIN2 (__90____29665), .Q
       (________29302));
  and2s1 _______505505(.DIN1 (____9___29551), .DIN2 (________29300), .Q
       (________29301));
  nnd2s1 _______505506(.DIN1 (________28620), .DIN2 (__9990), .Q
       (________29299));
  or2s1 _____505507(.DIN1 (__9__0__30291), .DIN2 (________29297), .Q
       (________29298));
  nnd2s1 _____9_505508(.DIN1 (_____9__29295), .DIN2 (___9____28691), .Q
       (_____0__29296));
  nor2s1 _____9_505509(.DIN1 (___9____28695), .DIN2 (________27149), .Q
       (________29294));
  xor2s1 ____0__505510(.DIN1 (___0_0___40566), .DIN2
       (__________________________________9__________), .Q
       (________29292));
  nor2s1 ____99_505511(.DIN1 (________26312), .DIN2 (________29241), .Q
       (________29291));
  xor2s1 _____0_505512(.DIN1 (_________36087), .DIN2 (___00____39929),
       .Q (________29290));
  nor2s1 ____99_505513(.DIN1 (__999___30539), .DIN2 (______0__41120),
       .Q (________29289));
  nor2s1 ____505514(.DIN1 (________28566), .DIN2 (___0_____31229), .Q
       (_____0__29288));
  nnd2s1 ____9_505515(.DIN1 (____0___28559), .DIN2 (________27528), .Q
       (____09__29287));
  nnd2s1 ____9__505516(.DIN1 (____0___28557), .DIN2 (____0___29285), .Q
       (____0___29286));
  nnd2s1 ____9__505517(.DIN1 (____0___29280), .DIN2 (____0___29283), .Q
       (____0___29284));
  nnd2s1 ____9__505518(.DIN1 (________28498), .DIN2 (_____9__28360), .Q
       (____0___29282));
  nnd2s1 ____9__505519(.DIN1 (____0___29280), .DIN2 (________27509), .Q
       (____0___29281));
  hi1s1 _______505520(.DIN (____99__29278), .Q (____00__29279));
  nnd2s1 _______505521(.DIN1 (____9___28549), .DIN2 (___0_____40602),
       .Q (____9___29276));
  nnd2s1 _______505522(.DIN1 (________28545), .DIN2 (______9__22030),
       .Q (____9___29275));
  nnd2s1 _______505523(.DIN1 (____9___29273), .DIN2 (___0__0__40581),
       .Q (____9___29274));
  nor2s1 _______505524(.DIN1 (__9__0__30120), .DIN2 (_____9__28529), .Q
       (_____9__29271));
  or2s1 _______505525(.DIN1 (________29269), .DIN2 (________29268), .Q
       (________29270));
  nnd2s1 _____0_505526(.DIN1 (____0___29280), .DIN2 (____0___27305), .Q
       (________29267));
  nor2s1 _______505527(.DIN1 (____9___28192), .DIN2 (________28521), .Q
       (________29266));
  or2s1 _______505528(.DIN1 (________29264), .DIN2 (____9___28552), .Q
       (________29265));
  nor2s1 _______505529(.DIN1 (_____0__29262), .DIN2 (_____9__28501), .Q
       (________29263));
  nnd2s1 _______505530(.DIN1 (_____0__28520), .DIN2 (____0___27483), .Q
       (_____9__29261));
  nor2s1 _______505531(.DIN1 (__90____29663), .DIN2 (________29259), .Q
       (________29260));
  nnd2s1 ______505532(.DIN1 (________29172), .DIN2 (____0___28382), .Q
       (________29258));
  or2s1 _______505533(.DIN1 (________29256), .DIN2 (________28516), .Q
       (________29257));
  nor2s1 _______505534(.DIN1 (___9____29615), .DIN2 (____00__29194), .Q
       (________29255));
  and2s1 _______505535(.DIN1 (_____0__28511), .DIN2 (________29253), .Q
       (________29254));
  nor2s1 _______505536(.DIN1 (__9_____29742), .DIN2 (________29251), .Q
       (_____9__29252));
  or2s1 _______505537(.DIN1 (________29249), .DIN2 (_________41122), .Q
       (________29250));
  nnd2s1 _______505538(.DIN1 (____0___29280), .DIN2 (________27314), .Q
       (________29248));
  nnd2s1 _______505539(.DIN1 (________29259), .DIN2 (________29246), .Q
       (________29247));
  and2s1 _______505540(.DIN1 (_____9__28510), .DIN2 (________29361), .Q
       (________29245));
  nor2s1 _____9_505541(.DIN1 (___9_9__26929), .DIN2 (________28524), .Q
       (_____9__29244));
  nor2s1 _____9_505542(.DIN1 (________29242), .DIN2 (________29241), .Q
       (________29243));
  nnd2s1 _____0_505543(.DIN1 (____0___29198), .DIN2 (________28388), .Q
       (________29240));
  and2s1 _____505544(.DIN1 (________29323), .DIN2 (________29238), .Q
       (________29239));
  nor2s1 _______505545(.DIN1 (________29236), .DIN2 (________28503), .Q
       (________29237));
  nnd2s1 _______505546(.DIN1 (________29323), .DIN2 (___9____28703), .Q
       (_____0__29235));
  nor2s1 ______505547(.DIN1 (________29233), .DIN2 (________28568), .Q
       (_____9__29234));
  and2s1 _______505548(.DIN1 (________28512), .DIN2 (________29231), .Q
       (________29232));
  nor2s1 _______505549(.DIN1 (________28604), .DIN2 (__9_____29862), .Q
       (________29230));
  nor2s1 _______505550(.DIN1 (________27616), .DIN2 (________28515), .Q
       (________29228));
  or2s1 _____9_505551(.DIN1 (________29225), .DIN2 (_________41124), .Q
       (________29226));
  nnd2s1 _____505552(.DIN1 (____0___28554), .DIN2 (________29223), .Q
       (________29224));
  nor2s1 _______505553(.DIN1 (________29221), .DIN2 (________29220), .Q
       (________29222));
  nor2s1 ____9__505554(.DIN1 (________28522), .DIN2 (_____9__29218), .Q
       (_____0__29219));
  nnd2s1 ____9__505555(.DIN1 (________29323), .DIN2 (___0____27872), .Q
       (________29215));
  nnd2s1 _______505556(.DIN1 (________28499), .DIN2 (_____0__29213), .Q
       (________29214));
  nnd2s1 _______505557(.DIN1 (________28506), .DIN2 (___0____26095), .Q
       (________29212));
  nor2s1 _______505558(.DIN1 (________29210), .DIN2 (________28496), .Q
       (________29211));
  nor2s1 _____505559(.DIN1 (________29208), .DIN2 (________29241), .Q
       (________29209));
  nnd2s1 _____9_505560(.DIN1 (________28539), .DIN2 (________27505), .Q
       (________29207));
  or2s1 _____9_505561(.DIN1 (________27429), .DIN2 (________29205), .Q
       (________29206));
  or2s1 _____9_505562(.DIN1 (_____9__27185), .DIN2 (________29241), .Q
       (_____0__29204));
  or2s1 _____9_505563(.DIN1 (____0___29202), .DIN2 (_____0___41114), .Q
       (____09__29203));
  nor2s1 _______505564(.DIN1 (____0___29200), .DIN2 (________28544), .Q
       (____0___29201));
  nnd2s1 _______505565(.DIN1 (____0___29198), .DIN2 (________28163), .Q
       (____0___29199));
  nor2s1 _______505566(.DIN1 (________27540), .DIN2 (________29241), .Q
       (____0___29197));
  nnd2s1 _______505567(.DIN1 (____0___29280), .DIN2 (___0____26978), .Q
       (____0___29196));
  or2s1 _______505568(.DIN1 (__9__9__29743), .DIN2 (____00__29194), .Q
       (____0___29195));
  nor2s1 _______505569(.DIN1 (________27169), .DIN2 (________29178), .Q
       (____99__29193));
  nor2s1 _______505570(.DIN1 (____0_9__31542), .DIN2 (________29268),
       .Q (____9___29192));
  or2s1 _______505571(.DIN1 (____9___29190), .DIN2 (________29241), .Q
       (____9___29191));
  or2s1 ______505572(.DIN1 (____0___28295), .DIN2 (________28542), .Q
       (____9___29189));
  nnd2s1 _______505573(.DIN1 (____0___29280), .DIN2 (________28212), .Q
       (____9___29188));
  nnd2s1 _______505574(.DIN1 (________28877), .DIN2 (____0___28475), .Q
       (____9___29187));
  and2s1 ____90_505575(.DIN1 (_____0__28890), .DIN2 (___9____28709), .Q
       (____9___29186));
  or2s1 ____9__505576(.DIN1 (___9____29608), .DIN2 (________28536), .Q
       (____90__29185));
  nor2s1 ____9__505577(.DIN1 (___9_0__27786), .DIN2 (________29183), .Q
       (_____9__29184));
  nor2s1 ____9_505578(.DIN1 (________29181), .DIN2 (________29241), .Q
       (________29182));
  nnd2s1 ____9__505579(.DIN1 (________29323), .DIN2 (________27328), .Q
       (________29180));
  nor2s1 ____9_505580(.DIN1 (___0____27877), .DIN2 (________29178), .Q
       (________29179));
  nor2s1 _____9_505581(.DIN1 (___0_____31262), .DIN2 (________28629),
       .Q (__9_____29876));
  hi1s1 ______505582(.DIN (________29177), .Q (__9_0___29805));
  nnd2s1 _____9_505583(.DIN1 (________28531), .DIN2 (________29176), .Q
       (__9_9___29799));
  or2s1 _______505584(.DIN1 (__9__9__30225), .DIN2 (____9___29273), .Q
       (_________38534));
  nor2s1 _______505585(.DIN1 (___0_), .DIN2 (________28579), .Q
       (__9_____29959));
  nnd2s1 ____0__505586(.DIN1 (_____0__28562), .DIN2 (_____0__29175), .Q
       (__9_____29731));
  nnd2s1 _______505587(.DIN1 (___9____28660), .DIN2 (________28270), .Q
       (__9_____29851));
  or2s1 ______505588(.DIN1 (_____9__29174), .DIN2 (___9____28686), .Q
       (__9_____29847));
  nnd2s1 _______505589(.DIN1 (_____9__28862), .DIN2 (__9__9__30056), .Q
       (__9__0__29926));
  or2s1 _______505590(.DIN1 (________29173), .DIN2 (________28851), .Q
       (__9_____29857));
  or2s1 _______505591(.DIN1 (____0____31545), .DIN2 (___9____28671), .Q
       (__9_____29835));
  nor2s1 _____0_505592(.DIN1 (______0__31950), .DIN2 (____9___28641),
       .Q (__9__9__29859));
  and2s1 ____0__505593(.DIN1 (________28564), .DIN2 (_________33695),
       .Q (______0__32646));
  and2s1 ____0__505594(.DIN1 (________29172), .DIN2 (________29171), .Q
       (__9__0__29832));
  nnd2s1 _____0_505595(.DIN1 (___9_0__28664), .DIN2 (________28260), .Q
       (____0____32548));
  nnd2s1 ____0_505596(.DIN1 (________28567), .DIN2 (_________33695), .Q
       (_____0___32583));
  nor2s1 ____0__505597(.DIN1 (_____9__27646), .DIN2 (________28540), .Q
       (__909___29718));
  nnd2s1 ____0__505598(.DIN1 (____0___29280), .DIN2 (________26359), .Q
       (_________31944));
  nor2s1 ____0__505599(.DIN1 (___0____27870), .DIN2 (________29241), .Q
       (_________32105));
  nnd2s1 ____0__505600(.DIN1 (____0___29280), .DIN2 (________29170), .Q
       (_________31873));
  hi1s1 ______505601(.DIN (______0__36766), .Q (__9_____29739));
  nor2s1 ____0_505602(.DIN1 (________29169), .DIN2 (________29168), .Q
       (______9__35773));
  nor2s1 _______505603(.DIN1 (_________31673), .DIN2 (___9____28715),
       .Q (__9_9___29893));
  and2s1 _____9_505604(.DIN1 (________28569), .DIN2 (______9__33037),
       .Q (__9_____30259));
  nnd2s1 _______505605(.DIN1 (________28867), .DIN2 (____0____31579),
       .Q (__9__0__30438));
  hi1s1 ______505606(.DIN (_________37223), .Q (__9_____29756));
  nnd2s1 ____0__505607(.DIN1 (____00___31507), .DIN2 (________29395),
       .Q (___0_____31132));
  hi1s1 _______505608(.DIN (_________34136), .Q (_________34225));
  dffacs1 _________________________________________0_____505609(.CLRB
       (reset), .CLK (clk), .DIN (___9_0__28689), .Q
       (_____________________________________0_______21759));
  dffacs1 _______________________________________________505610(.CLRB
       (reset), .CLK (clk), .DIN (________28563), .Q
       (__________________________________________________________________21986));
  nnd2s1 _______505611(.DIN1 (________29166), .DIN2 (___0_0__27009), .Q
       (________29167));
  nnd2s1 ____9__505612(.DIN1 (____9___28463), .DIN2 (____9___28464), .Q
       (_____0__29165));
  xor2s1 ____9__505613(.DIN1 (_____0__28118), .DIN2 (_____00__35736),
       .Q (_____9__29164));
  nnd2s1 _______505614(.DIN1 (________25331), .DIN2 (____9___28465), .Q
       (________29163));
  nor2s1 ____9__505615(.DIN1 (___0_____40585), .DIN2 (________25013),
       .Q (________29162));
  nnd2s1 ____9_505616(.DIN1 (_____0__28433), .DIN2 (____0___25679), .Q
       (________29161));
  nor2s1 ____9__505617(.DIN1 (________27171), .DIN2 (_____0__28404), .Q
       (________29160));
  nnd2s1 ____9_505618(.DIN1 (________28451), .DIN2 (________29158), .Q
       (________29159));
  nnd2s1 ____9__505619(.DIN1 (______________22109), .DIN2
       (___0_____40585), .Q (________29157));
  nor2s1 ____9__505620(.DIN1 (___0_____40585), .DIN2
       (______________22109), .Q (________29156));
  nnd2s1 ____9__505621(.DIN1 (________28409), .DIN2 (_________41196),
       .Q (_____0__29155));
  nor2s1 ____99_505622(.DIN1 (________22870), .DIN2 (________29153), .Q
       (________29154));
  nor2s1 ____0__505623(.DIN1 (_________33897), .DIN2 (________28431),
       .Q (________29152));
  nnd2s1 ____0__505624(.DIN1 (________28185), .DIN2 (________28416), .Q
       (________29151));
  nor2s1 ____0_505625(.DIN1 (________29149), .DIN2 (________28446), .Q
       (________29150));
  nor2s1 ____0__505626(.DIN1 (________28398), .DIN2 (_____0__28443), .Q
       (________29148));
  nor2s1 ____0_505627(.DIN1 (________28426), .DIN2 (________28303), .Q
       (________29147));
  nor2s1 ____0__505628(.DIN1 (________22957), .DIN2 (___0_____40400),
       .Q (_____0__29146));
  nnd2s1 ____0__505629(.DIN1 (_____9__28442), .DIN2 (__9_____30162), .Q
       (_____9__29145));
  nor2s1 ____0__505630(.DIN1 (__90____29663), .DIN2 (________28428), .Q
       (________29144));
  nor2s1 ____0__505631(.DIN1 (________29142), .DIN2 (________28430), .Q
       (________29143));
  nnd2s1 ____0__505632(.DIN1 (________28439), .DIN2 (________29140), .Q
       (________29141));
  nor2s1 ____0__505633(.DIN1 (____0____33491), .DIN2 (________28436),
       .Q (________29139));
  nor2s1 _______505634(.DIN1
       (__________________________________________0___21981), .DIN2
       (___0_____40400), .Q (________29138));
  nnd2s1 _______505635(.DIN1 (________28327), .DIN2 (________28177), .Q
       (________29137));
  and2s1 _______505636(.DIN1 (________28326), .DIN2 (__9__9__30063), .Q
       (_____0__29136));
  or2s1 _______505637(.DIN1 (_____9__28492), .DIN2 (________28868), .Q
       (_____9__29135));
  nor2s1 _____505638(.DIN1 (________28299), .DIN2 (_____9__28989), .Q
       (________29134));
  xnr2s1 _____0_505639(.DIN1
       (_____________________________________________21926), .DIN2
       (______________22106), .Q (________29133));
  xnr2s1 ______505640(.DIN1 (___0_____40433), .DIN2
       (_______________________________________________________________),
       .Q (________29132));
  xor2s1 ______505641(.DIN1
       (______________________________________________21931), .DIN2
       (___0_____40433), .Q (________29131));
  nnd2s1 _______505642(.DIN1 (_________41198), .DIN2 (________28418),
       .Q (________29130));
  xor2s1 _______505643(.DIN1 (________26455), .DIN2 (________27969), .Q
       (________29129));
  nor2s1 _______505644(.DIN1 (____9___23494), .DIN2 (___0_____40400),
       .Q (________29128));
  nor2s1 _______505645(.DIN1 (________27265), .DIN2 (________28449), .Q
       (_____0__29127));
  nnd2s1 ______505646(.DIN1 (____09__29106), .DIN2 (________28417), .Q
       (_____9__29126));
  nnd2s1 _______505647(.DIN1 (________28448), .DIN2 (____0___26593), .Q
       (________29125));
  and2s1 ______505648(.DIN1 (________29153), .DIN2 (________29123), .Q
       (________29124));
  nor2s1 _______505649(.DIN1 (________26795), .DIN2 (___9____28676), .Q
       (________29122));
  nor2s1 _______505650(.DIN1 (________28410), .DIN2 (___0_0__27894), .Q
       (________29121));
  nor2s1 _____9_505651(.DIN1 (________28450), .DIN2 (________29119), .Q
       (________29120));
  or2s1 _____0_505652(.DIN1 (_____0__29117), .DIN2 (____0___29372), .Q
       (________29118));
  nor2s1 _______505653(.DIN1 (________29115), .DIN2 (___9____28675), .Q
       (_____9__29116));
  or2s1 _______505654(.DIN1 (____0____32521), .DIN2 (________28301), .Q
       (________29114));
  nnd2s1 ______505655(.DIN1 (________28393), .DIN2 (________29112), .Q
       (________29113));
  nor2s1 ______505656(.DIN1 (________29110), .DIN2 (________28396), .Q
       (________29111));
  nnd2s1 _______505657(.DIN1 (______0__41130), .DIN2 (________29108),
       .Q (________29109));
  nnd2s1 _______505658(.DIN1 (____09__29106), .DIN2 (_____0__28414), .Q
       (_____0__29107));
  nor2s1 _______505659(.DIN1 (___9____28674), .DIN2 (____0___29104), .Q
       (____0___29105));
  nnd2s1 _______505660(.DIN1 (____0___29285), .DIN2 (____0___29101), .Q
       (____0___29103));
  and2s1 _______505661(.DIN1 (________29361), .DIN2 (____0___29101), .Q
       (____0___29102));
  nor2s1 ______505662(.DIN1 (___0____27846), .DIN2 (_____9__28403), .Q
       (____0___29100));
  nnd2s1 ______505663(.DIN1 (________28241), .DIN2 (_____0__27363), .Q
       (____0___29099));
  and2s1 _______505664(.DIN1 (____0___28208), .DIN2 (____9___28547), .Q
       (____0___29098));
  nnd2s1 _______505665(.DIN1 (________28391), .DIN2 (________27044), .Q
       (____00__29097));
  nor2s1 _______505666(.DIN1 (________28330), .DIN2 (_____9__27686), .Q
       (____99__29096));
  xor2s1 _____505667(.DIN1 (___0_____40596), .DIN2 (________28578), .Q
       (____9___29095));
  nnd2s1 ______505668(.DIN1 (_____0__28351), .DIN2 (___0____28793), .Q
       (____9___29094));
  nnd2s1 ______505669(.DIN1 (_____0__28385), .DIN2 (________29090), .Q
       (_____9__29091));
  nor2s1 _______505670(.DIN1 (________28311), .DIN2 (________28490), .Q
       (________29089));
  nnd2s1 ______505671(.DIN1 (________29086), .DIN2 (___0__0__40421), .Q
       (________29087));
  nnd2s1 ______505672(.DIN1 (________29084), .DIN2
       (______________________________________________21980), .Q
       (________29085));
  nor2s1 _______505673(.DIN1 (___0_99__40460), .DIN2 (____9___28287),
       .Q (_____0__29083));
  nnd2s1 _______505674(.DIN1 (________28347), .DIN2 (____9___26317), .Q
       (_____9__29082));
  nor2s1 _______505675(.DIN1 (________28365), .DIN2 (__999___30539), .Q
       (________29081));
  nnd2s1 _______505676(.DIN1 (________28224), .DIN2 (________29079), .Q
       (________29080));
  nor2s1 ______505677(.DIN1 (________28255), .DIN2 (__9_____30417), .Q
       (________29078));
  nnd2s1 _______505678(.DIN1 (________28974), .DIN2 (____00__26775), .Q
       (________29077));
  or2s1 _______505679(.DIN1 (_____0__28342), .DIN2 (___90___27749), .Q
       (________29076));
  or2s1 _____9_505680(.DIN1 (_____9__29074), .DIN2 (________28335), .Q
       (_____0__29075));
  nor2s1 _____9_505681(.DIN1 (________29072), .DIN2 (_____0__28333), .Q
       (________29073));
  nor2s1 _____505682(.DIN1 (________28271), .DIN2 (________24588), .Q
       (________29071));
  or2s1 _____0_505683(.DIN1 (________28331), .DIN2 (________27172), .Q
       (________29070));
  or2s1 _____0_505684(.DIN1 (________29068), .DIN2 (________28339), .Q
       (________29069));
  nnd2s1 _____505685(.DIN1 (________28249), .DIN2 (________29066), .Q
       (________29067));
  and2s1 ______505686(.DIN1 (________28251), .DIN2 (________27105), .Q
       (_____0__29065));
  nor2s1 _______505687(.DIN1 (________28319), .DIN2 (________27172), .Q
       (_____9__29064));
  nor2s1 _______505688(.DIN1 (___99___28734), .DIN2 (_____0__29046), .Q
       (________29063));
  nnd2s1 _______505689(.DIN1 (________28358), .DIN2 (___0____26981), .Q
       (________29062));
  nnd2s1 ______505690(.DIN1 (___0_____30783), .DIN2 (____0___26779), .Q
       (________29061));
  nnd2s1 ______505691(.DIN1 (____9___28374), .DIN2 (___90___28651), .Q
       (________29060));
  nnd2s1 _______505692(.DIN1 (_____9__28323), .DIN2 (________29537), .Q
       (________29059));
  nor2s1 _______505693(.DIN1 (___00___27831), .DIN2 (________28322), .Q
       (________29058));
  nor2s1 _______505694(.DIN1 (__9_____29783), .DIN2 (________29056), .Q
       (________29057));
  nnd2s1 _______505695(.DIN1 (________28352), .DIN2 (________27322), .Q
       (_____0__29055));
  nor2s1 _______505696(.DIN1 (________29053), .DIN2 (________28321), .Q
       (_____9__29054));
  nor2s1 _______505697(.DIN1 (________27639), .DIN2 (________29051), .Q
       (________29052));
  nor2s1 _______505698(.DIN1 (________29049), .DIN2 (_____0__28361), .Q
       (________29050));
  nnd2s1 ______505699(.DIN1 (___0_0___30748), .DIN2 (_____0__28314), .Q
       (________29048));
  nor2s1 _______505700(.DIN1 (________28497), .DIN2 (_____0__29046), .Q
       (________29047));
  or2s1 _______505701(.DIN1 (________27261), .DIN2 (_____9__28313), .Q
       (_____9__29045));
  nnd2s1 _______505702(.DIN1 (____90__28369), .DIN2 (________29043), .Q
       (________29044));
  nnd2s1 _______505703(.DIN1 (__9_9___30174), .DIN2 (________28312), .Q
       (________29042));
  or2s1 _______505704(.DIN1 (________29269), .DIN2 (________28996), .Q
       (________29041));
  or2s1 _______505705(.DIN1 (_________41136), .DIN2 (________29039), .Q
       (________29040));
  nnd2s1 _______505706(.DIN1 (________28489), .DIN2 (_____0__28247), .Q
       (________29038));
  or2s1 _______505707(.DIN1 (________28026), .DIN2 (____0___28379), .Q
       (_____9__29036));
  nnd2s1 ______505708(.DIN1 (____90__28191), .DIN2 (__9__0__30003), .Q
       (________29035));
  and2s1 _______505709(.DIN1 (____0___28381), .DIN2 (________29033), .Q
       (________29034));
  and2s1 _______505710(.DIN1 (____09__28384), .DIN2 (________29031), .Q
       (________29032));
  nor2s1 _____0_505711(.DIN1 (___9_9__27821), .DIN2 (________28861), .Q
       (________29030));
  nor2s1 ______505712(.DIN1 (________29233), .DIN2 (_____0__29028), .Q
       (________29029));
  nor2s1 _______505713(.DIN1 (________29026), .DIN2 (________28043), .Q
       (_____9__29027));
  nnd2s1 _______505714(.DIN1 (________28234), .DIN2 (___0_0___31119),
       .Q (________29025));
  nnd2s1 _______505715(.DIN1 (________28036), .DIN2 (________29023), .Q
       (________29024));
  and2s1 ______505716(.DIN1 (____00__28200), .DIN2 (_____9__28061), .Q
       (________29022));
  nnd2s1 _______505717(.DIN1 (________28459), .DIN2 (___9_0__27795), .Q
       (________29021));
  nor2s1 _______505718(.DIN1 (________25787), .DIN2 (________28422), .Q
       (________29020));
  or2s1 _______505719(.DIN1 (________27409), .DIN2 (_________41132), .Q
       (________29019));
  nnd2s1 _______505720(.DIN1 (___0_____31035), .DIN2 (________26806),
       .Q (____09__29018));
  nor2s1 _______505721(.DIN1 (________28387), .DIN2 (____0___29200), .Q
       (____0___29017));
  and2s1 ______505722(.DIN1 (________28253), .DIN2 (____0___29015), .Q
       (____0___29016));
  or2s1 _______505723(.DIN1 (____0___29013), .DIN2 (________28345), .Q
       (____0___29014));
  nor2s1 _____9_505724(.DIN1 (___0_____30760), .DIN2 (_____9__28413),
       .Q (____9___29365));
  nnd2s1 _______505725(.DIN1 (_____0__28453), .DIN2 (____0___29012), .Q
       (________29477));
  nor2s1 _______505726(.DIN1 (____0___29011), .DIN2 (________28438), .Q
       (________29494));
  nnd2s1 _____0_505727(.DIN1 (________28406), .DIN2 (_________31778),
       .Q (__90_0__29670));
  nnd2s1 _____505728(.DIN1 (________28458), .DIN2 (____0___29010), .Q
       (____9___29364));
  hi1s1 _______505729(.DIN
       (_________________________________________9___21929), .Q
       (__900___29641));
  nor2s1 _____9_505730(.DIN1 (____00__29009), .DIN2 (________28434), .Q
       (__90____29675));
  nnd2s1 ____9__505731(.DIN1 (____99__29008), .DIN2 (___0_____30709),
       .Q (___0_____31247));
  nnd2s1 _______505732(.DIN1 (________28435), .DIN2 (____9___29007), .Q
       (_________33030));
  nor2s1 ______505733(.DIN1 (____9___29006), .DIN2 (___0_____40400), .Q
       (___0_____40386));
  nor2s1 _______505734(.DIN1 (_____9__27176), .DIN2 (_____9__28394), .Q
       (__90____29701));
  nb1s1 _____9_505735(.DIN (____9___29005), .Q (_____9___34279));
  hi1s1 _____9_505736(.DIN (____9___29005), .Q (______0__33640));
  nor2s1 _______505737(.DIN1 (____00__26408), .DIN2 (________28437), .Q
       (_____9___38611));
  xnr2s1 _______505738(.DIN1
       (_____________________________________________21926), .DIN2
       (___0_90__40451), .Q (____9___29004));
  nnd2s1 _______505739(.DIN1 (____0___28926), .DIN2 (____9___29002), .Q
       (____9___29003));
  nor2s1 _____9_505740(.DIN1 (________28362), .DIN2 (________28048), .Q
       (____9___29001));
  nor2s1 _____0_505741(.DIN1 (____90__28999), .DIN2 (_____9__28998), .Q
       (____9___29000));
  or2s1 _______505742(.DIN1 (__9_____29742), .DIN2 (________28996), .Q
       (________28997));
  nor2s1 _______505743(.DIN1 (________28419), .DIN2 (________28994), .Q
       (________28995));
  nor2s1 _______505744(.DIN1 (__90____29663), .DIN2 (________28397), .Q
       (________28993));
  nor2s1 _______505745(.DIN1 (________28282), .DIN2 (___0____27866), .Q
       (________28992));
  nor2s1 _____9_505746(.DIN1 (____09__28931), .DIN2 (_____9__28989), .Q
       (_____0__28990));
  nnd2s1 _______505747(.DIN1 (_____0__28966), .DIN2 (________28987), .Q
       (________28988));
  nor2s1 ______505748(.DIN1 (__9__9__29935), .DIN2 (_____9__28284), .Q
       (________28986));
  nnd2s1 _______505749(.DIN1 (____9___28371), .DIN2
       (______________________________________________21931), .Q
       (________28985));
  nor2s1 _______505750(.DIN1 (________26710), .DIN2 (_____9__28180), .Q
       (________28984));
  nnd2s1 _______505751(.DIN1 (____0___28294), .DIN2 (___9____26935), .Q
       (________28983));
  nnd2s1 _______505752(.DIN1 (________28184), .DIN2 (________27553), .Q
       (_____0__28981));
  nnd2s1 _______505753(.DIN1 (_____9___32968), .DIN2 (________28188),
       .Q (________28978));
  nor2s1 _______505754(.DIN1 (________27608), .DIN2 (________28366), .Q
       (________28977));
  and2s1 ______505755(.DIN1 (__9_____29735), .DIN2 (__9_____30208), .Q
       (________28976));
  nnd2s1 _______505756(.DIN1 (________28974), .DIN2 (____0___28293), .Q
       (________28975));
  and2s1 _______505757(.DIN1 (_____9__28332), .DIN2 (_____9__28972), .Q
       (_____0__28973));
  nor2s1 ______505758(.DIN1 (____00__27300), .DIN2 (________28265), .Q
       (________28971));
  nnd2s1 _______505759(.DIN1 (________28254), .DIN2 (________28987), .Q
       (________28970));
  nor2s1 _____9_505760(.DIN1 (___0____26985), .DIN2 (________28968), .Q
       (________28969));
  nnd2s1 _____0_505761(.DIN1 (____0___28927), .DIN2 (___0____26994), .Q
       (________28967));
  nnd2s1 _____505762(.DIN1 (__9_____29735), .DIN2 (________27135), .Q
       (_____9__28965));
  nor2s1 _______505763(.DIN1 (___0____26987), .DIN2 (________28968), .Q
       (________28964));
  nnd2s1 ______505764(.DIN1 (_____9__28219), .DIN2 (___0____27840), .Q
       (________28963));
  or2s1 _______505765(.DIN1 (________26741), .DIN2 (________28961), .Q
       (________28962));
  nnd2s1 _______505766(.DIN1 (___0_____30783), .DIN2 (___9____26014),
       .Q (________28960));
  nor2s1 _______505767(.DIN1 (________28227), .DIN2 (________27496), .Q
       (________28959));
  nor2s1 _______505768(.DIN1 (__9_____29783), .DIN2 (________28957), .Q
       (________28958));
  nnd2s1 ______505769(.DIN1 (________27174), .DIN2 (________28955), .Q
       (_____9__28956));
  nnd2s1 _______505770(.DIN1 (_____9__29295), .DIN2 (________28262), .Q
       (________28954));
  and2s1 _______505771(.DIN1 (________28487), .DIN2 (________28952), .Q
       (________28953));
  and2s1 _______505772(.DIN1 (_____0__29495), .DIN2 (________28491), .Q
       (________28951));
  nor2s1 _______505773(.DIN1 (________28248), .DIN2 (__999___30539), .Q
       (________28950));
  nor2s1 _______505774(.DIN1 (________28239), .DIN2 (____90__27559), .Q
       (________28949));
  nor2s1 _______505775(.DIN1 (____90__24546), .DIN2 (_____9__28275), .Q
       (________28948));
  nor2s1 _______505776(.DIN1 (____9___28920), .DIN2 (________29051), .Q
       (_____0__28947));
  nor2s1 _______505777(.DIN1 (___9____26000), .DIN2 (_____0__29046), .Q
       (_____9__28946));
  nnd2s1 ______505778(.DIN1 (____0___29285), .DIN2 (_________41136), .Q
       (________28945));
  nnd2s1 _______505779(.DIN1 (__90____29661), .DIN2 (____9___28197), .Q
       (________28944));
  nor2s1 _______505780(.DIN1 (________28942), .DIN2 (_____0__29046), .Q
       (________28943));
  nor2s1 _______505781(.DIN1 (________27615), .DIN2 (________28226), .Q
       (_____0__28941));
  nor2s1 _______505782(.DIN1 (________28939), .DIN2 (________28165), .Q
       (_____9__28940));
  nor2s1 _______505783(.DIN1 (________28937), .DIN2 (________28325), .Q
       (________28938));
  and2s1 ____505784(.DIN1 (___0_____30783), .DIN2 (________28934), .Q
       (________28935));
  and2s1 ____90_505785(.DIN1 (________28274), .DIN2 (________29158), .Q
       (________28933));
  or2s1 ____90_505786(.DIN1 (____09__28931), .DIN2 (____0___28930), .Q
       (_____0__28932));
  and2s1 ____90_505787(.DIN1 (____09__28209), .DIN2 (__9_____29845), .Q
       (____0___28929));
  nnd2s1 ____9_505788(.DIN1 (____0___28927), .DIN2 (___9____28668), .Q
       (____0___28928));
  nnd2s1 ____9__505789(.DIN1 (_____9__28871), .DIN2 (___9____27820), .Q
       (____0___28925));
  nor2s1 ____9__505790(.DIN1 (___00____30630), .DIN2 (________28217),
       .Q (____00__28924));
  nor2s1 ____9__505791(.DIN1 (____9___28922), .DIN2 (________28968), .Q
       (____99__28923));
  nnd2s1 ____9__505792(.DIN1 (________28244), .DIN2 (____9___28920), .Q
       (____9___28921));
  nnd2s1 ____9_505793(.DIN1 (_____9__29295), .DIN2 (____0___28204), .Q
       (____9___28919));
  and2s1 ____9__505794(.DIN1 (________28359), .DIN2 (____9___28917), .Q
       (____9___28918));
  nor2s1 ____9__505795(.DIN1 (____0___28203), .DIN2 (____9___28915), .Q
       (____9___28916));
  nnd2s1 ____9__505796(.DIN1 (___0_____30783), .DIN2 (___0____27899),
       .Q (_____9__28914));
  and2s1 ____9__505797(.DIN1 (________29086), .DIN2 (____9___22446), .Q
       (________28913));
  and2s1 ____9__505798(.DIN1 (________28911), .DIN2 (___0____27004), .Q
       (________28912));
  or2s1 ____9__505799(.DIN1 (________28909), .DIN2 (________28911), .Q
       (________28910));
  nnd2s1 ____9__505800(.DIN1 (____0___28927), .DIN2 (________27492), .Q
       (________28908));
  nnd2s1 ____9_505801(.DIN1 (_____9__28237), .DIN2 (_____0__28608), .Q
       (________28907));
  or2s1 ____9__505802(.DIN1 (___9_9__28727), .DIN2 (_____9__28989), .Q
       (_____0__28906));
  nnd2s1 ____9_505803(.DIN1 (________28898), .DIN2 (____0___29285), .Q
       (_____9__28905));
  and2s1 ____9__505804(.DIN1 (________28356), .DIN2 (___009___30634),
       .Q (________28904));
  nnd2s1 ____9__505805(.DIN1 (________28215), .DIN2 (_____0__27411), .Q
       (________28903));
  nor2s1 ____9__505806(.DIN1 (________26345), .DIN2 (________29051), .Q
       (________28902));
  nnd2s1 ____99_505807(.DIN1 (________28240), .DIN2 (________28900), .Q
       (________28901));
  nor2s1 ____99_505808(.DIN1 (________27973), .DIN2 (________28898), .Q
       (________28899));
  xor2s1 ____00_505809(.DIN1 (________27612), .DIN2 (___0_____40534),
       .Q (_____0__28897));
  xor2s1 ____0_505810(.DIN1 (________27618), .DIN2 (______0__36697), .Q
       (_____9__28896));
  xor2s1 ____0__505811(.DIN1
       (_____________________________________________21787), .DIN2
       (________27618), .Q (________28894));
  and2s1 ____0__505812(.DIN1 (________28892), .DIN2 (________28891), .Q
       (________28893));
  and2s1 ______505813(.DIN1 (_____0__28174), .DIN2 (________28887), .Q
       (________28888));
  nnd2s1 _______505814(.DIN1 (________28279), .DIN2 (________28182), .Q
       (________28886));
  nnd2s1 _____9_505815(.DIN1 (________28172), .DIN2 (________29140), .Q
       (________28885));
  nnd2s1 _______505816(.DIN1 (_____9__28173), .DIN2 (__99__), .Q
       (________28884));
  xor2s1 ____0__505817(.DIN1 (________27618), .DIN2 (___99_0__39864),
       .Q (________28883));
  xor2s1 ____0__505818(.DIN1 (___0__9__40480), .DIN2 (________27618),
       .Q (________28882));
  nor2s1 _______505819(.DIN1 (________28183), .DIN2 (___9_9__27804), .Q
       (_____0__28881));
  nor2s1 _____505820(.DIN1 (________28879), .DIN2 (________28878), .Q
       (_____9__28880));
  nnd2s1 _____505821(.DIN1 (________29023), .DIN2 (________28876), .Q
       (__90____29651));
  nor2s1 ______505822(.DIN1 (________28875), .DIN2 (________28389), .Q
       (__90_9));
  nor2s1 _______505823(.DIN1 (___00____30587), .DIN2 (______0__41140),
       .Q (________29177));
  or2s1 _______505824(.DIN1 (________28874), .DIN2 (_____9__28989), .Q
       (________29505));
  or2s1 _____0_505825(.DIN1 (________27662), .DIN2 (______0__41140), .Q
       (________29499));
  nnd2s1 _______505826(.DIN1 (________28873), .DIN2 (_____0__28872), .Q
       (___900___38982));
  nor2s1 _______505827(.DIN1 (___00___26954), .DIN2 (________28961), .Q
       (____99__29278));
  nnd2s1 ____0__505828(.DIN1 (_____9__28871), .DIN2 (___0_0___30746),
       .Q (__9_____29834));
  nnd2s1 ____0__505829(.DIN1 (________28221), .DIN2 (________28870), .Q
       (___90___29559));
  nnd2s1 ____0__505830(.DIN1 (_____9__28546), .DIN2 (________26615), .Q
       (________29515));
  nnd2s1 ____0__505831(.DIN1 (________28218), .DIN2 (_________31781),
       .Q (________29216));
  nnd2s1 ______505832(.DIN1 (_________34531), .DIN2 (________28278), .Q
       (_________32688));
  nnd2s1 _______505833(.DIN1 (________28869), .DIN2 (___0____26977), .Q
       (________29293));
  nor2s1 _______505834(.DIN1 (___9____26945), .DIN2 (________28968), .Q
       (_____9___31690));
  nor2s1 ____0__505835(.DIN1 (________26830), .DIN2 (________28868), .Q
       (____9___29548));
  hi1s1 _______505836(.DIN (________28867), .Q (__9_____30303));
  nor2s1 ____0__505837(.DIN1 (________28866), .DIN2 (________28280), .Q
       (__9_9___29990));
  nor2s1 ____0__505838(.DIN1 (_________41291), .DIN2 (____0___28205),
       .Q (________29513));
  nor2s1 _______505839(.DIN1 (________28003), .DIN2 (_____9__28488), .Q
       (___9_9__29627));
  or2s1 ______505840(.DIN1 (___09____31429), .DIN2 (________28346), .Q
       (___999__29637));
  nor2s1 _______505841(.DIN1 (________28865), .DIN2 (________28864), .Q
       (_________38376));
  nor2s1 _______505842(.DIN1 (_________32658), .DIN2 (________28367),
       .Q (____9___29277));
  or2s1 ____0__505843(.DIN1 (___0_____31274), .DIN2 (_____9__28266), .Q
       (_________32982));
  nnd2s1 ____0_505844(.DIN1 (__9_____29735), .DIN2 (________25646), .Q
       (_____0___32577));
  nnd2s1 ____0_505845(.DIN1 (___0_____30783), .DIN2 (________26799), .Q
       (____0____32534));
  nor2s1 ____0__505846(.DIN1 (________28269), .DIN2 (__999___30539), .Q
       (_____00__33249));
  nor2s1 _______505847(.DIN1 (_____0__28863), .DIN2 (________28178), .Q
       (___0_____30870));
  hi1s1 _______505848(.DIN (_____9__28862), .Q (___9____29622));
  or2s1 ____0__505849(.DIN1 (____9___29190), .DIN2 (________28861), .Q
       (_____0___32676));
  or2s1 ____0__505850(.DIN1 (___0_9___40354), .DIN2 (________29084), .Q
       (___0_9___40358));
  dffacs1 _________________505851(.CLRB (reset), .CLK (clk), .DIN
       (________28340), .QN (______________22065));
  nor2s1 ____0__505852(.DIN1 (________28860), .DIN2 (_____0__28257), .Q
       (______0__36766));
  nor2s1 ____0__505853(.DIN1 (____0___23695), .DIN2 (________28355), .Q
       (_________37223));
  nnd2s1 ____0__505854(.DIN1 (________28258), .DIN2 (________26604), .Q
       (_________34136));
  or2s1 _______505855(.DIN1 (________28859), .DIN2 (________28353), .Q
       (_________37317));
  nor2s1 ______505856(.DIN1 (________28850), .DIN2 (____90__28101), .Q
       (________28858));
  nnd2s1 ____0__505857(.DIN1 (________28132), .DIN2 (____0___27035), .Q
       (________28856));
  nor2s1 ____0__505858(.DIN1 (________28135), .DIN2 (__9__0__30291), .Q
       (________28855));
  nnd2s1 _______505859(.DIN1 (________28852), .DIN2 (________27541), .Q
       (_____0__28854));
  nnd2s1 _______505860(.DIN1 (________28852), .DIN2 (____0___27926), .Q
       (_____9__28853));
  or2s1 _______505861(.DIN1 (________28850), .DIN2 (_____9__28127), .Q
       (________28851));
  hi1s1 _______505862(.DIN (________28848), .Q (________28849));
  hi1s1 _____505863(.DIN (____99__29008), .Q (________28847));
  and2s1 _______505864(.DIN1 (________28845), .DIN2 (___0_____30709),
       .Q (________28846));
  nor2s1 _______505865(.DIN1 (____9___28196), .DIN2 (____09__28843), .Q
       (_____0__28844));
  or2s1 _______505866(.DIN1 (________28866), .DIN2 (________28126), .Q
       (____0___28842));
  nnd2s1 _______505867(.DIN1 (__90____29661), .DIN2 (________28124), .Q
       (____0___28841));
  nnd2s1 _______505868(.DIN1 (________28420), .DIN2 (____0___28839), .Q
       (____0___28840));
  or2s1 ______505869(.DIN1 (___0____26979), .DIN2 (___0____28783), .Q
       (____0___28838));
  hi1s1 ______505870(.DIN (___0_____40400), .Q (____0___28837));
  nor2s1 _______505871(.DIN1 (___0_0__27018), .DIN2 (___9____28705), .Q
       (____0___28836));
  nnd2s1 _______505872(.DIN1 (____9___28469), .DIN2
       (_____________________________________________21973), .Q
       (____0___28835));
  nor2s1 _______505873(.DIN1
       (_____________________________________________21941), .DIN2
       (___0_____40115), .Q (____00__28834));
  nnd2s1 _______505874(.DIN1 (__9_____30019), .DIN2 (________27976), .Q
       (___099__28833));
  nnd2s1 ______505875(.DIN1 (____9___28551), .DIN2 (_____9__27940), .Q
       (___09___28832));
  nnd2s1 ______505876(.DIN1 (_____0__28042), .DIN2 (____990__33424), .Q
       (___09___28831));
  nor2s1 _______505877(.DIN1 (___09____31438), .DIN2 (___09___28829),
       .Q (___09___28830));
  nor2s1 _______505878(.DIN1 (____09__27215), .DIN2 (_____9__28004), .Q
       (___09___28828));
  nnd2s1 _______505879(.DIN1 (____0___28015), .DIN2 (clk), .Q
       (___09___28827));
  nnd2s1 _______505880(.DIN1 (________28099), .DIN2 (___09___28825), .Q
       (___09___28826));
  nnd2s1 _______505881(.DIN1 (________28095), .DIN2 (________27353), .Q
       (___0_9__28824));
  nnd2s1 _______505882(.DIN1 (________28093), .DIN2 (___0____28822), .Q
       (___0____28823));
  nor2s1 _______505883(.DIN1 (_____0__28082), .DIN2 (___0____28820), .Q
       (___0____28821));
  nnd2s1 _______505884(.DIN1 (________28092), .DIN2 (____990__33424),
       .Q (___0____28819));
  and2s1 ______505885(.DIN1 (___0____28817), .DIN2 (___9____28657), .Q
       (___0____28818));
  nnd2s1 _______505886(.DIN1 (___0____28790), .DIN2 (____0___27036), .Q
       (___0____28816));
  nnd2s1 _______505887(.DIN1 (________28085), .DIN2 (___0_9__28814), .Q
       (___0_0__28815));
  nor2s1 _______505888(.DIN1 (________28485), .DIN2 (________27947), .Q
       (___0____28813));
  and2s1 _______505889(.DIN1 (________28064), .DIN2 (___0____28811), .Q
       (___0____28812));
  nnd2s1 _______505890(.DIN1 (___0_9__27883), .DIN2 (_____0__27177), .Q
       (___0____28810));
  nnd2s1 _____505891(.DIN1 (________28079), .DIN2 (_________38856), .Q
       (___0____28809));
  nor2s1 _____9_505892(.DIN1 (_________32305), .DIN2 (________28075),
       .Q (___0____28808));
  or2s1 _____9_505893(.DIN1 (___0____28806), .DIN2 (________28073), .Q
       (___0____28807));
  nor2s1 _____9_505894(.DIN1 (_____9__28091), .DIN2 (___0_9__28804), .Q
       (___0_0__28805));
  and2s1 _____9_505895(.DIN1 (________28068), .DIN2 (_____0__27372), .Q
       (___0____28803));
  nnd2s1 _____9_505896(.DIN1 (________27990), .DIN2 (____9___28198), .Q
       (___0____28802));
  nnd2s1 _____9_505897(.DIN1 (__9_____29957), .DIN2 (_________41142),
       .Q (___0____28801));
  and2s1 _____0_505898(.DIN1 (________27959), .DIN2 (________26439), .Q
       (___0____28800));
  nor2s1 _____0_505899(.DIN1 (__9_____30335), .DIN2 (________28058), .Q
       (___0____28799));
  nor2s1 _____0_505900(.DIN1 (___0____28797), .DIN2 (________27172), .Q
       (___0____28798));
  nnd2s1 _____0_505901(.DIN1 (___0_____40115), .DIN2 (___9____26875),
       .Q (___0_0__28796));
  or2s1 _______505902(.DIN1 (_____9__28071), .DIN2 (___0____27908), .Q
       (___0_9__28795));
  nnd2s1 _______505903(.DIN1 (___9____28716), .DIN2 (___0____28793), .Q
       (___0____28794));
  nnd2s1 _______505904(.DIN1 (_____0__28052), .DIN2 (____990__33424),
       .Q (___0____28792));
  nor2s1 ______505905(.DIN1 (___0____28790), .DIN2 (________27172), .Q
       (___0____28791));
  and2s1 _______505906(.DIN1 (________28050), .DIN2 (___0____28788), .Q
       (___0____28789));
  nnd2s1 _______505907(.DIN1 (________28613), .DIN2 (_____9__26185), .Q
       (___0____28787));
  nnd2s1 _______505908(.DIN1 (___99___28732), .DIN2 (___90___25962), .Q
       (___0_0__28786));
  or2s1 _______505909(.DIN1 (___0____28784), .DIN2 (___0____28783), .Q
       (___0_9__28785));
  nnd2s1 _______505910(.DIN1 (__90_9__29717), .DIN2 (________26381), .Q
       (___0____28782));
  nnd2s1 _______505911(.DIN1 (________28055), .DIN2 (inData[10]), .Q
       (___0____28781));
  nor2s1 _______505912(.DIN1 (___0____28779), .DIN2 (________28037), .Q
       (___0____28780));
  or2s1 _______505913(.DIN1 (________28909), .DIN2 (________28035), .Q
       (___0____28778));
  nor2s1 ______505914(.DIN1 (________27081), .DIN2 (___0____28783), .Q
       (___0____28777));
  and2s1 _______505915(.DIN1 (_____9___33997), .DIN2 (_____9__29295),
       .Q (___0_0__28776));
  nor2s1 _______505916(.DIN1 (________26302), .DIN2 (_____9__28031), .Q
       (___0_9__28775));
  or2s1 _______505917(.DIN1 (______9__34266), .DIN2 (________27966), .Q
       (___0____28774));
  nnd2s1 ______505918(.DIN1 (________28086), .DIN2 (inData[16]), .Q
       (___0____28773));
  nor2s1 _______505919(.DIN1 (____9___27735), .DIN2 (____0___28558), .Q
       (___0____28772));
  nnd2s1 _______505920(.DIN1 (__90_9__29717), .DIN2 (_____0__28032), .Q
       (___0____28771));
  or2s1 _______505921(.DIN1 (________28589), .DIN2 (________28025), .Q
       (___0____28770));
  nor2s1 _______505922(.DIN1 (_____0__29037), .DIN2 (________28045), .Q
       (___0____28769));
  and2s1 _______505923(.DIN1 (____00__28108), .DIN2 (____99__25957), .Q
       (___0____28768));
  or2s1 ______505924(.DIN1 (__9__0__30093), .DIN2 (________28033), .Q
       (___0____28767));
  nor2s1 _____505925(.DIN1 (____0___28112), .DIN2 (___0_9__28765), .Q
       (___0_0__28766));
  nor2s1 _____9_505926(.DIN1 (________27961), .DIN2 (___0____28763), .Q
       (___0____28764));
  nnd2s1 _____9_505927(.DIN1 (___0____28761), .DIN2 (___90___27743), .Q
       (___0____28762));
  nnd2s1 _____9_505928(.DIN1 (____0___28018), .DIN2 (inData[24]), .Q
       (___0____28760));
  or2s1 _____505929(.DIN1 (___0____28758), .DIN2 (___0____28757), .Q
       (___0____28759));
  nnd2s1 _____0_505930(.DIN1 (____00__28376), .DIN2 (________27500), .Q
       (___0_0__28756));
  or2s1 _____0_505931(.DIN1 (___0____28754), .DIN2 (________28625), .Q
       (___0_9__28755));
  nor2s1 _____0_505932(.DIN1 (____00__28014), .DIN2 (__9_____30401), .Q
       (___0____28753));
  nor2s1 _____0_505933(.DIN1 (___0____28763), .DIN2 (________28166), .Q
       (___0____28752));
  or2s1 _____0_505934(.DIN1 (_________33551), .DIN2 (____9___28012), .Q
       (___0____28751));
  nor2s1 _____0_505935(.DIN1 (____9___28373), .DIN2 (________27970), .Q
       (___0____28750));
  nnd2s1 _______505936(.DIN1 (________28027), .DIN2 (___0____28748), .Q
       (___0____28749));
  nor2s1 _______505937(.DIN1 (________29500), .DIN2 (___9____28712), .Q
       (___0____28747));
  and2s1 _______505938(.DIN1 (________27952), .DIN2 (__9_____30096), .Q
       (___0_0__28746));
  nor2s1 _______505939(.DIN1 (___00___28744), .DIN2 (___990__28728), .Q
       (___009__28745));
  nor2s1 _______505940(.DIN1 (_____9__27426), .DIN2 (___00___28737), .Q
       (___00___28743));
  or2s1 _______505941(.DIN1 (___00___28741), .DIN2 (__9_0___30373), .Q
       (___00___28742));
  nnd2s1 _______505942(.DIN1 (________28141), .DIN2 (___0_09__30841),
       .Q (___00___28740));
  nnd2s1 _______505943(.DIN1 (________28080), .DIN2 (________27975), .Q
       (___00___28739));
  or2s1 _______505944(.DIN1 (________28000), .DIN2 (___00___28737), .Q
       (___00___28738));
  nor2s1 _______505945(.DIN1 (____9___28006), .DIN2 (________28233), .Q
       (___000__28736));
  or2s1 _______505946(.DIN1 (___99___28734), .DIN2 (___0____28783), .Q
       (___999__28735));
  and2s1 _______505947(.DIN1 (___99___28732), .DIN2 (___99___28731), .Q
       (___99___28733));
  nor2s1 _______505948(.DIN1 (___990__28728), .DIN2 (___9_9__28727), .Q
       (___99___28729));
  nnd2s1 _______505949(.DIN1 (____9___28102), .DIN2 (________29361), .Q
       (___9____28726));
  nnd2s1 ______505950(.DIN1 (___9____28670), .DIN2 (________27285), .Q
       (___9____28725));
  and2s1 _______505951(.DIN1 (__90_9__29717), .DIN2 (___9____28702), .Q
       (___9____28724));
  nnd2s1 _______505952(.DIN1 (____9___28288), .DIN2 (___9____28722), .Q
       (___9____28723));
  nor2s1 _______505953(.DIN1 (________28024), .DIN2 (____0___29200), .Q
       (___9____28721));
  nnd2s1 _______505954(.DIN1 (___9____28719), .DIN2 (___999__26050), .Q
       (___9____28720));
  or2s1 _______505955(.DIN1 (____9___28010), .DIN2 (_____9___33997), .Q
       (___9_0__28718));
  and2s1 _______505956(.DIN1 (___9____28716), .DIN2 (________28305), .Q
       (___9_9__28717));
  or2s1 _______505957(.DIN1 (__9_____30198), .DIN2 (_____0__28023), .Q
       (___9____28715));
  and2s1 _______505958(.DIN1 (___0____27879), .DIN2 (___00____30556),
       .Q (___9____28714));
  nor2s1 _______505959(.DIN1 (______0__31970), .DIN2 (___9____28712),
       .Q (___9____28713));
  nor2s1 _______505960(.DIN1 (________28076), .DIN2 (________29415), .Q
       (___9____28711));
  nnd2s1 _______505961(.DIN1 (___9____28709), .DIN2 (____9___28470), .Q
       (___9____28710));
  and2s1 _______505962(.DIN1 (________28078), .DIN2 (________28612), .Q
       (___9_0__28708));
  and2s1 _______505963(.DIN1 (___0_____30961), .DIN2 (________27418),
       .Q (___9_9__28707));
  nor2s1 ______505964(.DIN1 (________28090), .DIN2 (___9____28705), .Q
       (___9____28706));
  nor2s1 _____505965(.DIN1 (___9____28703), .DIN2 (___9____28702), .Q
       (___9____28704));
  nnd2s1 _____9_505966(.DIN1 (____9___28375), .DIN2 (________27439), .Q
       (___9____28701));
  nnd2s1 _____9_505967(.DIN1 (____9___28372), .DIN2 (_____9__27619), .Q
       (___9____28700));
  nor2s1 _____9_505968(.DIN1 (___9_0__28698), .DIN2 (________27979), .Q
       (___9____28699));
  and2s1 _____505969(.DIN1 (____9___28105), .DIN2 (___9____28696), .Q
       (___9____28697));
  nor2s1 ______505970(.DIN1 (___00____30605), .DIN2 (________27936), .Q
       (___9____28695));
  nnd2s1 _______505971(.DIN1 (___9____28692), .DIN2 (___0____27871), .Q
       (___9____28694));
  nnd2s1 _______505972(.DIN1 (___9____28692), .DIN2 (___0_0__26967), .Q
       (___9____28693));
  nnd2s1 _______505973(.DIN1 (____9___28011), .DIN2 (____09__26598), .Q
       (___9____28691));
  and2s1 _______505974(.DIN1 (__9_____30349), .DIN2 (________28300), .Q
       (___9____28690));
  nnd2s1 ______505975(.DIN1 (____0___27929), .DIN2 (_____9__27046), .Q
       (___9_0__28689));
  nnd2s1 ______505976(.DIN1 (__9_9___30270), .DIN2 (____0___27927), .Q
       (___9_9__28688));
  or2s1 _______505977(.DIN1 (_________41285), .DIN2 (_____0__27968), .Q
       (___9____28687));
  nnd2s1 _______505978(.DIN1 (____0___28110), .DIN2 (_____0__28181), .Q
       (___9____28686));
  nnd2s1 _______505979(.DIN1 (___9____28692), .DIN2 (________26668), .Q
       (___9____28685));
  nnd2s1 ______505980(.DIN1 (____09__29106), .DIN2 (________27944), .Q
       (___9____28684));
  nnd2s1 _______505981(.DIN1
       (_____________________________________________21926), .DIN2
       (______________22106), .Q (___9____28683));
  nnd2s1 _____0_505982(.DIN1 (________27988), .DIN2 (inData[6]), .Q
       (___9____28682));
  or2s1 _____0_505983(.DIN1 (_________32750), .DIN2 (________27963), .Q
       (___9_0__28681));
  or2s1 _____0_505984(.DIN1 (___9____28679), .DIN2 (____9___28009), .Q
       (___9_9__28680));
  nnd2s1 _____0_505985(.DIN1 (________28028), .DIN2 (inData[14]), .Q
       (___9____28678));
  hi1s1 _______505986(.DIN (___9____28676), .Q (___9____28677));
  nnd2s1 _______505987(.DIN1 (________27938), .DIN2 (____990__33424),
       .Q (___9_0__28673));
  xor2s1 _______505988(.DIN1
       (_____________________________________________21899), .DIN2
       (___0_____40439), .Q (___9_9__28672));
  nnd2s1 ______505989(.DIN1 (___9____28670), .DIN2 (_________31678), .Q
       (___9____28671));
  nor2s1 _______505990(.DIN1 (_____9__28636), .DIN2 (___9____28668), .Q
       (___9____28669));
  nnd2s1 _______505991(.DIN1 (__90_9__29717), .DIN2 (________26646), .Q
       (___9____28666));
  nnd2s1 _______505992(.DIN1 (___9____28692), .DIN2 (________27202), .Q
       (___9____28665));
  nnd2s1 _______505993(.DIN1 (________27993), .DIN2 (_________32836),
       .Q (___9_0__28664));
  nnd2s1 _______505994(.DIN1 (___9____28662), .DIN2 (inData[12]), .Q
       (___9_9__28663));
  nnd2s1 _______505995(.DIN1 (________28049), .DIN2 (inData[8]), .Q
       (___9____28661));
  nnd2s1 ______505996(.DIN1 (________27444), .DIN2 (____0___27928), .Q
       (___9____28660));
  nor2s1 _____9_505997(.DIN1 (___0____26113), .DIN2 (___0____27886), .Q
       (___9____28659));
  and2s1 _____9_505998(.DIN1 (_____0__28072), .DIN2 (___9____28657), .Q
       (___9____28658));
  nnd2s1 _____505999(.DIN1 (_____9__27957), .DIN2 (_____9__26747), .Q
       (___9____28656));
  nnd2s1 _____0_506000(.DIN1 (____0___29285), .DIN2 (________27953), .Q
       (___909__28654));
  xor2s1 _______506001(.DIN1 (________27445), .DIN2 (_________33321),
       .Q (____9___29005));
  nnd2s1 _______506002(.DIN1 (____0___27930), .DIN2 (___90___28653), .Q
       (________29450));
  nor2s1 _______506003(.DIN1 (___90___28652), .DIN2 (________28065), .Q
       (________29447));
  nnd2s1 _______506004(.DIN1 (________28098), .DIN2 (________29031), .Q
       (________29321));
  nnd2s1 _______506005(.DIN1 (________27942), .DIN2 (____9___29463), .Q
       (____0___29467));
  nnd2s1 _______506006(.DIN1 (____0___28021), .DIN2 (___90___28651), .Q
       (________29349));
  nor2s1 _______506007(.DIN1 (___99___25116), .DIN2 (________28067), .Q
       (________29420));
  or2s1 ______506008(.DIN1 (___09_9__31446), .DIN2 (________27933), .Q
       (__90____29653));
  nor2s1 _____0_506009(.DIN1 (___00___27830), .DIN2 (________27948), .Q
       (_________32347));
  nnd2s1 _____0_506010(.DIN1 (________28054), .DIN2 (___90___28650), .Q
       (____9___29092));
  and2s1 _____0_506011(.DIN1 (________28088), .DIN2 (_________31973),
       .Q (____09__29377));
  or2s1 _____0_506012(.DIN1 (____9___27738), .DIN2 (___0____27852), .Q
       (___0_____31010));
  and2s1 ______506013(.DIN1 (________28059), .DIN2 (___90___28649), .Q
       (________29452));
  or2s1 ______506014(.DIN1 (_____9___31789), .DIN2 (________28134), .Q
       (________29490));
  nor2s1 _______506015(.DIN1 (________25559), .DIN2 (___0_0__27884), .Q
       (____0____35363));
  dffacs1 _____________________________________________9_506016(.CLRB
       (reset), .CLK (clk), .DIN (________28056), .Q
       (_________________________________________9___21929));
  nnd2s1 ______506017(.DIN1 (___0_____40115), .DIN2 (___90___28648), .Q
       (___9_____39494));
  dffacs1 ________________________________________________506018(.CLRB
       (reset), .CLK (clk), .DIN (________28069), .Q
       (______________________________________________21904));
  and2s1 ____9__506019(.DIN1 (_____0___36015), .DIN2 (_________32663),
       .Q (______9__32949));
  nnd2s1 _______506020(.DIN1 (__9_____30423), .DIN2 (___0____27900), .Q
       (___90___28647));
  nor2s1 _______506021(.DIN1 (_____9__27977), .DIN2 (__90____29663), .Q
       (___900__28646));
  or2s1 ______506022(.DIN1 (____9___28644), .DIN2 (___0_0__27855), .Q
       (____99__28645));
  nor2s1 _______506023(.DIN1 (________27313), .DIN2 (___0____28783), .Q
       (____9___28643));
  or2s1 _______506024(.DIN1 (___0_90__31108), .DIN2 (___0____27904), .Q
       (____9___28641));
  nor2s1 ______506025(.DIN1 (________28038), .DIN2 (________29119), .Q
       (____9___28640));
  nor2s1 _______506026(.DIN1 (________22486), .DIN2 (___9____28662), .Q
       (____9___28639));
  nnd2s1 _______506027(.DIN1 (___9____28692), .DIN2 (________26343), .Q
       (____9___28638));
  nnd2s1 _______506028(.DIN1 (___9____28692), .DIN2 (_____9__28636), .Q
       (____90__28637));
  nor2s1 ______506029(.DIN1 (________28634), .DIN2 (____0___29104), .Q
       (________28635));
  nnd2s1 _______506030(.DIN1 (__9990), .DIN2 (___0____27898), .Q
       (________28633));
  and2s1 _______506031(.DIN1 (________28631), .DIN2 (____90__27472), .Q
       (________28632));
  nor2s1 ______506032(.DIN1 (________27997), .DIN2 (___0_9__28804), .Q
       (________28630));
  nnd2s1 _____9_506033(.DIN1 (____0___28113), .DIN2 (________28628), .Q
       (________28629));
  or2s1 _____9_506034(.DIN1 (_____9__28626), .DIN2 (___0____28783), .Q
       (_____0__28627));
  nor2s1 _____9_506035(.DIN1 (_________31667), .DIN2 (________28047),
       .Q (________28624));
  nor2s1 _____9_506036(.DIN1 (________27995), .DIN2 (________27149), .Q
       (________28623));
  nnd2s1 ____90_506037(.DIN1 (________29361), .DIN2 (________28121), .Q
       (________28622));
  or2s1 ____90_506038(.DIN1 (________27721), .DIN2 (________28857), .Q
       (________28621));
  nnd2s1 ____9__506039(.DIN1 (___0_9__27893), .DIN2 (________27256), .Q
       (________28620));
  or2s1 ____9__506040(.DIN1 (__9_0___29726), .DIN2 (________28002), .Q
       (________28619));
  nnd2s1 ____9__506041(.DIN1 (_____9__28617), .DIN2
       (__________________________________________________________________21990),
       .Q (_____0__28618));
  nnd2s1 ____9__506042(.DIN1 (________23845), .DIN2 (________27981), .Q
       (________28616));
  nor2s1 ____9__506043(.DIN1 (_________34167), .DIN2 (___9____28662),
       .Q (________28615));
  nnd2s1 ____9__506044(.DIN1 (________28613), .DIN2 (________28612), .Q
       (________28614));
  nor2s1 ____9_506045(.DIN1 (________28534), .DIN2 (________28610), .Q
       (________28611));
  nnd2s1 ____9__506046(.DIN1 (_____0__28608), .DIN2 (____0___28297), .Q
       (________28609));
  nor2s1 ____9__506047(.DIN1 (________27984), .DIN2 (_____0__27941), .Q
       (_____9__28607));
  and2s1 ____9__506048(.DIN1 (_____0__27950), .DIN2 (________28605), .Q
       (________28606));
  and2s1 ____9__506049(.DIN1 (_____9__28041), .DIN2 (____9___29463), .Q
       (________28604));
  and2s1 ____9_506050(.DIN1 (________28602), .DIN2 (___0____27842), .Q
       (________28603));
  or2s1 ____9__506051(.DIN1 (________28600), .DIN2 (___0____27895), .Q
       (________28601));
  nor2s1 ____9__506052(.DIN1 (________28164), .DIN2 (_________41168),
       .Q (________28599));
  nnd2s1 ____9__506053(.DIN1 (___0_____31078), .DIN2 (________28597),
       .Q (_____9__28598));
  nnd2s1 ____9_506054(.DIN1 (___0_0__27875), .DIN2 (________24879), .Q
       (________28595));
  nor2s1 ____9__506055(.DIN1 (_____0__28210), .DIN2 (___0____28783), .Q
       (________28594));
  nnd2s1 ____9_506056(.DIN1 (________28592), .DIN2 (_____0__28591), .Q
       (________28593));
  or2s1 ____9__506057(.DIN1 (________28589), .DIN2 (___0____27907), .Q
       (_____9__28590));
  or2s1 ____9_506058(.DIN1 (___9_9__27813), .DIN2 (________28587), .Q
       (________28588));
  nnd2s1 ____9__506059(.DIN1 (____09__27931), .DIN2 (________28585), .Q
       (________28586));
  nor2s1 ____9__506060(.DIN1 (________28583), .DIN2 (___0____28783), .Q
       (________28584));
  nnd2s1 ____9__506061(.DIN1 (___0____27891), .DIN2 (___0____27901), .Q
       (________28582));
  nnd2s1 ____9_506062(.DIN1 (__9_9___30174), .DIN2 (____0___28115), .Q
       (_____0__28581));
  nnd2s1 ____9__506063(.DIN1 (___9____28692), .DIN2 (___9_0__26901), .Q
       (_____9__28580));
  nor2s1 ____9__506064(.DIN1 (_______22180), .DIN2 (________28578), .Q
       (________28579));
  or2s1 ____9__506065(.DIN1 (_________41172), .DIN2 (___0____28783), .Q
       (________28577));
  nor2s1 ____99_506066(.DIN1 (__9_0___29995), .DIN2 (____00__28291), .Q
       (________28576));
  and2s1 ____99_506067(.DIN1 (________28123), .DIN2 (__9_____30332), .Q
       (________28575));
  and2s1 ____99_506068(.DIN1 (___9____28692), .DIN2 (________28573), .Q
       (________28574));
  nnd2s1 ____506069(.DIN1 (________27994), .DIN2 (________27946), .Q
       (________28572));
  nor2s1 ____90_506070(.DIN1 (________28077), .DIN2 (_____9__28570), .Q
       (_____0__28571));
  hi1s1 _______506071(.DIN (_________33175), .Q (________28569));
  or2s1 _______506072(.DIN1 (__9_____30098), .DIN2 (___0_9__27874), .Q
       (________28568));
  nnd2s1 _______506073(.DIN1 (_________32266), .DIN2 (_____9__26314),
       .Q (________28567));
  nnd2s1 _______506074(.DIN1 (________27539), .DIN2 (___0____27867), .Q
       (________28566));
  xor2s1 ____0__506075(.DIN1 (___0_____40527), .DIN2 (___9_0___39077),
       .Q (________28565));
  nnd2s1 _______506076(.DIN1 (_________32266), .DIN2 (________26334),
       .Q (________28564));
  nnd2s1 ______506077(.DIN1 (___0_0__27865), .DIN2 (___9_____39548), .Q
       (________28563));
  nor2s1 ______506078(.DIN1 (_____9__29174), .DIN2 (___0____27859), .Q
       (_____0__28562));
  xor2s1 ____0_506079(.DIN1 (____09__23890), .DIN2
       (__________________________________9__________), .Q
       (____09__28561));
  nor2s1 _______506080(.DIN1 (__9__9__29935), .DIN2 (___0_9__27854), .Q
       (____0___28560));
  nnd2s1 _______506081(.DIN1 (____0___28558), .DIN2 (__9_____30423), .Q
       (____0___28559));
  nnd2s1 _____506082(.DIN1 (________29525), .DIN2 (_____0__27490), .Q
       (____0___28557));
  xor2s1 ____0_506083(.DIN1
       (_____________________________________________21875), .DIN2
       (__________________________________9__________), .Q
       (____0___28556));
  xor2s1 ____0__506084(.DIN1 (_________37864), .DIN2 (_____0___32287),
       .Q (____0___28555));
  nor2s1 _______506085(.DIN1 (___9____27775), .DIN2 (_________41152),
       .Q (____0___28554));
  nnd2s1 _______506086(.DIN1
       (_________________________________________________________________________________________22089),
       .DIN2 (_________41367), .Q (____9___28553));
  nnd2s1 _______506087(.DIN1 (____9___28551), .DIN2 (____9___28550), .Q
       (____9___28552));
  hi1s1 ____0__506088(.DIN (____9___28548), .Q (____9___28549));
  hi1s1 ____0__506089(.DIN (___0_____40320), .Q (________28545));
  and2s1 _______506090(.DIN1 (___0_0__27845), .DIN2 (________28543), .Q
       (________28544));
  nor2s1 _____506091(.DIN1 (________28541), .DIN2 (________28175), .Q
       (________28542));
  hi1s1 ____09_506092(.DIN (___0_____30783), .Q (________28540));
  and2s1 _____0_506093(.DIN1 (_____0__28538), .DIN2 (________27203), .Q
       (________28539));
  or2s1 _______506094(.DIN1 (________28535), .DIN2 (________28534), .Q
       (________28536));
  nnd2s1 ______506095(.DIN1 (_____0___35741), .DIN2 (_________22033),
       .Q (________28532));
  and2s1 _______506096(.DIN1 (________27971), .DIN2 (_____0__28530), .Q
       (________28531));
  nnd2s1 ______506097(.DIN1 (________28528), .DIN2 (____9___29002), .Q
       (_____9__28529));
  nor2s1 _______506098(.DIN1 (________28509), .DIN2 (________27544), .Q
       (________28527));
  or2s1 _____9_506099(.DIN1 (________26445), .DIN2 (________28525), .Q
       (________28526));
  nnd2s1 _____9_506100(.DIN1 (________28176), .DIN2 (________28523), .Q
       (________28524));
  nnd2s1 _____0_506101(.DIN1 (____9___28551), .DIN2 (________27666), .Q
       (________28522));
  nor2s1 _____0_506102(.DIN1 (________28444), .DIN2 (___9____27816), .Q
       (________28521));
  nor2s1 _______506103(.DIN1 (____9___27566), .DIN2 (_________41158),
       .Q (_____0__28520));
  nnd2s1 _______506104(.DIN1 (________28513), .DIN2 (___0____22302), .Q
       (________28518));
  and2s1 ______506105(.DIN1 (___0_0__27836), .DIN2 (__9_____30314), .Q
       (________28517));
  nnd2s1 _______506106(.DIN1 (_____0__28538), .DIN2 (________28001), .Q
       (________28516));
  nnd2s1 _______506107(.DIN1 (____9___28642), .DIN2 (____9___27297), .Q
       (________28515));
  nnd2s1 ______506108(.DIN1 (________28513), .DIN2 (_______22206), .Q
       (________28514));
  and2s1 _______506109(.DIN1 (___00___27829), .DIN2 (__9__9__30319), .Q
       (________28512));
  nor2s1 _______506110(.DIN1 (________27325), .DIN2 (________28179), .Q
       (_____0__28511));
  nnd2s1 _______506111(.DIN1 (_________32692), .DIN2 (________28509),
       .Q (_____9__28510));
  and2s1 _______506112(.DIN1 (_____0___35741), .DIN2
       (_____________________________________9______21877), .Q
       (________28508));
  nor2s1 _____9_506113(.DIN1 (________26612), .DIN2 (___9____27818), .Q
       (________28506));
  or2s1 _____0_506114(.DIN1 (___0_____40592), .DIN2 (_____0___35741),
       .Q (________28505));
  and2s1 _____506115(.DIN1 (__9_____30306), .DIN2 (___0____27850), .Q
       (________28504));
  or2s1 _______506116(.DIN1 (_____0__28502), .DIN2 (____0___28478), .Q
       (________28503));
  or2s1 _______506117(.DIN1 (________28500), .DIN2 (___9____27812), .Q
       (_____9__28501));
  nor2s1 _____9_506118(.DIN1 (__9_9___30449), .DIN2 (________28156), .Q
       (________28499));
  and2s1 _______506119(.DIN1 (___9____27817), .DIN2 (________28497), .Q
       (________28498));
  nnd2s1 _______506120(.DIN1 (___0____27857), .DIN2 (________28495), .Q
       (________28496));
  nnd2s1 _______506121(.DIN1 (____09__29106), .DIN2 (___0_9__27844), .Q
       (________28494));
  nnd2s1 _______506122(.DIN1 (___00___27834), .DIN2 (inData[22]), .Q
       (________28493));
  nor2s1 ____00_506123(.DIN1 (__9_00__30272), .DIN2 (________28486), .Q
       (________28980));
  or2s1 ____00_506124(.DIN1 (________28485), .DIN2 (___0____27890), .Q
       (________29307));
  nnd2s1 ______506125(.DIN1 (___990__27822), .DIN2 (________28484), .Q
       (________29251));
  nor2s1 _______506126(.DIN1 (___0_0___40462), .DIN2 (________27612),
       .Q (________29220));
  and2s1 _______506127(.DIN1 (________27612), .DIN2 (___0_0___40462),
       .Q (________29221));
  nnd2s1 _______506128(.DIN1 (________28483), .DIN2 (________27155), .Q
       (________29205));
  nor2s1 ______506129(.DIN1 (________28344), .DIN2 (_________41158), .Q
       (________28877));
  and2s1 _______506130(.DIN1 (______9__33037), .DIN2 (________27579),
       .Q (______0__32744));
  and2s1 _______506131(.DIN1 (___9____27815), .DIN2 (_____9___34752),
       .Q (_________32349));
  and2s1 _______506132(.DIN1 (________28482), .DIN2 (___9____27808), .Q
       (_________33026));
  and2s1 ____506133(.DIN1 (_____0__27987), .DIN2 (_____0__28481), .Q
       (________29297));
  nor2s1 ______506134(.DIN1 (________28089), .DIN2 (___00___27827), .Q
       (________28867));
  xor2s1 ____0__506135(.DIN1
       (__________________________________9__________), .DIN2
       (_________37867), .Q (______0__35957));
  nor2s1 ____0__506136(.DIN1 (_________41273), .DIN2 (___0____27903),
       .Q (_____9__28862));
  nnd2s1 ____0__506137(.DIN1 (________28083), .DIN2 (___0____27888), .Q
       (___0_____30697));
  and2s1 ____0__506138(.DIN1 (_____0__27958), .DIN2 (___0_____30805),
       .Q (________29338));
  nnd2s1 ____0__506139(.DIN1 (____9___28289), .DIN2 (____09__28480), .Q
       (_____9__29334));
  or2s1 ____0__506140(.DIN1 (____0___28479), .DIN2 (________28096), .Q
       (____0___29471));
  xor2s1 ____0__506141(.DIN1
       (_________________________________________9_), .DIN2
       (__________________________________9__________), .Q
       (________28979));
  nnd2s1 ____0__506142(.DIN1 (____0___28114), .DIN2 (________27468), .Q
       (________29300));
  nor2s1 ____0__506143(.DIN1 (_________31762), .DIN2 (___0____27882),
       .Q (________29342));
  or2s1 ____0__506144(.DIN1 (____0___28479), .DIN2 (___0____27905), .Q
       (________29313));
  or2s1 _____9_506145(.DIN1 (_____0___31604), .DIN2 (__9__9__30337), .Q
       (________29183));
  nor2s1 _____0_506146(.DIN1 (________26333), .DIN2 (____0___28478), .Q
       (____0___29198));
  nor2s1 ______506147(.DIN1 (__9_____29870), .DIN2 (__9__9__30337), .Q
       (_____0__28890));
  nnd2s1 ______506148(.DIN1 (___9____27807), .DIN2 (__9_____30024), .Q
       (________29178));
  and2s1 _______506149(.DIN1 (_____0__27524), .DIN2 (____0___28477), .Q
       (__99____30490));
  nor2s1 _______506150(.DIN1 (_________37789), .DIN2 (________27618),
       .Q (________29168));
  or2s1 _______506151(.DIN1 (____0___28476), .DIN2 (___0____27841), .Q
       (_____0___32777));
  nnd2s1 ______506152(.DIN1 (____0___28475), .DIN2 (________28585), .Q
       (____00__29194));
  nor2s1 _______506153(.DIN1 (__909___29719), .DIN2 (____0___28558), .Q
       (________29172));
  nor2s1 _______506154(.DIN1 (_________37867), .DIN2 (_________41367),
       .Q (________29497));
  nor2s1 _______506155(.DIN1 (________28171), .DIN2 (___9____27811), .Q
       (________29259));
  or2s1 _______506156(.DIN1 (____0___28474), .DIN2 (____0___28473), .Q
       (________29268));
  nor2s1 _______506157(.DIN1 (___0_0___40463), .DIN2 (________27618),
       .Q (____9___29273));
  nnd2s1 _______506158(.DIN1 (________28513), .DIN2 (________28151), .Q
       (___9909__39806));
  nnd2s1 _______506159(.DIN1 (___0_____31204), .DIN2 (____0____31581),
       .Q (__9_0___29897));
  nor2s1 ______506160(.DIN1 (________28937), .DIN2 (___9____27810), .Q
       (___0_____30719));
  nnd2s1 ____0__506161(.DIN1 (___9____28692), .DIN2 (____0___28472), .Q
       (______9__32330));
  and2s1 _____506162(.DIN1 (________28482), .DIN2 (___0____27838), .Q
       (______0__33028));
  and2s1 _______506163(.DIN1 (________27618), .DIN2 (___0_0___40463),
       .Q (__9__9__30225));
  nnd2s1 _______506164(.DIN1 (_________41367), .DIN2 (_________37867),
       .Q (____09___35375));
  nor2s1 _____9_506165(.DIN1 (____00__28471), .DIN2 (_____0___35741),
       .Q (______0__35784));
  and2s1 _______506166(.DIN1 (_____9__27471), .DIN2 (________28044), .Q
       (____9____32439));
  and2s1 _____9_506167(.DIN1 (____9___28470), .DIN2 (____0___26145), .Q
       (____00___31507));
  dffacs1 _______________________________________________506168(.CLRB
       (reset), .CLK (clk), .DIN (_____9__28051), .QN
       (_____________________________________________21924));
  nnd2s1 ____0_506169(.DIN1 (________27943), .DIN2 (____9___28469), .Q
       (___0_____40166));
  hi1s1 ____09_506170(.DIN (________28968), .Q (________29323));
  hi1s1 ____09_506171(.DIN (_____0__29046), .Q (____0___29280));
  hi1s1 ____506172(.DIN (_____9__28871), .Q (________29241));
  xor2s1 ____9__506173(.DIN1 (___0__0__40413), .DIN2 (________28140),
       .Q (____9___28468));
  nor2s1 _______506174(.DIN1 (____9___28466), .DIN2 (________27581), .Q
       (____9___28467));
  xnr2s1 _______506175(.DIN1
       (_____________________________________0___0_), .DIN2
       (_____________________________________________21795), .Q
       (____9___28465));
  nnd2s1 _______506176(.DIN1 (_____0__28306), .DIN2 (___0_____30709),
       .Q (____9___28464));
  nnd2s1 _______506177(.DIN1 (________27603), .DIN2 (___9_9__26882), .Q
       (____9___28463));
  nor2s1 _______506178(.DIN1 (___9____26881), .DIN2 (________27603), .Q
       (____90__28462));
  nor2s1 _______506179(.DIN1 (___0__9__40590), .DIN2 (________27644),
       .Q (_____9__28461));
  nnd2s1 _______506180(.DIN1 (___0_____40326), .DIN2 (________22563),
       .Q (________28460));
  nor2s1 ______506181(.DIN1 (________29225), .DIN2 (____9___27648), .Q
       (________28459));
  nor2s1 _______506182(.DIN1 (________28457), .DIN2 (________28456), .Q
       (________28458));
  nor2s1 _______506183(.DIN1 (inData[11]), .DIN2 (______0__35537), .Q
       (________28455));
  nor2s1 ______506184(.DIN1 (________28860), .DIN2 (___90___27748), .Q
       (_____0__28453));
  nnd2s1 _______506185(.DIN1 (________25513), .DIN2 (___900__27742), .Q
       (_____9__28452));
  and2s1 ______506186(.DIN1 (____0___27306), .DIN2 (__9_____29941), .Q
       (________28451));
  nor2s1 _____506187(.DIN1 (_____9__28081), .DIN2 (________27599), .Q
       (________28450));
  or2s1 _____0_506188(.DIN1 (__9__9__30010), .DIN2 (___9____27756), .Q
       (________28449));
  and2s1 ______506189(.DIN1 (___90___27746), .DIN2 (________28447), .Q
       (________28448));
  nnd2s1 _______506190(.DIN1 (________28445), .DIN2 (________28444), .Q
       (________28446));
  and2s1 ______506191(.DIN1 (___9_____39219), .DIN2 (___0__0__40599),
       .Q (_____0__28443));
  nor2s1 _______506192(.DIN1 (________28441), .DIN2 (________28427), .Q
       (_____9__28442));
  nor2s1 _______506193(.DIN1 (inData[10]), .DIN2 (______0__35537), .Q
       (________28440));
  nor2s1 ______506194(.DIN1 (________27600), .DIN2 (________27513), .Q
       (________28439));
  nnd2s1 _______506195(.DIN1 (_________41166), .DIN2 (___009___30634),
       .Q (________28438));
  nnd2s1 _____9_506196(.DIN1 (___9____27753), .DIN2 (________24049), .Q
       (________28437));
  nnd2s1 _____9_506197(.DIN1 (________27698), .DIN2 (___9____29597), .Q
       (________28436));
  nor2s1 _____506198(.DIN1 (________28070), .DIN2 (_____0__27696), .Q
       (________28435));
  nnd2s1 _______506199(.DIN1 (________27727), .DIN2 (_____9__27967), .Q
       (________28434));
  nnd2s1 _______506200(.DIN1 (________27729), .DIN2 (clk), .Q
       (_____0__28433));
  nor2s1 _______506201(.DIN1 (_____0__28298), .DIN2 (__9_____30417), .Q
       (_____9__28432));
  nor2s1 _______506202(.DIN1 (____0____32541), .DIN2 (____9___27739),
       .Q (________28431));
  nnd2s1 _______506203(.DIN1 (_________41166), .DIN2 (________27690),
       .Q (________28430));
  and2s1 _______506204(.DIN1 (______0__35537), .DIN2 (____99__22938),
       .Q (________28429));
  nor2s1 ______506205(.DIN1 (___0_____31262), .DIN2 (________28427), .Q
       (________28428));
  nor2s1 ______506206(.DIN1
       (______________________________________________21955), .DIN2
       (___9_____39219), .Q (________28426));
  nor2s1 _______506207(.DIN1 (_____0__28424), .DIN2 (_____9__28423), .Q
       (________28425));
  nnd2s1 _____0_506208(.DIN1 (________27534), .DIN2 (________24902), .Q
       (________28422));
  hi1s1 _______506209(.DIN (________28420), .Q (________28421));
  xor2s1 _______506210(.DIN1 (__________0_), .DIN2 (___0_9___40452), .Q
       (________28419));
  and2s1 _______506211(.DIN1 (________27678), .DIN2 (__9__9__29779), .Q
       (________28418));
  nnd2s1 _____9_506212(.DIN1 (________27682), .DIN2 (__9_99__29992), .Q
       (________28417));
  nnd2s1 _______506213(.DIN1 (__90____29661), .DIN2 (_________41162),
       .Q (________28416));
  nor2s1 _______506214(.DIN1 (____0___24275), .DIN2 (___9_____39219),
       .Q (________28415));
  nnd2s1 _______506215(.DIN1 (________27596), .DIN2 (_____0__29175), .Q
       (_____0__28414));
  or2s1 ______506216(.DIN1 (________27220), .DIN2 (________28412), .Q
       (_____9__28413));
  nnd2s1 _______506217(.DIN1 (________28412), .DIN2 (__9990), .Q
       (________28411));
  nor2s1 _______506218(.DIN1 (________27693), .DIN2 (________29119), .Q
       (________28410));
  and2s1 _______506219(.DIN1 (________28408), .DIN2 (________28407), .Q
       (________28409));
  nor2s1 _______506220(.DIN1 (___0_____30764), .DIN2 (________27689),
       .Q (________28406));
  nnd2s1 _____506221(.DIN1 (___0_____40222), .DIN2 (________27685), .Q
       (________28405));
  or2s1 _____9_506222(.DIN1 (___9____29571), .DIN2 (________27684), .Q
       (_____0__28404));
  nor2s1 _____9_506223(.DIN1 (________27679), .DIN2 (________27149), .Q
       (_____9__28403));
  nor2s1 _____506224(.DIN1 (_____0__27677), .DIN2 (________27697), .Q
       (________28402));
  nnd2s1 ____9__506225(.DIN1 (________27152), .DIN2 (________27702), .Q
       (________28401));
  or2s1 ____9__506226(.DIN1 (_____9__27601), .DIN2 (________28399), .Q
       (________28400));
  nor2s1 ____9__506227(.DIN1 (___9____23205), .DIN2 (___9_____39219),
       .Q (________28398));
  and2s1 ____9__506228(.DIN1 (___0____27876), .DIN2 (________28628), .Q
       (________28397));
  nnd2s1 ____9__506229(.DIN1 (_____0__28395), .DIN2 (________29311), .Q
       (________28396));
  nnd2s1 ____9__506230(.DIN1 (___90___27750), .DIN2 (________28454), .Q
       (_____9__28394));
  nor2s1 ____9__506231(.DIN1 (________28392), .DIN2 (________27595), .Q
       (________28393));
  nnd2s1 _____506232(.DIN1 (________28390), .DIN2 (______0___22057), .Q
       (________28391));
  nnd2s1 _____9_506233(.DIN1 (____09__27659), .DIN2 (________26263), .Q
       (________28389));
  nor2s1 _____9_506234(.DIN1 (________25933), .DIN2 (_____9__27558), .Q
       (________28388));
  and2s1 _____9_506235(.DIN1 (____99__27653), .DIN2 (________28386), .Q
       (________28387));
  and2s1 _______506236(.DIN1 (___9____27760), .DIN2 (________28507), .Q
       (_____0__28385));
  and2s1 _______506237(.DIN1 (____0___28383), .DIN2 (____0___28382), .Q
       (____09__28384));
  nor2s1 ______506238(.DIN1 (____0___28380), .DIN2 (____9___28194), .Q
       (____0___28381));
  nnd2s1 _______506239(.DIN1 (________28155), .DIN2 (___0_____30807),
       .Q (____0___28379));
  nnd2s1 _______506240(.DIN1 (____0___28377), .DIN2 (________29537), .Q
       (____0___28378));
  hi1s1 ____0__506241(.DIN (____9___28373), .Q (____9___28374));
  hi1s1 ____0_506242(.DIN (___0_____40433), .Q (____9___28371));
  nnd2s1 _______506243(.DIN1 (________27249), .DIN2 (________27546), .Q
       (____9___28370));
  nor2s1 _______506244(.DIN1 (_____9__28368), .DIN2 (____00__27480), .Q
       (____90__28369));
  or2s1 _____0_506245(.DIN1 (___0_90__31108), .DIN2 (____9___27563), .Q
       (________28367));
  nnd2s1 _____0_506246(.DIN1 (____09__27577), .DIN2 (________29108), .Q
       (________28366));
  and2s1 _____0_506247(.DIN1 (________27588), .DIN2 (________28364), .Q
       (________28365));
  nnd2s1 _____506248(.DIN1 (________27152), .DIN2 (___9____26886), .Q
       (________28363));
  nor2s1 _______506249(.DIN1 (_________33321), .DIN2 (________23892),
       .Q (________28362));
  nnd2s1 _______506250(.DIN1 (________28264), .DIN2 (_____9__28360), .Q
       (_____0__28361));
  nor2s1 _______506251(.DIN1 (________26602), .DIN2 (________28357), .Q
       (________28359));
  nor2s1 _______506252(.DIN1 (____0___27570), .DIN2 (________28357), .Q
       (________28358));
  nor2s1 ______506253(.DIN1 (__9_0___29904), .DIN2 (________28236), .Q
       (________28356));
  nor2s1 ______506254(.DIN1 (____0___26324), .DIN2 (________27625), .Q
       (________28355));
  nor2s1 _______506255(.DIN1 (___0_99__40460), .DIN2 (____990__33424),
       .Q (________28354));
  nnd2s1 _______506256(.DIN1 (_____9__28256), .DIN2 (________23575), .Q
       (________28353));
  nor2s1 _______506257(.DIN1 (____99__27299), .DIN2 (____9___27562), .Q
       (________28352));
  and2s1 _______506258(.DIN1 (_____9__28350), .DIN2 (________28304), .Q
       (_____0__28351));
  nnd2s1 _______506259(.DIN1 (____90__27472), .DIN2 (________27310), .Q
       (________28349));
  nnd2s1 _______506260(.DIN1 (____00__27569), .DIN2 (inData[10]), .Q
       (________28348));
  nor2s1 _______506261(.DIN1 (____0___26687), .DIN2 (________27629), .Q
       (________28347));
  nnd2s1 ______506262(.DIN1 (________27631), .DIN2 (_________32260), .Q
       (________28346));
  or2s1 _______506263(.DIN1 (________28344), .DIN2 (________28343), .Q
       (________28345));
  nor2s1 ______506264(.DIN1 (_________41164), .DIN2 (___0_9__28804), .Q
       (_____0__28342));
  nor2s1 _______506265(.DIN1 (___0_00__40461), .DIN2
       (__________________________________9__________), .Q
       (_____9__28341));
  nnd2s1 _______506266(.DIN1 (________27632), .DIN2 (________26703), .Q
       (________28340));
  nnd2s1 _______506267(.DIN1 (_____9__27667), .DIN2 (_____0__27687), .Q
       (________28339));
  nor2s1 ______506268(.DIN1 (________28337), .DIN2 (___99___27823), .Q
       (________28338));
  nor2s1 _______506269(.DIN1 (________26536), .DIN2 (___0_9__28804), .Q
       (________28336));
  or2s1 ______506270(.DIN1 (________26816), .DIN2 (________28334), .Q
       (________28335));
  nnd2s1 _______506271(.DIN1 (________27580), .DIN2 (________29112), .Q
       (_____0__28333));
  nnd2s1 _______506272(.DIN1 (_________35859), .DIN2
       (_____________________________________________21897), .Q
       (_____9__28332));
  nor2s1 _____9_506273(.DIN1 (________28063), .DIN2 (______0__41170),
       .Q (________28331));
  nor2s1 _____0_506274(.DIN1 (_____9__29455), .DIN2 (___0_9__28804), .Q
       (________28330));
  nor2s1 _______506275(.DIN1 (________27423), .DIN2 (___09___28829), .Q
       (________28329));
  nnd2s1 _______506276(.DIN1
       (__________________________________9__________), .DIN2
       (_________________________________________9_), .Q
       (________28328));
  nor2s1 ______506277(.DIN1 (________27715), .DIN2 (________27663), .Q
       (________28327));
  and2s1 ______506278(.DIN1 (__9_____30035), .DIN2 (________28307), .Q
       (________28326));
  or2s1 _______506279(.DIN1 (______0__41160), .DIN2 (__9_____29883), .Q
       (________28325));
  and2s1 _______506280(.DIN1
       (__________________________________9__________), .DIN2
       (___0_00__40461), .Q (_____0__28324));
  nnd2s1 _______506281(.DIN1 (_________31778), .DIN2 (________27719),
       .Q (_____9__28323));
  nor2s1 ______506282(.DIN1 (__9__9__29935), .DIN2 (________27725), .Q
       (________28322));
  nnd2s1 _______506283(.DIN1 (________28320), .DIN2 (________28316), .Q
       (________28321));
  nor2s1 _______506284(.DIN1 (________28318), .DIN2 (________27525), .Q
       (________28319));
  nor2s1 ______506285(.DIN1 (________28316), .DIN2 (____0___28295), .Q
       (________28317));
  nor2s1 _______506286(.DIN1 (_____0__27345), .DIN2 (___9_9__27794), .Q
       (________28315));
  nnd2s1 _______506287(.DIN1 (________27671), .DIN2 (____0___29010), .Q
       (_____0__28314));
  nnd2s1 _______506288(.DIN1 (________27516), .DIN2 (________27282), .Q
       (_____9__28313));
  or2s1 _______506289(.DIN1 (________28311), .DIN2 (________27502), .Q
       (________28312));
  xor2s1 ____9_506290(.DIN1 (________27226), .DIN2 (________22511), .Q
       (___9_9__29601));
  hi1s1 ____09_506291(.DIN (___9____28692), .Q (________28861));
  nor2s1 _______506292(.DIN1 (_____9__27195), .DIN2 (___0_9___31405),
       .Q (____0___28926));
  nnd2s1 _______506293(.DIN1 (________27716), .DIN2 (________27286), .Q
       (___9____29584));
  nor2s1 ____0__506294(.DIN1 (____9___26677), .DIN2 (_____9__27695), .Q
       (___9____28674));
  nor2s1 ____0_506295(.DIN1 (__9_____30260), .DIN2 (__9__9__30262), .Q
       (__9_9___29801));
  and2s1 ____0_506296(.DIN1 (________27683), .DIN2 (__9_9___30267), .Q
       (_____0__29117));
  nnd2s1 ____0__506297(.DIN1 (________27692), .DIN2 (__9_____30162), .Q
       (___9____28675));
  and2s1 ____00_506298(.DIN1 (________27688), .DIN2 (________28309), .Q
       (______9__31660));
  nnd2s1 ____00_506299(.DIN1 (_____9__27705), .DIN2 (________28308), .Q
       (___9____28676));
  nnd2s1 ____506300(.DIN1 (________27680), .DIN2 (_____9___31697), .Q
       (____0___29101));
  nor2s1 _______506301(.DIN1 (___0_____31274), .DIN2 (________27643),
       .Q (_____9__28546));
  nor2s1 _______506302(.DIN1 (___0_0___40464), .DIN2
       (__________________________________9__________), .Q
       (________28865));
  nor2s1 _______506303(.DIN1 (___0_____30709), .DIN2 (________27603),
       .Q (________28848));
  and2s1 _______506304(.DIN1
       (__________________________________9__________), .DIN2
       (_________________________________________9___21861), .Q
       (_____9__28998));
  nnd2s1 _______506305(.DIN1 (___0_____40326), .DIN2 (___0_____40415),
       .Q (____9___28548));
  or2s1 _______506306(.DIN1 (____0___25866), .DIN2 (___0_9___31405), .Q
       (________28868));
  and2s1 _______506307(.DIN1 (________28307), .DIN2 (___0__0__31168),
       .Q (________29166));
  and2s1 _______506308(.DIN1
       (__________________________________9__________), .DIN2
       (___0_0___40464), .Q (________28864));
  nor2s1 _______506309(.DIN1
       (_________________________________________9___21861), .DIN2
       (_________38280), .Q (____90__28999));
  or2s1 _______506310(.DIN1
       (_________________________________________0___21862), .DIN2
       (_________38280), .Q (_____0__28872));
  nor2s1 _______506311(.DIN1 (__9_____30198), .DIN2 (__9_____29870), .Q
       (____9___28547));
  nnd2s1 _______506312(.DIN1
       (__________________________________9__________), .DIN2
       (_________________________________________0___21862), .Q
       (________28873));
  dffacs2 _________________506313(.CLRB (reset), .CLK (clk), .DIN
       (________27622), .Q (______________22066));
  nor2s1 _______506314(.DIN1 (________22537), .DIN2 (_____0__28306), .Q
       (____99__29008));
  nnd2s1 ____0__506315(.DIN1 (________27152), .DIN2 (_________41168),
       .Q (__9_09__30281));
  nor2s1 ____0__506316(.DIN1 (________27700), .DIN2 (________27699), .Q
       (________29153));
  dffacs1 _______________________________________________506317(.CLRB
       (reset), .CLK (clk), .DIN (________27641), .Q (___0_____40423));
  nnd2s1 _______506318(.DIN1 (________28305), .DIN2 (________28304), .Q
       (________28961));
  dffacs1 ______________________________________506319(.CLRB (reset),
       .CLK (clk), .DIN (___90___27745), .Q (___0_____40585));
  hi1s1 ____09_506320(.DIN (__90_9__29717), .Q (________29051));
  hi1s1 ____09_506321(.DIN (___0_____30961), .Q (__9_____29735));
  dffacs1 ______________________________________________0_506322(.CLRB
       (reset), .CLK (clk), .DIN (________27675), .Q
       (__________________________________________________________________21983));
  nor2s1 ______506323(.DIN1 (____9___27298), .DIN2 (____9___27736), .Q
       (___0_____40400));
  and2s1 _______506324(.DIN1 (___9_____39219), .DIN2
       (_________________________________________9___21943), .Q
       (________28303));
  nnd2s1 _______506325(.DIN1 (____9___27733), .DIN2 (________29537), .Q
       (________28302));
  nnd2s1 ____506326(.DIN1 (________27691), .DIN2 (________27701), .Q
       (________28301));
  nnd2s1 ______506327(.DIN1 (_____0__28298), .DIN2 (________27274), .Q
       (________28299));
  dffacs1 _______________506328(.CLRB (reset), .CLK (clk), .DIN
       (_____0__28306), .Q (outData[2]));
  nor2s1 _______506329(.DIN1 (_____9__29425), .DIN2 (____0___28295), .Q
       (____0___28296));
  and2s1 _______506330(.DIN1 (_____0__27593), .DIN2 (____0___28293), .Q
       (____0___28294));
  hi1s1 _______506331(.DIN (____9___28286), .Q (____9___28287));
  nor2s1 _______506332(.DIN1 (____0___27210), .DIN2 (________28283), .Q
       (_____9__28284));
  nor2s1 _______506333(.DIN1 (________28281), .DIN2 (____0___28295), .Q
       (________28282));
  hi1s1 _______506334(.DIN (____0____31556), .Q (________28280));
  or2s1 _______506335(.DIN1 (________28320), .DIN2 (____0___28295), .Q
       (________28279));
  nnd2s1 _____0_506336(.DIN1 (________27152), .DIN2 (________28277), .Q
       (________28278));
  or2s1 ______506337(.DIN1 (___0__0__40581), .DIN2
       (__________________________________9__________), .Q
       (_____0__28276));
  and2s1 _______506338(.DIN1 (_________34796), .DIN2 (_________33321),
       .Q (_____9__28275));
  nor2s1 _______506339(.DIN1 (___9____26927), .DIN2 (_____9__27713), .Q
       (________28274));
  nor2s1 _______506340(.DIN1 (________27447), .DIN2 (____0___28295), .Q
       (________28273));
  nnd2s1 _______506341(.DIN1 (____9___27567), .DIN2 (__9990), .Q
       (________28272));
  nor2s1 _______506342(.DIN1
       (__________________________________9__________), .DIN2
       (_________38164), .Q (________28271));
  nnd2s1 _______506343(.DIN1 (_________33321), .DIN2
       (______________22065), .Q (________28270));
  nor2s1 _______506344(.DIN1 (__9__0__30394), .DIN2 (________28268), .Q
       (________28269));
  nor2s1 _____9_506345(.DIN1 (________26291), .DIN2 (____9___27565), .Q
       (________28267));
  nnd2s1 _____0_506346(.DIN1 (_________41174), .DIN2 (__90_9__29688),
       .Q (_____9__28266));
  nnd2s1 _____0_506347(.DIN1 (________28264), .DIN2 (________26755), .Q
       (________28265));
  nor2s1 ______506348(.DIN1 (____9___27561), .DIN2 (____0___28295), .Q
       (________28263));
  nnd2s1 _______506349(.DIN1 (________27555), .DIN2 (________28261), .Q
       (________28262));
  nnd2s1 ______506350(.DIN1 (_____9__29314), .DIN2 (_________41176), .Q
       (________28260));
  nor2s1 _______506351(.DIN1 (_____0__22578), .DIN2 (___0_____40100),
       .Q (________28259));
  nor2s1 _______506352(.DIN1 (___0____26078), .DIN2 (____9___27650), .Q
       (________28258));
  nnd2s1 _______506353(.DIN1 (_____9__28256), .DIN2 (________26532), .Q
       (_____0__28257));
  nor2s1 _______506354(.DIN1 (____9____32449), .DIN2 (_____9__27722),
       .Q (________28255));
  and2s1 _______506355(.DIN1 (________27548), .DIN2 (__9__0__30130), .Q
       (________28254));
  and2s1 _______506356(.DIN1 (________27634), .DIN2 (________28252), .Q
       (________28253));
  nor2s1 _______506357(.DIN1 (________27956), .DIN2 (________28250), .Q
       (________28251));
  nor2s1 _______506358(.DIN1 (____99__26863), .DIN2 (________28334), .Q
       (________28249));
  and2s1 _______506359(.DIN1 (_____0__28247), .DIN2 (_____9__28246), .Q
       (________28248));
  nor2s1 _______506360(.DIN1 (___0____26968), .DIN2 (___0_9__28804), .Q
       (________28245));
  nor2s1 _______506361(.DIN1 (___9_0__26883), .DIN2 (____0___27572), .Q
       (________28244));
  nor2s1 _______506362(.DIN1 (________27556), .DIN2 (____0___29200), .Q
       (________28243));
  nor2s1 _______506363(.DIN1 (____9___25956), .DIN2 (____0___27575), .Q
       (________28241));
  nor2s1 ______506364(.DIN1 (________28268), .DIN2 (________27531), .Q
       (________28240));
  nor2s1 _______506365(.DIN1 (_____9__27523), .DIN2 (___0_____31336),
       .Q (________28239));
  nor2s1 _______506366(.DIN1 (_____0__27515), .DIN2 (__9_____30417), .Q
       (_____0__28238));
  nor2s1 _______506367(.DIN1 (________28236), .DIN2 (________28213), .Q
       (_____9__28237));
  nor2s1 _______506368(.DIN1 (________27536), .DIN2 (__9_____30417), .Q
       (________28235));
  nor2s1 _______506369(.DIN1 (________26749), .DIN2 (________28233), .Q
       (________28234));
  nnd2s1 _______506370(.DIN1 (_________38280), .DIN2 (_________37789),
       .Q (________28232));
  nor2s1 _______506371(.DIN1 (________28230), .DIN2 (________27172), .Q
       (________28231));
  nnd2s1 _______506372(.DIN1
       (__________________________________9__________), .DIN2
       (____99___36174), .Q (_____0__28229));
  nor2s1 _______506373(.DIN1 (____99___36174), .DIN2
       (__________________________________9__________), .Q
       (_____9__28228));
  nor2s1 _____506374(.DIN1 (________27235), .DIN2 (___09___28829), .Q
       (________28227));
  or2s1 _____9_506375(.DIN1 (________28170), .DIN2 (________28225), .Q
       (________28226));
  nor2s1 _____9_506376(.DIN1 (________28223), .DIN2 (________27661), .Q
       (________28224));
  nnd2s1 _____9_506377(.DIN1 (___0__0__40413), .DIN2 (_________33321),
       .Q (________28222));
  and2s1 _____0_506378(.DIN1 (________27517), .DIN2 (_____9___32965),
       .Q (________28221));
  nor2s1 _____0_506379(.DIN1 (________27275), .DIN2 (__9_____30417), .Q
       (_____0__28220));
  or2s1 _____0_506380(.DIN1 (________27991), .DIN2 (_________32692), .Q
       (_____9__28219));
  and2s1 _____0_506381(.DIN1 (__99____30468), .DIN2 (________27252), .Q
       (________28218));
  or2s1 _______506382(.DIN1 (________28216), .DIN2 (________27557), .Q
       (________28217));
  nor2s1 _______506383(.DIN1 (____0___25771), .DIN2 (________27630), .Q
       (________28215));
  nnd2s1 _______506384(.DIN1 (________28213), .DIN2 (____09__29106), .Q
       (________28214));
  nnd2s1 _______506385(.DIN1 (________28211), .DIN2 (_____0__28210), .Q
       (________28212));
  nor2s1 _______506386(.DIN1 (________28874), .DIN2 (________28159), .Q
       (____09__28209));
  nor2s1 _______506387(.DIN1 (____0___28207), .DIN2 (____0___28206), .Q
       (____0___28208));
  or2s1 _______506388(.DIN1 (________28600), .DIN2 (________27621), .Q
       (____0___28205));
  nnd2s1 _______506389(.DIN1 (________27586), .DIN2 (_________31731),
       .Q (____0___28204));
  or2s1 _______506390(.DIN1 (____0___28202), .DIN2 (____0___28201), .Q
       (____0___28203));
  or2s1 _______506391(.DIN1 (________28386), .DIN2 (____0___28295), .Q
       (____00__28200));
  or2s1 _______506392(.DIN1 (____9___28198), .DIN2 (___09___28829), .Q
       (____99__28199));
  or2s1 _______506393(.DIN1 (____9___28196), .DIN2 (_____9__27542), .Q
       (____9___28197));
  nnd2s1 _______506394(.DIN1 (____9___28194), .DIN2 (____0___29285), .Q
       (____9___28195));
  nor2s1 _______506395(.DIN1 (________27530), .DIN2 (__9__0__30291), .Q
       (____9___28193));
  and2s1 ______506396(.DIN1 (_____9__28368), .DIN2 (________29537), .Q
       (____9___28192));
  nor2s1 _______506397(.DIN1 (____0___27571), .DIN2 (________27519), .Q
       (____90__28191));
  nor2s1 _____9_506398(.DIN1 (________28189), .DIN2 (____0___28295), .Q
       (_____9__28190));
  nnd2s1 _____9_506399(.DIN1 (_____9__27471), .DIN2 (________28187), .Q
       (________28188));
  nnd2s1 ______506400(.DIN1 (____90__27472), .DIN2 (________28936), .Q
       (________28186));
  nnd2s1 _______506401(.DIN1 (____90__27472), .DIN2 (________28541), .Q
       (________28185));
  nnd2s1 _______506402(.DIN1 (________27152), .DIN2 (____00__29009), .Q
       (________28184));
  nor2s1 ______506403(.DIN1 (___0_____31182), .DIN2 (____0___28295), .Q
       (________28183));
  or2s1 _______506404(.DIN1 (_____0__28181), .DIN2 (__9_____30417), .Q
       (________28182));
  or2s1 _______506405(.DIN1 (___9____29606), .DIN2 (_____9__27506), .Q
       (_____9__28180));
  hi1s1 _______506406(.DIN (________28177), .Q (________28178));
  nor2s1 ____0__506407(.DIN1 (________27497), .DIN2 (________28337), .Q
       (_____0__28174));
  nor2s1 ____9__506408(.DIN1 (___9____26944), .DIN2 (_____0__27499), .Q
       (_____9__28173));
  nor2s1 _______506409(.DIN1 (________28171), .DIN2 (________28170), .Q
       (________28172));
  nor2s1 _______506410(.DIN1 (________27491), .DIN2 (________28268), .Q
       (________28489));
  nor2s1 _______506411(.DIN1 (___9____26924), .DIN2 (_____0__27637), .Q
       (________28957));
  nor2s1 ______506412(.DIN1 (_____9__28167), .DIN2 (___0_9__28804), .Q
       (___0_____31092));
  nor2s1 _____506413(.DIN1 (___09___27919), .DIN2 (________27503), .Q
       (________28869));
  or2s1 _______506414(.DIN1 (________29142), .DIN2 (__9_____29908), .Q
       (________28878));
  hi1s1 _______506415(.DIN (________28166), .Q (___9____29590));
  hi1s1 _______506416(.DIN (________28164), .Q (________28955));
  nnd2s1 _______506417(.DIN1 (_____0__27543), .DIN2 (____09___31598),
       .Q (________29026));
  nnd2s1 _______506418(.DIN1 (________28150), .DIN2 (________27417), .Q
       (_____0__29028));
  nor2s1 _______506419(.DIN1 (_____9__28147), .DIN2 (____0___27481), .Q
       (________28487));
  nor2s1 _______506420(.DIN1
       (_________________________________________________________________________________________22089),
       .DIN2 (__________________________________9__________), .Q
       (________29169));
  nor2s1 _______506421(.DIN1 (_________33321), .DIN2 (_________35622),
       .Q (________28939));
  nnd2s1 _______506422(.DIN1 (________28163), .DIN2 (________27425), .Q
       (_____9__28488));
  nnd2s1 _______506423(.DIN1 (_________33321), .DIN2
       (______________22066), .Q (________28892));
  and2s1 ______506424(.DIN1 (________27508), .DIN2 (________28162), .Q
       (________28974));
  or2s1 _______506425(.DIN1 (________28161), .DIN2 (________27230), .Q
       (______9__32703));
  or2s1 _______506426(.DIN1 (________28160), .DIN2 (________28159), .Q
       (____0___28930));
  nor2s1 _______506427(.DIN1 (___0_____31073), .DIN2 (________27590),
       .Q (________28491));
  hi1s1 _______506428(.DIN (_____0__28158), .Q (_____9__29218));
  hi1s1 _______506429(.DIN (_____9__28157), .Q (__9_____29979));
  hi1s1 _______506430(.DIN (________28156), .Q (_____0__28966));
  nnd2s1 _______506431(.DIN1 (________28155), .DIN2 (________28154), .Q
       (________28996));
  nnd2s1 _____506432(.DIN1 (____99__27568), .DIN2 (________27521), .Q
       (_____0___32780));
  nnd2s1 _____0_506433(.DIN1 (________27514), .DIN2 (__9_____30024), .Q
       (________28490));
  nor2s1 _____9_506434(.DIN1 (____0___29283), .DIN2 (________27510), .Q
       (________28942));
  nnd2s1 _______506435(.DIN1 (____0___27123), .DIN2 (___00____30606),
       .Q (_____9__28492));
  or2s1 _______506436(.DIN1 (________28149), .DIN2 (_____9___34186), .Q
       (________28898));
  hi1s1 ____09_506437(.DIN (___0____28783), .Q (____0___28927));
  and2s1 ______506438(.DIN1 (________28145), .DIN2 (________28152), .Q
       (___0_____31035));
  nor2s1 _______506439(.DIN1 (________28151), .DIN2 (___0_____40100),
       .Q (________29086));
  nnd2s1 _______506440(.DIN1 (________28150), .DIN2 (____0____31566),
       .Q (__9_____30039));
  nnd2s1 _______506441(.DIN1 (________27624), .DIN2 (________27288), .Q
       (________29084));
  or2s1 _______506442(.DIN1 (________28149), .DIN2 (____9___28194), .Q
       (________28911));
  nnd2s1 _______506443(.DIN1 (____90__27472), .DIN2 (_________32815),
       .Q (_________32649));
  nnd2s1 _______506444(.DIN1 (________27152), .DIN2 (____9___28196), .Q
       (___0_____30752));
  and2s1 _______506445(.DIN1 (________27623), .DIN2 (___0_____30943),
       .Q (___0_____30844));
  nor2s1 _______506446(.DIN1 (_____0__28148), .DIN2 (_____9__28147), .Q
       (________29056));
  nnd2s1 ______506447(.DIN1 (___0_____40326), .DIN2 (________28146), .Q
       (___0_____40320));
  and2s1 _____9_506448(.DIN1 (________28145), .DIN2 (___0_____31040),
       .Q (________29023));
  nnd2s1 _______506449(.DIN1 (________28143), .DIN2 (___09___27913), .Q
       (_____9__28871));
  hi1s1 _______506450(.DIN (_____0___35741), .Q (_________35718));
  dffacs1 _______________________________________________506451(.CLRB
       (reset), .CLK (clk), .DIN (________27635), .Q
       (_____________________________________________21953));
  dffacs1 ______________________________________506452(.CLRB (reset),
       .CLK (clk), .DIN (___90___27747), .QN (_____________22088));
  hi1s1 _______506453(.DIN (______0__36598), .Q (_________33924));
  or2s1 ______506454(.DIN1 (___0_____31073), .DIN2 (________29519), .Q
       (_____9__28989));
  nnd2s1 _______506455(.DIN1 (________28144), .DIN2 (inData[21]), .Q
       (_____0__29046));
  dffacs1 _________________________________________0_____506456(.CLRB
       (reset), .CLK (clk), .DIN (____9___27740), .Q (___0_____40573));
  nor2s1 _______506457(.DIN1 (_____0__27578), .DIN2 (____0___28295), .Q
       (_________33175));
  dffacs1 _______________________________________________506458(.CLRB
       (reset), .CLK (clk), .DIN (_____9__27628), .Q
       (_______________________________________________________________0__22010));
  nor2s1 _______506459(.DIN1 (___0_9__27911), .DIN2 (________28144), .Q
       (________28968));
  nnd2s1 ______506460(.DIN1 (________27717), .DIN2 (____0___26409), .Q
       (_________36087));
  dffacs1 _________________506461(.CLRB (reset), .CLK (clk), .DIN
       (________27645), .QN (______________22064));
  nor2s1 _______506462(.DIN1 (inData[21]), .DIN2 (________28143), .Q
       (___0_____30783));
  nnd2s1 _____9_506463(.DIN1 (______________22068), .DIN2
       (______9__32959), .Q (________28142));
  or2s1 _____0_506464(.DIN1 (___0_____40598), .DIN2 (________28140), .Q
       (________28141));
  nnd2s1 _____0_506465(.DIN1 (________28140), .DIN2 (___0_____40598),
       .Q (________28139));
  nor2s1 _______506466(.DIN1 (______9__32959), .DIN2 (________28140),
       .Q (_____0__28138));
  and2s1 _____9_506467(.DIN1 (________28140), .DIN2 (______9__32959),
       .Q (_____9__28137));
  nnd2s1 _______506468(.DIN1 (________27465), .DIN2 (inData[16]), .Q
       (________28136));
  nor2s1 _______506469(.DIN1 (___090___31413), .DIN2 (___9____27802),
       .Q (________28135));
  nnd2s1 _______506470(.DIN1 (________28133), .DIN2 (________26434), .Q
       (________28134));
  nor2s1 _____9_506471(.DIN1 (________28131), .DIN2 (________27455), .Q
       (________28132));
  nnd2s1 _______506472(.DIN1 (________27464), .DIN2 (________26376), .Q
       (________28130));
  nnd2s1 _______506473(.DIN1 (________27708), .DIN2 (_____0__28128), .Q
       (________28129));
  nnd2s1 _____9_506474(.DIN1 (____99__27479), .DIN2 (_____0__27231), .Q
       (_____9__28127));
  or2s1 ____9_506475(.DIN1 (________27454), .DIN2 (________28125), .Q
       (________28126));
  or2s1 ____9__506476(.DIN1 (____9___28196), .DIN2 (_____0__27453), .Q
       (________28124));
  and2s1 _____9_506477(.DIN1 (________27247), .DIN2 (________28122), .Q
       (________28123));
  nnd2s1 ______506478(.DIN1 (________28605), .DIN2 (________27159), .Q
       (________28121));
  xor2s1 ____00_506479(.DIN1
       (____________________________________________21818), .DIN2
       (_________35622), .Q (________28120));
  xor2s1 ____0_506480(.DIN1 (___0_9__25193), .DIN2 (_________34141), .Q
       (________28119));
  xor2s1 ____0__506481(.DIN1 (____0___25863), .DIN2 (_________34141),
       .Q (_____0__28118));
  nnd2s1 ____0_506482(.DIN1 (____0___28116), .DIN2 (___9____26879), .Q
       (____09__28117));
  or2s1 _______506483(.DIN1 (________27248), .DIN2 (____0___28111), .Q
       (____0___28115));
  and2s1 ______506484(.DIN1 (__9_9___30267), .DIN2 (________26640), .Q
       (____0___28114));
  nor2s1 _____0_506485(.DIN1 (____0___28112), .DIN2 (____0___28111), .Q
       (____0___28113));
  and2s1 _____0_506486(.DIN1 (_____0__27435), .DIN2 (____0___28109), .Q
       (____0___28110));
  and2s1 _______506487(.DIN1 (____99__28107), .DIN2 (___9____27781), .Q
       (____00__28108));
  nor2s1 _______506488(.DIN1 (______22139), .DIN2 (_____9___41202), .Q
       (____9___28106));
  nor2s1 _______506489(.DIN1 (________27323), .DIN2 (_____0__27507), .Q
       (____9___28105));
  nnd2s1 _______506490(.DIN1 (_____9__29314), .DIN2 (____9___28103), .Q
       (____9___28104));
  nnd2s1 _______506491(.DIN1 (_____9__27949), .DIN2 (_____9___31697),
       .Q (____9___28102));
  nnd2s1 _______506492(.DIN1 (____00__27392), .DIN2 (_____9__28100), .Q
       (____90__28101));
  nor2s1 ______506493(.DIN1 (____0___27484), .DIN2 (________27413), .Q
       (________28099));
  nor2s1 _______506494(.DIN1 (________27229), .DIN2 (________27587), .Q
       (________28098));
  nor2s1 _______506495(.DIN1 (________27373), .DIN2 (____0___29372), .Q
       (________28097));
  nnd2s1 _______506496(.DIN1 (____0___27399), .DIN2 (____9___29463), .Q
       (________28096));
  nor2s1 ______506497(.DIN1 (________28094), .DIN2 (____0___27655), .Q
       (________28095));
  nor2s1 _______506498(.DIN1 (________27355), .DIN2 (________27449), .Q
       (________28093));
  nnd2s1 _______506499(.DIN1 (____0___27395), .DIN2 (inData[22]), .Q
       (________28092));
  nor2s1 _______506500(.DIN1 (___0_____31198), .DIN2 (________27935),
       .Q (_____9__28091));
  or2s1 _______506501(.DIN1 (____0___26144), .DIN2 (________28089), .Q
       (________28090));
  nor2s1 ______506502(.DIN1 (__9_____30430), .DIN2 (________27271), .Q
       (________28088));
  nor2s1 _______506503(.DIN1 (____0___26506), .DIN2 (____0___29104), .Q
       (________28087));
  nor2s1 _______506504(.DIN1 (____09__26417), .DIN2 (________27332), .Q
       (________28086));
  and2s1 _______506505(.DIN1 (____9___27388), .DIN2 (________28084), .Q
       (________28085));
  nnd2s1 _______506506(.DIN1 (________28592), .DIN2 (____9___27118), .Q
       (________28083));
  nor2s1 _______506507(.DIN1 (_____9__28081), .DIN2 (____9___27385), .Q
       (_____0__28082));
  nor2s1 _______506508(.DIN1 (____9___27292), .DIN2 (__9_0___29904), .Q
       (________28080));
  nor2s1 _______506509(.DIN1 (________26459), .DIN2 (_____9__27381), .Q
       (________28079));
  nor2s1 _______506510(.DIN1 (_____0__27714), .DIN2 (________28077), .Q
       (________28078));
  nnd2s1 _______506511(.DIN1 (________27352), .DIN2 (________29501), .Q
       (________28076));
  nnd2s1 _______506512(.DIN1 (________27379), .DIN2 (________28074), .Q
       (________28075));
  nnd2s1 _______506513(.DIN1 (________27375), .DIN2 (___9____26904), .Q
       (________28073));
  and2s1 _______506514(.DIN1 (___9_0__27777), .DIN2 (_____9__29455), .Q
       (_____0__28072));
  and2s1 _______506515(.DIN1 (________28592), .DIN2 (________28070), .Q
       (_____9__28071));
  nnd2s1 ______506516(.DIN1 (_____9__27371), .DIN2 (________26562), .Q
       (________28069));
  nor2s1 _____506517(.DIN1 (___9____26018), .DIN2 (_________41186), .Q
       (________28068));
  nnd2s1 _____9_506518(.DIN1 (________28066), .DIN2 (________27999), .Q
       (________28067));
  nnd2s1 _____9_506519(.DIN1 (________27356), .DIN2 (___0____28822), .Q
       (________28065));
  nor2s1 _____506520(.DIN1 (________28063), .DIN2 (________28053), .Q
       (________28064));
  nor2s1 _____506521(.DIN1 (______0___22056), .DIN2 (________27617), .Q
       (_____0__28062));
  nnd2s1 _____0_506522(.DIN1 (_____9__29295), .DIN2 (________28060), .Q
       (_____9__28061));
  and2s1 _____0_506523(.DIN1 (________27364), .DIN2 (___0____28822), .Q
       (________28059));
  or2s1 _____0_506524(.DIN1 (________28057), .DIN2 (______0__41190), .Q
       (________28058));
  or2s1 _____0_506525(.DIN1 (_____0__25796), .DIN2 (_________41184), .Q
       (________28056));
  nor2s1 _____0_506526(.DIN1 (___0____24243), .DIN2 (____0___28016), .Q
       (________28055));
  nor2s1 ______506527(.DIN1 (________27627), .DIN2 (________28053), .Q
       (________28054));
  nnd2s1 _______506528(.DIN1 (________27412), .DIN2 (inData[12]), .Q
       (_____0__28052));
  nnd2s1 _______506529(.DIN1 (________27361), .DIN2 (________26560), .Q
       (_____9__28051));
  nor2s1 _______506530(.DIN1 (_____0__29305), .DIN2 (________27380), .Q
       (________28050));
  nnd2s1 _______506531(.DIN1 (________27348), .DIN2 (________27347), .Q
       (________28049));
  nor2s1 _______506532(.DIN1 (______________22068), .DIN2
       (________24818), .Q (________28048));
  or2s1 _______506533(.DIN1 (________28046), .DIN2 (________27331), .Q
       (________28047));
  or2s1 _______506534(.DIN1 (________28044), .DIN2 (________28043), .Q
       (________28045));
  nnd2s1 _______506535(.DIN1 (________27937), .DIN2 (___0__22157), .Q
       (_____0__28042));
  and2s1 _______506536(.DIN1 (________27407), .DIN2 (________28040), .Q
       (_____9__28041));
  nor2s1 _______506537(.DIN1 (__________0_), .DIN2 (________27071), .Q
       (________28039));
  nor2s1 _______506538(.DIN1 (_____9__28081), .DIN2 (____9___27384), .Q
       (________28038));
  nnd2s1 ______506539(.DIN1 (____0___27397), .DIN2 (_________41238), .Q
       (________28037));
  and2s1 _______506540(.DIN1 (________27321), .DIN2 (________27416), .Q
       (________28036));
  nnd2s1 _______506541(.DIN1 (________27346), .DIN2 (________28034), .Q
       (________28035));
  or2s1 ______506542(.DIN1 (_____0__28032), .DIN2 (________27319), .Q
       (________28033));
  nnd2s1 _______506543(.DIN1 (________28030), .DIN2 (________28029), .Q
       (_____9__28031));
  nnd2s1 _______506544(.DIN1 (_____0__27327), .DIN2 (_____9__27316), .Q
       (________28028));
  nor2s1 _______506545(.DIN1 (________28026), .DIN2 (___0____27896), .Q
       (________28027));
  nnd2s1 _______506546(.DIN1 (_________41192), .DIN2 (________29253),
       .Q (________28025));
  nor2s1 _______506547(.DIN1 (________27154), .DIN2 (________28060), .Q
       (________28024));
  nnd2s1 _______506548(.DIN1 (____09__28022), .DIN2 (________26607), .Q
       (_____0__28023));
  and2s1 ______506549(.DIN1 (____0___28020), .DIN2 (____0___28109), .Q
       (____0___28021));
  nnd2s1 _______506550(.DIN1 (_____9__29295), .DIN2 (___09___27914), .Q
       (____0___28019));
  nor2s1 ______506551(.DIN1 (____0___28017), .DIN2 (____0___28016), .Q
       (____0___28018));
  nor2s1 _____506552(.DIN1 (______9__37555), .DIN2 (________27403), .Q
       (____0___28015));
  nor2s1 _____9_506553(.DIN1 (____99__28013), .DIN2 (_____9__26757), .Q
       (____00__28014));
  or2s1 _____9_506554(.DIN1 (___00____30625), .DIN2 (_____0__27308), .Q
       (____9___28012));
  nor2s1 _____9_506555(.DIN1 (____9___28010), .DIN2 (________27312), .Q
       (____9___28011));
  nnd2s1 _____0_506556(.DIN1 (_____9__27410), .DIN2 (___0____26108), .Q
       (____9___28009));
  or2s1 _____0_506557(.DIN1 (________26198), .DIN2 (____9___28007), .Q
       (____9___28008));
  nnd2s1 _____0_506558(.DIN1 (_____9___41204), .DIN2 (________27440),
       .Q (____9___28006));
  and2s1 _______506559(.DIN1 (____09__29106), .DIN2 (________27350), .Q
       (____90__28005));
  or2s1 _______506560(.DIN1 (________28003), .DIN2 (___9____27755), .Q
       (_____9__28004));
  nnd2s1 _______506561(.DIN1 (________28001), .DIN2 (________27338), .Q
       (________28002));
  nnd2s1 _______506562(.DIN1 (________27999), .DIN2 (_____0__26438), .Q
       (________28000));
  nor2s1 _______506563(.DIN1 (________27239), .DIN2 (____0___29372), .Q
       (________27998));
  nor2s1 _______506564(.DIN1 (____9___26859), .DIN2 (_________41194),
       .Q (________27997));
  nor2s1 _______506565(.DIN1 (________27341), .DIN2 (____99__28013), .Q
       (________27995));
  nnd2s1 ______506566(.DIN1 (________27993), .DIN2 (____9___27389), .Q
       (________27994));
  nor2s1 _______506567(.DIN1 (________28605), .DIN2 (________27991), .Q
       (________27992));
  and2s1 _______506568(.DIN1 (________27406), .DIN2 (________27989), .Q
       (________27990));
  nor2s1 ______506569(.DIN1 (________27055), .DIN2 (_________33650), .Q
       (________27988));
  nor2s1 ______506570(.DIN1 (_____9__27986), .DIN2 (________27985), .Q
       (_____0__27987));
  nnd2s1 _______506571(.DIN1 (________27405), .DIN2 (___0____27885), .Q
       (________27984));
  or2s1 _______506572(.DIN1 (________27982), .DIN2 (___9____27799), .Q
       (________27983));
  nnd2s1 _______506573(.DIN1 (________27460), .DIN2 (inData[26]), .Q
       (________27981));
  nnd2s1 _______506574(.DIN1 (________27151), .DIN2 (_____0__27139), .Q
       (________27980));
  nnd2s1 _______506575(.DIN1 (_____0__27978), .DIN2 (____9___26585), .Q
       (________27979));
  and2s1 ______506576(.DIN1 (________27972), .DIN2 (________29246), .Q
       (_____9__27977));
  nnd2s1 _______506577(.DIN1 (________27424), .DIN2 (________27975), .Q
       (________27976));
  nor2s1 _______506578(.DIN1 (________27469), .DIN2 (________29119), .Q
       (________27974));
  nnd2s1 ______506579(.DIN1 (________27972), .DIN2 (____09__27489), .Q
       (________27973));
  nor2s1 _______506580(.DIN1 (________27970), .DIN2 (________27281), .Q
       (________27971));
  nnd2s1 _______506581(.DIN1 (__________0_), .DIN2
       (______________22103), .Q (________27969));
  nnd2s1 _______506582(.DIN1 (________27357), .DIN2 (_____9__27967), .Q
       (_____0__27968));
  nnd2s1 _______506583(.DIN1 (________27438), .DIN2 (_____90__33327),
       .Q (________27966));
  nnd2s1 _______506584(.DIN1 (________27945), .DIN2 (________27964), .Q
       (________27965));
  or2s1 _______506585(.DIN1 (________27264), .DIN2 (________27962), .Q
       (________27963));
  nnd2s1 _______506586(.DIN1 (________27535), .DIN2 (________27960), .Q
       (________27961));
  nor2s1 _____506587(.DIN1 (____9___26322), .DIN2 (________27955), .Q
       (________27959));
  nor2s1 _____0_506588(.DIN1 (________27277), .DIN2 (____0___28380), .Q
       (_____0__27958));
  nor2s1 _____0_506589(.DIN1 (________27956), .DIN2 (________27955), .Q
       (_____9__27957));
  nnd2s1 _____506590(.DIN1 (________27253), .DIN2 (_________31879), .Q
       (________27953));
  nor2s1 _____9_506591(.DIN1 (________26631), .DIN2 (__9_____29745), .Q
       (________27952));
  and2s1 _____9_506592(.DIN1 (_____9__27949), .DIN2 (________27532), .Q
       (_____0__27950));
  nor2s1 _____9_506593(.DIN1 (________27273), .DIN2 (________27153), .Q
       (________27948));
  nnd2s1 _____9_506594(.DIN1 (____9___27387), .DIN2 (____0___27398), .Q
       (________27947));
  nnd2s1 _____506595(.DIN1 (________27945), .DIN2 (___9_0__28655), .Q
       (________27946));
  hi1s1 _______506596(.DIN (_____0__28395), .Q (________27944));
  hi1s1 _______506597(.DIN (___0_____40156), .Q (________27943));
  nor2s1 _______506598(.DIN1 (________29088), .DIN2 (_____0__27941), .Q
       (________27942));
  nor2s1 ______506599(.DIN1 (________27939), .DIN2 (________27254), .Q
       (_____9__27940));
  nnd2s1 _______506600(.DIN1 (________27937), .DIN2 (inData[10]), .Q
       (________27938));
  nnd2s1 _______506601(.DIN1 (________27459), .DIN2 (________27493), .Q
       (________27936));
  nor2s1 _______506602(.DIN1 (_________31655), .DIN2 (____0___29104),
       .Q (________27934));
  or2s1 _______506603(.DIN1 (_____0__27932), .DIN2 (____9___27206), .Q
       (________27933));
  nor2s1 _______506604(.DIN1 (____0___28202), .DIN2 (________27592), .Q
       (____09__27931));
  nor2s1 ______506605(.DIN1 (________28485), .DIN2 (_____9__27240), .Q
       (____0___27930));
  or2s1 _______506606(.DIN1 (___0____22328), .DIN2 (____0___28016), .Q
       (____0___27929));
  nnd2s1 _______506607(.DIN1 (______________22068), .DIN2
       (_________32611), .Q (____0___27928));
  nnd2s1 ______506608(.DIN1 (________27589), .DIN2 (_____9__27434), .Q
       (____0___27927));
  nor2s1 _______506609(.DIN1 (________29173), .DIN2 (________27368), .Q
       (________28300));
  hi1s1 _______506610(.DIN (_____0__28306), .Q (________28845));
  xor2s1 ____00_506611(.DIN1 (________22371), .DIN2 (_________38155),
       .Q (________28420));
  nnd2s1 ____00_506612(.DIN1 (________27456), .DIN2 (____0___27926), .Q
       (____09__28843));
  or2s1 ______506613(.DIN1 (___0_____31191), .DIN2 (________27334), .Q
       (_____9__28570));
  nnd2s1 _______506614(.DIN1 (___0_____30771), .DIN2 (________25563),
       .Q (___00___28737));
  or2s1 _______506615(.DIN1 (_____9__26838), .DIN2 (____9_0__33415), .Q
       (___9_9__28727));
  or2s1 _______506616(.DIN1 (____0___27925), .DIN2 (____09__27307), .Q
       (___9____28668));
  nor2s1 _______506617(.DIN1 (________27433), .DIN2 (__9_____29881), .Q
       (___9____28670));
  nnd2s1 _______506618(.DIN1 (____0___27304), .DIN2 (___00___27828), .Q
       (___0____28757));
  nor2s1 ______506619(.DIN1 (____0___27924), .DIN2 (________27607), .Q
       (____00__28376));
  nor2s1 _______506620(.DIN1 (_________32058), .DIN2 (________27258),
       .Q (____9___28375));
  nnd2s1 _______506621(.DIN1
       (_____________________________________________21896), .DIN2
       (____0___27923), .Q (_____9__28972));
  nnd2s1 _______506622(.DIN1 (____00__27654), .DIN2 (________29331), .Q
       (____9___28373));
  and2s1 _______506623(.DIN1 (____9___27390), .DIN2 (________28230), .Q
       (___0____28817));
  nor2s1 ______506624(.DIN1 (___090___31413), .DIN2 (________27470), .Q
       (____9___28644));
  nnd2s1 _______506625(.DIN1 (________27606), .DIN2 (____00__27922), .Q
       (_____9__29386));
  nor2s1 _______506626(.DIN1 (__9_0___29724), .DIN2 (_____0__27336), .Q
       (___99___28732));
  and2s1 ______506627(.DIN1 (____0____31579), .DIN2 (________27267), .Q
       (___9____28709));
  nor2s1 _______506628(.DIN1 (___9____27771), .DIN2 (________27414), .Q
       (___0____28797));
  nor2s1 ______506629(.DIN1 (___099__27921), .DIN2 (________27337), .Q
       (____9___28372));
  nnd2s1 _______506630(.DIN1 (________27262), .DIN2 (___09___27920), .Q
       (___990__28728));
  nnd2s1 _______506631(.DIN1 (________27343), .DIN2 (_____9___31891),
       .Q (___9____29573));
  nor2s1 ______506632(.DIN1 (___09___27919), .DIN2 (___09___27918), .Q
       (_________33032));
  nor2s1 _______506633(.DIN1 (___09___27917), .DIN2 (________27431), .Q
       (___09____31438));
  nnd2s1 _____9_506634(.DIN1 (________28066), .DIN2 (________26752), .Q
       (__9__9__30444));
  nor2s1 _______506635(.DIN1 (___09___27916), .DIN2 (____0___29104), .Q
       (_________32344));
  or2s1 _____9_506636(.DIN1 (___09___27915), .DIN2 (___09___27914), .Q
       (_____9___33997));
  xor2s1 _______506637(.DIN1 (________27144), .DIN2 (________22537), .Q
       (_____0___36015));
  hi1s1 ____506638(.DIN (______0__35537), .Q (___9____28662));
  dffacs1 ________________________________________________506639(.CLRB
       (reset), .CLK (clk), .DIN (________27342), .Q
       (__________________________________________________________________21990));
  nor2s1 _____0_506640(.DIN1 (________28600), .DIN2 (__9_9___29892), .Q
       (______0__32108));
  nnd2s1 _____506641(.DIN1 (________27993), .DIN2 (________29431), .Q
       (_________34163));
  dffacs1 _______________________________________________506642(.CLRB
       (reset), .CLK (clk), .DIN (_____0__27354), .Q
       (_____________________________________________21926));
  hi1s1 ____09_506643(.DIN (___9_____39219), .Q (___0_____40115));
  dffacs1 ______________________________________________0_506644(.CLRB
       (reset), .CLK (clk), .DIN (________27360), .Q (___0_____40433));
  nnd2s1 ______506645(.DIN1 (___090__27912), .DIN2 (___09___27913), .Q
       (__90_9__29717));
  nnd2s1 _______506646(.DIN1 (___0____27910), .DIN2 (inData[21]), .Q
       (___0_____30961));
  nor2s1 _______506647(.DIN1 (inData[21]), .DIN2 (___090__27912), .Q
       (___9____28692));
  nor2s1 _______506648(.DIN1 (___0_9__27911), .DIN2 (___0____27910), .Q
       (___0____28783));
  nor2s1 _____9_506649(.DIN1 (________27238), .DIN2 (__9_____29827), .Q
       (___0____27909));
  nor2s1 _____0_506650(.DIN1 (____0___26783), .DIN2 (________29119), .Q
       (___0____27908));
  or2s1 _____0_506651(.DIN1 (___9____27797), .DIN2 (___0____27906), .Q
       (___0____27907));
  nnd2s1 ______506652(.DIN1 (________27272), .DIN2 (____9___29007), .Q
       (___0____27905));
  nnd2s1 _______506653(.DIN1 (________27467), .DIN2 (____0____31517),
       .Q (___0____27904));
  nnd2s1 _______506654(.DIN1 (________28585), .DIN2 (__9_____29873), .Q
       (___0____27903));
  nnd2s1 _______506655(.DIN1 (________28592), .DIN2 (___0_____31274),
       .Q (___0_9__27902));
  nnd2s1 _______506656(.DIN1 (________27993), .DIN2 (_________32305),
       .Q (___0____27901));
  or2s1 _______506657(.DIN1 (________29529), .DIN2 (_____9__27462), .Q
       (___0____27900));
  nnd2s1 ______506658(.DIN1 (________27268), .DIN2 (___0_____31151), .Q
       (___0____27899));
  or2s1 ______506659(.DIN1 (___0____27897), .DIN2 (___0____27896), .Q
       (___0____27898));
  nnd2s1 _______506660(.DIN1 (___0____27843), .DIN2 (________27068), .Q
       (___0____27895));
  nor2s1 _______506661(.DIN1 (____9___26678), .DIN2 (____0___29104), .Q
       (___0_0__27894));
  and2s1 _______506662(.DIN1 (___0____27892), .DIN2 (_____0__29213), .Q
       (___0_9__27893));
  nnd2s1 _______506663(.DIN1 (________28592), .DIN2 (____0___28479), .Q
       (___0____27891));
  nnd2s1 ______506664(.DIN1 (________27237), .DIN2 (___0____27889), .Q
       (___0____27890));
  nnd2s1 ______506665(.DIN1 (________27993), .DIN2 (________26726), .Q
       (___0____27888));
  nor2s1 _______506666(.DIN1 (____9___26495), .DIN2 (____0___29104), .Q
       (___0____27887));
  nnd2s1 ______506667(.DIN1 (___0____27885), .DIN2 (____9___27386), .Q
       (___0____27886));
  nnd2s1 ______506668(.DIN1 (_________41188), .DIN2 (___09___28825), .Q
       (___0_0__27884));
  nor2s1 _______506669(.DIN1 (________27664), .DIN2 (________27351), .Q
       (___0_9__27883));
  or2s1 _______506670(.DIN1 (______0__31950), .DIN2 (_____9__27250), .Q
       (___0____27882));
  and2s1 _______506671(.DIN1 (________28592), .DIN2 (___0_____30695),
       .Q (___0____27881));
  nor2s1 ______506672(.DIN1 (___0____27878), .DIN2 (_____90__41200), .Q
       (___0____27879));
  hi1s1 _______506673(.DIN (___0____27876), .Q (___0____27877));
  nor2s1 _______506674(.DIN1 (__9_0___29724), .DIN2 (________27263), .Q
       (___0_0__27875));
  or2s1 ______506675(.DIN1 (___0____27873), .DIN2 (_____0__27216), .Q
       (___0_9__27874));
  or2s1 ______506676(.DIN1 (________28046), .DIN2 (_____0__27196), .Q
       (___0____27872));
  nnd2s1 _______506677(.DIN1 (____9___27205), .DIN2 (___0____27870), .Q
       (___0____27871));
  nnd2s1 _______506678(.DIN1 (_____9__29295), .DIN2 (___0____27868), .Q
       (___0____27869));
  nnd2s1 _______506679(.DIN1 (________29361), .DIN2 (______0__41250),
       .Q (___0____27867));
  and2s1 _____0_506680(.DIN1 (__90____29661), .DIN2 (________29142), .Q
       (___0____27866));
  nor2s1 _____0_506681(.DIN1 (___09___25216), .DIN2 (________27188), .Q
       (___0_0__27865));
  nnd2s1 _____9_506682(.DIN1 (_____9__29295), .DIN2 (___0____27863), .Q
       (___0_9__27864));
  nor2s1 _____9_506683(.DIN1 (_____0__28481), .DIN2 (___0_0__27855), .Q
       (___0____27862));
  nnd2s1 _____9_506684(.DIN1 (__9990), .DIN2 (___0____27860), .Q
       (___0____27861));
  nnd2s1 _____506685(.DIN1 (____9___27476), .DIN2 (___0____27858), .Q
       (___0____27859));
  nor2s1 _______506686(.DIN1 (________27638), .DIN2 (____0___27211), .Q
       (___0____27857));
  nor2s1 ______506687(.DIN1 (____09___31598), .DIN2 (___0_0__27855), .Q
       (___0____27856));
  and2s1 _______506688(.DIN1 (___0____27892), .DIN2 (___0____27853), .Q
       (___0_9__27854));
  and2s1 _______506689(.DIN1 (________27151), .DIN2 (___0____27851), .Q
       (___0____27852));
  nor2s1 _______506690(.DIN1 (________27225), .DIN2 (___0____27849), .Q
       (___0____27850));
  or2s1 _______506691(.DIN1 (___0____27847), .DIN2 (________27991), .Q
       (___0____27848));
  nor2s1 ______506692(.DIN1 (____0___27213), .DIN2 (___0_0__27855), .Q
       (___0____27846));
  and2s1 _______506693(.DIN1 (________28320), .DIN2 (_____0__26728), .Q
       (___0_0__27845));
  nnd2s1 _______506694(.DIN1 (___0____27843), .DIN2 (___0____27842), .Q
       (___0_9__27844));
  nor2s1 _______506695(.DIN1 (________28628), .DIN2 (__9_____29827), .Q
       (___0____27841));
  nnd2s1 _______506696(.DIN1 (________29537), .DIN2 (_____0__28148), .Q
       (___0____27840));
  or2s1 _______506697(.DIN1 (___0_____31078), .DIN2 (___0_0__27855), .Q
       (___0____27839));
  nnd2s1 _____506698(.DIN1 (__9_____30019), .DIN2 (________28160), .Q
       (___0____27838));
  nor2s1 ______506699(.DIN1 (___9____27792), .DIN2 (__9_____29783), .Q
       (___0____27837));
  nor2s1 _______506700(.DIN1 (________29409), .DIN2 (___009__27835), .Q
       (___0_0__27836));
  nor2s1 _______506701(.DIN1 (________24880), .DIN2 (________27189), .Q
       (___00___27834));
  nor2s1 _______506702(.DIN1 (____0___27926), .DIN2 (___0_0__27855), .Q
       (___00___27833));
  nnd2s1 ______506703(.DIN1 (________29537), .DIN2 (________27547), .Q
       (___00___27832));
  and2s1 _______506704(.DIN1 (________29537), .DIN2 (__909___29719), .Q
       (___00___27831));
  nor2s1 _______506705(.DIN1 (________28305), .DIN2 (________27149), .Q
       (___00___27830));
  and2s1 _______506706(.DIN1 (________27193), .DIN2 (___00___27828), .Q
       (___00___27829));
  hi1s1 ______506707(.DIN (___00____30606), .Q (___00___27827));
  and2s1 ____0__506708(.DIN1 (________29361), .DIN2 (________27074), .Q
       (___99___27825));
  hi1s1 _____506709(.DIN (____0___28201), .Q (___990__27822));
  nor2s1 ____0__506710(.DIN1 (___9____27820), .DIN2 (________27184), .Q
       (___9_9__27821));
  hi1s1 _____0_506711(.DIN (___0_____40439), .Q (___9____27819));
  or2s1 ____0__506712(.DIN1 (________26548), .DIN2 (___9_9__27785), .Q
       (___9____27818));
  nor2s1 ____0__506713(.DIN1 (________27511), .DIN2 (________27200), .Q
       (___9____27817));
  nor2s1 ____0__506714(.DIN1 (________26212), .DIN2 (________27151), .Q
       (___9____27816));
  nnd2s1 ____9__506715(.DIN1 (________29361), .DIN2 (________27073), .Q
       (___9____27815));
  and2s1 ____9__506716(.DIN1 (___9____28696), .DIN2 (___9____25972), .Q
       (___9____27814));
  nnd2s1 ____9__506717(.DIN1 (________27191), .DIN2 (___0____26061), .Q
       (___9____27812));
  nnd2s1 ____90_506718(.DIN1 (________27501), .DIN2 (________28484), .Q
       (___9____27811));
  or2s1 _____9_506719(.DIN1 (________27939), .DIN2 (___9____27765), .Q
       (___9____27810));
  nnd2s1 _______506720(.DIN1 (__9_9___30270), .DIN2 (________26606), .Q
       (___9____27808));
  and2s1 _______506721(.DIN1 (___9____27806), .DIN2 (___9_0__27805), .Q
       (___9____27807));
  and2s1 _______506722(.DIN1 (_____9__29295), .DIN2 (___9____27803), .Q
       (___9_9__27804));
  nor2s1 _______506723(.DIN1 (____0___26597), .DIN2 (____9___29093), .Q
       (____9___28288));
  nor2s1 _____0_506724(.DIN1 (___9____27801), .DIN2 (___9____27802), .Q
       (________28852));
  nor2s1 ______506725(.DIN1 (___9____27801), .DIN2 (________27224), .Q
       (________28597));
  nnd2s1 ______506726(.DIN1 (____9___27473), .DIN2 (________29311), .Q
       (___00___28741));
  nor2s1 _______506727(.DIN1 (___9____27800), .DIN2 (___9____27799), .Q
       (________28613));
  or2s1 _______506728(.DIN1 (___9____27798), .DIN2 (___9____27797), .Q
       (________28625));
  or2s1 _______506729(.DIN1 (_____0___34102), .DIN2 (________27234), .Q
       (___9____28712));
  and2s1 _______506730(.DIN1 (________27584), .DIN2 (___9____27796), .Q
       (___9____28719));
  nnd2s1 ______506731(.DIN1 (________27349), .DIN2 (___9_0__27795), .Q
       (___9____28702));
  dffacs1 _________________________________________0____506732(.CLRB
       (reset), .CLK (clk), .DIN (________27376), .QN
       (_____________________________________0____));
  hi1s1 _____0_506733(.DIN (___9_9__27794), .Q (________28509));
  nnd2s1 ____0__506734(.DIN1 (________29361), .DIN2 (___9____27793), .Q
       (___0____28761));
  nnd2s1 ____0__506735(.DIN1 (___9____27806), .DIN2 (________28444), .Q
       (_____0__28168));
  nor2s1 ____0_506736(.DIN1 (___0_0___30746), .DIN2 (________27187), .Q
       (________29242));
  nnd2s1 ____0__506737(.DIN1 (___9____27792), .DIN2 (________27718), .Q
       (____0___28473));
  and2s1 ____506738(.DIN1 (___9____27791), .DIN2 (_____9___31694), .Q
       (________28483));
  nor2s1 ____09_506739(.DIN1 (___9_9__26939), .DIN2 (________29264), .Q
       (________28169));
  nnd2s1 ____09_506740(.DIN1 (____9___27207), .DIN2 (___0_____30789),
       .Q (____0___28478));
  nor2s1 _____0_506741(.DIN1 (________29229), .DIN2 (__9_____30260), .Q
       (________28528));
  nor2s1 _____0_506742(.DIN1 (________27194), .DIN2 (___0____26964), .Q
       (____9___28470));
  or2s1 _______506743(.DIN1 (___9____27790), .DIN2 (________27198), .Q
       (________28525));
  nnd2s1 _______506744(.DIN1 (____0___27485), .DIN2 (________29428), .Q
       (________28156));
  nnd2s1 _____506745(.DIN1 (__90____29661), .DIN2 (________29359), .Q
       (_____9__28157));
  nor2s1 _____0_506746(.DIN1 (___9____27789), .DIN2 (___9____27788), .Q
       (_____0__28158));
  nnd2s1 _______506747(.DIN1 (___9____27787), .DIN2 (________26723), .Q
       (________28179));
  nor2s1 _______506748(.DIN1 (___9_0__27786), .DIN2 (________27219), .Q
       (________28177));
  nor2s1 _______506749(.DIN1 (________27175), .DIN2 (___9_9__27785), .Q
       (________28176));
  nor2s1 _______506750(.DIN1 (_________41273), .DIN2 (________27218),
       .Q (____0___28475));
  nnd2s1 _______506751(.DIN1 (________28320), .DIN2 (________28261), .Q
       (________28175));
  nnd2s1 ______506752(.DIN1 (____09__29106), .DIN2 (__9_____29766), .Q
       (____0___28477));
  hi1s1 _______506753(.DIN (________28268), .Q (__9__0__30216));
  and2s1 _______506754(.DIN1 (__9990), .DIN2 (________29319), .Q
       (____0___28476));
  nor2s1 _______506755(.DIN1 (________26842), .DIN2 (___9____27788), .Q
       (__9_____29748));
  xnr2s1 ______506756(.DIN1 (______0__35711), .DIN2 (___0____26988), .Q
       (________28578));
  nnd2s1 _______506757(.DIN1 (____0___27486), .DIN2 (___9____27784), .Q
       (________28534));
  or2s1 _______506758(.DIN1 (___9____27783), .DIN2 (________29508), .Q
       (___0_9__28765));
  nnd2s1 _______506759(.DIN1 (________27960), .DIN2 (________25730), .Q
       (________28164));
  nnd2s1 _______506760(.DIN1 (________27366), .DIN2 (___9____27782), .Q
       (________28587));
  nor2s1 _______506761(.DIN1 (______________22068), .DIN2
       (_____9___38610), .Q (________28165));
  nnd2s1 _______506762(.DIN1 (___9____27781), .DIN2 (____0___29010), .Q
       (____0___28292));
  nnd2s1 ______506763(.DIN1 (___9____27779), .DIN2 (________29498), .Q
       (____00__28291));
  nnd2s1 _______506764(.DIN1 (________27146), .DIN2 (_____0__28608), .Q
       (________28166));
  nor2s1 _____506765(.DIN1 (___9_9__26919), .DIN2 (___9____27780), .Q
       (____0___28297));
  nnd2s1 _______506766(.DIN1 (___9____27779), .DIN2 (___9____27778), .Q
       (________28610));
  nor2s1 _______506767(.DIN1 (_____9___41301), .DIN2 (________27257),
       .Q (____90__28285));
  and2s1 _______506768(.DIN1 (___9_0__27777), .DIN2 (___0_0__26960), .Q
       (___0____28790));
  nnd2s1 ______506769(.DIN1 (________27232), .DIN2 (________25745), .Q
       (____9___28469));
  nor2s1 _______506770(.DIN1 (____0___22451), .DIN2 (_________33650),
       .Q (____9___28286));
  nnd2s1 ______506771(.DIN1 (___0____23297), .DIN2
       (______________22068), .Q (________28891));
  nor2s1 _______506772(.DIN1 (___9_9__27776), .DIN2 (_________41182),
       .Q (________28634));
  nnd2s1 _______506773(.DIN1 (_____0__27241), .DIN2 (___0_____31173),
       .Q (___9____28705));
  nnd2s1 _______506774(.DIN1 (___0_____30771), .DIN2 (________26751),
       .Q (___9____28679));
  nor2s1 _______506775(.DIN1 (___099__27921), .DIN2 (________27255), .Q
       (________28602));
  nor2s1 _______506776(.DIN1 (________27041), .DIN2 (___09____31480),
       .Q (____9___28289));
  nnd2s1 _______506777(.DIN1 (________27340), .DIN2 (___0_____31362),
       .Q (________28486));
  nor2s1 _______506778(.DIN1 (___0_9__25174), .DIN2 (___9____27775), .Q
       (____9___28290));
  or2s1 _____0_506779(.DIN1 (____9___28010), .DIN2 (_____0__27585), .Q
       (________28631));
  or2s1 _____0_506780(.DIN1 (___9____27774), .DIN2 (________27244), .Q
       (_____0__28591));
  nnd2s1 _____9_506781(.DIN1 (________27245), .DIN2 (___9____27773), .Q
       (___9____28667));
  nor2s1 _______506782(.DIN1 (____9___23592), .DIN2 (________27422), .Q
       (_________36713));
  nnd2s1 _______506783(.DIN1 (__9_____29845), .DIN2 (________27975), .Q
       (________28857));
  nor2s1 _______506784(.DIN1 (___9____27772), .DIN2 (________27420), .Q
       (____0____31556));
  or2s1 _______506785(.DIN1 (____0____31545), .DIN2 (________27430), .Q
       (___0_____31223));
  or2s1 _______506786(.DIN1 (___9____27771), .DIN2 (________27461), .Q
       (_________32836));
  nor2s1 _______506787(.DIN1 (___099__27921), .DIN2 (________27428), .Q
       (___9____28716));
  hi1s1 ______506788(.DIN (___0_____40100), .Q (________28513));
  hi1s1 _______506789(.DIN (__9_0___29729), .Q (____0___28558));
  nor2s1 _______506790(.DIN1 (___9____27781), .DIN2 (__9__9__29935), .Q
       (_________33002));
  hi1s1 ______506791(.DIN (___9____27770), .Q (________28987));
  and2s1 _______506792(.DIN1 (_____9___41204), .DIN2 (___9____25976),
       .Q (__9_____30306));
  nnd2s1 _______506793(.DIN1 (__9__0__30196), .DIN2 (___9____26918), .Q
       (__9__9__30073));
  and2s1 _______506794(.DIN1 (___9____27769), .DIN2 (________29384), .Q
       (_____0__28538));
  nor2s1 _______506795(.DIN1 (______9__32852), .DIN2 (___009__27835),
       .Q (____9___28642));
  or2s1 _______506796(.DIN1 (___0____28793), .DIN2 (________27149), .Q
       (_____9___32968));
  nor2s1 _____0_506797(.DIN1 (___9_0__27768), .DIN2 (___0_0__27855), .Q
       (_________32854));
  nnd2s1 _____0_506798(.DIN1 (__9990), .DIN2 (___099___31496), .Q
       (___09____31472));
  nnd2s1 _____0_506799(.DIN1 (____0___27212), .DIN2 (________26426), .Q
       (___0_09__30651));
  nnd2s1 _______506800(.DIN1 (________29537), .DIN2 (___9_9__27767), .Q
       (_________33096));
  nnd2s1 _____0_506801(.DIN1 (__9_9___30270), .DIN2 (___90___26867), .Q
       (________28482));
  nor2s1 ______506802(.DIN1 (___9____27766), .DIN2 (___0_0__27855), .Q
       (_________33143));
  nor2s1 _______506803(.DIN1 (____0____31547), .DIN2 (___9____27765),
       .Q (____9___28551));
  and2s1 _______506804(.DIN1 (___0____27847), .DIN2 (________28034), .Q
       (________29525));
  or2s1 _______506805(.DIN1 (___9____27764), .DIN2 (___0_0__27855), .Q
       (_________34531));
  or2s1 _______506806(.DIN1 (_____0__26518), .DIN2 (___0_0__27855), .Q
       (______9__33037));
  nnd2s1 _______506807(.DIN1 (____09__28480), .DIN2 (____0___27209), .Q
       (__9__9__30337));
  and2s1 _______506808(.DIN1 (__9_____30423), .DIN2 (______0__32214),
       .Q (______0__33008));
  ib1s1 _______506809(.DIN
       (__________________________________9__________), .Q
       (________27618));
  nor2s1 _______506810(.DIN1 (___0_____31381), .DIN2 (________27227),
       .Q (___0_____31204));
  and2s1 _______506811(.DIN1 (____09__28022), .DIN2 (___9____27763), .Q
       (___0_99__30832));
  hi1s1 _______506812(.DIN (______9__32753), .Q (_____90__32273));
  dffacs1 ________________________________________________506813(.CLRB
       (reset), .CLK (clk), .DIN (________27370), .Q
       (______________________________________________21905));
  dffacs1 _________________________________________0_____506814(.CLRB
       (reset), .CLK (clk), .DIN (________27404), .Q (___0_____40575));
  hi1s1 _______506815(.DIN
       (__________________________________9__________), .Q
       (________27612));
  dffacs1 ________________________________________________506816(.CLRB
       (reset), .CLK (clk), .DIN (________27276), .Q
       (__________________________________________________________________21985));
  hi1s1 _______506817(.DIN
       (__________________________________9__________), .Q
       (_________41367));
  nnd2s1 ______506818(.DIN1 (________29361), .DIN2 (___9____27762), .Q
       (_________33128));
  dffacs1 ______________________________________________0_506819(.CLRB
       (reset), .CLK (clk), .DIN (________27359), .QN
       (__________________________________________0___21935));
  dffacs1 ________________________________________________506820(.CLRB
       (reset), .CLK (clk), .DIN (________27330), .Q
       (______________________________________________21930));
  nor2s1 _______506821(.DIN1 (___0____25171), .DIN2 (________27437), .Q
       (______0__36598));
  hi1s1 _______506822(.DIN (______0__32253), .Q (_________32266));
  nor2s1 _____9_506823(.DIN1 (________23082), .DIN2 (________27182), .Q
       (_____0___35741));
  xnr2s1 _____9_506824(.DIN1
       (______________________________________________21958), .DIN2
       (_________38869), .Q (___9_9__27761));
  and2s1 ____00_506825(.DIN1 (____90__27647), .DIN2 (___0____26995), .Q
       (___9____27760));
  xor2s1 ____0__506826(.DIN1 (___9____27758), .DIN2 (___9____26874), .Q
       (___9____27759));
  xnr2s1 ____0__506827(.DIN1
       (_____________________________________________21799), .DIN2
       (___9__9__39731), .Q (___9____27757));
  or2s1 ______506828(.DIN1 (___9____27755), .DIN2 (___9____27754), .Q
       (___9____27756));
  nor2s1 _______506829(.DIN1 (_____0__23368), .DIN2 (_____0__27047), .Q
       (___9____27753));
  nor2s1 _______506830(.DIN1 (________22665), .DIN2 (__99____30514), .Q
       (___9_0__27752));
  and2s1 _______506831(.DIN1 (________27059), .DIN2 (________27602), .Q
       (___909__27751));
  nor2s1 _______506832(.DIN1 (____09__27128), .DIN2 (________27130), .Q
       (___90___27750));
  nor2s1 _______506833(.DIN1 (____9___27383), .DIN2 (___0____28820), .Q
       (___90___27749));
  nnd2s1 _______506834(.DIN1 (_____0__27129), .DIN2 (________28454), .Q
       (___90___27748));
  nnd2s1 _______506835(.DIN1 (____0___27124), .DIN2 (________25844), .Q
       (___90___27747));
  and2s1 ______506836(.DIN1 (____9___27120), .DIN2 (________27365), .Q
       (___90___27746));
  nnd2s1 _______506837(.DIN1 (____0___27125), .DIN2 (________25793), .Q
       (___90___27745));
  nnd2s1 _____9_506838(.DIN1 (____9___29551), .DIN2 (________26790), .Q
       (___90___27744));
  nnd2s1 _____506839(.DIN1 (__9_9___30174), .DIN2 (____0___28112), .Q
       (___90___27743));
  nnd2s1 _______506840(.DIN1 (____99__27741), .DIN2 (________27064), .Q
       (___900__27742));
  nnd2s1 _______506841(.DIN1 (________27045), .DIN2 (______9__35683),
       .Q (____9___27740));
  nnd2s1 _______506842(.DIN1 (___0_____30888), .DIN2 (________26624),
       .Q (____9___27739));
  nor2s1 _______506843(.DIN1 (____9___27115), .DIN2 (__9__9__29935), .Q
       (____9___27738));
  and2s1 _______506844(.DIN1 (_________34141), .DIN2 (________), .Q
       (____9___27737));
  nnd2s1 ______506845(.DIN1 (________27109), .DIN2 (____9___27649), .Q
       (____9___27736));
  nnd2s1 _______506846(.DIN1 (___0_____30805), .DIN2 (_____9__27636),
       .Q (____9___27735));
  nnd2s1 _______506847(.DIN1 (____0_0__37159), .DIN2 (________27133),
       .Q (____9___27734));
  nnd2s1 _______506848(.DIN1 (_________31778), .DIN2 (________27107),
       .Q (____9___27733));
  or2s1 _______506849(.DIN1 (________), .DIN2 (_________34141), .Q
       (____90__27732));
  or2s1 _______506850(.DIN1 (____0_0__32557), .DIN2 (________27106), .Q
       (_____9__27731));
  nnd2s1 _____9_506851(.DIN1 (___9____26908), .DIN2 (___0_____40515),
       .Q (________27730));
  nor2s1 _____506852(.DIN1 (________27065), .DIN2 (__90_9__29708), .Q
       (________27729));
  nor2s1 _____0_506853(.DIN1 (___0_____40515), .DIN2 (___9____26908),
       .Q (________27728));
  and2s1 _____0_506854(.DIN1 (________27726), .DIN2 (________27707), .Q
       (________27727));
  nor2s1 ____00_506855(.DIN1 (________27724), .DIN2 (_____0__27723), .Q
       (________27725));
  or2s1 ____99_506856(.DIN1 (________27721), .DIN2 (________27720), .Q
       (_____9__27722));
  and2s1 ____9__506857(.DIN1 (________28154), .DIN2 (________27718), .Q
       (________27719));
  nor2s1 ____9__506858(.DIN1 (____9___26316), .DIN2 (____0___27032), .Q
       (________27717));
  nor2s1 ____9_506859(.DIN1 (________27715), .DIN2 (_____0__27714), .Q
       (________27716));
  nnd2s1 ____9__506860(.DIN1 (________27712), .DIN2 (________27711), .Q
       (_____9__27713));
  and2s1 ____9__506861(.DIN1 (_____0__27085), .DIN2 (________27709), .Q
       (________27710));
  or2s1 ______506862(.DIN1 (________27962), .DIN2 (________27703), .Q
       (_____0__27706));
  nor2s1 ______506863(.DIN1 (________27704), .DIN2 (________27703), .Q
       (_____9__27705));
  nnd2s1 ______506864(.DIN1 (_________33931), .DIN2 (________27701), .Q
       (________27702));
  nor2s1 _____0_506865(.DIN1 (_____0__26211), .DIN2 (_________38650),
       .Q (________27700));
  and2s1 _____0_506866(.DIN1 (________26719), .DIN2 (_________38650),
       .Q (________27699));
  nor2s1 _____0_506867(.DIN1 (_____9__25900), .DIN2 (_____0___41216),
       .Q (________27698));
  nor2s1 _______506868(.DIN1 (___0____27889), .DIN2 (__9_____29862), .Q
       (________27697));
  nnd2s1 _______506869(.DIN1 (________27140), .DIN2 (____90__27382), .Q
       (_____0__27696));
  nnd2s1 ______506870(.DIN1 (________27048), .DIN2 (________27694), .Q
       (_____9__27695));
  nor2s1 ______506871(.DIN1 (___00___26955), .DIN2 (_____9__27222), .Q
       (________27693));
  nor2s1 _______506872(.DIN1 (________28171), .DIN2 (________28225), .Q
       (________27692));
  and2s1 _______506873(.DIN1 (__9_____30322), .DIN2 (________27690), .Q
       (________27691));
  nnd2s1 _______506874(.DIN1 (___0_____30805), .DIN2 (________26653),
       .Q (________27689));
  or2s1 _______506875(.DIN1 (_____0__27687), .DIN2 (____0___29372), .Q
       (________27688));
  nor2s1 ______506876(.DIN1 (____9___26862), .DIN2 (____0___29372), .Q
       (_____9__27686));
  nor2s1 _______506877(.DIN1 (________22520), .DIN2 (________27604), .Q
       (________27685));
  or2s1 _____0_506878(.DIN1 (___0____26971), .DIN2 (________27704), .Q
       (________27684));
  nor2s1 _____506879(.DIN1 (____09__26507), .DIN2 (________27704), .Q
       (________27683));
  nor2s1 _______506880(.DIN1 (____0___29374), .DIN2 (________27681), .Q
       (________27682));
  and2s1 _______506881(.DIN1 (____0___27034), .DIN2 (________28034), .Q
       (________27680));
  nor2s1 _______506882(.DIN1 (________27681), .DIN2 (________27069), .Q
       (________27679));
  nor2s1 _______506883(.DIN1 (________27221), .DIN2 (_____0__27057), .Q
       (________27678));
  nor2s1 _______506884(.DIN1 (________29066), .DIN2 (____0___29372), .Q
       (_____0__27677));
  xor2s1 _______506885(.DIN1
       (_____________________________________________21783), .DIN2
       (______0__34517), .Q (_____9__27676));
  or2s1 ____9_506886(.DIN1 (________27101), .DIN2 (________27674), .Q
       (________27675));
  xor2s1 _______506887(.DIN1
       (__________________________________________), .DIN2
       (___9_0___39709), .Q (________27673));
  xor2s1 _______506888(.DIN1 (____0___22553), .DIN2 (_________41252),
       .Q (________27672));
  nor2s1 ____9__506889(.DIN1 (_____9___41301), .DIN2 (________27670),
       .Q (________27671));
  xor2s1 _____9_506890(.DIN1
       (_____________________________________________21924), .DIN2
       (____9____38007), .Q (________27669));
  xor2s1 _____506891(.DIN1 (___9_____39511), .DIN2 (_____9___36360), .Q
       (________27668));
  and2s1 ____9_506892(.DIN1 (_____0__27093), .DIN2 (________26802), .Q
       (_____9__27667));
  nor2s1 ____9__506893(.DIN1 (________27665), .DIN2 (________27664), .Q
       (________27666));
  or2s1 ____9__506894(.DIN1 (________27662), .DIN2 (________26850), .Q
       (________27663));
  nnd2s1 ____9_506895(.DIN1 (____99__27208), .DIN2 (________27660), .Q
       (________27661));
  nor2s1 ____0__506896(.DIN1 (___9____25980), .DIN2 (____0___27658), .Q
       (____09__27659));
  nor2s1 ____0__506897(.DIN1 (____9___27293), .DIN2 (__9_____30401), .Q
       (____0___27656));
  hi1s1 _____9_506898(.DIN (___09___27914), .Q (____99__27653));
  nnd2s1 ____9__506899(.DIN1 (___99___26950), .DIN2 (inData[18]), .Q
       (____9___27652));
  nnd2s1 ____90_506900(.DIN1 (___0____26963), .DIN2 (____9___27649), .Q
       (____9___27650));
  nnd2s1 ____0_506901(.DIN1 (____90__27647), .DIN2 (_____9__27646), .Q
       (____9___27648));
  nnd2s1 ____90_506902(.DIN1 (___0____26970), .DIN2 (________26621), .Q
       (________27645));
  hi1s1 ______506903(.DIN (__________0_), .Q (________27644));
  nnd2s1 ____0__506904(.DIN1 (________27090), .DIN2 (___0_9__27017), .Q
       (________27643));
  nnd2s1 ____0__506905(.DIN1 (___0____27003), .DIN2 (inData[4]), .Q
       (________27642));
  nnd2s1 ____0__506906(.DIN1 (________27640), .DIN2 (____90__27113), .Q
       (________27641));
  nor2s1 ____0_506907(.DIN1 (________27638), .DIN2 (___0____26997), .Q
       (________27639));
  nnd2s1 ____0__506908(.DIN1 (_____9__27636), .DIN2 (________26716), .Q
       (_____0__27637));
  or2s1 ____0__506909(.DIN1 (_____9__26379), .DIN2 (________27078), .Q
       (________27635));
  and2s1 ____0__506910(.DIN1 (________27633), .DIN2 (________27415), .Q
       (________27634));
  nnd2s1 ____90_506911(.DIN1 (________27097), .DIN2 (inData[28]), .Q
       (________27632));
  nor2s1 ____90_506912(.DIN1 (________26451), .DIN2 (____9___29458), .Q
       (________27631));
  nnd2s1 ____0_506913(.DIN1 (_________41224), .DIN2 (________25807), .Q
       (________27630));
  nnd2s1 _____9_506914(.DIN1 (_________41224), .DIN2 (_____0__24516),
       .Q (________27629));
  nnd2s1 ____506915(.DIN1 (________27640), .DIN2 (________27143), .Q
       (_____9__27628));
  nnd2s1 _______506916(.DIN1 (___99___26951), .DIN2 (inData[22]), .Q
       (________27626));
  nor2s1 ______506917(.DIN1 (_____0__26528), .DIN2 (______0__41220), .Q
       (________27625));
  nor2s1 _______506918(.DIN1 (________26470), .DIN2 (___0____27025), .Q
       (________27624));
  and2s1 ______506919(.DIN1 (___0____26972), .DIN2 (___0_____31297), .Q
       (________27623));
  nnd2s1 _______506920(.DIN1 (________27083), .DIN2 (________26713), .Q
       (________27622));
  nnd2s1 _____9_506921(.DIN1 (_____0__27620), .DIN2 (_____9__27619), .Q
       (________27621));
  nnd2s1 ______506922(.DIN1 (_____9__29314), .DIN2 (___0_____31274), .Q
       (________28309));
  hi1s1 _____0_506923(.DIN (_____0__29495), .Q (________28159));
  hi1s1 _____0_506924(.DIN (___090__27912), .Q (________28144));
  hi1s1 _____0_506925(.DIN (___0____27910), .Q (________28143));
  hi1s1 _____9_506926(.DIN (________27617), .Q (________28390));
  or2s1 ____0__506927(.DIN1 (________27616), .DIN2 (____0___27487), .Q
       (________28875));
  nor2s1 _______506928(.DIN1 (________27615), .DIN2 (___0____26992), .Q
       (________28445));
  nnd2s1 _______506929(.DIN1 (________27614), .DIN2 (________27613), .Q
       (__9_____30109));
  nor2s1 _______506930(.DIN1 (____00___31509), .DIN2 (________28311),
       .Q (___0____27876));
  nor2s1 _____0_506931(.DIN1 (___9____29571), .DIN2 (____0___27037), .Q
       (________28407));
  nor2s1 ____0__506932(.DIN1 (___9_0__27805), .DIN2 (__90____29663), .Q
       (________28161));
  xor2s1 _______506933(.DIN1 (___0____22335), .DIN2 (_________41252),
       .Q (_____9__28423));
  nnd2s1 ____0__506934(.DIN1 (___9____26906), .DIN2 (________26308), .Q
       (______9__32733));
  and2s1 ____0_506935(.DIN1 (_________41222), .DIN2 (________27611), .Q
       (________28163));
  nor2s1 ______506936(.DIN1 (___9_9__26948), .DIN2 (___09___27918), .Q
       (____0____32550));
  nnd2s1 _______506937(.DIN1 (________27142), .DIN2 (_____0__26758), .Q
       (___0_____30939));
  nnd2s1 _______506938(.DIN1 (_____0__27610), .DIN2 (_____9__27609), .Q
       (________28427));
  or2s1 ______506939(.DIN1 (________28909), .DIN2 (____9___27114), .Q
       (________28456));
  and2s1 _______506940(.DIN1 (________27050), .DIN2 (__99____30533), .Q
       (_____0__28298));
  nor2s1 ____0__506941(.DIN1 (________24801), .DIN2 (___0____27024), .Q
       (________29223));
  or2s1 _______506942(.DIN1 (________25741), .DIN2 (________27982), .Q
       (__9_____30071));
  nor2s1 _______506943(.DIN1 (___9____27800), .DIN2 (________27051), .Q
       (__9_99__29895));
  hi1s1 _____0_506944(.DIN (________27607), .Q (____0____31577));
  and2s1 ______506945(.DIN1 (___0_____31362), .DIN2 (___0____26116), .Q
       (__9_____29843));
  nor2s1 _______506946(.DIN1 (________29531), .DIN2 (________27681), .Q
       (_____0__28395));
  nnd2s1 ______506947(.DIN1 (_____0__29213), .DIN2 (___0____27012), .Q
       (________28412));
  nor2s1 _______506948(.DIN1 (_________31906), .DIN2 (____09__27038),
       .Q (__9_____29941));
  hi1s1 _____0_506949(.DIN (________27606), .Q (___0_9___31405));
  hi1s1 _______506950(.DIN (________27603), .Q (_____0__28306));
  nnd2s1 _______506951(.DIN1 (________27170), .DIN2 (___0_90__30919),
       .Q (___0_____30956));
  nnd2s1 _______506952(.DIN1 (________27605), .DIN2 (________27432), .Q
       (__9__9__30262));
  hi1s1 _______506953(.DIN
       (_____________________________________________21896), .Q
       (_________35859));
  hi1s1 _______506954(.DIN (___0_9___40354), .Q (___0_____40326));
  nnd2s1 _______506955(.DIN1 (___0_____40222), .DIN2 (________27604),
       .Q (___0__9__40232));
  dffacs1 ______________________________________________9_506956(.CLRB
       (reset), .CLK (clk), .DIN (________27145), .QN
       (__________________________________________9___21934));
  hi1s1 _______506957(.DIN (____9____33397), .Q (___9_0___39170));
  nor2s1 _______506958(.DIN1 (________27150), .DIN2 (____0___27127), .Q
       (___0_____40156));
  hi1s1 _______506959(.DIN (________27945), .Q (___0_9__28804));
  nor2s1 _______506960(.DIN1 (________26611), .DIN2 (____9___27116), .Q
       (___9_____39219));
  nnd2s1 _______506961(.DIN1 (________27131), .DIN2 (________27602), .Q
       (______0__35537));
  hi1s1 ____0__506962(.DIN
       (_____________________________________0___0_), .Q
       (_____9__27601));
  or2s1 _______506963(.DIN1 (_____9__27138), .DIN2 (________28225), .Q
       (________27600));
  nnd2s1 _____9_506964(.DIN1 (____9___27119), .DIN2 (________27598), .Q
       (________27599));
  nor2s1 _______506965(.DIN1 (____9____32424), .DIN2 (__9_____29862),
       .Q (________27597));
  nor2s1 ______506966(.DIN1 (________27458), .DIN2 (___0__9__31347), .Q
       (________27596));
  nnd2s1 _______506967(.DIN1 (_____0___41214), .DIN2 (____9___28198),
       .Q (________27595));
  nor2s1 _______506968(.DIN1 (__90_9__29688), .DIN2 (___0____28820), .Q
       (________27594));
  nor2s1 _______506969(.DIN1 (________26279), .DIN2 (___0____26990), .Q
       (_____0__27593));
  hi1s1 _____0_506970(.DIN (________27589), .Q (________27590));
  hi1s1 _______506971(.DIN (________27587), .Q (________27588));
  hi1s1 _______506972(.DIN (_____0__27585), .Q (________27586));
  nor2s1 ______506973(.DIN1 (__9_____30222), .DIN2 (________27582), .Q
       (________27583));
  nnd2s1 _______506974(.DIN1 (________27086), .DIN2 (___9_0__26013), .Q
       (________27581));
  nor2s1 _______506975(.DIN1 (___90___28652), .DIN2 (________27096), .Q
       (________27580));
  or2s1 _______506976(.DIN1 (_____0__27578), .DIN2 (____0___29200), .Q
       (________27579));
  nor2s1 _______506977(.DIN1 (___00___26958), .DIN2 (____0___27576), .Q
       (____09__27577));
  nnd2s1 _______506978(.DIN1 (___09____40685), .DIN2 (____9___27295),
       .Q (____0___27575));
  or2s1 _______506979(.DIN1 (____0___27573), .DIN2 (____0___29200), .Q
       (____0___27574));
  or2s1 ______506980(.DIN1 (____0___27571), .DIN2 (____0___27570), .Q
       (____0___27572));
  nnd2s1 _______506981(.DIN1 (_____0__27067), .DIN2 (_____0___41212),
       .Q (____00__27569));
  or2s1 _____9_506982(.DIN1 (___0__0__31003), .DIN2 (__999___30539), .Q
       (____99__27568));
  or2s1 _____9_506983(.DIN1 (____9___27566), .DIN2 (__9_9___30449), .Q
       (____9___27567));
  nnd2s1 _____0_506984(.DIN1 (___990__26949), .DIN2 (____9___27564), .Q
       (____9___27565));
  or2s1 _____0_506985(.DIN1 (________26152), .DIN2 (________28937), .Q
       (____9___27563));
  nnd2s1 _____0_506986(.DIN1 (________27518), .DIN2 (___9____26922), .Q
       (____9___27562));
  nor2s1 _____506987(.DIN1 (___9_9__26910), .DIN2 (____9___27560), .Q
       (____9___27561));
  nor2s1 ______506988(.DIN1 (________28900), .DIN2 (__9_____29783), .Q
       (____90__27559));
  nnd2s1 _______506989(.DIN1 (_________41222), .DIN2 (________26369),
       .Q (_____9__27558));
  or2s1 _______506990(.DIN1 (________27190), .DIN2 (___0____27906), .Q
       (________27557));
  nor2s1 _______506991(.DIN1 (________29053), .DIN2 (___0____26961), .Q
       (________27556));
  nor2s1 ______506992(.DIN1 (________28936), .DIN2 (____9___27560), .Q
       (________27555));
  or2s1 ______506993(.DIN1 (___900__29553), .DIN2 (__9_____30401), .Q
       (________27553));
  nor2s1 _______506994(.DIN1 (_____9__27551), .DIN2 (__9_____29783), .Q
       (_____0__27552));
  nor2s1 _______506995(.DIN1 (________27549), .DIN2 (__9_____30401), .Q
       (________27550));
  nor2s1 _______506996(.DIN1 (___9____26898), .DIN2 (________27547), .Q
       (________27548));
  or2s1 _______506997(.DIN1 (________27545), .DIN2 (________27544), .Q
       (________27546));
  nor2s1 _______506998(.DIN1 (___0____25141), .DIN2 (________28936), .Q
       (_____0__27543));
  nnd2s1 _______506999(.DIN1 (__9_____30322), .DIN2 (________27541), .Q
       (_____9__27542));
  nor2s1 ______507000(.DIN1 (_____9__27498), .DIN2 (_________41226), .Q
       (________27540));
  or2s1 _______507001(.DIN1 (________27538), .DIN2 (__999___30539), .Q
       (________27539));
  or2s1 _______507002(.DIN1 (___0_____30810), .DIN2 (__90____29663), .Q
       (________27537));
  and2s1 _______507003(.DIN1 (_____0__28181), .DIN2 (________27535), .Q
       (________27536));
  nor2s1 _______507004(.DIN1 (_____0__24307), .DIN2 (______0__41220),
       .Q (________27534));
  nor2s1 ______507005(.DIN1 (________27532), .DIN2 (________27544), .Q
       (_____9__27533));
  nnd2s1 _______507006(.DIN1 (___0_9__26976), .DIN2 (_____9__27551), .Q
       (________27531));
  nor2s1 _______507007(.DIN1 (___090___31413), .DIN2 (___9____26943),
       .Q (________27530));
  or2s1 _______507008(.DIN1 (__9__9__29935), .DIN2 (____99__28107), .Q
       (________27529));
  or2s1 ______507009(.DIN1 (________29533), .DIN2 (__90____29663), .Q
       (________27528));
  or2s1 _______507010(.DIN1 (________27526), .DIN2 (________27991), .Q
       (________27527));
  or2s1 _______507011(.DIN1 (________27964), .DIN2 (___0____26969), .Q
       (________27525));
  or2s1 _______507012(.DIN1 (_________31811), .DIN2 (__9_____30401), .Q
       (_____0__27524));
  nor2s1 _______507013(.DIN1 (________27522), .DIN2 (___9____26946), .Q
       (_____9__27523));
  nnd2s1 _______507014(.DIN1 (____9____33386), .DIN2 (____0___29285),
       .Q (________27521));
  or2s1 ______507015(.DIN1 (______0__41230), .DIN2 (________27664), .Q
       (________27520));
  nnd2s1 _____9_507016(.DIN1 (________27518), .DIN2 (___0____26996), .Q
       (________27519));
  nor2s1 _____9_507017(.DIN1 (________26475), .DIN2 (______0__32892),
       .Q (________27517));
  nor2s1 _____507018(.DIN1 (________27721), .DIN2 (________27049), .Q
       (________27516));
  and2s1 _____0_507019(.DIN1 (________27535), .DIN2 (________26154), .Q
       (_____0__27515));
  nor2s1 _______507020(.DIN1 (________27615), .DIN2 (________27513), .Q
       (________27514));
  or2s1 _______507021(.DIN1 (_________41226), .DIN2 (________27511), .Q
       (________27512));
  or2s1 _______507022(.DIN1 (____0___26325), .DIN2 (________27509), .Q
       (________27510));
  nor2s1 _______507023(.DIN1 (___9_0__25968), .DIN2 (_____0__27507), .Q
       (________27508));
  nnd2s1 _______507024(.DIN1 (___0____26986), .DIN2 (________27505), .Q
       (_____9__27506));
  hi1s1 ____0__507025(.DIN (_____9___41208), .Q (________27503));
  hi1s1 ____0__507026(.DIN (________27501), .Q (________27502));
  or2s1 _______507027(.DIN1 (_____9__27498), .DIN2 (_____0___41218), .Q
       (_____0__27499));
  nnd2s1 ______507028(.DIN1 (___0____26983), .DIN2 (____0___28293), .Q
       (________27497));
  nor2s1 _______507029(.DIN1 (________27089), .DIN2 (___0____28820), .Q
       (________27496));
  or2s1 ____0_507030(.DIN1 (_________32065), .DIN2 (___0____27000), .Q
       (________28250));
  nnd2s1 ____09_507031(.DIN1 (_____9__27636), .DIN2 (________27495), .Q
       (___99___27824));
  or2s1 ____507032(.DIN1 (_____9__27102), .DIN2 (___09____31478), .Q
       (________28236));
  and2s1 _______507033(.DIN1 (________28154), .DIN2 (________27494), .Q
       (_____0__28247));
  nnd2s1 _______507034(.DIN1 (_________31935), .DIN2 (________27493),
       .Q (________28213));
  nor2s1 _______507035(.DIN1 (___0____27022), .DIN2 (________27492), .Q
       (________28211));
  nor2s1 ______507036(.DIN1 (________27491), .DIN2 (________27178), .Q
       (____0___28383));
  nor2s1 _______507037(.DIN1 (_____0__26508), .DIN2 (________28187), .Q
       (________28304));
  and2s1 _______507038(.DIN1 (_____0__27490), .DIN2 (____09__27489), .Q
       (________28155));
  nnd2s1 _______507039(.DIN1 (_____9__28246), .DIN2 (___0____26086), .Q
       (_____9__28147));
  nnd2s1 ______507040(.DIN1 (___0_9___31403), .DIN2 (_________32022),
       .Q (____0___28207));
  nor2s1 _______507041(.DIN1 (____0___27488), .DIN2 (_____9__27204), .Q
       (________28150));
  nor2s1 _______507042(.DIN1 (______9__32852), .DIN2 (___0____26974),
       .Q (__9_____29911));
  nor2s1 _______507043(.DIN1 (___0____25136), .DIN2 (___0____26980), .Q
       (_________32218));
  or2s1 _____9_507044(.DIN1 (_________32056), .DIN2 (___9____26941), .Q
       (________28233));
  nor2s1 _____9_507045(.DIN1 (____0___27487), .DIN2 (________27284), .Q
       (___99___27826));
  nnd2s1 ______507046(.DIN1 (___090__27026), .DIN2 (________27545), .Q
       (___9_9__27794));
  nor2s1 _____0_507047(.DIN1 (___0____27863), .DIN2 (____9___27560), .Q
       (________28316));
  or2s1 _____0_507048(.DIN1 (__9__0__29916), .DIN2 (_____0__27507), .Q
       (________28357));
  hi1s1 ____0__507049(.DIN (____0___27486), .Q (________28170));
  hi1s1 ____0_507050(.DIN (____0___27485), .Q (________28283));
  nnd2s1 _____0_507051(.DIN1 (____9___27474), .DIN2
       (_____________________21741), .Q (________28307));
  nnd2s1 _____507052(.DIN1 (___0____27020), .DIN2 (___9_0__27795), .Q
       (___99___27823));
  hi1s1 _____507053(.DIN (_________32241), .Q (________28145));
  nor2s1 _______507054(.DIN1 (____0___27484), .DIN2 (_____9__27092), .Q
       (_____9__28256));
  nor2s1 ____0__507055(.DIN1 (___9____27820), .DIN2 (________27087), .Q
       (________28264));
  nnd2s1 ____0__507056(.DIN1 (___0____26973), .DIN2 (________25340), .Q
       (________29238));
  nnd2s1 _______507057(.DIN1 (____0___27483), .DIN2 (___0____27853), .Q
       (___9____27770));
  or2s1 _______507058(.DIN1 (____0___27482), .DIN2 (___0____26984), .Q
       (________29519));
  nor2s1 _______507059(.DIN1 (________27491), .DIN2 (____0___27481), .Q
       (__9_0___29729));
  dffacs1 ________________________________________________507060(.CLRB
       (reset), .CLK (clk), .DIN (_____9__27147), .QN
       (______________________________________________21933));
  nor2s1 _______507061(.DIN1 (________27724), .DIN2 (____00__27480), .Q
       (__9_____30325));
  and2s1 _______507062(.DIN1 (________28154), .DIN2 (________28952), .Q
       (________29031));
  nnd2s1 _______507063(.DIN1 (___09___27027), .DIN2 (___9_0__27805), .Q
       (____0___28201));
  nnd2s1 _______507064(.DIN1 (____0___28382), .DIN2 (________27495), .Q
       (____0___28377));
  nnd2s1 _______507065(.DIN1 (___0_____31078), .DIN2 (___0_____30676),
       .Q (__9_0___30373));
  or2s1 _______507066(.DIN1 (___9____27766), .DIN2 (__9__0__30291), .Q
       (_________33137));
  dffacs1 _______________________________________________507067(.CLRB
       (reset), .CLK (clk), .DIN (________27098), .Q (___0_____40439));
  nnd2s1 _______507068(.DIN1 (____99__27479), .DIN2 (_____9__28100), .Q
       (________28334));
  nnd2s1 ______507069(.DIN1 (___9____26906), .DIN2 (________28034), .Q
       (____9___28194));
  nnd2s1 _______507070(.DIN1 (___09____31469), .DIN2 (___9_0__26911),
       .Q (________28343));
  nnd2s1 _______507071(.DIN1 (____9___27478), .DIN2 (____9___27477), .Q
       (_____9__28368));
  nnd2s1 _______507072(.DIN1 (____0___29285), .DIN2 (_________33123),
       .Q (_________33193));
  hi1s1 ____0__507073(.DIN (____9___27476), .Q (__9_____29908));
  nor2s1 _______507074(.DIN1 (_____0__26738), .DIN2 (________27544), .Q
       (___0_____31229));
  nnd2s1 ______507075(.DIN1 (____0___29285), .DIN2 (____9___27475), .Q
       (_________32808));
  nnd2s1 _______507076(.DIN1 (________29171), .DIN2 (____9___27477), .Q
       (____9___28915));
  nor2s1 _______507077(.DIN1 (___0____27019), .DIN2 (_________31843),
       .Q (________28386));
  nor2s1 _______507078(.DIN1 (_____9__27066), .DIN2 (_________32748),
       .Q (__99____30468));
  and2s1 _______507079(.DIN1 (____9___27474), .DIN2 (____0___25502), .Q
       (__9_____29870));
  nnd2s1 _______507080(.DIN1 (____9___27474), .DIN2 (________26618), .Q
       (___00____30606));
  dffacs1 _______________________________________507081(.CLRB (reset),
       .CLK (clk), .DIN (___099__27030), .Q (______________22111));
  nnd2s1 ______507082(.DIN1 (___9____26906), .DIN2 (_________31879), .Q
       (_____9___34186));
  dffacs1 _______________________________________507083(.CLRB (reset),
       .CLK (clk), .DIN (________27095), .QN (___0_____40449));
  hi1s1 _______507084(.DIN (____9___27473), .Q (_________31836));
  nor2s1 ______507085(.DIN1 (______0__41250), .DIN2 (____9____33386),
       .Q (_________32692));
  dffacs1 _____________________________________0_(.CLRB (reset), .CLK
       (clk), .DIN (________27088), .QN (___0__9__40450));
  nnd2s1 _____507086(.DIN1 (___9____26906), .DIN2 (inData[17]), .Q
       (______0__32253));
  hi1s1 _______507087(.DIN (__90____29665), .Q (___09___28829));
  nnd2s1 ______507088(.DIN1 (___0____26962), .DIN2 (____9____32424), .Q
       (_____9___34752));
  nnd2s1 _______507089(.DIN1 (___9____26906), .DIN2 (________26638), .Q
       (_________33695));
  nnd2s1 _______507090(.DIN1 (_____9__28246), .DIN2 (________28952), .Q
       (________28268));
  dffacs1 ______________________________________507091(.CLRB (reset),
       .CLK (clk), .DIN (____0___27126), .Q (_____________22084));
  nnd2s1 _______507092(.DIN1 (___0____26975), .DIN2 (________25735), .Q
       (_________37864));
  nnd2s1 _____9_507093(.DIN1 (___0____26965), .DIN2 (________26575), .Q
       (______9__37429));
  hi1s1 ______507094(.DIN (_________33650), .Q (____990__33424));
  nor2s1 _____9_507095(.DIN1 (____99__26407), .DIN2 (________27062), .Q
       (___9_0___39077));
  hi1s1 _______507096(.DIN (____90__27472), .Q (____0___28295));
  hi1s1 _______507097(.DIN (________27618), .Q (_________38280));
  nor2s1 _______507098(.DIN1 (inData[17]), .DIN2 (____9____33386), .Q
       (______9__32753));
  nor2s1 _____9_507099(.DIN1 (________26450), .DIN2 (___99___26952), .Q
       (___0_____40100));
  hi1s1 _______507100(.DIN (__9_____30019), .Q (__9_____30417));
  or2s1 ____99_507101(.DIN1 (_____9__27452), .DIN2 (________26811), .Q
       (________27470));
  nor2s1 _____9_507102(.DIN1 (___0_____30695), .DIN2 (________26663),
       .Q (________27469));
  and2s1 _______507103(.DIN1 (___09____31443), .DIN2 (________26667),
       .Q (________27467));
  and2s1 _______507104(.DIN1 (____0____37165), .DIN2 (________22687),
       .Q (________27466));
  nnd2s1 _______507105(.DIN1 (________26721), .DIN2 (_____9__26537), .Q
       (________27465));
  nor2s1 ______507106(.DIN1 (________25661), .DIN2 (_____0__27463), .Q
       (________27464));
  nnd2s1 _______507107(.DIN1 (________29171), .DIN2 (________26277), .Q
       (_____9__27462));
  nnd2s1 _______507108(.DIN1 (_____9__27075), .DIN2 (___90___28650), .Q
       (________27461));
  nor2s1 _______507109(.DIN1 (________22876), .DIN2 (_____0__26692), .Q
       (________27460));
  nor2s1 _______507110(.DIN1 (_____0__27427), .DIN2 (________27458), .Q
       (________27459));
  nnd2s1 _______507111(.DIN1 (_____9___38610), .DIN2 (_________33973),
       .Q (________27457));
  nor2s1 ______507112(.DIN1 (________27608), .DIN2 (__9_____30312), .Q
       (________27456));
  or2s1 _______507113(.DIN1 (________27454), .DIN2 (__9_____30312), .Q
       (________27455));
  or2s1 _______507114(.DIN1 (_____9__27452), .DIN2 (_____9__27986), .Q
       (_____0__27453));
  xnr2s1 ______507115(.DIN1
       (_____________________________________________21809), .DIN2
       (____0_0__38064), .Q (________27451));
  xor2s1 ______507116(.DIN1
       (_____________________________________________21842), .DIN2
       (___9_____39738), .Q (________27450));
  nnd2s1 _______507117(.DIN1 (________27448), .DIN2 (_____0__26608), .Q
       (________27449));
  and2s1 _______507118(.DIN1 (________28543), .DIN2 (________27446), .Q
       (________27447));
  xor2s1 _____9_507119(.DIN1 (________27444), .DIN2 (_________32611),
       .Q (________27445));
  xor2s1 _____9_507120(.DIN1 (________22436), .DIN2 (_________38666),
       .Q (_____0__27443));
  xnr2s1 _____9_507121(.DIN1
       (_____________________________________0___0___21760), .DIN2
       (____0_9__36267), .Q (_____9__27442));
  xor2s1 _____0_507122(.DIN1 (_________36856), .DIN2 (_________38876),
       .Q (________27441));
  nor2s1 ______507123(.DIN1 (___0_____31242), .DIN2 (________26763), .Q
       (________27438));
  nnd2s1 _______507124(.DIN1 (____9___26768), .DIN2 (____0___24747), .Q
       (________27437));
  nnd2s1 _______507125(.DIN1 (_________41232), .DIN2 (inData[22]), .Q
       (________27436));
  and2s1 _______507126(.DIN1 (________27283), .DIN2 (_____9__27434), .Q
       (_____0__27435));
  hi1s1 _______507127(.DIN (________27432), .Q (________27433));
  nnd2s1 _______507128(.DIN1 (________26659), .DIN2 (________28596), .Q
       (________27431));
  or2s1 _______507129(.DIN1 (________27429), .DIN2 (__9_____29881), .Q
       (________27430));
  or2s1 ______507130(.DIN1 (________28044), .DIN2 (_____0__27427), .Q
       (________27428));
  nnd2s1 _______507131(.DIN1 (________27425), .DIN2 (___0____27023), .Q
       (_____9__27426));
  nor2s1 _______507132(.DIN1 (___09____31478), .DIN2 (_____0__26839),
       .Q (________27424));
  and2s1 _______507133(.DIN1 (________26661), .DIN2 (________28596), .Q
       (________27423));
  nnd2s1 _______507134(.DIN1 (____0___26688), .DIN2 (________27421), .Q
       (________27422));
  nnd2s1 _______507135(.DIN1 (___09____31461), .DIN2 (________26745),
       .Q (________27420));
  nnd2s1 _______507136(.DIN1 (________26723), .DIN2
       (_____________________________________9_____), .Q
       (________27418));
  and2s1 _______507137(.DIN1 (________27416), .DIN2 (________27415), .Q
       (________27417));
  or2s1 _______507138(.DIN1 (____99__26774), .DIN2 (______9__33267), .Q
       (________27414));
  nnd2s1 _______507139(.DIN1 (________26825), .DIN2 (________25551), .Q
       (________27413));
  nor2s1 ______507140(.DIN1 (___0_____40620), .DIN2 (____0___27394), .Q
       (________27412));
  nor2s1 _____9_507141(.DIN1 (___9____26934), .DIN2 (________27409), .Q
       (_____9__27410));
  nor2s1 _____9_507142(.DIN1 (________28860), .DIN2 (_____9__26847), .Q
       (________27408));
  nor2s1 _____9_507143(.DIN1 (___0_0__26102), .DIN2 (________26623), .Q
       (________27407));
  and2s1 _____507144(.DIN1 (________27405), .DIN2 (___9____26903), .Q
       (________27406));
  nnd2s1 ____507145(.DIN1 (_____90__35555), .DIN2 (________26791), .Q
       (________27404));
  nnd2s1 ____90_507146(.DIN1 (________27402), .DIN2
       (_____________22081), .Q (________27403));
  nnd2s1 ____90_507147(.DIN1 (____9___26766), .DIN2 (inData[6]), .Q
       (_____0__27401));
  nor2s1 ____507148(.DIN1 (inData[24]), .DIN2 (____0____37165), .Q
       (____09__27400));
  and2s1 ____9__507149(.DIN1 (___90___26866), .DIN2 (____0___27398), .Q
       (____0___27399));
  and2s1 ____9__507150(.DIN1 (___0____28788), .DIN2 (____0___27396), .Q
       (____0___27397));
  nor2s1 ____9__507151(.DIN1 (___0_99__40460), .DIN2 (____0___27394),
       .Q (____0___27395));
  nor2s1 ____9__507152(.DIN1 (___0_9__26091), .DIN2 (____99__27391), .Q
       (____00__27392));
  nor2s1 ____9__507153(.DIN1 (____9___27389), .DIN2 (____09__26691), .Q
       (____9___27390));
  nor2s1 ____9__507154(.DIN1 (___9____26897), .DIN2 (_________32701),
       .Q (____9___27388));
  and2s1 ____9__507155(.DIN1 (___9____26905), .DIN2 (____9___27386), .Q
       (____9___27387));
  nnd2s1 ____9__507156(.DIN1 (_________41244), .DIN2 (________28074),
       .Q (____9___27385));
  nnd2s1 ____9__507157(.DIN1 (____9___27383), .DIN2 (____90__27382), .Q
       (____9___27384));
  nnd2s1 ____9__507158(.DIN1 (________26801), .DIN2 (________25889), .Q
       (_____9__27381));
  nnd2s1 ____9__507159(.DIN1 (________26813), .DIN2 (___9____26900), .Q
       (________27380));
  nor2s1 ____9_507160(.DIN1 (________27378), .DIN2 (_____9__26803), .Q
       (________27379));
  or2s1 ____9_507161(.DIN1 (_____00__34847), .DIN2 (________26852), .Q
       (________27377));
  nnd2s1 ____9__507162(.DIN1 (______0__41240), .DIN2 (________24590),
       .Q (________27376));
  nor2s1 ____9__507163(.DIN1 (___9____26885), .DIN2 (_________41236),
       .Q (________27375));
  nnd2s1 ____9__507164(.DIN1 (________27324), .DIN2 (____9___25854), .Q
       (________27374));
  nor2s1 ____9__507165(.DIN1 (________28850), .DIN2 (_____9__29074), .Q
       (________27373));
  nnd2s1 ____9__507166(.DIN1 (________26836), .DIN2 (________26819), .Q
       (_____0__27372));
  nnd2s1 ____9__507167(.DIN1 (_____9__26672), .DIN2 (inData[24]), .Q
       (_____9__27371));
  or2s1 ____9_507168(.DIN1 (_____0__26203), .DIN2 (________26670), .Q
       (________27370));
  nnd2s1 ____9__507169(.DIN1 (________26792), .DIN2 (inData[26]), .Q
       (________27369));
  or2s1 ____9__507170(.DIN1 (_____9__26447), .DIN2 (_________41234), .Q
       (________27368));
  and2s1 ____9__507171(.DIN1 (____0____37165), .DIN2 (________22404),
       .Q (________27367));
  and2s1 ____9__507172(.DIN1 (__9_____29968), .DIN2 (__99____30506), .Q
       (________27366));
  and2s1 ____9__507173(.DIN1 (________27448), .DIN2 (_____0__27363), .Q
       (________27364));
  nnd2s1 ____9__507174(.DIN1 (____0_0__37159), .DIN2 (________22815),
       .Q (_____9__27362));
  nnd2s1 ____9__507175(.DIN1 (_____9__26821), .DIN2 (inData[10]), .Q
       (________27361));
  nnd2s1 ____9__507176(.DIN1 (________26697), .DIN2 (______0__37731),
       .Q (________27360));
  nnd2s1 ____9__507177(.DIN1 (____9___26771), .DIN2 (________26196), .Q
       (________27359));
  and2s1 ____9__507178(.DIN1 (___0_____40222), .DIN2 (_______22175), .Q
       (________27358));
  and2s1 ____9__507179(.DIN1 (_____0__26645), .DIN2 (___9____27764), .Q
       (________27357));
  nor2s1 ____9__507180(.DIN1 (________27355), .DIN2 (_________41236),
       .Q (________27356));
  nnd2s1 ____9_507181(.DIN1 (_________41228), .DIN2 (____99__25677), .Q
       (_____0__27354));
  and2s1 ____9__507182(.DIN1 (________26761), .DIN2 (________28523), .Q
       (________27352));
  nnd2s1 ____9__507183(.DIN1 (________27711), .DIN2 (____0___26780), .Q
       (________27351));
  nnd2s1 ____9__507184(.DIN1 (___900__29553), .DIN2 (________28122), .Q
       (________27350));
  nor2s1 ____9__507185(.DIN1 (________27638), .DIN2 (____0___26776), .Q
       (________27349));
  nnd2s1 ____9__507186(.DIN1 (_____9__27326), .DIN2
       (_____________________________________________21778), .Q
       (________27348));
  or2s1 ____99_507187(.DIN1
       (_____________________________________________21778), .DIN2
       (________27315), .Q (________27347));
  nor2s1 ____99_507188(.DIN1 (_____0__27345), .DIN2 (_____9__27344), .Q
       (________27346));
  and2s1 ____99_507189(.DIN1 (___00___26957), .DIN2 (________25541), .Q
       (________27343));
  nnd2s1 ____99_507190(.DIN1 (________26844), .DIN2 (__9_____29949), .Q
       (________27342));
  and2s1 ____99_507191(.DIN1 (_____9__26831), .DIN2 (________27339), .Q
       (________27340));
  and2s1 ____507192(.DIN1 (_____9__27335), .DIN2 (___0_9__26121), .Q
       (________27338));
  or2s1 ____00_507193(.DIN1 (________26740), .DIN2 (_____0__27427), .Q
       (________27337));
  nnd2s1 ____00_507194(.DIN1 (_____9___32673), .DIN2 (_____9__27335),
       .Q (_____0__27336));
  or2s1 ____00_507195(.DIN1 (________27333), .DIN2 (_____0__28863), .Q
       (________27334));
  nor2s1 ____00_507196(.DIN1 (________26820), .DIN2 (________26515), .Q
       (________27332));
  or2s1 ____00_507197(.DIN1 (__9_____30054), .DIN2 (____9___26861), .Q
       (________27331));
  nnd2s1 ____00_507198(.DIN1 (________26788), .DIN2 (________26166), .Q
       (________27330));
  and2s1 ____0__507199(.DIN1 (____0_0__37159), .DIN2 (___0_____40572),
       .Q (________27329));
  nnd2s1 ____0__507200(.DIN1 (___99___28731), .DIN2 (________25936), .Q
       (________27328));
  nnd2s1 ____0__507201(.DIN1 (_____9__27326), .DIN2 (____0____35320),
       .Q (_____0__27327));
  nnd2s1 ____0__507202(.DIN1 (________27324), .DIN2 (_____9__27056), .Q
       (________27325));
  nnd2s1 ____0__507203(.DIN1 (________27322), .DIN2 (___9____25969), .Q
       (________27323));
  nor2s1 ____0__507204(.DIN1 (________27320), .DIN2 (_____9__26793), .Q
       (________27321));
  nnd2s1 ____0__507205(.DIN1 (________26800), .DIN2 (___0____26982), .Q
       (________27319));
  nnd2s1 ____0_507206(.DIN1 (_____0__27317), .DIN2 (________23524), .Q
       (________27318));
  or2s1 ____0_507207(.DIN1 (____0____35320), .DIN2 (________27315), .Q
       (_____9__27316));
  nnd2s1 ____0__507208(.DIN1 (____0___26689), .DIN2 (________27313), .Q
       (________27314));
  nnd2s1 ____0__507209(.DIN1 (________27311), .DIN2 (_____0__27578), .Q
       (________27312));
  nnd2s1 ____0__507210(.DIN1 (_____0__26848), .DIN2 (________27446), .Q
       (________27310));
  or2s1 ____0_507211(.DIN1 (_________33986), .DIN2 (_____0__26785), .Q
       (_____0__27308));
  nnd2s1 ____0__507212(.DIN1 (_____9__28626), .DIN2 (____9___25954), .Q
       (____09__27307));
  and2s1 ____0__507213(.DIN1 (________27365), .DIN2 (________27168), .Q
       (____0___27306));
  nnd2s1 ____0__507214(.DIN1 (___0____27021), .DIN2 (________27313), .Q
       (____0___27305));
  nor2s1 ____0_507215(.DIN1 (____90__27290), .DIN2 (____0___27301), .Q
       (____0___27304));
  nnd2s1 ____0_507216(.DIN1 (____99__26498), .DIN2 (____09__26784), .Q
       (____0___27303));
  xor2s1 _______507217(.DIN1 (___09_), .DIN2 (___9_0___39624), .Q
       (________27708));
  nnd2s1 ____0__507218(.DIN1 (___90___26869), .DIN2 (________28074), .Q
       (____9___28103));
  nor2s1 ____0__507219(.DIN1 (__90____29692), .DIN2 (____9___27291), .Q
       (___0_9___31301));
  nor2s1 ____0__507220(.DIN1 (inData[21]), .DIN2 (___0900), .Q
       (___0_9__27911));
  nor2s1 ____0_507221(.DIN1 (________26750), .DIN2 (____0___27301), .Q
       (________27999));
  or2s1 ____0__507222(.DIN1 (_________34207), .DIN2 (________26630), .Q
       (____9___28007));
  nor2s1 ____0__507223(.DIN1 (____00__27300), .DIN2 (____99__27299), .Q
       (________28030));
  nor2s1 ____0__507224(.DIN1 (____9___27298), .DIN2 (________26817), .Q
       (____9___29006));
  nnd2s1 ____0__507225(.DIN1 (_________41246), .DIN2 (____9___27297),
       .Q (________27951));
  nor2s1 ____09_507226(.DIN1 (inData[31]), .DIN2 (_____9__26625), .Q
       (_________31648));
  and2s1 ____09_507227(.DIN1 (___9_9__26891), .DIN2 (_________33172),
       .Q (___0__9__30661));
  nnd2s1 ____09_507228(.DIN1 (____9___27296), .DIN2 (____9___27295), .Q
       (____0___27655));
  or2s1 ____09_507229(.DIN1 (________26383), .DIN2 (___0_____30866), .Q
       (___9____27797));
  nnd2s1 ____09_507230(.DIN1 (____9___27294), .DIN2 (___9____26896), .Q
       (________29039));
  nnd2s1 _____507231(.DIN1 (____9___27293), .DIN2 (___0____27858), .Q
       (________28043));
  nor2s1 _____0_507232(.DIN1 (________26753), .DIN2 (____9___27292), .Q
       (____00__27654));
  nor2s1 _____0_507233(.DIN1 (________27072), .DIN2 (____9___27291), .Q
       (_____9__27949));
  or2s1 _______507234(.DIN1 (___0____28758), .DIN2 (____90__27290), .Q
       (________28003));
  nnd2s1 ____0__507235(.DIN1 (________26837), .DIN2 (________28230), .Q
       (________28053));
  xor2s1 _______507236(.DIN1 (________22512), .DIN2 (_________36856),
       .Q (____0___28116));
  nnd2s1 ______507237(.DIN1 (____0_0__37159), .DIN2 (________22927), .Q
       (________27617));
  nnd2s1 ____0__507238(.DIN1 (__99____30480), .DIN2 (___0_____30676),
       .Q (___9____27780));
  nnd2s1 _______507239(.DIN1 (________27690), .DIN2 (_____9__27289), .Q
       (___9____27802));
  and2s1 _______507240(.DIN1 (___9____26893), .DIN2 (______0__31921),
       .Q (________28133));
  xor2s1 ____0__507241(.DIN1 (________26541), .DIN2 (___0____24250), .Q
       (________27603));
  nor2s1 ______507242(.DIN1 (_____9__27269), .DIN2 (___0____27878), .Q
       (________27606));
  nnd2s1 _______507243(.DIN1 (___0_____31297), .DIN2 (____9____32422),
       .Q (________27607));
  nnd2s1 ____0__507244(.DIN1 (________26723), .DIN2 (inData[21]), .Q
       (___09___27913));
  nnd2s1 _______507245(.DIN1 (_____0__27280), .DIN2 (________26702), .Q
       (________27945));
  nnd2s1 _______507246(.DIN1 (_____9__26856), .DIN2 (________27288), .Q
       (____00__28471));
  nnd2s1 ______507247(.DIN1 (______0__32205), .DIN2 (____00__27922), .Q
       (__9__0__30120));
  and2s1 _______507248(.DIN1 (________27287), .DIN2 (__9__0__29966), .Q
       (___9____28722));
  nor2s1 ______507249(.DIN1 (inData[16]), .DIN2 (___0900), .Q
       (___0____27910));
  nnd2s1 _______507250(.DIN1 (________26723), .DIN2 (inData[16]), .Q
       (___090__27912));
  nnd2s1 _______507251(.DIN1 (________27311), .DIN2 (________28543), .Q
       (________28060));
  or2s1 _______507252(.DIN1 (_____________________21745), .DIN2
       (____0___26781), .Q (____09__28022));
  nnd2s1 ______507253(.DIN1 (________26299), .DIN2 (___9____29578), .Q
       (____0____32532));
  nnd2s1 _______507254(.DIN1 (________27286), .DIN2 (___0_____30979),
       .Q (___0_____31191));
  nnd2s1 _______507255(.DIN1 (__9_____30423), .DIN2 (___9____26928), .Q
       (______9__32615));
  nor2s1 _____9_507256(.DIN1 (___9____23207), .DIN2 (____0___26778), .Q
       (____9____33397));
  nnd2s1 _______507257(.DIN1 (________26299), .DIN2 (___9____26878), .Q
       (_________32898));
  nnd2s1 _______507258(.DIN1 (________27285), .DIN2 (_____0___41313),
       .Q (________28077));
  nor2s1 ______507259(.DIN1 (________26805), .DIN2 (________27284), .Q
       (________28066));
  nor2s1 _______507260(.DIN1 (_____0__27260), .DIN2 (___00___28744), .Q
       (____0___28020));
  nnd2s1 _______507261(.DIN1 (________27311), .DIN2 (________28982), .Q
       (___09___27914));
  or2s1 _______507262(.DIN1 (___9____27809), .DIN2 (________26843), .Q
       (________29415));
  dffacs1 _____________________________________9_(.CLRB (reset), .CLK
       (clk), .DIN (________26827), .Q (______9__22017));
  nnd2s1 _______507263(.DIN1 (________27283), .DIN2 (________27975), .Q
       (____9_0__33415));
  dffacs1 _______________________________________________507264(.CLRB
       (reset), .CLK (clk), .DIN (____0___26777), .Q
       (_____________________________________________21896));
  nnd2s1 ______507265(.DIN1 (__9__0__29966), .DIN2 (_________31811), .Q
       (__9_9___29892));
  nnd2s1 _______507266(.DIN1 (_____0__28530), .DIN2 (________27282), .Q
       (__9_0___29904));
  nor2s1 _______507267(.DIN1 (_________41271), .DIN2 (________27720),
       .Q (_____0__29495));
  hi1s1 _______507268(.DIN (________27281), .Q (__9_____29845));
  hi1s1 ______507269(.DIN (____0___29372), .Q (__9_____29957));
  hi1s1 ______507270(.DIN (__9_____29862), .Q (__9_____30255));
  xor2s1 ____0__507271(.DIN1 (________26540), .DIN2 (_________38271),
       .Q (________28140));
  dffacs1 _____________________________________0_507272(.CLRB (reset),
       .CLK (clk), .DIN (________26808), .Q (__________0_));
  dffacs1 _________________________________________0___0_(.CLRB
       (reset), .CLK (clk), .DIN (___9____26887), .Q
       (_____________________________________0___0_));
  dffacs1 ______________________________________507273(.CLRB (reset),
       .CLK (clk), .DIN (________26818), .Q (___0_____40589));
  nnd2s1 _______507274(.DIN1 (________26854), .DIN2 (________25656), .Q
       (_________32241));
  hi1s1 _______507275(.DIN (_____9__29314), .Q (________29119));
  hi1s1 _______507276(.DIN (________27172), .Q (________27993));
  nnd2s1 _______507277(.DIN1 (_____0__27280), .DIN2 (___90___26865), .Q
       (__90____29665));
  hi1s1 _______507278(.DIN (____9___29551), .Q (____0___29104));
  hi1s1 _______507279(.DIN (__9__0__30291), .Q (__90____29661));
  nor2s1 _____9_507280(.DIN1 (________26643), .DIN2 (____9___26767), .Q
       (___0_9___40354));
  dffacs2 _________________507281(.CLRB (reset), .CLK (clk), .DIN
       (_____9__26654), .Q (______________22068));
  nnd2s1 _____507282(.DIN1 (_____9__26664), .DIN2 (inData[8]), .Q
       (_____9__27279));
  and2s1 _____0_507283(.DIN1 (__9_9___30174), .DIN2 (________27277), .Q
       (________27278));
  or2s1 _____0_507284(.DIN1 (________26762), .DIN2 (________27674), .Q
       (________27276));
  and2s1 _____0_507285(.DIN1 (________27274), .DIN2 (___90___28651), .Q
       (________27275));
  and2s1 ______507286(.DIN1 (_____0__28181), .DIN2 (_____0__28530), .Q
       (________27273));
  nor2s1 _______507287(.DIN1 (________27242), .DIN2 (_____9__26473), .Q
       (________27272));
  or2s1 _______507288(.DIN1 (_____0__27270), .DIN2 (_____9__27269), .Q
       (________27271));
  and2s1 _______507289(.DIN1 (________27322), .DIN2 (___9____26923), .Q
       (________27268));
  and2s1 ______507290(.DIN1 (________26641), .DIN2 (___090___31415), .Q
       (________27267));
  or2s1 _______507291(.DIN1 (__9_____30098), .DIN2 (________27265), .Q
       (________27266));
  nnd2s1 ______507292(.DIN1 (_____9__27084), .DIN2 (________26796), .Q
       (________27264));
  nnd2s1 _______507293(.DIN1 (________26628), .DIN2 (________26335), .Q
       (________27263));
  nor2s1 _______507294(.DIN1 (________27261), .DIN2 (_____0__27260), .Q
       (________27262));
  nor2s1 _______507295(.DIN1 (________28860), .DIN2 (________26828), .Q
       (________27259));
  or2s1 ______507296(.DIN1 (________28344), .DIN2 (_________41273), .Q
       (________27258));
  nnd2s1 _______507297(.DIN1 (________27256), .DIN2 (____0___26683), .Q
       (________27257));
  or2s1 _______507298(.DIN1 (________27246), .DIN2 (________27458), .Q
       (________27255));
  or2s1 _______507299(.DIN1 (__9_____30016), .DIN2 (________26815), .Q
       (________27254));
  nor2s1 _______507300(.DIN1 (____9___27475), .DIN2 (______0__41250),
       .Q (________27253));
  and2s1 _______507301(.DIN1 (_____0__27251), .DIN2 (_____0__26832), .Q
       (________27252));
  nnd2s1 _______507302(.DIN1 (____9___26858), .DIN2 (___0_____31391),
       .Q (_____9__27250));
  nnd2s1 _______507303(.DIN1 (__9_9___30174), .DIN2 (________27248), .Q
       (________27249));
  nor2s1 _______507304(.DIN1 (________27246), .DIN2 (______9__32117),
       .Q (________27247));
  and2s1 _____9_507305(.DIN1 (___9____26876), .DIN2 (_________32811),
       .Q (________27245));
  or2s1 _____507306(.DIN1 (________27243), .DIN2 (________27242), .Q
       (________27244));
  nnd2s1 _____0_507307(.DIN1 (________26786), .DIN2 (___9____26912), .Q
       (_____0__27241));
  nnd2s1 _____0_507308(.DIN1 (____9___26675), .DIN2 (________29112), .Q
       (_____9__27240));
  and2s1 _____0_507309(.DIN1 (____9___26681), .DIN2 (________27694), .Q
       (________27239));
  nor2s1 _____0_507310(.DIN1 (____0___26685), .DIN2 (__90____29692), .Q
       (________27238));
  and2s1 _____0_507311(.DIN1 (________27236), .DIN2 (________27235), .Q
       (________27237));
  or2s1 _____507312(.DIN1 (________25802), .DIN2 (___0_____30866), .Q
       (________27234));
  nnd2s1 _______507313(.DIN1 (__9_9___30174), .DIN2 (________29149), .Q
       (________27233));
  nor2s1 _______507314(.DIN1 (____9___27298), .DIN2 (_____0__26665), .Q
       (________27232));
  nor2s1 _______507315(.DIN1 (_________41297), .DIN2 (_________41234),
       .Q (_____0__27231));
  and2s1 _______507316(.DIN1 (__9_____30423), .DIN2 (________27229), .Q
       (________27230));
  xor2s1 ______507317(.DIN1 (___0_____40526), .DIN2 (___9_0___39705),
       .Q (________27228));
  hi1s1 ____0__507318(.DIN (___0_9___31403), .Q (________27227));
  xor2s1 ____0_507319(.DIN1 (_________35727), .DIN2 (________26542), .Q
       (________27226));
  or2s1 _______507320(.DIN1 (________27320), .DIN2 (________27160), .Q
       (________27225));
  hi1s1 _______507321(.DIN (________27707), .Q (________27224));
  and2s1 _____0_507322(.DIN1 (____0____37165), .DIN2 (________24036),
       .Q (________27223));
  nor2s1 _____0_507323(.DIN1 (____0___26590), .DIN2 (________26715), .Q
       (________27219));
  or2s1 ______507324(.DIN1 (____0___29013), .DIN2 (________27217), .Q
       (________27218));
  or2s1 _______507325(.DIN1 (____09__27215), .DIN2 (________29236), .Q
       (_____0__27216));
  nor2s1 _______507326(.DIN1 (_____9__27452), .DIN2 (___9____27772), .Q
       (____0___27213));
  nor2s1 _______507327(.DIN1 (________26433), .DIN2 (___0____26993), .Q
       (____0___27212));
  nnd2s1 _______507328(.DIN1 (________26722), .DIN2 (________29208), .Q
       (____0___27211));
  hi1s1 ____0_507329(.DIN (___09____31469), .Q (____0___27210));
  hi1s1 ____0__507330(.DIN (________29229), .Q (____0___27209));
  hi1s1 _____0_507331(.DIN (____0___27658), .Q (____9___27207));
  or2s1 _____507332(.DIN1 (________26287), .DIN2 (________27265), .Q
       (____9___27206));
  hi1s1 ____0__507333(.DIN (_________41226), .Q (____9___27205));
  nnd2s1 ______507334(.DIN1 (_____0__27186), .DIN2 (___9____25979), .Q
       (________27202));
  nnd2s1 _______507335(.DIN1 (________26699), .DIN2 (inData[18]), .Q
       (________27201));
  or2s1 _______507336(.DIN1 (_____0__26266), .DIN2 (________27199), .Q
       (________27200));
  or2s1 _______507337(.DIN1 (________25333), .DIN2 (________27221), .Q
       (________27198));
  nnd2s1 _______507338(.DIN1 (___9____26884), .DIN2 (________28887), .Q
       (________27197));
  or2s1 _____507339(.DIN1 (___0__0__31061), .DIN2 (________26709), .Q
       (_____0__27196));
  nor2s1 _____9_507340(.DIN1 (__________________0___21750), .DIN2
       (____9____32422), .Q (_____9__27195));
  nor2s1 _______507341(.DIN1 (_____________________21745), .DIN2
       (___9____26894), .Q (________27194));
  nor2s1 _______507342(.DIN1 (________27616), .DIN2 (________27192), .Q
       (________27193));
  nor2s1 _______507343(.DIN1 (________27190), .DIN2 (_________33664),
       .Q (________27191));
  nor2s1 _______507344(.DIN1 (____0___25313), .DIN2 (____9___26679), .Q
       (________27189));
  nnd2s1 _______507345(.DIN1 (________26648), .DIN2 (____0___25681), .Q
       (________27188));
  nnd2s1 _______507346(.DIN1 (_____0__27186), .DIN2 (_____9__27185), .Q
       (________27187));
  or2s1 _____9_507347(.DIN1 (________27183), .DIN2 (___9____26902), .Q
       (________27184));
  nnd2s1 _____0_507348(.DIN1 (________26712), .DIN2 (________23739), .Q
       (________27182));
  and2s1 _______507349(.DIN1 (________26299), .DIN2 (___0_9__27008), .Q
       (___09___27919));
  nnd2s1 _______507350(.DIN1 (___0_____31266), .DIN2 (_________32296),
       .Q (________27592));
  or2s1 _______507351(.DIN1 (________27181), .DIN2 (________26658), .Q
       (___9____27775));
  nnd2s1 _______507352(.DIN1 (________28242), .DIN2 (________25599), .Q
       (___9____27799));
  nor2s1 _______507353(.DIN1 (___0____27006), .DIN2 (_________31870),
       .Q (________27591));
  nor2s1 _______507354(.DIN1 (____9____32449), .DIN2 (_________31809),
       .Q (________27589));
  and2s1 _______507355(.DIN1 (___9____27778), .DIN2 (________27180), .Q
       (________27972));
  nnd2s1 _______507356(.DIN1 (________27538), .DIN2 (__99____30513), .Q
       (________27587));
  nor2s1 _______507357(.DIN1 (___0_____31198), .DIN2 (_____0__26636),
       .Q (___9_0__27777));
  and2s1 _______507358(.DIN1 (___0_____31096), .DIN2 (________27179),
       .Q (________29393));
  hi1s1 ____0__507359(.DIN (____9___27477), .Q (____0___28474));
  or2s1 ______507360(.DIN1 (_________41271), .DIN2 (________28160), .Q
       (________27970));
  hi1s1 ____0_507361(.DIN (________27178), .Q (___9____27792));
  nor2s1 _______507362(.DIN1 (__9_____29766), .DIN2 (______9__32117),
       .Q (____9___27473));
  nnd2s1 _______507363(.DIN1 (_____9__26700), .DIN2 (_____0__27177), .Q
       (________27955));
  nnd2s1 _______507364(.DIN1 (________26633), .DIN2 (____9_9__32410),
       .Q (___0____27880));
  nnd2s1 _______507365(.DIN1 (________28543), .DIN2 (________28281), .Q
       (_____0__27585));
  nnd2s1 _____9_507366(.DIN1 (________26841), .DIN2 (___0____27014), .Q
       (__9_9___30360));
  nor2s1 _____9_507367(.DIN1 (_________32071), .DIN2 (________26669),
       .Q (________27584));
  nor2s1 _____9_507368(.DIN1 (_____9__27176), .DIN2 (________26650), .Q
       (___9____29600));
  hi1s1 _______507369(.DIN (________27175), .Q (___9____27769));
  nnd2s1 _____9_507370(.DIN1 (________27180), .DIN2 (___9____26899), .Q
       (____0___28111));
  nor2s1 _____507371(.DIN1 (________26634), .DIN2 (______0__32351), .Q
       (_____0__27978));
  nnd2s1 _____0_507372(.DIN1 (________26652), .DIN2 (________29181), .Q
       (_____9__28636));
  hi1s1 ____0_507373(.DIN (________27174), .Q (________27985));
  hi1s1 _____0_507374(.DIN (________27173), .Q (___9____27765));
  nnd2s1 ______507375(.DIN1 (___9____26877), .DIN2 (___9_0__27768), .Q
       (________28125));
  nnd2s1 _______507376(.DIN1 (____0___29010), .DIN2 (________29033), .Q
       (___0____27896));
  and2s1 ______507377(.DIN1 (___0__9__31260), .DIN2 (____00__27922), .Q
       (___9____27791));
  nor2s1 _______507378(.DIN1 (_____________________21745), .DIN2
       (____9___26674), .Q (________28089));
  nor2s1 _______507379(.DIN1 (________27171), .DIN2 (________26851), .Q
       (___0____27885));
  hi1s1 _______507380(.DIN (________27149), .Q (_____9__27471));
  hi1s1 _______507381(.DIN (________27170), .Q (___0__9__31050));
  or2s1 ______507382(.DIN1 (____9___27389), .DIN2 (______9__33267), .Q
       (________27935));
  nor2s1 _______507383(.DIN1 (____00__22450), .DIN2 (____0___27394), .Q
       (________27937));
  nor2s1 _______507384(.DIN1 (_____9__27452), .DIN2 (________26754), .Q
       (____9___27476));
  nor2s1 _______507385(.DIN1 (________27169), .DIN2 (_____9__26708), .Q
       (____0___27486));
  nor2s1 ______507386(.DIN1 (________27220), .DIN2 (________27217), .Q
       (____0___27485));
  nor2s1 _____0_507387(.DIN1 (________28441), .DIN2 (________29115), .Q
       (________27501));
  nor2s1 _____9_507388(.DIN1 (________27164), .DIN2 (________28153), .Q
       (________27500));
  nnd2s1 _______507389(.DIN1 (________26711), .DIN2 (________29384), .Q
       (___9_9__27785));
  nor2s1 _______507390(.DIN1 (_________34207), .DIN2 (________28216),
       .Q (___9____27787));
  nnd2s1 _______507391(.DIN1 (________27168), .DIN2 (_____0__27167), .Q
       (___9_9__27813));
  and2s1 _______507392(.DIN1 (__9__0__29878), .DIN2 (_____0__29175), .Q
       (___0____27843));
  nor2s1 ______507393(.DIN1 (_____9___41301), .DIN2 (_____9__27166), .Q
       (__90____29657));
  nnd2s1 _____0_507394(.DIN1 (____9___28198), .DIN2 (_________41242),
       .Q (_________32750));
  nnd2s1 ______507395(.DIN1 (_________36521), .DIN2 (___90___26870), .Q
       (_________36621));
  dffacs1 ________________________________________________507396(.CLRB
       (reset), .CLK (clk), .DIN (___9____26889), .QN
       (_________________________________________________________________21991));
  or2s1 _______507397(.DIN1 (________27162), .DIN2 (___0_____40284), .Q
       (___0_____40294));
  nor2s1 _______507398(.DIN1 (____0___29013), .DIN2 (_____9__27166), .Q
       (__9__9__30056));
  or2s1 _______507399(.DIN1 (________28149), .DIN2 (________29149), .Q
       (____0___28380));
  nor2s1 ____9__507400(.DIN1 (___00____30625), .DIN2 (____9____32434),
       .Q (______0__31815));
  nor2s1 ____9__507401(.DIN1 (___9_9__25996), .DIN2 (________27192), .Q
       (__9__0__30196));
  nor2s1 ____9__507402(.DIN1 (________27165), .DIN2 (________27164), .Q
       (____9___29367));
  nnd2s1 ____9_507403(.DIN1 (________26619), .DIN2 (________27163), .Q
       (________29264));
  nnd2s1 _______507404(.DIN1 (__9_9___30174), .DIN2 (___9____29608), .Q
       (______9__32998));
  nnd2s1 ____0__507405(.DIN1 (_____0__27148), .DIN2 (________26707), .Q
       (____90__27472));
  nnd2s1 _______507406(.DIN1 (____9___27296), .DIN2 (________25570), .Q
       (_____0__27941));
  nnd2s1 _______507407(.DIN1 (__99____30533), .DIN2 (_____0__28530), .Q
       (________28874));
  or2s1 ______507408(.DIN1 (____9___26586), .DIN2 (________27458), .Q
       (____9___29093));
  dffacs1 _____________________________________________0_507409(.CLRB
       (reset), .CLK (clk), .DIN (________26798), .Q
       (_________________________________________0___21895));
  dffacs1 ________________________________________________507410(.CLRB
       (reset), .CLK (clk), .DIN (________26849), .Q (_________22023));
  nnd2s1 ______507411(.DIN1 (__9_9___30174), .DIN2 (___0____27015), .Q
       (____0____32499));
  hi1s1 _______507412(.DIN (________27513), .Q (___9____27806));
  nnd2s1 _______507413(.DIN1 (____9___26405), .DIN2 (________27162), .Q
       (___0_0___40281));
  or2s1 ______507414(.DIN1 (____0_0__31523), .DIN2 (________27160), .Q
       (___009__27835));
  hi1s1 ____0__507415(.DIN (____00___31511), .Q (___9____27788));
  nor2s1 _______507416(.DIN1 (_________41268), .DIN2 (____9___27292),
       .Q (_____0__28608));
  or2s1 _______507417(.DIN1 (___0_____31381), .DIN2 (________27164), .Q
       (___9____29580));
  and2s1 _______507418(.DIN1 (________26299), .DIN2 (_________31673),
       .Q (_________32746));
  and2s1 _______507419(.DIN1 (________27159), .DIN2 (________27526), .Q
       (___0____27847));
  nor2s1 ______507420(.DIN1 (___0_____31282), .DIN2 (________27217), .Q
       (___0____27892));
  and2s1 _______507421(.DIN1 (________26694), .DIN2 (____9___28920), .Q
       (___9____28696));
  nnd2s1 _______507422(.DIN1 (_________36521), .DIN2 (___90___26871),
       .Q (____0___28016));
  nor2s1 _______507423(.DIN1 (________27158), .DIN2 (_________31870),
       .Q (___9____27781));
  nor2s1 _______507424(.DIN1 (________28866), .DIN2 (________28879), .Q
       (________27960));
  nnd2s1 ______507425(.DIN1 (____09___31595), .DIN2 (________25941), .Q
       (___0_00__30642));
  nor2s1 _______507426(.DIN1 (________29149), .DIN2 (__90____29692), .Q
       (___9____27779));
  nnd2s1 _______507427(.DIN1 (______9__31688), .DIN2 (___0_____31385),
       .Q (__9_____29745));
  or2s1 _______507428(.DIN1 (________29529), .DIN2 (_____0__26718), .Q
       (______0__32214));
  or2s1 _______507429(.DIN1 (__9_00__29993), .DIN2 (______9__32117), .Q
       (____99__28013));
  and2s1 ______507430(.DIN1 (_____9___31891), .DIN2 (_____0__27157), .Q
       (____9___29002));
  nor2s1 _______507431(.DIN1 (___0____28779), .DIN2 (___0900), .Q
       (_____9___33329));
  and2s1 _______507432(.DIN1 (___0__9__31280), .DIN2 (___0_____31237),
       .Q (___0_____30771));
  nnd2s1 ______507433(.DIN1 (____0___29010), .DIN2 (________26696), .Q
       (________29508));
  or2s1 _______507434(.DIN1 (______9__37555), .DIN2 (________27402), .Q
       (______9__37652));
  nor2s1 _______507435(.DIN1 (_________33123), .DIN2 (______0__41250),
       .Q (________28605));
  nnd2s1 _______507436(.DIN1 (__9_____29775), .DIN2 (________28364), .Q
       (_________32602));
  nor2s1 _______507437(.DIN1 (_________41262), .DIN2 (________28344),
       .Q (________28585));
  dffacs1 _______________________________________507438(.CLRB (reset),
       .CLK (clk), .DIN (________26846), .Q (______________22108));
  nnd2s1 _______507439(.DIN1 (________27156), .DIN2 (________27155), .Q
       (__9_____30260));
  dffacs1 _____________________________________9_507440(.CLRB (reset),
       .CLK (clk), .DIN (________26833), .Q (__________9___22107));
  nnd2s1 _______507441(.DIN1 (__9_9___30451), .DIN2 (_________32022),
       .Q (___09____31480));
  dffacs1 _________________________________________0_____507442(.CLRB
       (reset), .CLK (clk), .DIN (___9_0__26892), .Q (___0_____40576));
  nor2s1 ______507443(.DIN1 (____9___26680), .DIN2 (____99__27391), .Q
       (__9_9___30267));
  nor2s1 ______507444(.DIN1 (________27154), .DIN2 (____9___28010), .Q
       (________28320));
  dffacs1 _______________________________________________507445(.CLRB
       (reset), .CLK (clk), .DIN (________26797), .Q
       (_____________________________________________21899));
  dffacs1 _______________________________________507446(.CLRB (reset),
       .CLK (clk), .DIN (____9___26769), .Q (______________22110));
  nor2s1 _____9_507447(.DIN1 (________27150), .DIN2 (_____9__26644), .Q
       (_________33650));
  hi1s1 _______507448(.DIN (___0____28820), .Q (________28592));
  hi1s1 _______507449(.DIN (__9_____30401), .Q (____09__29106));
  hi1s1 _______507450(.DIN (________27151), .Q (__9_____29827));
  hi1s1 ______507451(.DIN (________27153), .Q (__9_9___30270));
  nnd2s1 ____0__507452(.DIN1 (_____0__27148), .DIN2 (________26705), .Q
       (__9_____30019));
  hi1s1 _______507453(.DIN (________27152), .Q (___0_0__27855));
  hi1s1 _______507454(.DIN (____0___29200), .Q (_____9__29295));
  hi1s1 ______507455(.DIN (__999___30539), .Q (________29537));
  hi1s1 ______507456(.DIN (________27544), .Q (________29361));
  hi1s1 ______507457(.DIN (__9__9__29935), .Q (__9990));
  nnd2s1 _____9_507458(.DIN1 (________26567), .DIN2 (_____0__24373), .Q
       (_____9__27147));
  hi1s1 ____0__507459(.DIN (____9___28010), .Q (________27146));
  nnd2s1 _____507460(.DIN1 (________26569), .DIN2 (________24591), .Q
       (________27145));
  xor2s1 _____507461(.DIN1 (___________________), .DIN2
       (___0_____30709), .Q (________27144));
  nor2s1 _______507462(.DIN1 (________26252), .DIN2 (_____9__26389), .Q
       (________27143));
  nor2s1 _______507463(.DIN1 (________26436), .DIN2 (________27141), .Q
       (________27142));
  nor2s1 _______507464(.DIN1 (____99__26682), .DIN2 (____9___27117), .Q
       (________27140));
  or2s1 _______507465(.DIN1 (_____9__27138), .DIN2 (________27248), .Q
       (_____0__27139));
  nnd2s1 _______507466(.DIN1 (________26477), .DIN2 (inData[16]), .Q
       (________27137));
  nnd2s1 _______507467(.DIN1 (____9___26493), .DIN2 (inData[4]), .Q
       (________27136));
  nnd2s1 _______507468(.DIN1 (________26534), .DIN2 (____9___28922), .Q
       (________27135));
  nnd2s1 _______507469(.DIN1 (_____0__26538), .DIN2
       (_____________________________________________21940), .Q
       (________27134));
  nor2s1 _______507470(.DIN1
       (_____________________________________________21799), .DIN2
       (________26463), .Q (________27133));
  nor2s1 ______507471(.DIN1 (________23676), .DIN2 (___0_____40188), .Q
       (________27132));
  nor2s1 _____507472(.DIN1 (________28859), .DIN2 (________26533), .Q
       (________27131));
  or2s1 ____90_507473(.DIN1 (____0___27484), .DIN2 (____9___26318), .Q
       (________27130));
  nor2s1 ____9__507474(.DIN1 (____09__27128), .DIN2 (________26350), .Q
       (_____0__27129));
  nnd2s1 ____9__507475(.DIN1 (________26487), .DIN2 (________25813), .Q
       (____0___27127));
  nnd2s1 ____9__507476(.DIN1 (________26513), .DIN2 (_____0__24915), .Q
       (____0___27126));
  nor2s1 ____9__507477(.DIN1 (____0___25864), .DIN2 (________26512), .Q
       (____0___27125));
  nnd2s1 ____9__507478(.DIN1 (____9___26496), .DIN2 (inData[12]), .Q
       (____0___27124));
  nor2s1 ____9_507479(.DIN1 (_________41283), .DIN2 (____0___27122), .Q
       (____0___27123));
  nnd2s1 ____9__507480(.DIN1 (________26511), .DIN2 (inData[26]), .Q
       (____0___27121));
  nor2s1 ____9__507481(.DIN1 (___0____26090), .DIN2 (________26807), .Q
       (____9___27120));
  nor2s1 ____9__507482(.DIN1 (____9___27118), .DIN2 (____9___27117), .Q
       (____9___27119));
  nnd2s1 ____0__507483(.DIN1 (_____0__26474), .DIN2 (_____9__24059), .Q
       (____9___27116));
  nor2s1 ____0__507484(.DIN1 (________28026), .DIN2 (_____9___41301),
       .Q (____9___27115));
  or2s1 ____0_507485(.DIN1 (_________33123), .DIN2 (____9___27566), .Q
       (____9___27114));
  and2s1 _______507486(.DIN1 (________26572), .DIN2 (_____9__26255), .Q
       (____90__27113));
  nor2s1 ____0__507487(.DIN1 (___90), .DIN2 (___0_____40188), .Q
       (_____9__27112));
  nor2s1 ____0__507488(.DIN1 (________22500), .DIN2 (___0_____40188),
       .Q (________27111));
  nnd2s1 ____0__507489(.DIN1 (________26573), .DIN2 (___09___26137), .Q
       (________27110));
  nor2s1 ____0_507490(.DIN1 (___0____26064), .DIN2 (____0___26502), .Q
       (________27109));
  nnd2s1 ____0__507491(.DIN1 (_____9__26517), .DIN2 (_________36480),
       .Q (________27108));
  and2s1 ____0_507492(.DIN1 (___0_____30807), .DIN2 (__99____30513), .Q
       (________27107));
  nnd2s1 ____0__507493(.DIN1 (________26809), .DIN2 (________27105), .Q
       (________27106));
  nor2s1 ____0__507494(.DIN1 (______22163), .DIN2 (________27060), .Q
       (________27104));
  nor2s1 _______507495(.DIN1 (__9_____30208), .DIN2 (________27080), .Q
       (_____0__27103));
  or2s1 _______507496(.DIN1 (__9_____29750), .DIN2 (_________41271), .Q
       (_____9__27102));
  or2s1 _______507497(.DIN1 (________26396), .DIN2 (________26184), .Q
       (________27101));
  or2s1 _______507498(.DIN1
       (______________________________________0_______21890), .DIN2
       (________27099), .Q (________27100));
  nnd2s1 _______507499(.DIN1 (________26387), .DIN2 (___9_____39548),
       .Q (________27098));
  nor2s1 _______507500(.DIN1 (______9__32360), .DIN2 (________27082),
       .Q (________27097));
  nnd2s1 _______507501(.DIN1 (_____0__26276), .DIN2 (_____0__27363), .Q
       (________27096));
  nnd2s1 ______507502(.DIN1 (________26386), .DIN2 (________27094), .Q
       (________27095));
  nor2s1 _______507503(.DIN1 (___9____26926), .DIN2 (____9___26494), .Q
       (_____0__27093));
  or2s1 _______507504(.DIN1 (________25254), .DIN2 (_____0__26571), .Q
       (_____9__27092));
  nor2s1 _______507505(.DIN1 (___9____26938), .DIN2 (___0_9__26998), .Q
       (________27091));
  and2s1 _______507506(.DIN1 (________27089), .DIN2 (____9___25763), .Q
       (________27090));
  nnd2s1 _______507507(.DIN1 (____90__26400), .DIN2 (________27094), .Q
       (________27088));
  nnd2s1 _______507508(.DIN1 (____9___26401), .DIN2 (_________31933),
       .Q (________27087));
  nnd2s1 _______507509(.DIN1 (___9____26933), .DIN2
       (______________22066), .Q (________27086));
  and2s1 _____0_507510(.DIN1 (_____9__27084), .DIN2 (___0____26124), .Q
       (_____0__27085));
  or2s1 _______507511(.DIN1 (___0_____40479), .DIN2 (________27082), .Q
       (________27083));
  nor2s1 _______507512(.DIN1 (________27080), .DIN2 (________27079), .Q
       (________27081));
  and2s1 _______507513(.DIN1 (________27077), .DIN2 (________22369), .Q
       (________27078));
  nnd2s1 ______507514(.DIN1 (________26388), .DIN2 (inData[20]), .Q
       (________27076));
  or2s1 ______507515(.DIN1 (________27073), .DIN2 (________27072), .Q
       (________27074));
  nor2s1 ______507516(.DIN1
       (__________________________________________________________________21986),
       .DIN2 (________26552), .Q (________27070));
  hi1s1 _____507517(.DIN (________27068), .Q (________27069));
  or2s1 _______507518(.DIN1 (___________), .DIN2 (_____0__26363), .Q
       (_____0__27067));
  or2s1 _______507519(.DIN1 (___0_____30821), .DIN2 (________26375), .Q
       (_____9__27066));
  xor2s1 _______507520(.DIN1 (_________22016), .DIN2 (________27063),
       .Q (________27065));
  xnr2s1 ______507521(.DIN1 (_________22015), .DIN2 (________27063), .Q
       (________27064));
  nnd2s1 _______507522(.DIN1 (________26378), .DIN2 (________26257), .Q
       (________27062));
  nor2s1 _______507523(.DIN1 (________22759), .DIN2 (________27060), .Q
       (________27061));
  nor2s1 ______507524(.DIN1 (________27058), .DIN2 (________26479), .Q
       (________27059));
  nnd2s1 _______507525(.DIN1 (________26543), .DIN2 (_____9__27056), .Q
       (_____0__27057));
  nnd2s1 _______507526(.DIN1 (________27054), .DIN2 (________22409), .Q
       (________27055));
  nor2s1 _______507527(.DIN1 (_____9__22928), .DIN2 (________27052), .Q
       (________27053));
  or2s1 _____9_507528(.DIN1 (____0___26596), .DIN2 (_________32042), .Q
       (________27051));
  nor2s1 _______507529(.DIN1 (_________41271), .DIN2 (________27049),
       .Q (________27050));
  nor2s1 _______507530(.DIN1 (__9_____30400), .DIN2 (____9___26492), .Q
       (________27048));
  nnd2s1 _______507531(.DIN1 (________26544), .DIN2 (____09__23510), .Q
       (_____0__27047));
  nnd2s1 _______507532(.DIN1 (________27060), .DIN2 (_________37321),
       .Q (_____9__27046));
  nor2s1 _______507533(.DIN1 (________26347), .DIN2 (________26539), .Q
       (________27045));
  nnd2s1 ______507534(.DIN1 (________27052), .DIN2 (________27043), .Q
       (________27044));
  or2s1 _______507535(.DIN1 (________27040), .DIN2 (__9_____30432), .Q
       (________27041));
  or2s1 ______507536(.DIN1 (_________32065), .DIN2 (______0__31950), .Q
       (____09__27038));
  nnd2s1 _____9_507537(.DIN1 (____0___27036), .DIN2 (____0___26690), .Q
       (____0___27037));
  nor2s1 _______507538(.DIN1 (____9___27475), .DIN2 (_________33123),
       .Q (____0___27034));
  xor2s1 _______507539(.DIN1 (___0_____40536), .DIN2 (___0__9__40158),
       .Q (____0___27033));
  nnd2s1 _____9_507540(.DIN1 (_____0__26380), .DIN2 (_____9__23747), .Q
       (____0___27032));
  nnd2s1 _______507541(.DIN1 (________26480), .DIN2 (________26346), .Q
       (____00__27031));
  nnd2s1 _____9_507542(.DIN1 (_____0__26555), .DIN2 (________24612), .Q
       (___099__27030));
  or2s1 _____0_507543(.DIN1 (_________35587), .DIN2 (________26395), .Q
       (___09___27029));
  hi1s1 _____0_507544(.DIN (________28535), .Q (___09___27027));
  hi1s1 _____0_507545(.DIN (____9___27291), .Q (___090__27026));
  nnd2s1 _______507546(.DIN1 (____0___26327), .DIN2 (___0____25183), .Q
       (___0____27025));
  hi1s1 _____507547(.DIN (___0____27023), .Q (___0____27024));
  hi1s1 _____9_507548(.DIN (___0____27021), .Q (___0____27022));
  and2s1 ______507549(.DIN1 (__9_____30163), .DIN2 (________26391), .Q
       (___0____27020));
  hi1s1 ____0__507550(.DIN (____0___27573), .Q (___0____27019));
  nor2s1 _______507551(.DIN1 (____0____33496), .DIN2 (________26524),
       .Q (____0___27302));
  hi1s1 ____0_507552(.DIN (_________41246), .Q (___0____27849));
  nor2s1 _______507553(.DIN1 (_____0__26349), .DIN2 (___0_0__27018), .Q
       (________27170));
  nnd2s1 _______507554(.DIN1 (________26509), .DIN2 (___0____27842), .Q
       (________27341));
  hi1s1 _______507555(.DIN (______0__38770), .Q (_________36753));
  hi1s1 _______507556(.DIN (______9__31688), .Q (____0___27487));
  and2s1 _______507557(.DIN1 (___0____27889), .DIN2 (___0_9__27017), .Q
       (________28408));
  nnd2s1 ______507558(.DIN1 (________26468), .DIN2 (___0____27016), .Q
       (_____9__27222));
  nnd2s1 _______507559(.DIN1 (____0___26504), .DIN2 (__99____30516), .Q
       (___9____27754));
  nor2s1 ____0_507560(.DIN1 (_____90__41299), .DIN2 (_________41258),
       .Q (________27440));
  nnd2s1 _______507561(.DIN1 (_____9__26465), .DIN2 (________25544), .Q
       (______9__31910));
  nnd2s1 ____0__507562(.DIN1 (________26476), .DIN2 (___9____27773), .Q
       (__9_____29860));
  nor2s1 _______507563(.DIN1 (___9____26025), .DIN2 (________26471), .Q
       (________27604));
  nnd2s1 _______507564(.DIN1 (________26368), .DIN2 (____0___26147), .Q
       (________27509));
  dffacs2 __________________507565(.CLRB (reset), .CLK (clk), .DIN
       (________26460), .QN
       (__________________________________9__________));
  nnd2s1 _____9_507566(.DIN1 (___0____27005), .DIN2 (inData[28]), .Q
       (________27172));
  nor2s1 ____0__507567(.DIN1 (________27724), .DIN2 (___9____29615), .Q
       (________27439));
  nor2s1 _____0_507568(.DIN1 (___0____27015), .DIN2 (________28171), .Q
       (_____0__27610));
  nnd2s1 ______507569(.DIN1 (____0___26500), .DIN2 (___0____27014), .Q
       (__9_____30339));
  nnd2s1 ______507570(.DIN1 (___9____27763), .DIN2 (___090___31415), .Q
       (___9_0__28698));
  or2s1 _______507571(.DIN1 (___9_9__27776), .DIN2 (________26488), .Q
       (________27703));
  nnd2s1 ____9__507572(.DIN1 (________26549), .DIN2 (___0____27013), .Q
       (________27175));
  nor2s1 _______507573(.DIN1 (________28131), .DIN2 (________27608), .Q
       (________27707));
  nnd2s1 _______507574(.DIN1 (___0_____31162), .DIN2 (___0_____30917),
       .Q (________27664));
  hi1s1 _______507575(.DIN (__9__0__29966), .Q (___00____30605));
  or2s1 _______507576(.DIN1 (__9_____29742), .DIN2 (________27248), .Q
       (________28311));
  nnd2s1 _______507577(.DIN1 (________26724), .DIN2 (__9_____30162), .Q
       (____0___28112));
  nnd2s1 _____0_507578(.DIN1 (___0_____31006), .DIN2 (___9____26947),
       .Q (________27982));
  and2s1 _______507579(.DIN1 (____0___27483), .DIN2 (___0____27012), .Q
       (____99__28107));
  hi1s1 _______507580(.DIN (___0____27011), .Q (__9_____30380));
  hi1s1 _______507581(.DIN (___0____27010), .Q (_________33778));
  or2s1 ______507582(.DIN1 (____09__28931), .DIN2 (_____9__29174), .Q
       (________27721));
  nor2s1 _______507583(.DIN1 (________27040), .DIN2 (________26464), .Q
       (___0_____30793));
  nor2s1 _______507584(.DIN1 (___0_0__27009), .DIN2 (___0__9__30890),
       .Q (___09___27918));
  nor2s1 ______507585(.DIN1 (________28859), .DIN2 (________26529), .Q
       (__99____30514));
  or2s1 _______507586(.DIN1 (___0_9__27008), .DIN2 (__9_____30432), .Q
       (__9__0__29824));
  and2s1 _______507587(.DIN1 (___0_____30903), .DIN2 (___0__0__31168),
       .Q (___0_____31362));
  nor2s1 _______507588(.DIN1 (__9__9__30419), .DIN2 (___0__9__30813),
       .Q (___0_____30888));
  nor2s1 _______507589(.DIN1 (_____9__26527), .DIN2 (____0___27924), .Q
       (___0_____31175));
  and2s1 _______507590(.DIN1 (___9____27764), .DIN2 (___9____27766), .Q
       (_________33931));
  nnd2s1 _______507591(.DIN1 (___0____27007), .DIN2 (________25821), .Q
       (________27704));
  hi1s1 ______507592(.DIN (_____9___38610), .Q (_________35622));
  or2s1 _______507593(.DIN1 (___00_0__30612), .DIN2 (________27248), .Q
       (________28225));
  nor2s1 _______507594(.DIN1 (________28026), .DIN2 (___0____27006), .Q
       (_____0__29213));
  nor2s1 _______507595(.DIN1 (____0___26591), .DIN2 (__909___29719), .Q
       (___0_____30805));
  nor2s1 _______507596(.DIN1 (inData[28]), .DIN2 (_____0__27280), .Q
       (____9___29551));
  nnd2s1 _______507597(.DIN1 (___0____27858), .DIN2 (________26364), .Q
       (________27681));
  nor2s1 _______507598(.DIN1 (_____0__29037), .DIN2 (___9____26937), .Q
       (_________31935));
  nnd2s1 _______507599(.DIN1 (_____9__26202), .DIN2 (________27287), .Q
       (___0__9__31347));
  hi1s1 _______507600(.DIN (___0____27004), .Q (________27991));
  nor2s1 ______507601(.DIN1 (_____0__26701), .DIN2 (___0____27005), .Q
       (___0____28820));
  nnd2s1 _____507602(.DIN1 (_________41254), .DIN2 (________26576), .Q
       (_________38155));
  nor2s1 _______507603(.DIN1 (_________35587), .DIN2 (_____0__27280),
       .Q (_____9__29314));
  dffacs1 _________________________________________0____507604(.CLRB
       (reset), .CLK (clk), .DIN (____0___26505), .Q
       (_____________________________________0______21756));
  nnd2s1 _____9_507605(.DIN1 (_____9__26489), .DIN2 (_____9__23482), .Q
       (_________36871));
  nor2s1 _____9_507606(.DIN1 (___9____24144), .DIN2 (____90__26490), .Q
       (_________38650));
  hi1s1 _______507607(.DIN (__9_____30423), .Q (__9_____29783));
  nnd2s1 _____9_507608(.DIN1 (___0____27005), .DIN2 (_________35587),
       .Q (__9_____29862));
  nor2s1 _____9_507609(.DIN1 (___900__26864), .DIN2 (___0____27005), .Q
       (____0___29372));
  hi1s1 ______507610(.DIN (___0_____31336), .Q (___0_0___30748));
  nb1s1 _______507611(.DIN (___0____27004), .Q (____0___29285));
  and2s1 _______507612(.DIN1 (________27077), .DIN2 (________24053), .Q
       (___0____27003));
  nor2s1 ______507613(.DIN1
       (__________________________________________9___21977), .DIN2
       (___0_____40284), .Q (___0____27002));
  and2s1 ______507614(.DIN1 (________26377), .DIN2 (_____9___37002), .Q
       (___0____27001));
  or2s1 _______507615(.DIN1 (___0_0__26999), .DIN2 (___0_9__26998), .Q
       (___0____27000));
  nnd2s1 _______507616(.DIN1 (___0____26996), .DIN2 (___0____26995), .Q
       (___0____26997));
  or2s1 _______507617(.DIN1 (________29170), .DIN2 (________26393), .Q
       (___0____26994));
  nnd2s1 ____9_507618(.DIN1 (________29498), .DIN2 (_________41281), .Q
       (___0____26992));
  nor2s1 _______507619(.DIN1 (_____9__24973), .DIN2 (________27060), .Q
       (___0_9__26991));
  nnd2s1 _______507620(.DIN1 (___0____26989), .DIN2 (________26693), .Q
       (___0____26990));
  nor2s1 _______507621(.DIN1 (_____9__26220), .DIN2 (________26398), .Q
       (___0____26988));
  nor2s1 _____0_507622(.DIN1 (________29049), .DIN2 (__9_0___29724), .Q
       (___0____26987));
  and2s1 ____0__507623(.DIN1 (________29090), .DIN2 (___0____26985), .Q
       (___0____26986));
  hi1s1 ____0__507624(.DIN (________29523), .Q (___0____26984));
  and2s1 _______507625(.DIN1 (___0____26982), .DIN2 (___0____26981), .Q
       (___0____26983));
  or2s1 _______507626(.DIN1 (___9____27800), .DIN2 (____9___27294), .Q
       (___0____26980));
  nor2s1 ______507627(.DIN1 (___0____26978), .DIN2 (____0___26326), .Q
       (___0____26979));
  or2s1 _______507628(.DIN1 (___0_00__30740), .DIN2 (___0__9__30890),
       .Q (___0____26977));
  and2s1 _______507629(.DIN1 (____9___27478), .DIN2 (________27495), .Q
       (___0_9__26976));
  nor2s1 _____0_507630(.DIN1 (____0___25593), .DIN2 (____0___26328), .Q
       (___0____26975));
  nnd2s1 _____507631(.DIN1 (__99____30516), .DIN2 (___9____26915), .Q
       (___0____26974));
  nor2s1 _____9_507632(.DIN1 (________26336), .DIN2 (________28046), .Q
       (___0____26973));
  nnd2s1 _____9_507633(.DIN1 (____9___26584), .DIN2
       (__________________0___21750), .Q (___0____26972));
  nnd2s1 _____9_507634(.DIN1 (____00__26323), .DIN2 (________28040), .Q
       (___0____26971));
  or2s1 _____507635(.DIN1 (______________22065), .DIN2 (________27082),
       .Q (___0____26970));
  nnd2s1 _______507636(.DIN1 (___0____26968), .DIN2 (___0____26106), .Q
       (___0____26969));
  or2s1 _______507637(.DIN1 (________26651), .DIN2 (___0_9__26966), .Q
       (___0_0__26967));
  nor2s1 ______507638(.DIN1 (___0____23299), .DIN2 (____90__26315), .Q
       (___0____26965));
  nor2s1 _______507639(.DIN1 (________26431), .DIN2 (____9___26319), .Q
       (___0____26964));
  nor2s1 _______507640(.DIN1 (________24989), .DIN2 (________26384), .Q
       (___0____26963));
  nor2s1 ______507641(.DIN1 (_____0__26617), .DIN2 (____9___27294), .Q
       (___0____26962));
  nnd2s1 ______507642(.DIN1 (________27446), .DIN2 (________28189), .Q
       (___0____26961));
  nnd2s1 _______507643(.DIN1 (________27099), .DIN2 (___9____24105), .Q
       (___009__26959));
  nnd2s1 _______507644(.DIN1 (____0___26592), .DIN2 (___9____27766), .Q
       (___00___26958));
  hi1s1 ____0__507645(.DIN (_________41244), .Q (___00___26955));
  hi1s1 ____0__507646(.DIN (_____0__27620), .Q (___00___26954));
  and2s1 _______507647(.DIN1 (___9____26931), .DIN2 (_____0__29417), .Q
       (___99___26953));
  nnd2s1 ______507648(.DIN1 (________26338), .DIN2 (________25878), .Q
       (___99___26952));
  nor2s1 _______507649(.DIN1 (________22598), .DIN2 (________27082), .Q
       (___99___26951));
  nor2s1 _______507650(.DIN1 (____0___22551), .DIN2 (________27082), .Q
       (___99___26950));
  and2s1 ______507651(.DIN1 (________27416), .DIN2 (_____0__26371), .Q
       (___990__26949));
  nor2s1 _______507652(.DIN1 (___9____26947), .DIN2 (____0____32539),
       .Q (___9_9__26948));
  or2s1 _______507653(.DIN1 (____0___29013), .DIN2 (__9__9__29743), .Q
       (___9____26946));
  nor2s1 ____507654(.DIN1 (_________32001), .DIN2 (___9____26944), .Q
       (___9____26945));
  or2s1 _______507655(.DIN1 (____00__29009), .DIN2 (____0____32521), .Q
       (___9____26943));
  nnd2s1 _____0_507656(.DIN1 (________26756), .DIN2 (________29231), .Q
       (___9____26941));
  nnd2s1 _______507657(.DIN1 (________26579), .DIN2 (___009___30634),
       .Q (________27281));
  or2s1 _______507658(.DIN1 (____9___27475), .DIN2 (___9____27762), .Q
       (___9____27793));
  hi1s1 ____0__507659(.DIN (_________31778), .Q (____0___27481));
  hi1s1 ____0_507660(.DIN (_____9__27344), .Q (_____0__27490));
  nor2s1 _______507661(.DIN1 (___9_0__26940), .DIN2 (__9_00__29993), .Q
       (_____9__27619));
  or2s1 ____0__507662(.DIN1 (inData[14]), .DIN2 (_____0__27148), .Q
       (________27149));
  or2s1 _______507663(.DIN1 (________27158), .DIN2 (_________41262), .Q
       (________27670));
  nor2s1 ______507664(.DIN1 (___9_9__26939), .DIN2 (___9____26938), .Q
       (____99__27208));
  nor2s1 _____9_507665(.DIN1 (_________33580), .DIN2 (________26521),
       .Q (________27614));
  and2s1 _______507666(.DIN1 (___0_____31156), .DIN2 (________25517),
       .Q (_____0___31895));
  and2s1 ______507667(.DIN1 (________27611), .DIN2 (______0__32196), .Q
       (_____0__29407));
  nor2s1 _____507668(.DIN1 (____00__27300), .DIN2 (________26385), .Q
       (____90__27647));
  nnd2s1 _____9_507669(.DIN1 (________26566), .DIN2 (___0__0__31290),
       .Q (_____0__27714));
  and2s1 ____90_507670(.DIN1 (__99____30473), .DIN2 (___0____27014), .Q
       (________27712));
  nnd2s1 ____9__507671(.DIN1 (________26361), .DIN2 (________24909), .Q
       (________27173));
  nor2s1 _______507672(.DIN1 (_____9__26304), .DIN2 (___9____26944), .Q
       (________27203));
  nnd2s1 _______507673(.DIN1 (________29090), .DIN2 (___9____26936), .Q
       (____0___27570));
  nor2s1 _______507674(.DIN1 (__9_____29766), .DIN2 (___9____26937), .Q
       (________27549));
  and2s1 ______507675(.DIN1 (____9___28550), .DIN2 (___0__9__30671), .Q
       (___0_____30968));
  and2s1 _______507676(.DIN1 (___9____26936), .DIN2 (___9____26935), .Q
       (________27518));
  nor2s1 _______507677(.DIN1 (________25707), .DIN2 (___9____26934), .Q
       (___99___28730));
  nor2s1 ______507678(.DIN1 (______________22066), .DIN2
       (___9____26933), .Q (____9___28466));
  nor2s1 _______507679(.DIN1 (_____0__26448), .DIN2 (________26510), .Q
       (____99__27479));
  or2s1 _______507680(.DIN1 (_____0___31803), .DIN2 (________26565), .Q
       (________27662));
  nnd2s1 _____9_507681(.DIN1 (_________31973), .DIN2 (_____9__26554),
       .Q (____9___27651));
  nnd2s1 _____507682(.DIN1 (________27256), .DIN2 (___9____26932), .Q
       (_____0__27723));
  nor2s1 _____507683(.DIN1 (__99____30485), .DIN2 (___09_9__31446), .Q
       (________27633));
  nnd2s1 _____0_507684(.DIN1 (________26372), .DIN2 (____9___27564), .Q
       (_____9__27204));
  nnd2s1 _____0_507685(.DIN1 (________26352), .DIN2 (___0_____30979),
       .Q (____0___28206));
  nnd2s1 _____0_507686(.DIN1 (___9____26931), .DIN2 (_____90__32080),
       .Q (___9____27755));
  nor2s1 _______507687(.DIN1 (____0___27576), .DIN2 (____00__29009), .Q
       (________27174));
  nnd2s1 ______507688(.DIN1 (____9___27478), .DIN2 (________27494), .Q
       (________27178));
  nnd2s1 _____9_507689(.DIN1 (________26519), .DIN2
       (_____________________21745), .Q (________27432));
  nor2s1 _______507690(.DIN1 (___9_0__26930), .DIN2 (___9_9__26929), .Q
       (________28001));
  nor2s1 ____9__507691(.DIN1 (___90___25959), .DIN2 (___9____26928), .Q
       (____0___28382));
  nor2s1 ____9__507692(.DIN1 (___9____26895), .DIN2 (___9____26928), .Q
       (__9__0__30130));
  nnd2s1 ____9__507693(.DIN1 (________26356), .DIN2 (__9_____29981), .Q
       (____0_0__32557));
  nor2s1 ____0_507694(.DIN1 (__99_9__30508), .DIN2 (_____0__27148), .Q
       (________27152));
  nor2s1 ____9_507695(.DIN1 (___9____26927), .DIN2 (______0__41270), .Q
       (________29079));
  nnd2s1 ____9__507696(.DIN1 (__9__0__29760), .DIN2 (___0____25150), .Q
       (____0___27658));
  nor2s1 ____9_507697(.DIN1 (________26483), .DIN2 (___9____26926), .Q
       (_________31655));
  nnd2s1 ____9__507698(.DIN1 (________27256), .DIN2 (___9____26925), .Q
       (____00__27480));
  nor2s1 _______507699(.DIN1 (___9____26924), .DIN2 (__9_0___30179), .Q
       (________28537));
  nnd2s1 ____0_507700(.DIN1 (___9____26909), .DIN2 (__99_9__30508), .Q
       (________27153));
  nor2s1 _______507701(.DIN1 (___00___26054), .DIN2 (_________41266),
       .Q (________28187));
  nnd2s1 _______507702(.DIN1 (____9___27478), .DIN2 (____0___26414), .Q
       (________27547));
  hi1s1 ____0__507703(.DIN (________27975), .Q (_________31817));
  nnd2s1 _______507704(.DIN1 (____9___27294), .DIN2 (___0____26066), .Q
       (_____9___31886));
  nor2s1 _______507705(.DIN1 (_____9__29174), .DIN2 (________29217), .Q
       (________27535));
  nnd2s1 ______507706(.DIN1 (________26556), .DIN2 (___09_9__31426), .Q
       (___0____27906));
  and2s1 _______507707(.DIN1 (_____0__26332), .DIN2
       (__________________0___21750), .Q (____9___27474));
  hi1s1 ____0__507708(.DIN (_____9__27166), .Q (___0____27853));
  or2s1 ______507709(.DIN1 (___9____26917), .DIN2 (__9_0___30179), .Q
       (________29269));
  nnd2s1 _______507710(.DIN1 (___9____26923), .DIN2 (___9____26922), .Q
       (_____0__27507));
  and2s1 _______507711(.DIN1 (________27235), .DIN2 (________27089), .Q
       (__9_____30349));
  nnd2s1 ______507712(.DIN1 (____0___26330), .DIN2 (________23726), .Q
       (________27640));
  nnd2s1 _______507713(.DIN1 (___9____26921), .DIN2 (____09__28480), .Q
       (__990___30461));
  or2s1 _______507714(.DIN1 (___9_0__26920), .DIN2 (____9_0__33356), .Q
       (________29500));
  or2s1 _______507715(.DIN1 (___09___27915), .DIN2 (___9_9__26919), .Q
       (________28541));
  nnd2s1 _______507716(.DIN1 (________27446), .DIN2 (_________31731),
       .Q (_________31843));
  nnd2s1 ____9__507717(.DIN1 (___9____27784), .DIN2 (_________41281),
       .Q (________27513));
  nnd2s1 ______507718(.DIN1 (________26339), .DIN2 (________29066), .Q
       (________27962));
  hi1s1 ____507719(.DIN (___9____26918), .Q (__9_____30222));
  or2s1 _______507720(.DIN1 (________25628), .DIN2 (_________32658), .Q
       (__9_____29883));
  nor2s1 ____507721(.DIN1 (___9____26917), .DIN2 (___9____26928), .Q
       (_____9__27636));
  nnd2s1 ______507722(.DIN1 (____9___25675), .DIN2 (___9____26916), .Q
       (________28337));
  nnd2s1 ____9__507723(.DIN1 (____9___26403), .DIN2 (___0_____31391),
       .Q (____9___29458));
  nor2s1 ____0__507724(.DIN1 (inData[23]), .DIN2 (________26486), .Q
       (________27151));
  and2s1 ____9__507725(.DIN1 (__9__0__29760), .DIN2 (___9____26915), .Q
       (__9_____30096));
  or2s1 _____507726(.DIN1 (____9___26581), .DIN2 (_____9__26370), .Q
       (_____9__28246));
  dffacs1 _______________________________________507727(.CLRB (reset),
       .CLK (clk), .DIN (________26467), .Q (___0_____40445));
  hi1s1 ____0__507728(.DIN (________28900), .Q (___0_____30764));
  nor2s1 _______507729(.DIN1 (___0_____30801), .DIN2 (___9____26914),
       .Q (____9___27477));
  nor2s1 _______507730(.DIN1 (_________31783), .DIN2 (_________31955),
       .Q (___0__9__30851));
  hi1s1 ____09_507731(.DIN (_________41248), .Q (_________35867));
  nor2s1 ______507732(.DIN1 (________25392), .DIN2 (___9____26913), .Q
       (____00___31511));
  and2s1 ____9_507733(.DIN1 (___0_____31040), .DIN2 (__9_____29818), .Q
       (___0_0___31119));
  or2s1 ____9__507734(.DIN1 (_________33609), .DIN2 (__9_9___30362), .Q
       (______0__32892));
  nor2s1 _____0_507735(.DIN1 (____99__25767), .DIN2 (________27504), .Q
       (___0_____31173));
  nnd2s1 _____0_507736(.DIN1 (____0___26329), .DIN2 (________25925), .Q
       (___0_9___31403));
  nor2s1 _____0_507737(.DIN1 (___9____26912), .DIN2 (________26313), .Q
       (________29229));
  nor2s1 _____0_507738(.DIN1 (________28441), .DIN2 (________26348), .Q
       (________28628));
  and2s1 _______507739(.DIN1 (_________31738), .DIN2 (___0_____30810),
       .Q (________29246));
  nnd2s1 _____507740(.DIN1 (____9___26320), .DIN2 (________26814), .Q
       (________28937));
  or2s1 _______507741(.DIN1 (___0____27868), .DIN2 (_________32815), .Q
       (____9___27560));
  nor2s1 _______507742(.DIN1 (________29326), .DIN2 (________28277), .Q
       (__9_____30322));
  nnd2s1 ______507743(.DIN1 (____0___27483), .DIN2 (___9_0__26911), .Q
       (__9_9___30449));
  or2s1 _______507744(.DIN1 (___09___27915), .DIN2 (___9_9__26910), .Q
       (________28936));
  nnd2s1 ____0__507745(.DIN1 (___9____26907), .DIN2 (inData[23]), .Q
       (________27544));
  nnd2s1 _______507746(.DIN1 (__99____30465), .DIN2 (_________32140),
       .Q (_____9___33059));
  nor2s1 _______507747(.DIN1 (____0___26412), .DIN2 (____00__29009), .Q
       (___0_____31078));
  nnd2s1 _______507748(.DIN1 (________26310), .DIN2 (____9___23782), .Q
       (________28154));
  nnd2s1 _______507749(.DIN1 (___9____26932), .DIN2 (___0_____30679),
       .Q (___0_____30760));
  dffacs1 _____________________________________0_507750(.CLRB (reset),
       .CLK (clk), .DIN (_____9__26570), .QN (___0_____40446));
  nor2s1 _______507751(.DIN1 (___0____27860), .DIN2 (__9__9__29743), .Q
       (___09____31469));
  nnd2s1 ____0__507752(.DIN1 (___9____26909), .DIN2 (inData[14]), .Q
       (____0___29200));
  dffacs1 ________________9_507753(.CLRB (reset), .CLK (clk), .DIN
       (________26522), .QN
       (_________________________________________________________________________________________22089));
  hi1s1 _______507754(.DIN (___9____26908), .Q (_________34141));
  hi1s1 ______507755(.DIN (__9_9___30174), .Q (__90____29663));
  nor2s1 ____0__507756(.DIN1 (________26610), .DIN2 (___9____26907), .Q
       (__9__9__29935));
  nor2s1 ____0_507757(.DIN1 (________26706), .DIN2 (___9____26909), .Q
       (__9__0__30291));
  nor2s1 ____0__507758(.DIN1 (________26704), .DIN2 (___9____26909), .Q
       (__9_____30401));
  nor2s1 ____0__507759(.DIN1 (________26485), .DIN2 (________26609), .Q
       (__999___30539));
  hi1s1 ____09_507760(.DIN (___9____26906), .Q (____9____33386));
  and2s1 _______507761(.DIN1 (___9____26904), .DIN2 (___9____26903), .Q
       (___9____26905));
  or2s1 ____0__507762(.DIN1 (_____0__25596), .DIN2 (___9_0__26901), .Q
       (___9____26902));
  hi1s1 ____0__507763(.DIN (___9____26898), .Q (___9____26899));
  nnd2s1 ______507764(.DIN1 (____0___27396), .DIN2 (________26729), .Q
       (___9____26897));
  nor2s1 ______507765(.DIN1 (___9____26895), .DIN2 (_____9__27138), .Q
       (___9____26896));
  nnd2s1 _______507766(.DIN1 (____99__26588), .DIN2 (________26601), .Q
       (___9____26894));
  nor2s1 ____9__507767(.DIN1 (___0_____31129), .DIN2 (___9____27789),
       .Q (___9____26893));
  or2s1 ____9__507768(.DIN1 (_____9___35559), .DIN2 (________26160), .Q
       (___9_0__26892));
  nor2s1 _______507769(.DIN1 (________24893), .DIN2 (___9____26890), .Q
       (___9_9__26891));
  or2s1 ____9_507770(.DIN1 (________26183), .DIN2 (_________37837), .Q
       (___9____26889));
  nor2s1 ____9__507771(.DIN1 (_______22238), .DIN2 (________26720), .Q
       (___9____26888));
  nnd2s1 ____507772(.DIN1 (_____0__26186), .DIN2 (________25906), .Q
       (___9____26887));
  nnd2s1 ____0__507773(.DIN1 (________27726), .DIN2 (____0___27035), .Q
       (___9____26886));
  nor2s1 _____0_507774(.DIN1 (________26301), .DIN2 (___9_0__26883), .Q
       (___9____26884));
  nor2s1 ______507775(.DIN1 (_________32663), .DIN2 (___0_____30709),
       .Q (___9_9__26882));
  nor2s1 _______507776(.DIN1 (________22537), .DIN2 (___0_____30709),
       .Q (___9____26881));
  nor2s1 _______507777(.DIN1 (___9____26879), .DIN2 (____0___26411), .Q
       (___9____26880));
  nnd2s1 _____9_507778(.DIN1 (_____9___31694), .DIN2 (________26736),
       .Q (___9____26878));
  nor2s1 _______507779(.DIN1 (____9___28196), .DIN2 (________26730), .Q
       (___9____26877));
  and2s1 _______507780(.DIN1 (_________32720), .DIN2 (__9_____30239),
       .Q (___9____26876));
  nor2s1 _______507781(.DIN1
       (__________________________________________________________________22002),
       .DIN2 (___90___28648), .Q (___9____26875));
  xnr2s1 _______507782(.DIN1
       (____________________________________________21772), .DIN2
       (_________37884), .Q (___9____26874));
  xor2s1 _______507783(.DIN1
       (____________________________________________21833), .DIN2
       (_____9___41303), .Q (___9_0__26873));
  xor2s1 ______507784(.DIN1 (________25914), .DIN2
       (_______________22070), .Q (___909__26872));
  hi1s1 ____0__507785(.DIN (___90___26870), .Q (___90___26871));
  nor2s1 ______507786(.DIN1 (____9___25759), .DIN2 (____9___27118), .Q
       (___90___26869));
  nnd2s1 _______507787(.DIN1 (___90___26867), .DIN2 (______22152), .Q
       (___90___26868));
  nor2s1 _______507788(.DIN1 (________27355), .DIN2 (________29431), .Q
       (___90___26866));
  hi1s1 ____0__507789(.DIN (___900__26864), .Q (___90___26865));
  nnd2s1 _______507790(.DIN1 (_____0__26482), .DIN2 (____9___26862), .Q
       (____99__26863));
  nnd2s1 _______507791(.DIN1 (_____0__26626), .DIN2 (________26281), .Q
       (____9___26861));
  nor2s1 _______507792(.DIN1 (__________22059), .DIN2 (____09___37180),
       .Q (____9___26860));
  nnd2s1 ______507793(.DIN1 (___0____26128), .DIN2 (________25381), .Q
       (____9___26859));
  nor2s1 _______507794(.DIN1 (___0_____30882), .DIN2 (_________41287),
       .Q (____9___26858));
  nnd2s1 _______507795(.DIN1 (_____0__26822), .DIN2
       (_____________________________________9_____), .Q
       (____90__26857));
  nor2s1 _____0_507796(.DIN1 (________27150), .DIN2 (___9____26026), .Q
       (_____9__26856));
  and2s1 _______507797(.DIN1 (________26823), .DIN2 (________27071), .Q
       (________26855));
  nnd2s1 _______507798(.DIN1 (____00__26589), .DIN2 (_____0__24487), .Q
       (________26854));
  nor2s1 _______507799(.DIN1 (___0_9___40457), .DIN2 (______0__37929),
       .Q (________26853));
  nnd2s1 _______507800(.DIN1 (___9_9___39611), .DIN2
       (__________________________________________9___21918), .Q
       (________26852));
  or2s1 ______507801(.DIN1 (________27355), .DIN2 (___00___26058), .Q
       (________26851));
  and2s1 _____507802(.DIN1 (___00____30589), .DIN2 (___9____26912), .Q
       (________26850));
  or2s1 _____9_507803(.DIN1 (___0____26127), .DIN2 (________26250), .Q
       (________26849));
  nor2s1 _____9_507804(.DIN1 (___9____27803), .DIN2 (____0___29011), .Q
       (_____0__26848));
  nnd2s1 _____9_507805(.DIN1 (___09___28825), .DIN2 (________25808), .Q
       (_____9__26847));
  or2s1 _____507806(.DIN1 (____9___25673), .DIN2 (___9____26024), .Q
       (________26846));
  or2s1 _____507807(.DIN1
       (_____________________________________________21777), .DIN2
       (________26835), .Q (________26845));
  nor2s1 _____0_507808(.DIN1 (____99__26228), .DIN2 (________25849), .Q
       (________26844));
  or2s1 _____0_507809(.DIN1 (___0____26100), .DIN2 (________27511), .Q
       (________26843));
  nnd2s1 _____0_507810(.DIN1 (________26153), .DIN2 (___0_____30917),
       .Q (________26842));
  nor2s1 _______507811(.DIN1 (________26840), .DIN2 (________26452), .Q
       (________26841));
  or2s1 _______507812(.DIN1 (____0___27482), .DIN2 (_____9__26838), .Q
       (_____0__26839));
  nor2s1 _______507813(.DIN1 (____9___27389), .DIN2 (____9___26772), .Q
       (________26837));
  nnd2s1 _______507814(.DIN1 (________26835), .DIN2 (________26834), .Q
       (________26836));
  nnd2s1 _______507815(.DIN1 (___9____26022), .DIN2 (________25471), .Q
       (________26833));
  nor2s1 _______507816(.DIN1 (________26481), .DIN2 (________26830), .Q
       (_____9__26831));
  nor2s1 ______507817(.DIN1 (__9__), .DIN2 (___0____26076), .Q
       (________26829));
  nnd2s1 ______507818(.DIN1 (________28454), .DIN2 (____0___26232), .Q
       (________26828));
  nnd2s1 _______507819(.DIN1 (________26165), .DIN2 (________26826), .Q
       (________26827));
  nor2s1 _______507820(.DIN1 (________25390), .DIN2 (____0___26686), .Q
       (________26825));
  nor2s1 _______507821(.DIN1 (________26823), .DIN2 (_____0__26822), .Q
       (________26824));
  nor2s1 _______507822(.DIN1 (_________37424), .DIN2 (________26671),
       .Q (_____9__26821));
  nor2s1 _______507823(.DIN1 (________26819), .DIN2 (________26835), .Q
       (________26820));
  nnd2s1 _______507824(.DIN1 (____00__26229), .DIN2 (______0__36932),
       .Q (________26818));
  nnd2s1 ______507825(.DIN1 (___9____26038), .DIN2 (____09__25871), .Q
       (________26817));
  nnd2s1 ______507826(.DIN1 (___0____26070), .DIN2 (________26789), .Q
       (________26816));
  nnd2s1 _______507827(.DIN1 (________26743), .DIN2 (________26814), .Q
       (________26815));
  nor2s1 _______507828(.DIN1 (___9____26890), .DIN2 (___0____26126), .Q
       (________26813));
  nnd2s1 _______507829(.DIN1 (_____9__27289), .DIN2 (_____9__26285), .Q
       (________26811));
  nnd2s1 _______507830(.DIN1 (________26809), .DIN2 (________25731), .Q
       (________26810));
  or2s1 _______507831(.DIN1 (_____9__23539), .DIN2 (___9____26017), .Q
       (________26808));
  nor2s1 _______507832(.DIN1 (________26805), .DIN2 (_____0__26804), .Q
       (________26806));
  nnd2s1 _______507833(.DIN1 (________27709), .DIN2 (________26802), .Q
       (_____9__26803));
  or2s1 _______507834(.DIN1 (___0_____40624), .DIN2 (___9____26035), .Q
       (________26801));
  nor2s1 _______507835(.DIN1 (________26799), .DIN2 (________26759), .Q
       (________26800));
  nnd2s1 _______507836(.DIN1 (___9_9__25987), .DIN2 (____9___25403), .Q
       (________26798));
  or2s1 _______507837(.DIN1 (____0___25680), .DIN2 (_________41277), .Q
       (________26797));
  nor2s1 ______507838(.DIN1 (________26795), .DIN2 (________26725), .Q
       (________26796));
  nnd2s1 _______507839(.DIN1 (_________37538), .DIN2
       (______________________________________0_____), .Q
       (_____0__26794));
  nnd2s1 _______507840(.DIN1 (_____0__26748), .DIN2 (________25715), .Q
       (_____9__26793));
  nnd2s1 _______507841(.DIN1 (________26214), .DIN2 (________26205), .Q
       (________26792));
  and2s1 ______507842(.DIN1 (____0___26142), .DIN2 (________25874), .Q
       (________26791));
  nnd2s1 ______507843(.DIN1 (________26789), .DIN2 (________27694), .Q
       (________26790));
  or2s1 _______507844(.DIN1
       (_______________________________________________________________9__21995),
       .DIN2 (________26787), .Q (________26788));
  and2s1 _______507845(.DIN1 (________26175), .DIN2
       (______________________21751), .Q (________26786));
  or2s1 _____9_507846(.DIN1 (__9_____29932), .DIN2 (_____09__31999), .Q
       (_____0__26785));
  nnd2s1 _____9_507847(.DIN1 (____0___26237), .DIN2 (inData[8]), .Q
       (____09__26784));
  nor2s1 _____507848(.DIN1 (____0___26782), .DIN2 (________26253), .Q
       (____0___26783));
  nnd2s1 _____507849(.DIN1 (___9____26033), .DIN2 (___9_9__25977), .Q
       (____0___26781));
  and2s1 _____0_507850(.DIN1 (____9___26404), .DIN2 (________26373), .Q
       (____0___26780));
  nnd2s1 _____0_507851(.DIN1 (___0____26995), .DIN2 (________28495), .Q
       (____0___26779));
  nnd2s1 _____0_507852(.DIN1 (____9___26227), .DIN2 (________24037), .Q
       (____0___26778));
  nnd2s1 _______507853(.DIN1 (________26178), .DIN2 (________24963), .Q
       (____0___26777));
  nnd2s1 _______507854(.DIN1 (____00__26775), .DIN2 (_____0__26390), .Q
       (____0___26776));
  or2s1 _______507855(.DIN1 (____9___26773), .DIN2 (____9___26772), .Q
       (____99__26774));
  or2s1 _______507856(.DIN1 (____9___26770), .DIN2 (________26787), .Q
       (____9___26771));
  or2s1 _______507857(.DIN1 (________25482), .DIN2 (________26245), .Q
       (____9___26769));
  nor2s1 _______507858(.DIN1 (____0___26501), .DIN2 (________26215), .Q
       (____9___26768));
  nnd2s1 _______507859(.DIN1 (___9____26032), .DIN2 (____9___27649), .Q
       (____9___26767));
  nor2s1 _______507860(.DIN1 (___00___26056), .DIN2 (____9___26226), .Q
       (____9___26766));
  nnd2s1 _______507861(.DIN1 (______9__34050), .DIN2 (_________32298),
       .Q (________26763));
  nnd2s1 _______507862(.DIN1 (____0___26235), .DIN2 (___9____26029), .Q
       (________26762));
  nor2s1 _______507863(.DIN1 (________26760), .DIN2 (________26759), .Q
       (________26761));
  nnd2s1 _______507864(.DIN1 (___0____26074), .DIN2 (_____0__26758), .Q
       (________28223));
  hi1s1 _______507865(.DIN (________27248), .Q (_____9__27609));
  hi1s1 _______507866(.DIN (____9____38949), .Q (_____0__27317));
  hi1s1 _______507867(.DIN (__9_00__30177), .Q (_____0__27260));
  xor2s1 _____9_507868(.DIN1 (_____9__25917), .DIN2 (________25811), .Q
       (___9____26908));
  hi1s1 ____0__507869(.DIN (_____9__26757), .Q (_____9__28350));
  xor2s1 ______507870(.DIN1 (________23774), .DIN2 (_________37884), .Q
       (___0____27010));
  nnd2s1 _______507871(.DIN1 (___9_9__26040), .DIN2
       (_____________________21742), .Q (___00___26957));
  nor2s1 ______507872(.DIN1 (________29110), .DIN2 (___099__27921), .Q
       (________27068));
  xor2s1 ______507873(.DIN1 (________26516), .DIN2 (_____9___37002), .Q
       (_____0__27463));
  or2s1 _____0_507874(.DIN1 (___9____27772), .DIN2 (____0___27576), .Q
       (________27454));
  nor2s1 _____9_507875(.DIN1 (________26297), .DIN2 (_____9__26635), .Q
       (_____9__27075));
  hi1s1 ____9__507876(.DIN (________26756), .Q (________27160));
  nor2s1 _______507877(.DIN1 (___0____26109), .DIN2 (________26746), .Q
       (____90__27290));
  nnd2s1 _______507878(.DIN1 (____00__26775), .DIN2 (________26755), .Q
       (____99__27299));
  nor2s1 _______507879(.DIN1 (________29256), .DIN2 (___9____26009), .Q
       (_____9__27335));
  nor2s1 ______507880(.DIN1 (____0___29283), .DIN2 (____09__26148), .Q
       (___0____27021));
  nor2s1 _______507881(.DIN1 (_________32755), .DIN2 (________26179),
       .Q (____0___27393));
  nor2s1 _______507882(.DIN1 (_________41285), .DIN2 (________26754),
       .Q (________27541));
  nor2s1 _______507883(.DIN1 (________26174), .DIN2 (___0____26072), .Q
       (_____9__27269));
  nor2s1 _______507884(.DIN1 (________26753), .DIN2 (___00___28744), .Q
       (_____9__27434));
  nnd2s1 _______507885(.DIN1 (________26752), .DIN2 (________26264), .Q
       (_____0__28502));
  nor2s1 _______507886(.DIN1 (___9____24101), .DIN2 (___0____26076), .Q
       (___0_____40063));
  and2s1 _______507887(.DIN1 (___0__9__31299), .DIN2 (________26751),
       .Q (____0___29015));
  nnd2s1 _____9_507888(.DIN1 (________26169), .DIN2 (________24879), .Q
       (___9____28703));
  nor2s1 _____9_507889(.DIN1 (____9___24740), .DIN2 (________26750), .Q
       (___0____27023));
  nor2s1 _____9_507890(.DIN1 (________28500), .DIN2 (___9____25995), .Q
       (________27324));
  nnd2s1 _____9_507891(.DIN1 (____99__26498), .DIN2 (________26213), .Q
       (________27315));
  or2s1 _____9_507892(.DIN1 (________26657), .DIN2 (_____0__26804), .Q
       (________27409));
  nor2s1 _____507893(.DIN1 (________26204), .DIN2 (__9_____29754), .Q
       (________27286));
  nor2s1 ____507894(.DIN1 (________26241), .DIN2 (________26749), .Q
       (_____0__27419));
  nnd2s1 ____90_507895(.DIN1 (________26201), .DIN2 (___9____26912), .Q
       (________27285));
  and2s1 ____90_507896(.DIN1 (_____0__26748), .DIN2 (________25709), .Q
       (________27415));
  and2s1 ____90_507897(.DIN1 (_____9__26747), .DIN2 (__9_9___29986), .Q
       (_____0__27251));
  nor2s1 ____90_507898(.DIN1 (____0___26594), .DIN2 (________26746), .Q
       (____0___27301));
  nor2s1 ____9__507899(.DIN1 (____00__25497), .DIN2 (________29233), .Q
       (___0____27011));
  hi1s1 ____0__507900(.DIN (___9____26932), .Q (___9____27783));
  nor2s1 _______507901(.DIN1 (___0____27863), .DIN2 (____0___29011), .Q
       (____0___27573));
  hi1s1 ____0_507902(.DIN (________27180), .Q (________29115));
  nnd2s1 _______507903(.DIN1 (___0_0__26060), .DIN2
       (__________________0___21750), .Q (___0_____30894));
  nnd2s1 _______507904(.DIN1 (_____0__27687), .DIN2 (___9____25985), .Q
       (____99__27391));
  or2s1 _____0_507905(.DIN1 (__9_____30204), .DIN2 (___0____27873), .Q
       (________27192));
  hi1s1 ____0__507906(.DIN (________27054), .Q (____0___27394));
  hi1s1 ____0__507907(.DIN (____00___31509), .Q (__9_____29775));
  hi1s1 ____0__507908(.DIN (________26745), .Q (________28879));
  and2s1 _______507909(.DIN1 (_____9__27967), .DIN2 (____0___27035), .Q
       (________27690));
  nnd2s1 ____9_507910(.DIN1 (________26744), .DIN2 (___0_____31094), .Q
       (_____9__29074));
  and2s1 ____9__507911(.DIN1 (________26743), .DIN2 (________26742), .Q
       (________27711));
  nor2s1 ____9__507912(.DIN1 (_____0__26168), .DIN2 (________26759), .Q
       (___99___28731));
  nor2s1 ____9__507913(.DIN1 (___9____25983), .DIN2 (________26746), .Q
       (________27284));
  nor2s1 ____9__507914(.DIN1 (________26741), .DIN2 (________26740), .Q
       (___0____28793));
  nnd2s1 ____9__507915(.DIN1 (________26243), .DIN2 (_________31868),
       .Q (________27265));
  nor2s1 ____9_507916(.DIN1 (__909___29721), .DIN2 (___0_0___30649), .Q
       (________29379));
  nor2s1 ____9__507917(.DIN1 (________26739), .DIN2 (______9__34266),
       .Q (_________33020));
  nnd2s1 ____9__507918(.DIN1 (________26446), .DIN2 (_____0__26738), .Q
       (____9___27291));
  nnd2s1 ____9__507919(.DIN1 (________29043), .DIN2 (____0___26684), .Q
       (________28535));
  and2s1 ____9__507920(.DIN1 (___9____25993), .DIN2 (_____9__26737), .Q
       (__9_____29968));
  nor2s1 ____9__507921(.DIN1 (_____9___32184), .DIN2 (___9____26016),
       .Q (___0____28788));
  nnd2s1 ____9__507922(.DIN1 (________26435), .DIN2 (________27282), .Q
       (________27720));
  nor2s1 ____9__507923(.DIN1 (_____________________21690), .DIN2
       (_____0__26177), .Q (____9___27292));
  nor2s1 ____9__507924(.DIN1 (________28310), .DIN2 (________26353), .Q
       (__9_____29758));
  nor2s1 ____9_507925(.DIN1 (___0_0___31125), .DIN2 (________28153), .Q
       (________29389));
  nnd2s1 ____9__507926(.DIN1 (________26736), .DIN2 (________26735), .Q
       (___9____29578));
  nor2s1 ____9_507927(.DIN1 (________28392), .DIN2 (_____9__26427), .Q
       (____9___27296));
  nor2s1 ____9__507928(.DIN1 (________26734), .DIN2 (________26218), .Q
       (___00____30556));
  nor2s1 _______507929(.DIN1 (___00_0__30612), .DIN2 (__9_0___29995),
       .Q (___9____27778));
  or2s1 _____507930(.DIN1 (________26733), .DIN2 (__999___30543), .Q
       (____9____32434));
  nnd2s1 _____9_507931(.DIN1 (________26732), .DIN2 (____00__26140), .Q
       (________28160));
  or2s1 ____9__507932(.DIN1 (___900__25958), .DIN2 (___0____26075), .Q
       (__99____30480));
  nnd2s1 ____9_507933(.DIN1 (___0_9___40070), .DIN2 (________26731), .Q
       (___0__9__40048));
  or2s1 _______507934(.DIN1 (_________41285), .DIN2 (________26730), .Q
       (__9_____30312));
  or2s1 ____9__507935(.DIN1 (_____________________21744), .DIN2
       (_____0___31609), .Q (____0____31579));
  nnd2s1 ____9__507936(.DIN1 (________26729), .DIN2 (_________32696),
       .Q (___0_____30977));
  and2s1 ____9__507937(.DIN1 (________25654), .DIN2 (_____0__26728), .Q
       (________27311));
  and2s1 ____9__507938(.DIN1 (___0__9__31299), .DIN2 (_____9__26727),
       .Q (_____09__31612));
  or2s1 ____9__507939(.DIN1 (________26726), .DIN2 (________26725), .Q
       (______9__33267));
  hi1s1 ______507940(.DIN (________26724), .Q (________29149));
  and2s1 ____9_507941(.DIN1 (___99___29629), .DIN2 (__9_____29792), .Q
       (_________31781));
  hi1s1 _______507942(.DIN (___0_____40188), .Q (___0_____40222));
  nnd2s1 _____507943(.DIN1 (________26180), .DIN2 (________26577), .Q
       (_____9___38610));
  hi1s1 ______507944(.DIN (________26723), .Q (___0900));
  hi1s1 _______507945(.DIN (________27052), .Q (____0_0__37159));
  nor2s1 _____0_507946(.DIN1 (___9_0__26901), .DIN2 (________26298), .Q
       (________26722));
  or2s1 _______507947(.DIN1 (___0__0__40431), .DIN2 (________26720), .Q
       (________26721));
  nnd2s1 _______507948(.DIN1 (________26187), .DIN2 (________22592), .Q
       (________26719));
  nnd2s1 _______507949(.DIN1 (_____9__26717), .DIN2 (________26716), .Q
       (_____0__26718));
  nnd2s1 _____9_507950(.DIN1 (___0____26071), .DIN2
       (_____________________21745), .Q (________26715));
  hi1s1 ____0__507951(.DIN (___0_____30903), .Q (________26714));
  nnd2s1 _______507952(.DIN1 (____9____33350), .DIN2 (inData[6]), .Q
       (________26713));
  nnd2s1 ______507953(.DIN1 (___0____26065), .DIN2 (________25268), .Q
       (________26712));
  nor2s1 _______507954(.DIN1 (________26306), .DIN2 (________26710), .Q
       (________26711));
  nnd2s1 ____0__507955(.DIN1 (________26627), .DIN2 (___9____29574), .Q
       (________26709));
  hi1s1 ____99_507956(.DIN (________28444), .Q (_____9__26708));
  hi1s1 ____9__507957(.DIN (________26706), .Q (________26707));
  hi1s1 ____9__507958(.DIN (________26704), .Q (________26705));
  nnd2s1 _______507959(.DIN1 (____9____33350), .DIN2 (inData[4]), .Q
       (________26703));
  hi1s1 ____0__507960(.DIN (_____0__26701), .Q (________26702));
  hi1s1 ____0__507961(.DIN (__99____30492), .Q (_____9__26700));
  nor2s1 _____9_507962(.DIN1 (________26698), .DIN2 (___9_____39657),
       .Q (________26699));
  nor2s1 ______507963(.DIN1 (____0___26233), .DIN2 (________25698), .Q
       (________26697));
  hi1s1 _______507964(.DIN (___9____29615), .Q (________26696));
  nor2s1 _______507965(.DIN1 (________25722), .DIN2 (___9____26001), .Q
       (________26695));
  and2s1 ______507966(.DIN1 (________26693), .DIN2 (________28519), .Q
       (________26694));
  nnd2s1 ____09_507967(.DIN1 (________27063), .DIN2 (____9___26223), .Q
       (_____0__26692));
  nnd2s1 _____0_507968(.DIN1 (_____0__26547), .DIN2 (____0___26690), .Q
       (____09__26691));
  nor2s1 _______507969(.DIN1 (________29170), .DIN2 (________26367), .Q
       (____0___26689));
  nor2s1 _______507970(.DIN1 (____0___26687), .DIN2 (____0___26686), .Q
       (____0___26688));
  nnd2s1 _______507971(.DIN1 (___0____26084), .DIN2 (____0___26684), .Q
       (____0___26685));
  and2s1 _______507972(.DIN1 (____90__26580), .DIN2 (___0__0__31003),
       .Q (____0___26683));
  nor2s1 _______507973(.DIN1 (____9___26680), .DIN2 (________26639), .Q
       (____9___26681));
  and2s1 _______507974(.DIN1 (________26647), .DIN2
       (__________________________________________________________________21986),
       .Q (____9___26679));
  nor2s1 _______507975(.DIN1 (____9___26677), .DIN2 (____9___26676), .Q
       (____9___26678));
  nor2s1 ______507976(.DIN1 (________28392), .DIN2 (________26660), .Q
       (____9___26675));
  nnd2s1 _______507977(.DIN1 (_________41275), .DIN2 (____90__26673),
       .Q (____9___26674));
  nor2s1 _______507978(.DIN1 (_____9), .DIN2 (________26671), .Q
       (_____9__26672));
  nor2s1 _______507979(.DIN1 (___0____22351), .DIN2 (________26671), .Q
       (________26670));
  or2s1 ______507980(.DIN1 (________26553), .DIN2 (________26764), .Q
       (________26669));
  or2s1 _______507981(.DIN1 (________26337), .DIN2 (________28573), .Q
       (________26668));
  nor2s1 _______507982(.DIN1 (________26666), .DIN2 (_____0__26355), .Q
       (________26667));
  or2s1 _______507983(.DIN1 (_____9__26616), .DIN2 (________26172), .Q
       (_____0__26665));
  nor2s1 _______507984(.DIN1 (________22809), .DIN2 (___0_00__31023),
       .Q (_____9__26664));
  or2s1 _______507985(.DIN1 (____0___28479), .DIN2 (________26662), .Q
       (________26663));
  nor2s1 _______507986(.DIN1 (________26660), .DIN2 (________27042), .Q
       (________26661));
  and2s1 _______507987(.DIN1 (________27989), .DIN2 (__99_0__30469), .Q
       (________26659));
  or2s1 _______507988(.DIN1 (________26657), .DIN2 (________26656), .Q
       (________26658));
  nnd2s1 ______507989(.DIN1 (___99___26047), .DIN2 (inData[8]), .Q
       (_____0__26655));
  nnd2s1 _____9_507990(.DIN1 (________25609), .DIN2 (____0___26143), .Q
       (_____9__26654));
  nor2s1 _____9_507991(.DIN1 (___9____26924), .DIN2 (___9_9__27767), .Q
       (________26653));
  nor2s1 _____9_507992(.DIN1 (___9____27820), .DIN2 (________26651), .Q
       (________26652));
  nnd2s1 _____9_507993(.DIN1 (___09___28825), .DIN2 (_____0__26256), .Q
       (________26650));
  nnd2s1 _____507994(.DIN1 (___0_99__30926), .DIN2 (__9_____29737), .Q
       (________26649));
  nnd2s1 _____9_507995(.DIN1 (________26647), .DIN2
       (______________________________________0_______21893), .Q
       (________26648));
  nnd2s1 _____0_507996(.DIN1 (________29090), .DIN2 (___9_9__26012), .Q
       (________26646));
  nor2s1 _____0_507997(.DIN1 (____0___26595), .DIN2 (___9____27801), .Q
       (_____0__26645));
  or2s1 _____0_507998(.DIN1 (________26643), .DIN2 (___9_0__26031), .Q
       (_____9__26644));
  nnd2s1 _____0_507999(.DIN1 (___00___26057), .DIN2 (inData[28]), .Q
       (________26642));
  and2s1 ______508000(.DIN1 (________26564), .DIN2 (________27339), .Q
       (________26641));
  nor2s1 _______508001(.DIN1 (________29068), .DIN2 (________26639), .Q
       (________26640));
  and2s1 _______508002(.DIN1 (___9____27800), .DIN2 (________26637), .Q
       (________26638));
  or2s1 _______508003(.DIN1 (___9____27771), .DIN2 (_____9__26635), .Q
       (_____0__26636));
  nnd2s1 ______508004(.DIN1 (___0_____30997), .DIN2 (__9_0___29899), .Q
       (________26634));
  nor2s1 _______508005(.DIN1 (________26632), .DIN2 (________26631), .Q
       (________26633));
  nnd2s1 _______508006(.DIN1 (________26629), .DIN2 (________26600), .Q
       (________26630));
  and2s1 _______508007(.DIN1 (________26627), .DIN2 (_____0__26626), .Q
       (________26628));
  nnd2s1 _______508008(.DIN1 (______0__33736), .DIN2 (___0____26063),
       .Q (_____9__26625));
  and2s1 _______508009(.DIN1 (________27163), .DIN2 (___0_____30912),
       .Q (________26624));
  nnd2s1 _______508010(.DIN1 (________26622), .DIN2 (________26366), .Q
       (________26623));
  nnd2s1 _______508011(.DIN1 (____9____33350), .DIN2 (inData[3]), .Q
       (________26621));
  xor2s1 ______508012(.DIN1
       (_____________________________________0_______21758), .DIN2
       (_________36301), .Q (________26620));
  hi1s1 _______508013(.DIN (__900_), .Q (________26619));
  nnd2s1 _______508014(.DIN1 (___9____26007), .DIN2 (________26618), .Q
       (___0____26993));
  nnd2s1 _______508015(.DIN1 (___0_____30997), .DIN2 (_____0__26617),
       .Q (________27715));
  nor2s1 ______508016(.DIN1 (_____9__26616), .DIN2 (___9____26039), .Q
       (________27162));
  and2s1 _______508017(.DIN1 (________27989), .DIN2 (____9____32424),
       .Q (________27236));
  and2s1 ______508018(.DIN1 (________27526), .DIN2 (_________31879), .Q
       (________27532));
  nor2s1 _____9_508019(.DIN1 (____9___25765), .DIN2 (____9___26676), .Q
       (________27353));
  and2s1 _____9_508020(.DIN1 (_____0__28481), .DIN2 (________28189), .Q
       (_____9__29542));
  and2s1 _____9_508021(.DIN1 (________26615), .DIN2 (__90_9__29688), .Q
       (____9___27383));
  nnd2s1 _____0_508022(.DIN1 (_____9__26717), .DIN2 (_____9__25710), .Q
       (________27229));
  nnd2s1 _____508023(.DIN1 (___99___26046), .DIN2
       (_____________________21742), .Q (_____0__27157));
  nor2s1 _______508024(.DIN1 (___9_0__26940), .DIN2 (________29531), .Q
       (____9___27293));
  or2s1 _______508025(.DIN1 (________26284), .DIN2 (___9_0__26883), .Q
       (________27199));
  or2s1 _______508026(.DIN1 (________26614), .DIN2 (________26613), .Q
       (__9_____30441));
  or2s1 _______508027(.DIN1 (____0___25225), .DIN2 (________26612), .Q
       (________28991));
  nnd2s1 _______508028(.DIN1 (___9____26005), .DIN2 (________26611), .Q
       (________27159));
  hi1s1 ____0_508029(.DIN (________27446), .Q (________27154));
  or2s1 ____0__508030(.DIN1 (________26610), .DIN2 (________26609), .Q
       (___0____27004));
  nor2s1 _______508031(.DIN1 (_____9__27498), .DIN2 (________26311), .Q
       (_____0__27186));
  and2s1 _______508032(.DIN1 (_____0__26608), .DIN2 (________26622), .Q
       (________27405));
  or2s1 _______508033(.DIN1 (___00____30608), .DIN2 (_________41283),
       .Q (________27333));
  nor2s1 _______508034(.DIN1 (___09___26135), .DIN2 (________25725), .Q
       (_____9__27326));
  hi1s1 ______508035(.DIN (________26607), .Q (___0_0___30743));
  and2s1 ______508036(.DIN1 (________26732), .DIN2 (____0___26413), .Q
       (________27274));
  hi1s1 _______508037(.DIN (________26606), .Q (________27283));
  nnd2s1 _______508038(.DIN1 (________26578), .DIN2 (________25923), .Q
       (___9____26906));
  nor2s1 _____9_508039(.DIN1 (_________31866), .DIN2 (_________32142),
       .Q (___9____26918));
  nor2s1 _______508040(.DIN1 (________26605), .DIN2 (________26207), .Q
       (___00___26956));
  hi1s1 ____0_508041(.DIN (________27608), .Q (________27701));
  hi1s1 _______508042(.DIN (______0__36697), .Q (______0__34517));
  nor2s1 _______508043(.DIN1 (________25238), .DIN2 (___9_9__26929), .Q
       (_____9___32673));
  nor2s1 _______508044(.DIN1 (________26604), .DIN2 (___9_9__26030), .Q
       (_____9__27166));
  or2s1 _______508045(.DIN1 (________26614), .DIN2 (________26262), .Q
       (________27582));
  nor2s1 _____508046(.DIN1 (____0___26410), .DIN2 (________26248), .Q
       (_____9__27344));
  nnd2s1 ____9__508047(.DIN1 (_________36955), .DIN2 (________26170),
       .Q (_________37454));
  and2s1 _______508048(.DIN1 (_____9__26563), .DIN2 (________26603), .Q
       (________27448));
  nor2s1 _______508049(.DIN1 (____0___25589), .DIN2 (________27079), .Q
       (_____9__28626));
  nnd2s1 _______508050(.DIN1 (____90__27382), .DIN2 (________26164), .Q
       (________27242));
  hi1s1 _______508051(.DIN (_________37547), .Q (______9__37353));
  nor2s1 _______508052(.DIN1 (_____0__29534), .DIN2 (________26602), .Q
       (________27322));
  nor2s1 _______508053(.DIN1 (________27724), .DIN2 (________27158), .Q
       (________29033));
  nor2s1 _______508054(.DIN1 (___0_0__26999), .DIN2 (___9____25997), .Q
       (________27168));
  hi1s1 ____09_508055(.DIN (___00____39910), .Q (___9_0___39709));
  nnd2s1 _______508056(.DIN1 (___0____26068), .DIN2 (________26601), .Q
       (________27156));
  nnd2s1 _______508057(.DIN1 (________26751), .DIN2 (__9__0__30234), .Q
       (________29236));
  nnd2s1 _______508058(.DIN1 (___00___26052), .DIN2 (________25946), .Q
       (________27402));
  hi1s1 _______508059(.DIN (_____9___33155), .Q (___0_____31266));
  nnd2s1 ______508060(.DIN1 (________25236), .DIN2 (________26600), .Q
       (________28216));
  nnd2s1 _______508061(.DIN1 (_____0__26599), .DIN2 (______0__37929),
       .Q (____0____38104));
  nnd2s1 ______508062(.DIN1 (___9____26900), .DIN2 (________25372), .Q
       (_________33664));
  and2s1 _______508063(.DIN1 (___0__0__31003), .DIN2 (____9___26587),
       .Q (________27538));
  nnd2s1 _______508064(.DIN1 (__9_90__30169), .DIN2 (________25246), .Q
       (________27221));
  and2s1 _______508065(.DIN1 (____0____33459), .DIN2 (_________32104),
       .Q (__9__9__29779));
  hi1s1 ____00_508066(.DIN (___9____26937), .Q (__9__0__29878));
  hi1s1 ____0__508067(.DIN (_____09__31708), .Q (________27164));
  nor2s1 _______508068(.DIN1 (________26734), .DIN2 (____00___31505),
       .Q (__9_____30035));
  or2s1 _______508069(.DIN1 (___9____25998), .DIN2 (________27220), .Q
       (____0___28202));
  and2s1 _______508070(.DIN1 (________28261), .DIN2 (____09__26598), .Q
       (_____9__29425));
  nor2s1 ______508071(.DIN1 (________29110), .DIN2 (____0___26597), .Q
       (_____0__27620));
  or2s1 _______508072(.DIN1 (________26454), .DIN2 (________27246), .Q
       (_____0__27427));
  nor2s1 _______508073(.DIN1 (___0_____31073), .DIN2 (__9_____30142),
       .Q (___9____29592));
  nor2s1 _______508074(.DIN1 (________27040), .DIN2 (____0___26596), .Q
       (________28242));
  nor2s1 ____9__508075(.DIN1 (________23583), .DIN2 (_________37538),
       .Q (______0__38770));
  nor2s1 _______508076(.DIN1 (____0___26595), .DIN2 (___9____27803), .Q
       (___09____31461));
  or2s1 _______508077(.DIN1 (____0___26594), .DIN2 (________26197), .Q
       (___0__9__31280));
  nor2s1 _______508078(.DIN1 (___9____25974), .DIN2 (___9____26036), .Q
       (________28344));
  hi1s1 ____0__508079(.DIN (______0__32351), .Q (______0__32205));
  and2s1 _______508080(.DIN1 (________27163), .DIN2 (____0___26593), .Q
       (___0_____31096));
  hi1s1 ____0_508081(.DIN (____0___26592), .Q (_____9__27452));
  nnd2s1 ______508082(.DIN1 (________26443), .DIN2 (________28895), .Q
       (________27615));
  hi1s1 ____0__508083(.DIN (________29176), .Q (___09____31478));
  nnd2s1 _______508084(.DIN1 (________26357), .DIN2 (________29405), .Q
       (__9_____29881));
  hi1s1 ____0__508085(.DIN (________27522), .Q (__9900));
  nor2s1 _______508086(.DIN1 (________27261), .DIN2 (________26288), .Q
       (____0___28109));
  hi1s1 ____0_508087(.DIN (____0___26591), .Q (________28364));
  nor2s1 ______508088(.DIN1 (____0___26590), .DIN2 (_________31678), .Q
       (___0_____30656));
  nnd2s1 ____9__508089(.DIN1 (____00__26589), .DIN2 (________24304), .Q
       (______9__31688));
  nnd2s1 ______508090(.DIN1 (____99__26588), .DIN2 (________25797), .Q
       (___0__9__31260));
  nor2s1 _____9_508091(.DIN1 (________26419), .DIN2 (___00___26053), .Q
       (________27458));
  nor2s1 ______508092(.DIN1 (_____0__28148), .DIN2 (________26193), .Q
       (________28900));
  nnd2s1 _____9_508093(.DIN1 (________29311), .DIN2 (___0____27842), .Q
       (___0_____30669));
  nnd2s1 _______508094(.DIN1 (_____9__27967), .DIN2 (________26273), .Q
       (_____9__27986));
  nor2s1 _____9_508095(.DIN1 (___9_9__27767), .DIN2 (___9____26917), .Q
       (________29171));
  hi1s1 ____0_508096(.DIN (_________41268), .Q (__99____30533));
  nnd2s1 _____9_508097(.DIN1 (________27495), .DIN2 (____9___26587), .Q
       (____0_9__31542));
  nnd2s1 _____0_508098(.DIN1 (___00____30589), .DIN2
       (_____________________21745), .Q (___0_90__30919));
  nor2s1 _____0_508099(.DIN1 (___9_0__26940), .DIN2 (____9___26586), .Q
       (___900__29553));
  and2s1 _____0_508100(.DIN1 (____9___26585), .DIN2 (__9_____30241), .Q
       (____09___31595));
  hi1s1 _____9_508101(.DIN (____9___26584), .Q (____9____32422));
  hi1s1 _____0_508102(.DIN (___0____28748), .Q (________27217));
  dffacs1 _________________________________________0____508103(.CLRB
       (reset), .CLK (clk), .DIN (________26162), .QN (___0__9__40580));
  nnd2s1 ____99_508104(.DIN1 (________26150), .DIN2 (____9___26583), .Q
       (__9__0__29966));
  and2s1 _______508105(.DIN1 (________26251), .DIN2 (____9___26583), .Q
       (______9__32117));
  and2s1 _______508106(.DIN1 (________28261), .DIN2 (___0_____31182),
       .Q (________28543));
  nnd2s1 ____9_508107(.DIN1 (________25694), .DIN2 (____9___26582), .Q
       (___0_____30866));
  nnd2s1 ______508108(.DIN1 (___00___26055), .DIN2 (___9____25984), .Q
       (_____0__28530));
  nnd2s1 _______508109(.DIN1 (___9____26027), .DIN2 (___9_9__26020), .Q
       (_________32022));
  nor2s1 _______508110(.DIN1 (_____________________21742), .DIN2
       (___9_0__26021), .Q (____0____31545));
  nnd2s1 _______508111(.DIN1 (___099__26139), .DIN2
       (_____________________21691), .Q (________27975));
  nnd2s1 ____9__508112(.DIN1 (________26752), .DIN2 (_____9__24802), .Q
       (_________32130));
  hi1s1 _______508113(.DIN (___9____26916), .Q (_________31667));
  nnd2s1 _______508114(.DIN1 (_____9__26246), .DIN2 (________26429), .Q
       (________29523));
  nor2s1 _______508115(.DIN1 (________26280), .DIN2 (___9_9__26003), .Q
       (____9___28010));
  nor2s1 ____99_508116(.DIN1 (____9___26581), .DIN2 (______0__41279),
       .Q (__9__0__30394));
  nnd2s1 ____9__508117(.DIN1 (____90__26580), .DIN2 (________28484), .Q
       (___0_____31262));
  nnd2s1 ____508118(.DIN1 (________26206), .DIN2 (___99___24165), .Q
       (_________38242));
  hi1s1 ____0__508119(.DIN (________26579), .Q (____9____32449));
  nor2s1 _______508120(.DIN1 (_____0__25566), .DIN2 (________26191), .Q
       (___9__9__39731));
  nnd2s1 _______508121(.DIN1 (________26578), .DIN2 (_____0__25479), .Q
       (_________31778));
  nnd2s1 ____0__508122(.DIN1 (________26609), .DIN2 (inData[23]), .Q
       (___0_____31336));
  hi1s1 ____0_508123(.DIN (________27060), .Q (_________36521));
  nnd2s1 _______508124(.DIN1 (_____9__26176), .DIN2 (________24883), .Q
       (___9_____39511));
  nnd2s1 ____00_508125(.DIN1 (________26219), .DIN2 (________26577), .Q
       (_________38869));
  nnd2s1 ____00_508126(.DIN1 (________26200), .DIN2 (________26576), .Q
       (____90___36104));
  nor2s1 ______508127(.DIN1 (____9___26581), .DIN2 (___009__26059), .Q
       (_________31870));
  dffacs1 _______________0_(.CLRB (reset), .CLK (clk), .DIN
       (___9____26028), .Q (_________22038));
  nor2s1 ____00_508128(.DIN1 (________24609), .DIN2 (____9___26221), .Q
       (____9____38007));
  and2s1 ____0__508129(.DIN1 (____0___26230), .DIN2 (________26575), .Q
       (___909___39065));
  nnd2s1 ____0__508130(.DIN1 (________26574), .DIN2 (________26484), .Q
       (__9_9___30174));
  nor2s1 ____0__508131(.DIN1 (inData[23]), .DIN2 (________26574), .Q
       (__9_____30423));
  nnd2s1 ____0__508132(.DIN1 (___9____26015), .DIN2 (________27602), .Q
       (____0____37165));
  nnd2s1 _______508133(.DIN1 (________26514), .DIN2
       (_____________________________________________21777), .Q
       (________26573));
  nnd2s1 ______508134(.DIN1 (___00____39925), .DIN2 (___0_____40612),
       .Q (________26572));
  nor2s1 _____0_508135(.DIN1 (______22154), .DIN2 (________25916), .Q
       (_____0__26571));
  nnd2s1 _______508136(.DIN1 (____09__25777), .DIN2 (________26826), .Q
       (_____9__26570));
  nnd2s1 _______508137(.DIN1 (________26568), .DIN2
       (__________________________________________9___21918), .Q
       (________26569));
  nnd2s1 _______508138(.DIN1 (________26568), .DIN2
       (______________________________________________21915), .Q
       (________26567));
  hi1s1 ____00_508139(.DIN (___0_____31277), .Q (________26566));
  hi1s1 ____9__508140(.DIN (________26564), .Q (________26565));
  nnd2s1 ______508141(.DIN1 (________26559), .DIN2
       (______________________________________0_______21892), .Q
       (________26562));
  nnd2s1 _______508142(.DIN1 (________26559), .DIN2
       (_____________________________________________21907), .Q
       (________26560));
  nnd2s1 _______508143(.DIN1 (________26557), .DIN2
       (______________________________________________21980), .Q
       (________26558));
  hi1s1 _____9_508144(.DIN (___0__9__31147), .Q (________26556));
  nnd2s1 _______508145(.DIN1 (________26557), .DIN2
       (______________________________________________21979), .Q
       (_____0__26555));
  hi1s1 _______508146(.DIN (________26553), .Q (_____9__26554));
  or2s1 _______508147(.DIN1 (___0__9__40440), .DIN2 (___9____25971), .Q
       (________26552));
  nnd2s1 ____9__508148(.DIN1 (___9____27758), .DIN2
       (____________________________________________21772), .Q
       (________26551));
  or2s1 ____9__508149(.DIN1
       (____________________________________________21772), .DIN2
       (___9____27758), .Q (________26550));
  hi1s1 _______508150(.DIN (________26548), .Q (________26549));
  nor2s1 _______508151(.DIN1 (________26545), .DIN2 (________26360), .Q
       (_____9__26546));
  nnd2s1 _______508152(.DIN1 (________25887), .DIN2 (______22153), .Q
       (________26544));
  nor2s1 _______508153(.DIN1 (___9____25994), .DIN2 (________26472), .Q
       (________26543));
  xnr2s1 _______508154(.DIN1 (_________22038), .DIN2 (_________35523),
       .Q (________26542));
  xor2s1 _______508155(.DIN1 (___0____24251), .DIN2 (_________35523),
       .Q (________26541));
  xor2s1 ______508156(.DIN1 (________26209), .DIN2 (_____9__26210), .Q
       (________26540));
  nor2s1 _______508157(.DIN1 (___0_____40411), .DIN2 (____99__26498),
       .Q (________26539));
  hi1s1 _____9_508158(.DIN (_____9__26537), .Q (_____0__26538));
  nor2s1 _______508159(.DIN1 (___0_____31198), .DIN2 (________27627),
       .Q (________26536));
  nor2s1 _______508160(.DIN1 (___0_9___40455), .DIN2 (________26458),
       .Q (________26535));
  and2s1 _____9_508161(.DIN1 (________25835), .DIN2 (________28533), .Q
       (________26534));
  nnd2s1 _____9_508162(.DIN1 (___0____26073), .DIN2 (________26532), .Q
       (________26533));
  or2s1 _____9_508163(.DIN1 (________26530), .DIN2 (____0___25865), .Q
       (________26531));
  or2s1 _____9_508164(.DIN1 (_____0__26528), .DIN2 (________25788), .Q
       (________26529));
  nor2s1 _____0_508165(.DIN1 (________22397), .DIN2 (________25803), .Q
       (_____9__26527));
  nnd2s1 _____0_508166(.DIN1 (________25827), .DIN2 (________26525), .Q
       (________26526));
  nnd2s1 _______508167(.DIN1 (________25902), .DIN2 (________26523), .Q
       (________26524));
  or2s1 _______508168(.DIN1 (________24029), .DIN2 (________25877), .Q
       (________26522));
  nnd2s1 _______508169(.DIN1 (________26520), .DIN2 (____0___26593), .Q
       (________26521));
  nor2s1 ______508170(.DIN1 (___0____25163), .DIN2 (_____0__25842), .Q
       (________26519));
  nnd2s1 _______508171(.DIN1 (________26442), .DIN2 (___0____26077), .Q
       (_____0__26518));
  nor2s1 _______508172(.DIN1 (________26516), .DIN2 (_____9___37002),
       .Q (_____9__26517));
  and2s1 _______508173(.DIN1 (________26514), .DIN2 (________26819), .Q
       (________26515));
  nnd2s1 _______508174(.DIN1 (________25719), .DIN2 (inData[22]), .Q
       (________26513));
  and2s1 _______508175(.DIN1 (________25833), .DIN2
       (_____________22084), .Q (________26512));
  nor2s1 ______508176(.DIN1 (_____0___38616), .DIN2 (________25801), .Q
       (________26511));
  hi1s1 ____9_508177(.DIN (________28308), .Q (________26510));
  nor2s1 ______508178(.DIN1 (________26740), .DIN2 (_____0__26508), .Q
       (________26509));
  nnd2s1 ______508179(.DIN1 (____0___26506), .DIN2 (________26181), .Q
       (____09__26507));
  nnd2s1 _______508180(.DIN1 (________25692), .DIN2 (___09___23305), .Q
       (____0___26505));
  nor2s1 ______508181(.DIN1 (____0___26503), .DIN2 (_________32931), .Q
       (____0___26504));
  nnd2s1 _______508182(.DIN1 (_____9__25814), .DIN2 (________26171), .Q
       (____0___26502));
  nor2s1 _______508183(.DIN1 (________25374), .DIN2 (________26840), .Q
       (____0___26500));
  and2s1 _____9_508184(.DIN1 (____99__26498), .DIN2 (___0___22171), .Q
       (____00__26499));
  nor2s1 _____0_508185(.DIN1 (_______22184), .DIN2 (_________37834), .Q
       (____9___26497));
  nor2s1 _____0_508186(.DIN1 (________22504), .DIN2 (_________38638),
       .Q (____9___26496));
  nor2s1 _______508187(.DIN1 (____9___25766), .DIN2 (____9___26494), .Q
       (____9___26495));
  and2s1 _______508188(.DIN1 (_____9__26765), .DIN2 (________25839), .Q
       (____9___26493));
  nnd2s1 _______508189(.DIN1 (___09___27916), .DIN2 (____9___26491), .Q
       (____9___26492));
  nnd2s1 _______508190(.DIN1 (_____9__25841), .DIN2 (____09__24276), .Q
       (____90__26490));
  nor2s1 _______508191(.DIN1 (________23615), .DIN2 (_____0__25695), .Q
       (_____9__26489));
  nnd2s1 ______508192(.DIN1 (____0___26506), .DIN2 (_____0__26295), .Q
       (________26488));
  and2s1 _______508193(.DIN1 (________25904), .DIN2 (_____9__24914), .Q
       (________26487));
  hi1s1 _______508194(.DIN (________26609), .Q (________26486));
  hi1s1 _______508195(.DIN (________26484), .Q (________26485));
  hi1s1 _______508196(.DIN (_____0__26482), .Q (________26483));
  xor2s1 ____09_508197(.DIN1 (_______________22076), .DIN2
       (________25903), .Q (________26480));
  nnd2s1 _____0_508198(.DIN1 (________26532), .DIN2 (________25370), .Q
       (________26479));
  or2s1 _____0_508199(.DIN1 (____9___23130), .DIN2 (____9____34338), .Q
       (________26478));
  nor2s1 _____0_508200(.DIN1 (___09___23304), .DIN2 (____9____34338),
       .Q (________26477));
  nor2s1 _____508201(.DIN1 (___0____28754), .DIN2 (________26475), .Q
       (________26476));
  nor2s1 _______508202(.DIN1 (_____9__26616), .DIN2 (_____0__25872), .Q
       (_____0__26474));
  nnd2s1 ______508203(.DIN1 (________26453), .DIN2 (____9___25582), .Q
       (_____9__26473));
  or2s1 _______508204(.DIN1 (________26470), .DIN2 (________25879), .Q
       (________26471));
  and2s1 ______508205(.DIN1 (____99__26498), .DIN2 (________22600), .Q
       (________26469));
  nor2s1 _______508206(.DIN1 (____9___25760), .DIN2 (____99__26682), .Q
       (________26468));
  nnd2s1 _______508207(.DIN1 (____90__25852), .DIN2 (________26826), .Q
       (________26467));
  or2s1 _______508208(.DIN1 (_____9__25851), .DIN2 (_________34916), .Q
       (_____0__26466));
  nnd2s1 _______508209(.DIN1 (_____0__28481), .DIN2 (_________31749),
       .Q (_____9__26465));
  nor2s1 _____9_508210(.DIN1 (____09__26331), .DIN2 (________25798), .Q
       (________26464));
  nnd2s1 _____0_508211(.DIN1 (___0_0__26069), .DIN2 (___0__0__40571),
       .Q (________26463));
  nnd2s1 _______508212(.DIN1 (________25907), .DIN2 (_________33596),
       .Q (________26462));
  nnd2s1 _______508213(.DIN1 (________25922), .DIN2 (inData[26]), .Q
       (________26461));
  or2s1 _______508214(.DIN1 (________25895), .DIN2 (____0____38052), .Q
       (________26460));
  nor2s1 _______508215(.DIN1 (___9____26034), .DIN2 (________26458), .Q
       (________26459));
  xnr2s1 _______508216(.DIN1 (___0_____40573), .DIN2 (______0__35711),
       .Q (_____0__26457));
  xor2s1 ______508217(.DIN1
       (__________________________________________________________________22005),
       .DIN2 (____0____38091), .Q (_____9__26456));
  xnr2s1 _______508218(.DIN1 (___0_9___40452), .DIN2 (_________9_), .Q
       (________26455));
  nnd2s1 _____9_508219(.DIN1 (________26425), .DIN2 (________26259), .Q
       (________26745));
  xnr2s1 ______508220(.DIN1 (___0_9___40452), .DIN2 (___________), .Q
       (_________36317));
  nnd2s1 _______508221(.DIN1 (________28122), .DIN2 (__9_99__29992), .Q
       (_____9__26757));
  nnd2s1 _______508222(.DIN1 (_________41295), .DIN2 (________26258),
       .Q (____0___26592));
  hi1s1 ____0__508223(.DIN (___0990__31494), .Q (___9____26931));
  nor2s1 _____9_508224(.DIN1 (________26454), .DIN2 (____0___29374), .Q
       (________27954));
  nnd2s1 ______508225(.DIN1 (________26453), .DIN2 (________26163), .Q
       (____9___27117));
  hi1s1 ____0__508226(.DIN (__9_____30241), .Q (___09____31467));
  hi1s1 ____00_508227(.DIN (_____9__27551), .Q (___9____26914));
  hi1s1 _____9_508228(.DIN (________26574), .Q (___9____26907));
  hi1s1 ______508229(.DIN (________26452), .Q (________28447));
  hi1s1 _______508230(.DIN (___99___28734), .Q (________27080));
  nor2s1 _______508231(.DIN1 (inData[14]), .DIN2 (____0____32541), .Q
       (________26706));
  hi1s1 _____508232(.DIN (________26451), .Q (__9_____29976));
  hi1s1 _____0_508233(.DIN (________28982), .Q (___9_9__26919));
  nnd2s1 _______508234(.DIN1 (________26520), .DIN2 (________25239), .Q
       (________27141));
  nor2s1 _____9_508235(.DIN1 (________26449), .DIN2 (__9_____29932), .Q
       (________28889));
  and2s1 _______508236(.DIN1 (________25784), .DIN2 (________27694), .Q
       (____0___27036));
  nor2s1 ____90_508237(.DIN1 (________26217), .DIN2 (________26432), .Q
       (____0___27122));
  nor2s1 ____90_508238(.DIN1 (_____0__26448), .DIN2 (_____9__26447), .Q
       (___0____27007));
  hi1s1 _______508239(.DIN (________26446), .Q (________27073));
  nnd2s1 _____0_508240(.DIN1 (___0_00__31216), .DIN2 (________26374),
       .Q (________26807));
  nor2s1 ____9__508241(.DIN1 (_____), .DIN2 (________25812), .Q
       (________27444));
  or2s1 _______508242(.DIN1 (________26445), .DIN2 (________26444), .Q
       (___09___27028));
  hi1s1 ____9__508243(.DIN (________26443), .Q (___0____27851));
  hi1s1 ____0__508244(.DIN (__9_00__30272), .Q (________27155));
  nor2s1 _______508245(.DIN1 (inData[28]), .DIN2 (_________31809), .Q
       (_____0__26701));
  nor2s1 _______508246(.DIN1 (________26440), .DIN2 (________25606), .Q
       (___9_0__27786));
  nnd2s1 _____508247(.DIN1 (__9_____29873), .DIN2 (________29140), .Q
       (________28457));
  nnd2s1 _______508248(.DIN1 (________26442), .DIN2 (_____0__26418), .Q
       (________26579));
  nnd2s1 _______508249(.DIN1 (________29140), .DIN2 (________26420), .Q
       (___9____26898));
  nnd2s1 ____9_508250(.DIN1 (________25843), .DIN2 (________25829), .Q
       (________26724));
  nor2s1 _______508251(.DIN1 (________26441), .DIN2 (________25886), .Q
       (___0_0__27009));
  nor2s1 _______508252(.DIN1 (______0__35694), .DIN2 (________25779),
       .Q (___90___26870));
  or2s1 _______508253(.DIN1 (________28441), .DIN2 (__9_____29773), .Q
       (________27277));
  nor2s1 _______508254(.DIN1 (____9___25761), .DIN2 (_________31827),
       .Q (________27105));
  nor2s1 _______508255(.DIN1 (________26440), .DIN2 (________25894), .Q
       (___0_0__27018));
  nor2s1 _______508256(.DIN1 (___9____26019), .DIN2 (________25810), .Q
       (____0___26591));
  nnd2s1 ____9__508257(.DIN1 (________26439), .DIN2 (___909__25967), .Q
       (___0__9__30813));
  dffacs1 _________________________________________0____508258(.CLRB
       (reset), .CLK (clk), .DIN (_____0__25909), .QN (___0_____40578));
  nnd2s1 _____0_508259(.DIN1 (_____0__26438), .DIN2 (________25708), .Q
       (________27616));
  nor2s1 _______508260(.DIN1 (____09__28931), .DIN2 (________29217), .Q
       (________29176));
  nnd2s1 ______508261(.DIN1 (_________31725), .DIN2 (__9_____30058), .Q
       (________27522));
  nor2s1 _____0_508262(.DIN1 (_____9__26437), .DIN2 (________26436), .Q
       (___0__9__30880));
  nnd2s1 ______508263(.DIN1 (________25911), .DIN2 (________27288), .Q
       (________27054));
  nnd2s1 ____9__508264(.DIN1 (________26435), .DIN2 (_____9__27289), .Q
       (___0____28763));
  and2s1 ____9__508265(.DIN1 (________25693), .DIN2 (________26434), .Q
       (________27365));
  or2s1 _______508266(.DIN1 (________26433), .DIN2 (________26432), .Q
       (________27605));
  nor2s1 _______508267(.DIN1 (_________41291), .DIN2 (___0____27863),
       .Q (_________31953));
  nnd2s1 _______508268(.DIN1 (________25545), .DIN2 (___90___28651), .Q
       (________27049));
  nor2s1 ____9__508269(.DIN1 (________26431), .DIN2 (_____9__25908), .Q
       (_____0__28863));
  nnd2s1 _______508270(.DIN1 (____999__33432), .DIN2 (________26430),
       .Q (___00____30630));
  or2s1 _______508271(.DIN1 (____0____33465), .DIN2 (____0___25776), .Q
       (_________32701));
  nnd2s1 ____9_508272(.DIN1 (_____0__25824), .DIN2 (________26429), .Q
       (________27287));
  nnd2s1 ____0__508273(.DIN1 (________25893), .DIN2
       (____0________________21664), .Q (________26723));
  nnd2s1 ____9__508274(.DIN1 (____99__26498), .DIN2 (____0___26236), .Q
       (______9__35683));
  nor2s1 ____9__508275(.DIN1 (___9____25992), .DIN2 (_____0__26428), .Q
       (_____9___32868));
  nor2s1 ____9_508276(.DIN1 (__________________0___21750), .DIN2
       (________25789), .Q (____0___27924));
  hi1s1 _______508277(.DIN (_________31731), .Q (___0____27868));
  hi1s1 _______508278(.DIN (___090___31413), .Q (___9_0__27768));
  hi1s1 _____9_508279(.DIN (_____9__26427), .Q (_____0__27363));
  nnd2s1 _______508280(.DIN1 (________29341), .DIN2 (_____0__26286), .Q
       (__99____30492));
  hi1s1 _______508281(.DIN (_________37538), .Q (________27099));
  hi1s1 _____0_508282(.DIN (________29326), .Q (________29108));
  hi1s1 ____0_508283(.DIN (_____0__29175), .Q (__9_00__29993));
  nor2s1 ____9__508284(.DIN1 (inData[23]), .DIN2 (_________31809), .Q
       (___0____27005));
  nnd2s1 _______508285(.DIN1 (________25645), .DIN2 (____0___26415), .Q
       (___0__0__31168));
  nor2s1 ____508286(.DIN1 (______0__35694), .DIN2 (________25848), .Q
       (________27052));
  nnd2s1 _______508287(.DIN1 (________25913), .DIN2 (________26426), .Q
       (___0_____30903));
  and2s1 ____9__508288(.DIN1 (________27494), .DIN2 (____9___26587), .Q
       (___0_____30807));
  nnd2s1 ____9_508289(.DIN1 (________26425), .DIN2 (___09___24263), .Q
       (___0____27858));
  and2s1 ____9_508290(.DIN1 (__9_9___29991), .DIN2 (________26426), .Q
       (__9_____30198));
  nor2s1 _______508291(.DIN1 (________26424), .DIN2 (________26423), .Q
       (____9____33393));
  nor2s1 ____9__508292(.DIN1 (________25756), .DIN2 (____0___25870), .Q
       (________28026));
  and2s1 ______508293(.DIN1 (________26422), .DIN2 (___90___28651), .Q
       (_____0__28181));
  nor2s1 _______508294(.DIN1 (________27169), .DIN2 (_____9__27138), .Q
       (________29498));
  and2s1 _______508295(.DIN1 (___0_00__30740), .DIN2 (________25697),
       .Q (___0_____30654));
  or2s1 _____9_508296(.DIN1 (_____________________21745), .DIN2
       (________28612), .Q (__9_9___30451));
  nor2s1 _____9_508297(.DIN1 (________26421), .DIN2 (________26432), .Q
       (__9_____30432));
  nnd2s1 ____9__508298(.DIN1 (________25545), .DIN2 (inData[23]), .Q
       (_____0__27280));
  nnd2s1 _____508299(.DIN1 (________25816), .DIN2 (________26601), .Q
       (___0_____31297));
  nnd2s1 _______508300(.DIN1 (________26420), .DIN2 (________29533), .Q
       (________28171));
  or2s1 ____9__508301(.DIN1 (________26419), .DIN2 (____9___25858), .Q
       (___9____27764));
  nnd2s1 ____9__508302(.DIN1 (____99__25861), .DIN2 (_____0__26418), .Q
       (__9_00__30177));
  nor2s1 ____9__508303(.DIN1 (________26309), .DIN2 (____0___26416), .Q
       (___9____29615));
  nnd2s1 ____9__508304(.DIN1 (____09__26417), .DIN2 (____0___26141), .Q
       (_____90__35555));
  nor2s1 _______508305(.DIN1 (________24877), .DIN2 (________25847), .Q
       (________27060));
  nor2s1 _______508306(.DIN1 (_____0__26247), .DIN2 (____0___26416), .Q
       (__9_____29742));
  and2s1 _______508307(.DIN1 (________25883), .DIN2
       (_____________________21678), .Q (______0__31950));
  nor2s1 ____99_508308(.DIN1 (___9_9___39339), .DIN2 (________25836),
       .Q (____9____38949));
  nnd2s1 ____99_508309(.DIN1 (___0____26103), .DIN2 (________29428), .Q
       (_____9___33155));
  nnd2s1 ____9__508310(.DIN1 (________25799), .DIN2 (____0___26415), .Q
       (_____9___31891));
  and2s1 _______508311(.DIN1 (__9_9___29991), .DIN2
       (_____________________21742), .Q (_________32042));
  hi1s1 ____0__508312(.DIN (____0___26414), .Q (__909___29719));
  hi1s1 ____0__508313(.DIN (____0___26413), .Q (_____9__29174));
  nnd2s1 ____9__508314(.DIN1 (________26274), .DIN2 (________26269), .Q
       (________27256));
  nor2s1 _______508315(.DIN1 (________26307), .DIN2 (____9___25859), .Q
       (________27608));
  nor2s1 ____508316(.DIN1 (____0________________21716), .DIN2
       (________25791), .Q (_________33123));
  hi1s1 ____0__508317(.DIN (________26299), .Q (___0__9__30890));
  hi1s1 ______508318(.DIN (____0___26412), .Q (____09___31598));
  hi1s1 ____09_508319(.DIN (____0___26411), .Q (_________36856));
  nnd2s1 _______508320(.DIN1 (____0___25867), .DIN2 (____9___26406), .Q
       (_________38666));
  nor2s1 ____99_508321(.DIN1 (____0___26410), .DIN2 (________25830), .Q
       (________27248));
  nnd2s1 ____508322(.DIN1 (________25873), .DIN2 (___0____26125), .Q
       (______0__36697));
  nnd2s1 ______508323(.DIN1 (________25921), .DIN2 (____0___26409), .Q
       (___00____39910));
  nnd2s1 ____00_508324(.DIN1 (________25890), .DIN2 (________25600), .Q
       (____0_9__36267));
  or2s1 _______508325(.DIN1 (____00__26408), .DIN2 (_____9__25720), .Q
       (___9_____39738));
  nor2s1 ____00_508326(.DIN1 (____99__26407), .DIN2 (_____9__25703), .Q
       (___9_0___39624));
  nnd2s1 ____00_508327(.DIN1 (________25809), .DIN2 (____9___26406), .Q
       (_________38463));
  nor2s1 ____0_508328(.DIN1 (________26450), .DIN2 (________25875), .Q
       (___0_____40188));
  dffacs1 __________________508329(.CLRB (reset), .CLK (clk), .DIN
       (________25782), .QN (_______________22075));
  hi1s1 ____0__508330(.DIN (____9___26405), .Q (___0_____40284));
  nor2s1 _______508331(.DIN1 (___0_____30882), .DIN2 (____9___26402),
       .Q (____9___26403));
  and2s1 ______508332(.DIN1 (________25616), .DIN2 (________25935), .Q
       (____9___26401));
  and2s1 _____9_508333(.DIN1 (________25666), .DIN2 (____9___25400), .Q
       (____90__26400));
  nor2s1 _____9_508334(.DIN1 (___0_____40447), .DIN2 (________26557),
       .Q (_____9__26399));
  nor2s1 _____9_508335(.DIN1 (___9____25063), .DIN2 (_________36301),
       .Q (________26398));
  nor2s1 ______508336(.DIN1 (___0_____40448), .DIN2 (________26557), .Q
       (________26397));
  nor2s1 _______508337(.DIN1 (________22507), .DIN2 (________26559), .Q
       (________26396));
  nnd2s1 _______508338(.DIN1 (________26394), .DIN2 (____9___23126), .Q
       (________26395));
  or2s1 _______508339(.DIN1 (____0___27925), .DIN2 (________26392), .Q
       (________26393));
  and2s1 _______508340(.DIN1 (_____0__26390), .DIN2 (________28495), .Q
       (________26391));
  nor2s1 _______508341(.DIN1 (___0_0__22297), .DIN2 (___00____39925),
       .Q (_____9__26389));
  nor2s1 _______508342(.DIN1 (___0_____40534), .DIN2 (_____0__26341),
       .Q (________26388));
  nor2s1 _______508343(.DIN1 (____0___25684), .DIN2 (____9___25304), .Q
       (________26387));
  and2s1 ______508344(.DIN1 (_____9__25603), .DIN2 (____9___25401), .Q
       (________26386));
  nnd2s1 _______508345(.DIN1 (________26344), .DIN2 (__99__), .Q
       (________26385));
  nnd2s1 _____9_508346(.DIN1 (____9___25674), .DIN2 (________23648), .Q
       (________26384));
  or2s1 _____9_508347(.DIN1 (__99____30487), .DIN2 (________26382), .Q
       (________26383));
  nnd2s1 _____0_508348(.DIN1 (_____9__28360), .DIN2 (_____0__26390), .Q
       (________26381));
  nor2s1 _____0_508349(.DIN1 (________23566), .DIN2 (________25658), .Q
       (_____0__26380));
  and2s1 _____508350(.DIN1 (___00____39925), .DIN2 (___0__0__40431), .Q
       (_____9__26379));
  nor2s1 _______508351(.DIN1 (________23519), .DIN2 (________25655), .Q
       (________26378));
  nnd2s1 _______508352(.DIN1 (________26376), .DIN2 (_____0__25520), .Q
       (________26377));
  nnd2s1 _______508353(.DIN1 (________26374), .DIN2 (________26373), .Q
       (________26375));
  and2s1 ______508354(.DIN1 (____9___25672), .DIN2 (_____0__26371), .Q
       (________26372));
  nnd2s1 _______508355(.DIN1 (________25621), .DIN2 (___0____26099), .Q
       (_____9__26370));
  hi1s1 ____9__508356(.DIN (________26367), .Q (________26368));
  nnd2s1 _______508357(.DIN1 (________26394), .DIN2 (________22723), .Q
       (________26365));
  hi1s1 ____0__508358(.DIN (________28600), .Q (________26364));
  hi1s1 _______508359(.DIN (_____0__26822), .Q (_____0__26363));
  or2s1 ______508360(.DIN1 (__99____30501), .DIN2 (_____0__25786), .Q
       (_____9__26362));
  nnd2s1 _______508361(.DIN1 (____9___26321), .DIN2 (____0___25411), .Q
       (________26361));
  dffacs1 _______________508362(.CLRB (reset), .CLK (clk), .DIN
       (________26360), .Q (outData[1]));
  or2s1 ___9___508363(.DIN1 (________27554), .DIN2 (____0___29283), .Q
       (________26359));
  hi1s1 ____9_508364(.DIN (_____0__26355), .Q (________26356));
  nor2s1 _______508365(.DIN1 (inData[5]), .DIN2 (________26261), .Q
       (_____9__26354));
  hi1s1 ____99_508366(.DIN (________26830), .Q (________26352));
  xor2s1 _______508367(.DIN1 (___0___22273), .DIN2 (_________37614), .Q
       (________26351));
  nnd2s1 _______508368(.DIN1 (___90___25960), .DIN2 (_____0__27411), .Q
       (________26350));
  hi1s1 ____0__508369(.DIN (_________31973), .Q (_____0__26349));
  hi1s1 ____0__508370(.DIN (___0_____30810), .Q (________26348));
  and2s1 _______508371(.DIN1 (____99__26498), .DIN2 (___00___23222), .Q
       (________26347));
  and2s1 ____09_508372(.DIN1 (____90__29272), .DIN2 (________26344), .Q
       (________26345));
  nnd2s1 ____09_508373(.DIN1 (___0____26982), .DIN2 (____0___25223), .Q
       (________26343));
  or2s1 _____0_508374(.DIN1 (_____9__22528), .DIN2 (_____0__26341), .Q
       (________26342));
  or2s1 _____0_508375(.DIN1 (________22428), .DIN2 (_____0__26341), .Q
       (_____9__26340));
  and2s1 _____0_508376(.DIN1 (________26271), .DIN2 (_____9__27996), .Q
       (________26339));
  nnd2s1 _______508377(.DIN1 (________25611), .DIN2 (____0___25314), .Q
       (________26338));
  nnd2s1 _______508378(.DIN1 (________26335), .DIN2 (________26282), .Q
       (________26336));
  or2s1 ______508379(.DIN1 (_________31942), .DIN2 (________26333), .Q
       (________26334));
  nor2s1 _______508380(.DIN1 (____09__26331), .DIN2 (________25639), .Q
       (_____0__26332));
  nor2s1 _______508381(.DIN1 (________23642), .DIN2 (___00____39925),
       .Q (____0___26330));
  nor2s1 _______508382(.DIN1 (___0____25204), .DIN2 (___9____26006), .Q
       (____0___26329));
  nnd2s1 _______508383(.DIN1 (____9___26406), .DIN2 (________25637), .Q
       (____0___26328));
  nor2s1 _______508384(.DIN1 (____9___23783), .DIN2 (________25652), .Q
       (____0___26327));
  or2s1 ______508385(.DIN1 (___0____26117), .DIN2 (____0___26325), .Q
       (____0___26326));
  nor2s1 _______508386(.DIN1 (______22154), .DIN2 (_____9__27176), .Q
       (____0___26324));
  nor2s1 ______508387(.DIN1 (___0_0__26122), .DIN2 (_________41297), .Q
       (____00__26323));
  nor2s1 ______508388(.DIN1 (____0___25412), .DIN2 (____9___26321), .Q
       (____9___26322));
  or2s1 _______508389(.DIN1 (_____9__25378), .DIN2 (____9___26321), .Q
       (____9___26320));
  nnd2s1 _______508390(.DIN1 (_____0__25633), .DIN2 (___0____25161), .Q
       (____9___26319));
  nnd2s1 _______508391(.DIN1 (________25905), .DIN2 (____9___26317), .Q
       (____9___26318));
  nnd2s1 _____9_508392(.DIN1 (_____0__25651), .DIN2 (________25702), .Q
       (____90__26315));
  nnd2s1 _____9_508393(.DIN1 (___0_____31084), .DIN2 (________25713),
       .Q (_____9__26314));
  nnd2s1 _____508394(.DIN1 (_________41293), .DIN2 (____0___26415), .Q
       (________26313));
  nor2s1 _____0_508395(.DIN1 (_____0__26305), .DIN2 (________26311), .Q
       (________26312));
  nor2s1 _______508396(.DIN1 (________26309), .DIN2 (_____9__25669), .Q
       (________26310));
  and2s1 ______508397(.DIN1 (_____0__26617), .DIN2 (________26637), .Q
       (________26308));
  nnd2s1 _______508398(.DIN1 (_____9__27185), .DIN2 (________29208), .Q
       (___0_9__26966));
  nnd2s1 _______508399(.DIN1 (________25818), .DIN2
       (_________________0___21740), .Q (________26607));
  nor2s1 _______508400(.DIN1 (________24897), .DIN2 (________26632), .Q
       (____9___27297));
  nor2s1 _______508401(.DIN1 (________26307), .DIN2 (_____9__25659), .Q
       (________26606));
  hi1s1 ____0__508402(.DIN (___9_9___39611), .Q (___9_9___39610));
  nnd2s1 _______508403(.DIN1 (________25820), .DIN2 (____0___26231), .Q
       (__9_9___29989));
  nor2s1 _______508404(.DIN1 (_________35587), .DIN2 (_________31809),
       .Q (___900__26864));
  hi1s1 ____99_508405(.DIN (____0___26595), .Q (________29511));
  or2s1 ___9__508406(.DIN1 (________26306), .DIN2 (________26283), .Q
       (___9_0__26930));
  hi1s1 ____00_508407(.DIN (______0__33984), .Q (____0____33487));
  nor2s1 ___9___508408(.DIN1 (_____0__26305), .DIN2 (_____9__26304), .Q
       (___0____26989));
  nor2s1 ___9___508409(.DIN1 (_________32001), .DIN2 (________26303),
       .Q (___0____26985));
  and2s1 _______508410(.DIN1 (___0____26119), .DIN2 (___90___28650), .Q
       (___0_0__26960));
  nor2s1 ____9_508411(.DIN1 (___9____26912), .DIN2 (________25638), .Q
       (____9___26584));
  nnd2s1 _______508412(.DIN1 (________25629), .DIN2 (_____0__26832), .Q
       (________27956));
  hi1s1 _______508413(.DIN (________26302), .Q (___0____26981));
  hi1s1 ____0__508414(.DIN (________28189), .Q (___9_9__26910));
  hi1s1 _______508415(.DIN (________26301), .Q (___0____26996));
  nor2s1 _______508416(.DIN1 (___0_____31088), .DIN2 (________25716),
       .Q (________26756));
  nnd2s1 ______508417(.DIN1 (_________36928), .DIN2 (______9__32959),
       .Q (___9____26933));
  nor2s1 ______508418(.DIN1 (________26300), .DIN2 (____0___27571), .Q
       (___9____26923));
  hi1s1 ___9___508419(.DIN (________26298), .Q (___9____26935));
  or2s1 ______508420(.DIN1 (________29210), .DIN2 (____0___26325), .Q
       (________27492));
  nor2s1 _______508421(.DIN1 (________26726), .DIN2 (________26297), .Q
       (___0____26968));
  nnd2s1 _______508422(.DIN1 (___09____31487), .DIN2 (_____9__26265),
       .Q (____09__27215));
  hi1s1 ____0_508423(.DIN (________29531), .Q (________27493));
  nor2s1 _______508424(.DIN1 (__99_9__30508), .DIN2 (____0____32541),
       .Q (________26704));
  nor2s1 ______508425(.DIN1 (________26296), .DIN2 (_____9__25891), .Q
       (________27425));
  nor2s1 _______508426(.DIN1 (_________32305), .DIN2 (________26297),
       .Q (_____9__28167));
  nor2s1 ______508427(.DIN1 (________25631), .DIN2 (________26333), .Q
       (________28252));
  nor2s1 ______508428(.DIN1 (________25294), .DIN2 (____9___26321), .Q
       (___9____26913));
  nor2s1 _______508429(.DIN1 (________25607), .DIN2 (_____9__25650), .Q
       (___0_9__26998));
  or2s1 _______508430(.DIN1 (________27665), .DIN2 (________25608), .Q
       (___9_9__26939));
  nnd2s1 ______508431(.DIN1 (________27468), .DIN2 (_____0__26295), .Q
       (___9____26926));
  and2s1 _______508432(.DIN1 (________29309), .DIN2 (________28162), .Q
       (___9____26936));
  or2s1 _______508433(.DIN1 (________27181), .DIN2 (____00___33437), .Q
       (___9____26934));
  nor2s1 _____0_508434(.DIN1 (_____9__26294), .DIN2 (________26293), .Q
       (________29253));
  or2s1 _____9_508435(.DIN1 (____0_0__31523), .DIN2 (__9_____30115), .Q
       (________27320));
  nor2s1 _____9_508436(.DIN1 (________23643), .DIN2 (___00____39925),
       .Q (________27077));
  nor2s1 _____508437(.DIN1 (_____9__28081), .DIN2 (____0___26782), .Q
       (________27089));
  nnd2s1 _______508438(.DIN1 (___0_9__26111), .DIN2 (________26292), .Q
       (_____0__29305));
  nor2s1 _______508439(.DIN1 (_____9__24705), .DIN2 (________25718), .Q
       (________27504));
  nnd2s1 _______508440(.DIN1 (____0____32541), .DIN2 (________24879),
       .Q (______0__32980));
  or2s1 _______508441(.DIN1 (_____0__25918), .DIN2 (________26382), .Q
       (____9_0__33356));
  nor2s1 _______508442(.DIN1 (___0____26105), .DIN2 (________26559), .Q
       (________27674));
  or2s1 _______508443(.DIN1 (________26291), .DIN2 (_________31942), .Q
       (__9__9__30010));
  nor2s1 ______508444(.DIN1 (______0__31903), .DIN2 (________25643), .Q
       (____0___28293));
  or2s1 _______508445(.DIN1 (____0___25227), .DIN2 (________26290), .Q
       (__9_9___30362));
  and2s1 _______508446(.DIN1 (___09_9__31426), .DIN2 (____0___25775),
       .Q (____9____32417));
  nor2s1 _______508447(.DIN1 (___9____25970), .DIN2 (____0____32541),
       .Q (__99____30473));
  or2s1 ______508448(.DIN1 (_____9__25728), .DIN2 (___9_0__26004), .Q
       (___9____27784));
  nor2s1 _____0_508449(.DIN1 (__99____30485), .DIN2 (________26632), .Q
       (__9_____30314));
  nor2s1 _______508450(.DIN1 (________25617), .DIN2 (________28589), .Q
       (____0____32516));
  nor2s1 ______508451(.DIN1 (____9___27389), .DIN2 (________28485), .Q
       (_____9__27084));
  nnd2s1 _______508452(.DIN1 (_____0__25623), .DIN2 (________25569), .Q
       (___9____27763));
  and2s1 _______508453(.DIN1 (________26742), .DIN2 (________25627), .Q
       (____9___28550));
  hi1s1 ____508454(.DIN (_________41287), .Q (___0_____31162));
  nor2s1 _______508455(.DIN1 (________26289), .DIN2 (____0___26325), .Q
       (________28497));
  hi1s1 ____00_508456(.DIN (________26288), .Q (________29331));
  nnd2s1 _______508457(.DIN1 (___0__0__30787), .DIN2 (________25624),
       .Q (____000__31503));
  nor2s1 ______508458(.DIN1 (___0__0__30872), .DIN2 (________26287), .Q
       (________27416));
  nnd2s1 _______508459(.DIN1 (________26242), .DIN2 (_____0__27177), .Q
       (__900_));
  nnd2s1 _______508460(.DIN1 (_____0__26286), .DIN2 (_____0__26758), .Q
       (___0_9___31015));
  hi1s1 ____99_508461(.DIN (_____9__26285), .Q (________28277));
  nnd2s1 _______508462(.DIN1 (________25919), .DIN2 (________25920), .Q
       (________28305));
  nor2s1 ____9__508463(.DIN1 (________26284), .DIN2 (________26283), .Q
       (________28523));
  dffacs1 ______________________________________508464(.CLRB (reset),
       .CLK (clk), .DIN (________25837), .Q (_____________22079));
  nnd2s1 _______508465(.DIN1 (________26282), .DIN2 (________26281), .Q
       (___9____26944));
  nor2s1 _______508466(.DIN1 (________26280), .DIN2 (________25636), .Q
       (___9____26937));
  nnd2s1 _______508467(.DIN1 (________25714), .DIN2 (________27545), .Q
       (___9____27762));
  or2s1 ___9___508468(.DIN1 (________26279), .DIN2 (________26303), .Q
       (________29049));
  nnd2s1 ____9__508469(.DIN1 (________25689), .DIN2 (____0___26146), .Q
       (___0____28748));
  nnd2s1 _______508470(.DIN1 (_____0__25604), .DIN2 (________26272), .Q
       (_____09__31708));
  hi1s1 ____0__508471(.DIN (_____9___31697), .Q (________28149));
  and2s1 _______508472(.DIN1 (________26442), .DIN2 (________26429), .Q
       (________28044));
  nnd2s1 _______508473(.DIN1 (________25828), .DIN2 (________26426), .Q
       (___0_____31006));
  nnd2s1 ___90_508474(.DIN1 (________26270), .DIN2 (___0____25172), .Q
       (___9____26916));
  hi1s1 ____99_508475(.DIN (________26278), .Q (__99____30465));
  hi1s1 ____00_508476(.DIN (________26277), .Q (________27491));
  hi1s1 ____0__508477(.DIN (___0_____31282), .Q (___0_____30679));
  hi1s1 ____0__508478(.DIN (____0___29011), .Q (________28281));
  hi1s1 ____0_508479(.DIN (____9___26586), .Q (__9_____30332));
  hi1s1 ______508480(.DIN (__9_____29777), .Q (___0_____31151));
  nnd2s1 _______508481(.DIN1 (________25615), .DIN2 (________26611), .Q
       (________28444));
  hi1s1 ____0__508482(.DIN (________26749), .Q (__99____30516));
  and2s1 _____0_508483(.DIN1 (_____0__26276), .DIN2 (________28040), .Q
       (___0____27889));
  hi1s1 ____0__508484(.DIN (_____9__26275), .Q (___0_____31237));
  nnd2s1 _______508485(.DIN1 (________26274), .DIN2 (________26267), .Q
       (____0___27483));
  or2s1 _______508486(.DIN1 (____9___25860), .DIN2 (________25724), .Q
       (___0_____31156));
  hi1s1 ____508487(.DIN (________26273), .Q (________29142));
  nnd2s1 _______508488(.DIN1 (________26268), .DIN2 (________25282), .Q
       (________27180));
  nor2s1 _______508489(.DIN1 (________25391), .DIN2 (____9___26321), .Q
       (_________32748));
  nnd2s1 _____508490(.DIN1 (________25619), .DIN2 (________26272), .Q
       (____09__28480));
  or2s1 _____508491(.DIN1 (____00___33437), .DIN2 (________26333), .Q
       (__9_____30098));
  nnd2s1 _____0_508492(.DIN1 (________28230), .DIN2 (________26271), .Q
       (________27964));
  nor2s1 _____0_508493(.DIN1 (____09__24848), .DIN2 (________27190), .Q
       (______0__33727));
  hi1s1 ____0__508494(.DIN (_________31879), .Q (________28909));
  nnd2s1 ______508495(.DIN1 (________25649), .DIN2
       (_____________________21736), .Q (__9__0__29760));
  nnd2s1 ____90_508496(.DIN1 (________25544), .DIN2 (inData[19]), .Q
       (_____0__27148));
  nnd2s1 ____90_508497(.DIN1 (________25705), .DIN2 (____00__24746), .Q
       (___0_____31040));
  or2s1 _______508498(.DIN1 (________25699), .DIN2 (____0___27214), .Q
       (___00_9__30621));
  nnd2s1 ___9__508499(.DIN1 (________26270), .DIN2 (________25380), .Q
       (_________31933));
  nnd2s1 _______508500(.DIN1 (_____0__25642), .DIN2 (________26269), .Q
       (___9____26932));
  nor2s1 _______508501(.DIN1 (__________________0___21750), .DIN2
       (________25888), .Q (______0__32351));
  nor2s1 _______508502(.DIN1 (inData[19]), .DIN2 (____0____32541), .Q
       (___9____26909));
  hi1s1 _____0_508503(.DIN (___0____27015), .Q (_________31738));
  hi1s1 _______508504(.DIN (___0____27860), .Q (_________32296));
  nor2s1 _____9_508505(.DIN1 (____9___25955), .DIN2 (________25691), .Q
       (___9____26928));
  nnd2s1 _______508506(.DIN1 (________25618), .DIN2
       (_____________________21742), .Q (___0__0__31290));
  dffacs1 _________________________________________0____508507(.CLRB
       (reset), .CLK (clk), .DIN (_____9__25805), .Q
       (_____________________________________0______21755));
  nor2s1 _______508508(.DIN1 (____9___26581), .DIN2 (________25826), .Q
       (____00___31509));
  nnd2s1 _______508509(.DIN1 (________26268), .DIN2 (________26267), .Q
       (____9___27294));
  nor2s1 _______508510(.DIN1 (____9___25952), .DIN2 (_____0__26266), .Q
       (__9_____30163));
  nor2s1 ____9__508511(.DIN1 (___0_0__25135), .DIN2 (____9___26321), .Q
       (_________32658));
  dffacs1 ________________0_508512(.CLRB (reset), .CLK (clk), .DIN
       (_____0__25704), .QN
       (______________________________________________________________________________________0__22093));
  nnd2s1 _______508513(.DIN1 (_____9__26265), .DIN2 (________26264), .Q
       (___09_9__31446));
  nnd2s1 ____9__508514(.DIN1 (____9___25671), .DIN2 (____9___25404), .Q
       (__9_____30024));
  nor2s1 _______508515(.DIN1 (___0____26083), .DIN2 (________25635), .Q
       (__9_0___30179));
  nor2s1 ______508516(.DIN1 (________26604), .DIN2 (________25641), .Q
       (__9__9__29743));
  nnd2s1 _______508517(.DIN1 (________25664), .DIN2 (________26269), .Q
       (____9___27478));
  hi1s1 ___9__508518(.DIN (________26263), .Q (_________31955));
  hi1s1 ___9___508519(.DIN (________26262), .Q (______0__32196));
  nnd2s1 _______508520(.DIN1 (________26261), .DIN2 (________26260), .Q
       (________27082));
  nnd2s1 _____9_508521(.DIN1 (________25625), .DIN2 (________26259), .Q
       (________27446));
  nor2s1 _______508522(.DIN1 (___9____24134), .DIN2 (_____0__25832), .Q
       (____0_0__38064));
  and2s1 _______508523(.DIN1 (________25885), .DIN2 (________26258), .Q
       (____00__29009));
  hi1s1 ____0__508524(.DIN (____0____32543), .Q (____0____32539));
  and2s1 ____9__508525(.DIN1 (________25667), .DIN2 (________26257), .Q
       (___9_0___39705));
  dffacs1 __________________508526(.CLRB (reset), .CLK (clk), .DIN
       (________25780), .QN (_______________22077));
  nor2s1 ____9_508527(.DIN1 (___9____23175), .DIN2 (________25610), .Q
       (_________37547));
  nor2s1 ______508528(.DIN1 (____09__27128), .DIN2 (________25819), .Q
       (_____0__26256));
  nnd2s1 ______508529(.DIN1 (________26254), .DIN2 (________24004), .Q
       (_____9__26255));
  nnd2s1 _______508530(.DIN1 (____9___29007), .DIN2 (________27598), .Q
       (________26253));
  nor2s1 _______508531(.DIN1
       (_____________________________________________21940), .DIN2
       (________26254), .Q (________26252));
  nor2s1 ____0__508532(.DIN1 (_____0__26149), .DIN2 (________25524), .Q
       (________26251));
  nor2s1 ______508533(.DIN1 (________24039), .DIN2 (________26249), .Q
       (________26250));
  or2s1 _______508534(.DIN1 (_____0__26247), .DIN2 (________25273), .Q
       (________26248));
  and2s1 ______508535(.DIN1 (___9____26002), .DIN2 (________25751), .Q
       (_____9__26246));
  nor2s1 _____0_508536(.DIN1 (___0_____40414), .DIN2 (___0_____40380),
       .Q (________26245));
  nnd2s1 _______508537(.DIN1 (______0__37345), .DIN2 (_____9__23386),
       .Q (________26244));
  and2s1 _______508538(.DIN1 (___0_____31385), .DIN2 (__9__9__30319),
       .Q (________26243));
  nnd2s1 _______508539(.DIN1 (________26240), .DIN2 (________26239), .Q
       (________26241));
  nor2s1 _______508540(.DIN1 (____9__22224), .DIN2 (____99___37096), .Q
       (____09__26238));
  nor2s1 ______508541(.DIN1 (___0_____40573), .DIN2 (____0___26236), .Q
       (____0___26237));
  or2s1 _______508542(.DIN1
       (______________________________________0_______21893), .DIN2
       (____0___26234), .Q (____0___26235));
  and2s1 _______508543(.DIN1 (___0_____30688), .DIN2
       (__________________________________________0_), .Q
       (____0___26233));
  and2s1 _______508544(.DIN1 (____0___26231), .DIN2 (________25350), .Q
       (____0___26232));
  and2s1 _______508545(.DIN1 (________25530), .DIN2 (________23541), .Q
       (____0___26230));
  nor2s1 _______508546(.DIN1 (____9___24926), .DIN2 (________25542), .Q
       (____00__26229));
  and2s1 ______508547(.DIN1 (__9_9___29888), .DIN2
       (______________________________________0_______21891), .Q
       (____99__26228));
  nor2s1 _______508548(.DIN1 (_____9__22998), .DIN2 (________25463), .Q
       (____9___26227));
  nor2s1 _______508549(.DIN1 (_____0___41311), .DIN2 (____0___25504),
       .Q (____9___26226));
  nnd2s1 _____0_508550(.DIN1 (_________38435), .DIN2 (____00__22644),
       .Q (____9___26225));
  and2s1 _____0_508551(.DIN1 (_________38435), .DIN2
       (_____________________________________________21783), .Q
       (____9___26224));
  or2s1 _____0_508552(.DIN1 (______________22104), .DIN2
       (______________________________________________21932), .Q
       (____9___26223));
  or2s1 _____508553(.DIN1 (________23610), .DIN2 (________25509), .Q
       (____9___26221));
  nor2s1 _____9_508554(.DIN1 (___0____24252), .DIN2 (_____9__25546), .Q
       (_____9__26220));
  nor2s1 _____9_508555(.DIN1 (_____9__25478), .DIN2 (___0____24244), .Q
       (________26219));
  nor2s1 _____508556(.DIN1 (________26217), .DIN2 (________25934), .Q
       (________26218));
  xor2s1 ______508557(.DIN1 (_________37245), .DIN2 (_____09__35744),
       .Q (________26216));
  or2s1 _______508558(.DIN1 (________26199), .DIN2 (________25433), .Q
       (________26215));
  nnd2s1 ______508559(.DIN1 (____0___25410), .DIN2 (________24431), .Q
       (________26214));
  nor2s1 ______508560(.DIN1 (________22424), .DIN2 (____0___26236), .Q
       (________26213));
  and2s1 _______508561(.DIN1 (____9____32424), .DIN2 (___0__0__40431),
       .Q (________26212));
  nnd2s1 _____508562(.DIN1 (_____9__26210), .DIN2 (________26209), .Q
       (_____0__26211));
  and2s1 _______508563(.DIN1 (___0_9___40452), .DIN2 (___________), .Q
       (________26208));
  or2s1 _______508564(.DIN1 (_________31958), .DIN2 (________25465), .Q
       (________26207));
  nor2s1 ______508565(.DIN1 (___0____23247), .DIN2 (________25486), .Q
       (________26206));
  nnd2s1 _______508566(.DIN1 (________25422), .DIN2
       (______________________________________0___9_), .Q
       (________26205));
  nor2s1 _______508567(.DIN1 (_____________________21742), .DIN2
       (____9___25303), .Q (________26204));
  nor2s1 _______508568(.DIN1 (___0__9__40440), .DIN2 (____0___26234),
       .Q (_____0__26203));
  hi1s1 _____508569(.DIN (____0___29374), .Q (_____9__26202));
  nor2s1 ______508570(.DIN1 (_____9__25632), .DIN2 (________26173), .Q
       (________26201));
  nor2s1 _______508571(.DIN1 (________26199), .DIN2 (___0_0__25194), .Q
       (________26200));
  nnd2s1 _______508572(.DIN1 (____9___25950), .DIN2 (_____9__25368), .Q
       (________26197));
  nnd2s1 ______508573(.DIN1 (________26249), .DIN2
       (__________________________________________0___21919), .Q
       (________26196));
  and2s1 _______508574(.DIN1 (___00_0__39902), .DIN2 (________23371),
       .Q (_____0__26195));
  nor2s1 _______508575(.DIN1 (___0_____40436), .DIN2 (____90__25576),
       .Q (_____9__26194));
  hi1s1 _____0_508576(.DIN (__99____30513), .Q (________26193));
  and2s1 _______508577(.DIN1 (___00_0__39902), .DIN2 (___09___22359),
       .Q (________26192));
  nnd2s1 _____0_508578(.DIN1 (________25237), .DIN2 (___0____24232), .Q
       (________26191));
  nnd2s1 ______508579(.DIN1 (________26188), .DIN2 (________24984), .Q
       (________26189));
  or2s1 _______508580(.DIN1 (____99__23038), .DIN2 (_____9__26210), .Q
       (________26187));
  or2s1 _______508581(.DIN1
       (___________________________________________), .DIN2
       (________28399), .Q (_____0__26186));
  nnd2s1 _______508582(.DIN1 (___0____26085), .DIN2 (____90__26673), .Q
       (_____9__26185));
  nor2s1 _______508583(.DIN1 (________22611), .DIN2 (____0___26234), .Q
       (________26184));
  or2s1 _____9_508584(.DIN1 (________25485), .DIN2 (_____9__25424), .Q
       (________26183));
  or2s1 _______508585(.DIN1 (___0_____40576), .DIN2 (________28399), .Q
       (________26182));
  nor2s1 _______508586(.DIN1 (_____0__25445), .DIN2 (________23990), .Q
       (________26180));
  nnd2s1 _______508587(.DIN1 (___0____27014), .DIN2 (_____9__25757), .Q
       (________26179));
  nnd2s1 _______508588(.DIN1 (_____9__25388), .DIN2 (inData[28]), .Q
       (________26178));
  nnd2s1 _______508589(.DIN1 (________25382), .DIN2 (________23801), .Q
       (_____0__26177));
  nor2s1 _______508590(.DIN1 (________23840), .DIN2 (________25532), .Q
       (_____9__26176));
  nor2s1 _______508591(.DIN1 (________26174), .DIN2 (________26173), .Q
       (________26175));
  nnd2s1 _____0_508592(.DIN1 (________25449), .DIN2 (________26171), .Q
       (________26172));
  nor2s1 _____0_508593(.DIN1 (________24415), .DIN2 (________25292), .Q
       (________26170));
  nor2s1 _____0_508594(.DIN1 (_____0__26168), .DIN2 (__9_____30054), .Q
       (________26169));
  nor2s1 _____0_508595(.DIN1 (________25432), .DIN2 (_________38249),
       .Q (_____9__26167));
  nnd2s1 _____0_508596(.DIN1 (________26249), .DIN2
       (______________________________________________21911), .Q
       (________26166));
  and2s1 _____9_508597(.DIN1 (___9____25049), .DIN2 (________25473), .Q
       (________26165));
  and2s1 ______508598(.DIN1 (____9___25764), .DIN2 (________26163), .Q
       (________26164));
  or2s1 _______508599(.DIN1 (______0__34259), .DIN2 (________25427), .Q
       (________26162));
  or2s1 _______508600(.DIN1 (___0_9___40452), .DIN2 (___________), .Q
       (________26161));
  nnd2s1 _______508601(.DIN1 (________25429), .DIN2 (________25385), .Q
       (________26160));
  xor2s1 _______508602(.DIN1
       (____________________________________________21820), .DIN2
       (_________37202), .Q (_____0__26159));
  xnr2s1 _______508603(.DIN1
       (_________________________________________0___21856), .DIN2
       (___9_____39554), .Q (_____9__26158));
  xor2s1 _______508604(.DIN1 (___0__0__40571), .DIN2 (________22381),
       .Q (________26157));
  xnr2s1 _______508605(.DIN1 (______0_), .DIN2 (_____09__35744), .Q
       (________26156));
  xor2s1 _______508606(.DIN1 (___9_____39773), .DIN2 (_________38860),
       .Q (________26155));
  hi1s1 ____0__508607(.DIN (___0_____31073), .Q (________26154));
  nor2s1 _______508608(.DIN1 (__9__9__30419), .DIN2 (________25341), .Q
       (________26153));
  nnd2s1 _______508609(.DIN1 (___0_0__26082), .DIN2 (________26151), .Q
       (________26152));
  nor2s1 ______508610(.DIN1 (_____0__26149), .DIN2 (_____0__25528), .Q
       (________26150));
  nnd2s1 _______508611(.DIN1 (___9____25973), .DIN2 (____0___26147), .Q
       (____09__26148));
  hi1s1 _______508612(.DIN (____0___26144), .Q (____0___26145));
  or2s1 _______508613(.DIN1 (________26530), .DIN2 (________25423), .Q
       (____0___26143));
  nnd2s1 ______508614(.DIN1 (____0___26141), .DIN2 (___0_99__40560), .Q
       (____0___26142));
  hi1s1 _____508615(.DIN (__9_____29750), .Q (____00__26140));
  nor2s1 _______508616(.DIN1 (________24762), .DIN2 (____0___25505), .Q
       (___099__26139));
  nnd2s1 _______508617(.DIN1 (___0_____30688), .DIN2
       (______________________________________________21912), .Q
       (___09___26138));
  nnd2s1 _______508618(.DIN1 (____0___26141), .DIN2 (________25850), .Q
       (___09___26137));
  nnd2s1 _______508619(.DIN1 (____0____37139), .DIN2 (__________22061),
       .Q (___09___26136));
  or2s1 _______508620(.DIN1 (___0__9__40540), .DIN2 (____0___26236), .Q
       (___09___26135));
  and2s1 _______508621(.DIN1 (___00____30587), .DIN2 (_____9__22633),
       .Q (___09___26134));
  nnd2s1 _______508622(.DIN1 (___9____26023), .DIN2
       (______________22110), .Q (___09___26133));
  or2s1 ______508623(.DIN1 (___0_____40617), .DIN2 (____0___26234), .Q
       (___090__26132));
  nnd2s1 _______508624(.DIN1 (___0____26097), .DIN2
       (_____________________________________9_______21883), .Q
       (___0_9__26131));
  nnd2s1 _______508625(.DIN1 (__9_9___29888), .DIN2 (___0__0__40619),
       .Q (___0____26130));
  nnd2s1 _______508626(.DIN1 (__9_9___29888), .DIN2
       (______________________________________0___9_), .Q
       (___0____26129));
  nnd2s1 _______508627(.DIN1 (________25939), .DIN2
       (_________________________________________9___21861), .Q
       (___0____26128));
  and2s1 _______508628(.DIN1 (________26249), .DIN2
       (______________________________________________21916), .Q
       (___0____26127));
  and2s1 _______508629(.DIN1 (____9___26491), .DIN2 (___0_0__25165), .Q
       (________26744));
  hi1s1 _____508630(.DIN (_________31725), .Q (___0____27897));
  hi1s1 _____9_508631(.DIN (________26435), .Q (_____9__26838));
  hi1s1 _______508632(.DIN (___0____26126), .Q (________27309));
  nnd2s1 ______508633(.DIN1 (_____9__25444), .DIN2 (___0____26125), .Q
       (____0___26411));
  nnd2s1 _______508634(.DIN1 (___0____26124), .DIN2 (________24823), .Q
       (_____9__26427));
  nnd2s1 _______508635(.DIN1 (__99____30506), .DIN2 (___0____26123), .Q
       (________26452));
  nnd2s1 _____0_508636(.DIN1 (____9___25307), .DIN2 (________26611), .Q
       (________26446));
  nnd2s1 _____9_508637(.DIN1 (____9____32424), .DIN2 (inData[23]), .Q
       (________26484));
  nor2s1 _____9_508638(.DIN1 (________23438), .DIN2 (________25289), .Q
       (________26578));
  nor2s1 _____9_508639(.DIN1 (inData[23]), .DIN2 (___0____25136), .Q
       (________26610));
  nor2s1 _____9_508640(.DIN1 (________23555), .DIN2 (___0____26104), .Q
       (________27165));
  nnd2s1 _______508641(.DIN1 (____0___25312), .DIN2 (________26611), .Q
       (________26443));
  nor2s1 _____508642(.DIN1 (_____________________21736), .DIN2
       (________25232), .Q (____00__26589));
  nor2s1 _______508643(.DIN1 (___0_0__26122), .DIN2 (________28063), .Q
       (_____0__26547));
  nnd2s1 _______508644(.DIN1 (________25439), .DIN2
       (_________________9___21749), .Q (___9____27796));
  nnd2s1 ____9__508645(.DIN1 (___09___25218), .DIN2 (______9__32019),
       .Q (________26451));
  nor2s1 _______508646(.DIN1 (________28070), .DIN2 (___9____27774), .Q
       (________26615));
  nnd2s1 ______508647(.DIN1 (___0____25200), .DIN2 (___0_9__26121), .Q
       (________26548));
  nnd2s1 _______508648(.DIN1 (____9___25491), .DIN2 (___0____26120), .Q
       (________26720));
  nor2s1 _______508649(.DIN1 (______________22066), .DIN2
       (________25241), .Q (____0___27657));
  nnd2s1 _______508650(.DIN1 (________25447), .DIN2 (___0____26120), .Q
       (_____9__26537));
  nor2s1 _______508651(.DIN1 (______________________21753), .DIN2
       (___0_9__26101), .Q (________26553));
  nnd2s1 _______508652(.DIN1 (___0____26119), .DIN2 (___0____26107), .Q
       (____9___26772));
  nor2s1 _______508653(.DIN1 (___0____26089), .DIN2 (___9____25982), .Q
       (________26750));
  nor2s1 ______508654(.DIN1 (________29068), .DIN2 (____9___25762), .Q
       (_____0__26482));
  hi1s1 _______508655(.DIN (___0____26118), .Q (________26743));
  hi1s1 ______508656(.DIN (___9____26925), .Q (___9____26895));
  and2s1 ______508657(.DIN1 (________26603), .DIN2 (____0___24847), .Q
       (___9____26903));
  nor2s1 _______508658(.DIN1 (_____9__24525), .DIN2 (_____0__25507), .Q
       (________27429));
  nnd2s1 _______508659(.DIN1 (___0____28811), .DIN2 (_____9__25747), .Q
       (________26725));
  nor2s1 _______508660(.DIN1 (___0____26117), .DIN2 (________26289), .Q
       (___0____28784));
  and2s1 _______508661(.DIN1 (________26434), .DIN2 (______0__31921),
       .Q (________27660));
  nnd2s1 _______508662(.DIN1 (____0___26141), .DIN2 (___0_____40574),
       .Q (________26834));
  nnd2s1 _______508663(.DIN1 (____00__25222), .DIN2 (___99___26049), .Q
       (________26357));
  hi1s1 ____0__508664(.DIN (_________31827), .Q (________27613));
  nor2s1 _______508665(.DIN1 (____0___26590), .DIN2 (___0____26116), .Q
       (________26481));
  hi1s1 ____0_508666(.DIN (__9_____29773), .Q (____90__26580));
  nor2s1 _______508667(.DIN1 (___0____26115), .DIN2 (________29173), .Q
       (________26789));
  hi1s1 _______508668(.DIN (_____0__28481), .Q (________26754));
  hi1s1 ____0__508669(.DIN (____0____37113), .Q (____9_0__36107));
  or2s1 ______508670(.DIN1 (________25783), .DIN2 (________29072), .Q
       (________26660));
  nnd2s1 ______508671(.DIN1 (________25521), .DIN2 (________25362), .Q
       (____9___26582));
  nor2s1 _______508672(.DIN1 (________25736), .DIN2 (___0____26114), .Q
       (________26366));
  nor2s1 _______508673(.DIN1 (___0____26113), .DIN2 (___0_0__26112), .Q
       (_____9__26563));
  nnd2s1 _______508674(.DIN1 (___0_____30684), .DIN2 (___0_9___31214),
       .Q (_____0__26355));
  and2s1 _______508675(.DIN1 (___0_9__26111), .DIN2 (___0____26110), .Q
       (________26729));
  nor2s1 _______508676(.DIN1 (________28057), .DIN2 (_____0__25778), .Q
       (_____9__26747));
  nor2s1 _____508677(.DIN1 (________29336), .DIN2 (___9____25091), .Q
       (_____0__26748));
  nor2s1 _______508678(.DIN1 (___0_____31140), .DIN2 (________26296),
       .Q (________26358));
  nnd2s1 _______508679(.DIN1 (________25516), .DIN2 (_____9__27996), .Q
       (________26662));
  nor2s1 _____0_508680(.DIN1 (___0____26109), .DIN2 (___0____26088), .Q
       (___0____28758));
  hi1s1 ____0__508681(.DIN (___9____26921), .Q (_____0___31604));
  nnd2s1 _______508682(.DIN1 (________25233), .DIN2 (___0____26108), .Q
       (________26749));
  nor2s1 ______508683(.DIN1 (___0____26113), .DIN2 (____9___25577), .Q
       (________26622));
  nnd2s1 _______508684(.DIN1 (___00_0__39902), .DIN2 (_____0__25319),
       .Q (___9_____39644));
  hi1s1 ____0_508685(.DIN (__909___29721), .Q (___0_____31394));
  nnd2s1 _______508686(.DIN1 (___0____26107), .DIN2 (___0____26106), .Q
       (_____9__26635));
  nnd2s1 _______508687(.DIN1 (____0___26234), .DIN2 (___0____26105), .Q
       (________26671));
  nor2s1 _______508688(.DIN1 (________26440), .DIN2 (___0____26104), .Q
       (________26830));
  nnd2s1 _______508689(.DIN1 (_____0__25435), .DIN2 (______22153), .Q
       (__9_____29792));
  nnd2s1 _______508690(.DIN1 (________25436), .DIN2 (________26426), .Q
       (________29405));
  nor2s1 _______508691(.DIN1 (___0__0__31080), .DIN2 (________25487),
       .Q (________27611));
  hi1s1 ____00_508692(.DIN (___0____26103), .Q (____9___27566));
  nor2s1 _______508693(.DIN1 (________24605), .DIN2 (_____9__25488), .Q
       (________26752));
  nor2s1 _______508694(.DIN1 (__9__0__29916), .DIN2 (________29225), .Q
       (____00__26775));
  nor2s1 _______508695(.DIN1 (__909___29720), .DIN2 (___0_0__26102), .Q
       (____9___27295));
  nor2s1 ______508696(.DIN1 (___0____26080), .DIN2 (___0_9__26101), .Q
       (__9_____30430));
  nor2s1 ______508697(.DIN1 (___0____26100), .DIN2 (___9____26011), .Q
       (___0____26995));
  nnd2s1 _______508698(.DIN1 (________25253), .DIN2 (___0____26099), .Q
       (_____9__26717));
  nor2s1 _______508699(.DIN1 (________24791), .DIN2 (________25451), .Q
       (___0____27878));
  or2s1 ______508700(.DIN1 (___0____26098), .DIN2 (___0____26097), .Q
       (_________38856));
  or2s1 _____0_508701(.DIN1 (________28070), .DIN2 (___0____26096), .Q
       (____9___27118));
  nnd2s1 _______508702(.DIN1 (___0____26095), .DIN2 (__9_____29771), .Q
       (________26759));
  nor2s1 _______508703(.DIN1 (____0___24936), .DIN2 (___9____26037), .Q
       (___90___28648));
  nnd2s1 _______508704(.DIN1 (_____0___33721), .DIN2 (___0_9__28814),
       .Q (___9____26890));
  nnd2s1 _______508705(.DIN1 (____0___25414), .DIN2 (________25750), .Q
       (________27282));
  nor2s1 _______508706(.DIN1 (___0____26100), .DIN2 (________29225), .Q
       (__9__0__30003));
  nnd2s1 _______508707(.DIN1 (__9_____29921), .DIN2 (___0____26094), .Q
       (______0__31970));
  nor2s1 ______508708(.DIN1 (________25553), .DIN2 (____9___25492), .Q
       (________26730));
  and2s1 ____9__508709(.DIN1 (___0____25209), .DIN2
       (_____________________21678), .Q (___9____27789));
  nnd2s1 ______508710(.DIN1 (___0_____40380), .DIN2 (________23749), .Q
       (___0__9__40392));
  nnd2s1 _______508711(.DIN1 (___0_9__28814), .DIN2 (________26523), .Q
       (_________33849));
  nnd2s1 ______508712(.DIN1 (________29066), .DIN2 (____9___26491), .Q
       (________26639));
  nor2s1 _______508713(.DIN1 (________25518), .DIN2 (__99____30463), .Q
       (________26809));
  nnd2s1 _______508714(.DIN1 (____9____32424), .DIN2 (___0____25196),
       .Q (________27042));
  nnd2s1 _______508715(.DIN1 (________29441), .DIN2 (___0____25189), .Q
       (___0_____30986));
  nnd2s1 _______508716(.DIN1 (___0____26093), .DIN2 (___0_0__26092), .Q
       (________26656));
  nor2s1 _____9_508717(.DIN1 (________27071), .DIN2 (___90___25961), .Q
       (_____0__26822));
  nnd2s1 _____508718(.DIN1 (____0___26141), .DIN2 (____9____35264), .Q
       (________26835));
  nor2s1 _____0_508719(.DIN1 (___0_9__26091), .DIN2 (__9_____30400), .Q
       (________28308));
  nor2s1 _______508720(.DIN1 (_________33553), .DIN2 (________25755),
       .Q (_________32298));
  nnd2s1 ______508721(.DIN1 (_________31868), .DIN2 (________26239), .Q
       (_____0__26804));
  or2s1 _______508722(.DIN1 (____9___25581), .DIN2 (__9_9___29888), .Q
       (___0_00__31023));
  nnd2s1 _______508723(.DIN1 (__90____29672), .DIN2 (___0____26062), .Q
       (___9____27798));
  and2s1 _______508724(.DIN1 (_____0__27039), .DIN2 (____0____31527),
       .Q (_________32720));
  or2s1 _______508725(.DIN1 (_____________________21683), .DIN2
       (________25297), .Q (________27163));
  or2s1 ____90_508726(.DIN1 (____0____________9___21722), .DIN2
       (________26249), .Q (________26787));
  nor2s1 ____9__508727(.DIN1 (___9____27801), .DIN2 (____0___27576), .Q
       (________27726));
  nor2s1 ____9__508728(.DIN1 (___0_0__25145), .DIN2 (___0____26090), .Q
       (___09____31443));
  nor2s1 ____508729(.DIN1 (__99____30487), .DIN2 (___0____28754), .Q
       (_________33934));
  nnd2s1 _____508730(.DIN1 (________25462), .DIN2 (_____0__25349), .Q
       (________28859));
  nor2s1 _____9_508731(.DIN1 (___0____26089), .DIN2 (___0____26088), .Q
       (___0_9___31111));
  nor2s1 _____9_508732(.DIN1 (________25510), .DIN2 (________25940), .Q
       (___9____27803));
  nor2s1 _____508733(.DIN1 (___0____26087), .DIN2 (________25441), .Q
       (___00___28744));
  hi1s1 _____0_508734(.DIN (___0____26086), .Q (________29529));
  nor2s1 _______508735(.DIN1 (____9___24928), .DIN2 (________26173), .Q
       (___00____30589));
  nor2s1 _____9_508736(.DIN1 (________26739), .DIN2 (____0____31589),
       .Q (______9__34050));
  nor2s1 ____90_508737(.DIN1 (________26174), .DIN2 (____09__25416), .Q
       (___0_0___30649));
  nor2s1 ______508738(.DIN1 (________28063), .DIN2 (____9___26773), .Q
       (_____9__29455));
  nnd2s1 ______508739(.DIN1 (___0____26085), .DIN2 (________25508), .Q
       (___0_____30997));
  hi1s1 ____0__508740(.DIN (___0____26084), .Q (___00_0__30612));
  nor2s1 ____9__508741(.DIN1 (___0____26083), .DIN2 (____99__25406), .Q
       (___0____27860));
  nnd2s1 _____0_508742(.DIN1 (___0_0__26082), .DIN2 (___0_9__26081), .Q
       (__9_0___30274));
  nor2s1 _____9_508743(.DIN1 (________26309), .DIN2 (________25456), .Q
       (________27158));
  nor2s1 _______508744(.DIN1 (inData[3]), .DIN2 (___0____25136), .Q
       (________26609));
  nor2s1 _______508745(.DIN1 (___0____26080), .DIN2 (________25817), .Q
       (___0_0___31125));
  nnd2s1 ______508746(.DIN1 (_____99__33716), .DIN2 (___0____26079), .Q
       (______9__34266));
  nnd2s1 _______508747(.DIN1 (________25468), .DIN2 (___0____26078), .Q
       (___9_0__27805));
  nor2s1 ______508748(.DIN1 (_____________________21691), .DIN2
       (________25428), .Q (___099__27921));
  hi1s1 ____0_508749(.DIN (_________37893), .Q (_________37616));
  hi1s1 ____508750(.DIN (___9____27758), .Q (_________34026));
  nnd2s1 _______508751(.DIN1 (________25266), .DIN2 (___0____26077), .Q
       (________28189));
  or2s1 _______508752(.DIN1 (___0____26087), .DIN2 (_____0__25928), .Q
       (___009___30634));
  nnd2s1 _______508753(.DIN1 (________25286), .DIN2 (____0___25774), .Q
       (________28261));
  nnd2s1 _______508754(.DIN1 (_________34243), .DIN2 (________28084),
       .Q (_________33551));
  nnd2s1 _______508755(.DIN1 (____9___25493), .DIN2
       (_____________________21742), .Q (_____9___31694));
  hi1s1 _______508756(.DIN (_________37834), .Q (______0__37929));
  hi1s1 ____0__508757(.DIN (___0____26076), .Q (___0_9___40070));
  hi1s1 ____09_508758(.DIN (________26360), .Q (___0_____30709));
  hi1s1 _______508759(.DIN (________26425), .Q (___0____26075));
  hi1s1 _______508760(.DIN (________26840), .Q (___0____26074));
  or2s1 _____9_508761(.DIN1 (________25644), .DIN2 (_____9__25460), .Q
       (___0____26072));
  nor2s1 ___9___508762(.DIN1 (________22853), .DIN2 (___0____25205), .Q
       (___0____26071));
  nor2s1 ___9__508763(.DIN1 (___0____26067), .DIN2 (___0_9__25202), .Q
       (___0____26068));
  hi1s1 ____0__508764(.DIN (____9___27475), .Q (___0____26066));
  or2s1 ___9___508765(.DIN1 (___0____26064), .DIN2 (________25476), .Q
       (___0____26065));
  and2s1 ____0_508766(.DIN1 (___0____26062), .DIN2 (___0____26061), .Q
       (___0____26063));
  nor2s1 ____0_508767(.DIN1 (___99___26045), .DIN2 (____0___25503), .Q
       (___0_0__26060));
  nnd2s1 ____0__508768(.DIN1 (________25418), .DIN2 (________25634), .Q
       (___009__26059));
  or2s1 ____0__508769(.DIN1 (___9____25981), .DIN2 (___90___28652), .Q
       (___00___26058));
  nor2s1 ____0__508770(.DIN1 (___00___26056), .DIN2 (________25255), .Q
       (___00___26057));
  nor2s1 ____0_508771(.DIN1 (___00___26054), .DIN2 (________25533), .Q
       (___00___26055));
  or2s1 ____0__508772(.DIN1 (_____9__25823), .DIN2 (________25269), .Q
       (___00___26053));
  and2s1 ____09_508773(.DIN1 (________25234), .DIN2 (_________33686),
       .Q (___00___26052));
  nor2s1 ____09_508774(.DIN1 (___90___23138), .DIN2 (___0_____30688),
       .Q (___000__26051));
  nnd2s1 ____09_508775(.DIN1 (________25717), .DIN2 (___99___26049), .Q
       (___999__26050));
  nor2s1 ____09_508776(.DIN1 (___9____23185), .DIN2 (___0_____30688),
       .Q (___99___26048));
  nnd2s1 _____0_508777(.DIN1 (____0___25408), .DIN2 (_____9__24811), .Q
       (___99___26047));
  nor2s1 ______508778(.DIN1 (___99___26045), .DIN2 (_____0__25453), .Q
       (___99___26046));
  or2s1 _______508779(.DIN1 (___99___26043), .DIN2 (____9___26222), .Q
       (___99___26044));
  nnd2s1 _______508780(.DIN1 (___0____28811), .DIN2 (________25342), .Q
       (___99___26042));
  nnd2s1 _______508781(.DIN1 (___9_____39206), .DIN2 (_____0__22605),
       .Q (___990__26041));
  nor2s1 _______508782(.DIN1 (___99___26045), .DIN2 (___09___25215), .Q
       (___9_9__26040));
  nnd2s1 _______508783(.DIN1 (____9___25495), .DIN2 (________24519), .Q
       (___9____26039));
  nor2s1 _______508784(.DIN1 (________24861), .DIN2 (___9____26037), .Q
       (___9____26038));
  nnd2s1 _______508785(.DIN1 (________25477), .DIN2 (________23072), .Q
       (___9____26036));
  nor2s1 _______508786(.DIN1 (___9____26034), .DIN2 (___0____26097), .Q
       (___9____26035));
  nor2s1 _______508787(.DIN1 (___0____26080), .DIN2 (________25457), .Q
       (___9____26033));
  nor2s1 ______508788(.DIN1 (___0____26064), .DIN2 (________25299), .Q
       (___9____26032));
  nnd2s1 _______508789(.DIN1 (________25384), .DIN2 (________23927), .Q
       (___9_0__26031));
  nnd2s1 _______508790(.DIN1 (________25258), .DIN2 (________25931), .Q
       (___9_9__26030));
  nnd2s1 _______508791(.DIN1 (____0___26234), .DIN2 (________22993), .Q
       (___9____26029));
  nnd2s1 _______508792(.DIN1 (________25298), .DIN2 (____0_0__34423),
       .Q (___9____26028));
  nor2s1 _______508793(.DIN1 (___0____25210), .DIN2 (___099__25221), .Q
       (___9____26027));
  or2s1 _______508794(.DIN1 (___9____26025), .DIN2 (________25386), .Q
       (___9____26026));
  and2s1 ______508795(.DIN1 (___9____26023), .DIN2 (___0____22295), .Q
       (___9____26024));
  nnd2s1 ______508796(.DIN1 (___9____26023), .DIN2 (_____0__22509), .Q
       (___9____26022));
  nnd2s1 _______508797(.DIN1 (___0____25211), .DIN2 (___9_9__26020), .Q
       (___9_0__26021));
  nor2s1 _______508798(.DIN1 (_________36762), .DIN2 (____0___26141),
       .Q (___9____26018));
  nor2s1 _______508799(.DIN1 (___0_9___40452), .DIN2 (________28994),
       .Q (___9____26017));
  nnd2s1 _______508800(.DIN1 (_____9___32965), .DIN2 (________28084),
       .Q (___9____26016));
  and2s1 _____9_508801(.DIN1 (____0___26231), .DIN2 (________24444), .Q
       (___9____26015));
  or2s1 _____0_508802(.DIN1 (_____0__29534), .DIN2 (________26300), .Q
       (___9____26014));
  nnd2s1 _____0_508803(.DIN1 (___9_____39206), .DIN2 (___0__0__40413),
       .Q (___9_0__26013));
  nor2s1 _____0_508804(.DIN1 (___9____26011), .DIN2 (___9____26010), .Q
       (___9_9__26012));
  nnd2s1 ___9___508805(.DIN1 (___90___25963), .DIN2 (___90___25964), .Q
       (___9____26009));
  xor2s1 _______508806(.DIN1 (___0_____40519), .DIN2 (___9_____39542),
       .Q (___9____26008));
  hi1s1 ___9_0_508807(.DIN (___9____26006), .Q (___9____26007));
  hi1s1 ___909_508808(.DIN (___9_0__26004), .Q (___9____26005));
  nnd2s1 _______508809(.DIN1 (___9____26002), .DIN2 (___9_0__25095), .Q
       (___9_9__26003));
  nor2s1 _______508810(.DIN1 (______9__22026), .DIN2 (___0_9__25212),
       .Q (___9____26001));
  nor2s1 _______508811(.DIN1 (___9____25999), .DIN2 (___0____26117), .Q
       (___9____26000));
  hi1s1 _______508812(.DIN (__9_____29873), .Q (___9____25998));
  hi1s1 ______508813(.DIN (_________32239), .Q (___9____25997));
  or2s1 _______508814(.DIN1 (___9____25994), .DIN2 (_____0__25901), .Q
       (___9____25995));
  hi1s1 _______508815(.DIN (___9____25992), .Q (___9____25993));
  xor2s1 _______508816(.DIN1 (______0___22057), .DIN2 (_________35526),
       .Q (___9____25991));
  nnd2s1 _______508817(.DIN1 (_________38435), .DIN2 (___9____23179),
       .Q (___9____25990));
  nor2s1 ___9___508818(.DIN1 (____99___36174), .DIN2 (___9_0__25988),
       .Q (___9____25989));
  nnd2s1 _______508819(.DIN1 (_____0__25262), .DIN2 (inData[4]), .Q
       (___9_9__25987));
  or2s1 _______508820(.DIN1 (________25430), .DIN2 (_________35186), .Q
       (___9____25986));
  hi1s1 ___9___508821(.DIN (_________41297), .Q (___9____25985));
  nnd2s1 ____9__508822(.DIN1 (___90___25965), .DIN2 (__9__0__30206), .Q
       (________26302));
  nnd2s1 _______508823(.DIN1 (___0_____31084), .DIN2 (_________41321),
       .Q (________26278));
  nnd2s1 _____9_508824(.DIN1 (____0___25228), .DIN2 (___9____25984), .Q
       (_____9__26285));
  nnd2s1 _____508825(.DIN1 (____9___25305), .DIN2 (________25825), .Q
       (________26277));
  nor2s1 _______508826(.DIN1 (________25929), .DIN2 (________25540), .Q
       (________26288));
  nnd2s1 _______508827(.DIN1 (______0__41366), .DIN2 (___90___25030),
       .Q (________26273));
  nor2s1 _______508828(.DIN1 (___9____25983), .DIN2 (___9____25982), .Q
       (_____9__26275));
  nor2s1 _____9_508829(.DIN1 (___0____26114), .DIN2 (___09___27917), .Q
       (____9___27386));
  hi1s1 ___9___508830(.DIN (________26344), .Q (_________31668));
  or2s1 _____9_508831(.DIN1 (___9____25981), .DIN2 (___09___27917), .Q
       (___9____26885));
  or2s1 _____9_508832(.DIN1 (___9____25980), .DIN2 (________25242), .Q
       (________26631));
  nnd2s1 _______508833(.DIN1 (________25924), .DIN2 (____90__25758), .Q
       (____0___26414));
  nnd2s1 _______508834(.DIN1 (____9___25301), .DIN2 (___0____26077), .Q
       (____0___26413));
  nnd2s1 _______508835(.DIN1 (________25601), .DIN2 (___9____25979), .Q
       (____0___28472));
  nor2s1 _______508836(.DIN1 (____9___25490), .DIN2 (___9_0__25978), .Q
       (___90___26867));
  nnd2s1 _______508837(.DIN1 (________25265), .DIN2 (___9_9__25977), .Q
       (________26736));
  nnd2s1 _______508838(.DIN1 (_____0___41317), .DIN2 (________25942),
       .Q (________26564));
  nnd2s1 _______508839(.DIN1 (___9____25976), .DIN2 (___9____25975), .Q
       (________26353));
  nnd2s1 _____0_508840(.DIN1 (________25264), .DIN2 (___9____25974), .Q
       (____9___26405));
  nnd2s1 _______508841(.DIN1 (____9___25951), .DIN2 (____9___25953), .Q
       (________26651));
  nnd2s1 _______508842(.DIN1 (___9____25973), .DIN2 (___9____25972), .Q
       (________26367));
  hi1s1 ______508843(.DIN (___9____25971), .Q (________26647));
  nnd2s1 _______508844(.DIN1 (________25277), .DIN2 (___0____26078), .Q
       (____0___26684));
  nor2s1 ______508845(.DIN1 (___9____25970), .DIN2 (___9____26927), .Q
       (____9___26404));
  nor2s1 _______508846(.DIN1 (___0__0__31080), .DIN2 (___0____25151),
       .Q (________26369));
  nnd2s1 _______508847(.DIN1 (___90___28649), .DIN2 (____9____32424),
       .Q (___0____28806));
  nor2s1 _______508848(.DIN1 (________26280), .DIN2 (________25245), .Q
       (________26741));
  or2s1 ______508849(.DIN1 (________25744), .DIN2 (___0____26104), .Q
       (____9___26585));
  nnd2s1 ____90_508850(.DIN1 (___9____25969), .DIN2 (_____9__27646), .Q
       (________26301));
  nnd2s1 _____9_508851(.DIN1 (________25446), .DIN2 (_____0__26418), .Q
       (_____0__26728));
  nor2s1 ______508852(.DIN1 (________29249), .DIN2 (_____0__26168), .Q
       (_____0__26626));
  or2s1 _______508853(.DIN1 (___9_0__25968), .DIN2 (___9____29606), .Q
       (________26602));
  hi1s1 ___9___508854(.DIN (________27468), .Q (____9___26677));
  nnd2s1 _______508855(.DIN1 (__90_9__29688), .DIN2 (_____9__24584), .Q
       (________27243));
  nnd2s1 ______508856(.DIN1 (___909__25967), .DIN2 (_____9__26737), .Q
       (__99____30525));
  hi1s1 ___9___508857(.DIN (_________32078), .Q (________26613));
  hi1s1 ___9___508858(.DIN (_________32755), .Q (________27179));
  hi1s1 _____508859(.DIN (___09___27920), .Q (________26753));
  and2s1 _______508860(.DIN1 (______0__41319), .DIN2 (___9____25062),
       .Q (________26629));
  nor2s1 _____0_508861(.DIN1 (________25737), .DIN2 (___0_0__26112), .Q
       (___9____26904));
  hi1s1 ____0__508862(.DIN (________28034), .Q (________27072));
  hi1s1 ____9__508863(.DIN (___90___25966), .Q (____0___26596));
  hi1s1 ____0__508864(.DIN (________28122), .Q (____0___26597));
  and2s1 ___9___508865(.DIN1 (___90___25965), .DIN2 (_____9__27646), .Q
       (________26693));
  nor2s1 ___9___508866(.DIN1 (____0___26590), .DIN2 (___0____25201), .Q
       (____99__26588));
  and2s1 ___9___508867(.DIN1 (___0____26095), .DIN2 (___0_____30958),
       .Q (________26627));
  nnd2s1 ___9___508868(.DIN1 (________25945), .DIN2 (________25355), .Q
       (________26600));
  nnd2s1 ___9___508869(.DIN1 (___0__9__30984), .DIN2 (___90___25964),
       .Q (________26612));
  nnd2s1 ___9__508870(.DIN1 (___90___25963), .DIN2 (___90___25962), .Q
       (________26710));
  nnd2s1 ___9_9_508871(.DIN1 (________25943), .DIN2 (___9_0__27795), .Q
       (________26298));
  nor2s1 _______508872(.DIN1
       (_____________________________________9_____), .DIN2
       (___90___25961), .Q (________26823));
  hi1s1 ____508873(.DIN (___90___25960), .Q (____0___26686));
  hi1s1 _______508874(.DIN (___90___25959), .Q (________27718));
  nor2s1 ___9__508875(.DIN1 (_____0__25556), .DIN2 (____0___25317), .Q
       (________26262));
  nnd2s1 ___9_9_508876(.DIN1 (________25450), .DIN2 (________24710), .Q
       (________26263));
  hi1s1 ___9___508877(.DIN (________27554), .Q (_____0__28210));
  nor2s1 ____9__508878(.DIN1 (___900__25958), .DIN2 (____0___25501), .Q
       (____0___26412));
  hi1s1 ____99_508879(.DIN (____99__25957), .Q (___0____27006));
  hi1s1 ____9__508880(.DIN (____9___25956), .Q (_____0__26608));
  nnd2s1 _______508881(.DIN1 (________25396), .DIN2 (____0___26415), .Q
       (________26735));
  nnd2s1 _______508882(.DIN1 (__90____29672), .DIN2 (________26523), .Q
       (______0__33984));
  nor2s1 _____9_508883(.DIN1 (________24659), .DIN2 (___0____25192), .Q
       (____0___27488));
  nor2s1 ____9__508884(.DIN1 (____9___25955), .DIN2 (_____0__25470), .Q
       (___0____27015));
  and2s1 ____9__508885(.DIN1 (____9___25954), .DIN2 (____9___25953), .Q
       (________29501));
  nor2s1 ____9__508886(.DIN1 (_____9__25575), .DIN2 (_________38177),
       .Q (______9__38245));
  nor2s1 ____9__508887(.DIN1 (____9___25952), .DIN2 (____00__27300), .Q
       (________28887));
  or2s1 ______508888(.DIN1 (________25263), .DIN2 (_________32903), .Q
       (___0_09__31127));
  nor2s1 ___90__508889(.DIN1 (________25571), .DIN2 (____0___25773), .Q
       (__9_____29777));
  nnd2s1 _______508890(.DIN1 (____0___25311), .DIN2 (________24798), .Q
       (___9_9__26929));
  nnd2s1 ____9__508891(.DIN1 (______________22104), .DIN2
       (______________________________________________21932), .Q
       (________27063));
  nnd2s1 _____0_508892(.DIN1 (_________33570), .DIN2 (___0090__30632),
       .Q (_____09__31999));
  hi1s1 ___9___508893(.DIN (_____0__27167), .Q (___09____31429));
  hi1s1 ___9___508894(.DIN (_____90__41299), .Q (____0____31566));
  nnd2s1 _____0_508895(.DIN1 (____9___25951), .DIN2 (___9____25979), .Q
       (________28573));
  hi1s1 ___9___508896(.DIN (_____0__27932), .Q (________26751));
  hi1s1 ___9__508897(.DIN (___9____26947), .Q (___00____30608));
  nnd2s1 _____0_508898(.DIN1 (____9___25950), .DIN2 (________25352), .Q
       (________26746));
  nnd2s1 _____0_508899(.DIN1 (_________38435), .DIN2 (____9___25949),
       .Q (____09___37180));
  nor2s1 ______508900(.DIN1 (___09___25214), .DIN2 (________27171), .Q
       (________27235));
  hi1s1 ___9___508901(.DIN (_____9__26727), .Q (_________31846));
  nor2s1 _______508902(.DIN1 (________25467), .DIN2 (________25295), .Q
       (___99___29629));
  nor2s1 ______508903(.DIN1 (___0____26117), .DIN2 (____0___27925), .Q
       (___99___28734));
  nor2s1 _______508904(.DIN1 (____90__25948), .DIN2 (________25240), .Q
       (____0___27396));
  nnd2s1 ____90_508905(.DIN1 (____9____32424), .DIN2 (inData[3]), .Q
       (________26574));
  nor2s1 _______508906(.DIN1 (___900__25958), .DIN2 (________25244), .Q
       (____9___26586));
  nor2s1 ______508907(.DIN1 (________25626), .DIN2 (____0____31591), .Q
       (________29158));
  nor2s1 _______508908(.DIN1 (___090__25213), .DIN2 (_____9__25947), .Q
       (________27709));
  nnd2s1 _______508909(.DIN1 (________25293), .DIN2 (___0____26077), .Q
       (________26732));
  and2s1 _______508910(.DIN1 (____9___25302), .DIN2 (___0____26077), .Q
       (________27246));
  nnd2s1 _______508911(.DIN1 (________28507), .DIN2 (________28533), .Q
       (________27511));
  and2s1 ___9___508912(.DIN1 (________25484), .DIN2 (________25944), .Q
       (__999___30543));
  nnd2s1 _______508913(.DIN1 (________25706), .DIN2 (____9___26862), .Q
       (____9___26676));
  nor2s1 ___9___508914(.DIN1 (___0____25188), .DIN2 (________25946), .Q
       (__9_____30204));
  nnd2s1 ___9__508915(.DIN1 (________25945), .DIN2 (________25944), .Q
       (___9____26900));
  nnd2s1 ___9___508916(.DIN1 (___9_____39743), .DIN2 (________23959),
       .Q (___9_____39657));
  nnd2s1 ___9___508917(.DIN1 (________25945), .DIN2 (________25373), .Q
       (__9_90__30169));
  nnd2s1 ___9___508918(.DIN1 (____9___25953), .DIN2 (____0___24752), .Q
       (___9_0__26901));
  nnd2s1 ___9___508919(.DIN1 (____9___28917), .DIN2 (________25943), .Q
       (___9_0__26883));
  nor2s1 _____508920(.DIN1 (inData[31]), .DIN2 (___99___25116), .Q
       (________26299));
  nnd2s1 ______508921(.DIN1 (________25296), .DIN2 (________25942), .Q
       (________29395));
  or2s1 _______508922(.DIN1 (___0____25153), .DIN2 (________29170), .Q
       (________27079));
  nnd2s1 _______508923(.DIN1 (________25567), .DIN2 (___0_9___31214),
       .Q (__9_____30016));
  hi1s1 ____99_508924(.DIN (________25941), .Q (____00___31505));
  nor2s1 _______508925(.DIN1 (_____9__25280), .DIN2 (________25940), .Q
       (____0___26595));
  hi1s1 ____0__508926(.DIN (________26422), .Q (__9_____30142));
  hi1s1 ____0__508927(.DIN (___9_0__26911), .Q (________29319));
  nor2s1 ____9__508928(.DIN1 (________24703), .DIN2 (___0____25191), .Q
       (_____9__27498));
  nnd2s1 ____9__508929(.DIN1 (________25511), .DIN2 (___0____26077), .Q
       (________28982));
  hi1s1 ____0__508930(.DIN (________29053), .Q (___0_____31182));
  hi1s1 ____0__508931(.DIN (____0___27926), .Q (___9____27772));
  and2s1 _____9_508932(.DIN1 (________25419), .DIN2 (___0____26078), .Q
       (___9_9__27767));
  nor2s1 _____9_508933(.DIN1 (____0___26590), .DIN2 (________25288), .Q
       (_____0___31803));
  nor2s1 ______508934(.DIN1 (___99___26045), .DIN2 (________25274), .Q
       (__9_00__30272));
  nor2s1 _____9_508935(.DIN1 (__9__9__29751), .DIN2 (_____0__27270), .Q
       (____0____31581));
  nor2s1 _______508936(.DIN1 (________27288), .DIN2 (________25284), .Q
       (___0_____31282));
  or2s1 _____508937(.DIN1 (________28318), .DIN2 (________25939), .Q
       (________29431));
  and2s1 ____9__508938(.DIN1 (___0__0__30787), .DIN2 (________26240),
       .Q (___0_99__30926));
  nor2s1 ____9_508939(.DIN1 (____0___26409), .DIN2 (____9___25399), .Q
       (________29326));
  nnd2s1 ______508940(.DIN1 (_____0__25938), .DIN2 (_____0__24849), .Q
       (_________33986));
  nnd2s1 ____9__508941(.DIN1 (_____9__25937), .DIN2 (________25454), .Q
       (__9_____30208));
  nnd2s1 ____9_508942(.DIN1 (________25936), .DIN2 (________25935), .Q
       (________28046));
  nor2s1 _______508943(.DIN1 (________26421), .DIN2 (________25934), .Q
       (___0_____31277));
  nor2s1 _______508944(.DIN1 (________26433), .DIN2 (________25934), .Q
       (________28153));
  nnd2s1 _______508945(.DIN1 (_____9__25290), .DIN2 (________26426), .Q
       (___0_____30943));
  nor2s1 ____90_508946(.DIN1 (________25933), .DIN2 (____9___29544), .Q
       (___0__9__31299));
  nor2s1 ___9___508947(.DIN1 (___0____25207), .DIN2 (___9_0__25978), .Q
       (_________32815));
  or2s1 ____508948(.DIN1 (___0_____31345), .DIN2 (________25932), .Q
       (________29233));
  nnd2s1 _______508949(.DIN1 (____0___25226), .DIN2 (___9____26912), .Q
       (_________31678));
  nnd2s1 _______508950(.DIN1 (_____9__25261), .DIN2 (________25931), .Q
       (_____9__27551));
  nnd2s1 _______508951(.DIN1 (________25598), .DIN2 (___0____26061), .Q
       (____0____33491));
  nnd2s1 ______508952(.DIN1 (_____0__25291), .DIN2
       (_____________________21744), .Q (__9_____30241));
  or2s1 _______508953(.DIN1 (________26174), .DIN2 (_____9__25452), .Q
       (_____0___31609));
  nnd2s1 ____90_508954(.DIN1 (_____0__25281), .DIN2 (________23449), .Q
       (___0_____30676));
  nnd2s1 _______508955(.DIN1 (________25630), .DIN2 (____0____31554),
       .Q (___0990__31494));
  nor2s1 _______508956(.DIN1 (_____9__25947), .DIN2 (___9____25088), .Q
       (________27989));
  hi1s1 ____0__508957(.DIN (_________41291), .Q (___0____27842));
  nnd2s1 ____9__508958(.DIN1 (___9____25090), .DIN2 (___0____26094), .Q
       (___0__9__31147));
  nnd2s1 _______508959(.DIN1 (____0___25499), .DIN2 (___9____25984), .Q
       (_____9__27967));
  nnd2s1 ___9___508960(.DIN1 (________25945), .DIN2 (___0____25176), .Q
       (____0____33459));
  nor2s1 ____9__508961(.DIN1 (_____0__25461), .DIN2 (________27058), .Q
       (___09___28825));
  nnd2s1 ____9_508962(.DIN1 (________25442), .DIN2 (________26611), .Q
       (________27495));
  nnd2s1 ____9__508963(.DIN1 (_________38435), .DIN2 (________25930),
       .Q (_________38550));
  nnd2s1 _____9_508964(.DIN1 (___0____25195), .DIN2 (___0____26077), .Q
       (_____0__29175));
  nnd2s1 _____9_508965(.DIN1 (________25279), .DIN2 (___0____26078), .Q
       (_____9___31697));
  nor2s1 _____9_508966(.DIN1 (________25929), .DIN2 (_____0__25928), .Q
       (____0___29011));
  dffacs1 _________________________________________0_____508967(.CLRB
       (reset), .CLK (clk), .DIN (___09___25217), .Q (___0_0___40567));
  nor2s1 _______508968(.DIN1 (________25440), .DIN2 (________25383), .Q
       (________29531));
  hi1s1 _______508969(.DIN (_____0__26617), .Q (___9____27800));
  nor2s1 _______508970(.DIN1 (_____9__25927), .DIN2 (________25421), .Q
       (___9_9___39611));
  nor2s1 _______508971(.DIN1 (___9_0__25068), .DIN2 (____99__25309), .Q
       (________28600));
  nnd2s1 _______508972(.DIN1 (___0____25197), .DIN2 (________25749), .Q
       (___0_____30810));
  nor2s1 _______508973(.DIN1 (_____0__26247), .DIN2 (________25459), .Q
       (__9_0___29995));
  nnd2s1 _______508974(.DIN1 (___09___25220), .DIN2 (________25740), .Q
       (___0__0__31003));
  hi1s1 ___9___508975(.DIN (________25926), .Q (_________31866));
  nnd2s1 ______508976(.DIN1 (____09__25230), .DIN2 (________25925), .Q
       (_________31973));
  nor2s1 _______508977(.DIN1 (_____________________21691), .DIN2
       (________25256), .Q (________29359));
  nnd2s1 ______508978(.DIN1 (________25543), .DIN2 (_____0__25748), .Q
       (________29311));
  hi1s1 ____0__508979(.DIN (___0__9__40098), .Q (___0__9__40158));
  nnd2s1 ____9__508980(.DIN1 (________25481), .DIN2 (____90__25489), .Q
       (_________31731));
  nor2s1 ____9__508981(.DIN1 (________26280), .DIN2 (________25474), .Q
       (___090___31413));
  nor2s1 ____9_508982(.DIN1 (________24279), .DIN2 (________25420), .Q
       (_________37538));
  hi1s1 ___9_9_508983(.DIN (_________31715), .Q (_____9___32376));
  hi1s1 ___9_508984(.DIN (________26261), .Q (____9____33350));
  hi1s1 ___9_9_508985(.DIN (______0__34524), .Q (_________33897));
  nnd2s1 ____9__508986(.DIN1 (________25924), .DIN2 (________23915), .Q
       (____0___29010));
  hi1s1 ______508987(.DIN (______0__41289), .Q (___90____39008));
  nnd2s1 _____508988(.DIN1 (________25287), .DIN2 (________25923), .Q
       (_________31879));
  hi1s1 ____0__508989(.DIN (___0____27012), .Q (_________32058));
  nor2s1 ______508990(.DIN1 (_____9__25019), .DIN2 (________25884), .Q
       (____0____32521));
  nnd2s1 ____9__508991(.DIN1 (________25480), .DIN2 (____9___27298), .Q
       (__9_____30162));
  nor2s1 _____0_508992(.DIN1 (_________32159), .DIN2 (___99___25116),
       .Q (____0____32543));
  nnd2s1 _______508993(.DIN1 (________24919), .DIN2 (________24511), .Q
       (________25922));
  nor2s1 ____09_508994(.DIN1 (________25007), .DIN2 (________25920), .Q
       (________25921));
  nor2s1 _____9_508995(.DIN1 (________23563), .DIN2 (________25723), .Q
       (________25919));
  hi1s1 ___9__508996(.DIN (____9_0__32391), .Q (_____0__25918));
  xor2s1 _______508997(.DIN1 (________22576), .DIN2 (_________38871),
       .Q (_____9__25917));
  nor2s1 _____0_508998(.DIN1 (________24718), .DIN2 (____9___24831), .Q
       (________25916));
  xor2s1 _______508999(.DIN1 (___0_____40487), .DIN2 (_________38573),
       .Q (________25915));
  xor2s1 _______509000(.DIN1 (_________41341), .DIN2 (_____0___32287),
       .Q (________25914));
  nor2s1 _______509001(.DIN1 (_____9__25555), .DIN2 (_____0__25815), .Q
       (________25913));
  nnd2s1 _______509002(.DIN1 (____9___24933), .DIN2 (____9____38898),
       .Q (________25912));
  and2s1 _____509003(.DIN1 (_____0__24991), .DIN2 (____0___26410), .Q
       (________25911));
  and2s1 _______509004(.DIN1 (___9_____39539), .DIN2
       (_____________________________________________21810), .Q
       (________25910));
  nnd2s1 _____9_509005(.DIN1 (_________35435), .DIN2 (_________33973),
       .Q (_____0__25909));
  nnd2s1 ______509006(.DIN1 (___9_9__25077), .DIN2 (___9_9__25977), .Q
       (_____9__25908));
  nnd2s1 _______509007(.DIN1 (________25525), .DIN2 (____00__22549), .Q
       (________25907));
  nnd2s1 _______509008(.DIN1 (_________35186), .DIN2
       (_________________________________________________________________________________________22090),
       .Q (________25906));
  nor2s1 ______509009(.DIN1 (_____9__23665), .DIN2 (____0___25770), .Q
       (________25905));
  nnd2s1 _______509010(.DIN1 (________24862), .DIN2
       (____0_______________), .Q (________25904));
  nor2s1 _______509011(.DIN1 (_____0__25901), .DIN2 (_____9__25900), .Q
       (________25902));
  or2s1 _______509012(.DIN1 (________25898), .DIN2 (________25897), .Q
       (________25899));
  or2s1 _______509013(.DIN1 (____0___24273), .DIN2 (_____0___34932), .Q
       (________25896));
  nnd2s1 _______509014(.DIN1 (___9____25050), .DIN2 (___9____25042), .Q
       (________25895));
  nnd2s1 _______509015(.DIN1 (___9____25061), .DIN2 (________22694), .Q
       (________25894));
  nor2s1 _______509016(.DIN1 (___999), .DIN2 (____9___24930), .Q
       (________25893));
  xor2s1 _______509017(.DIN1 (_____9___36721), .DIN2 (_____9___38412),
       .Q (_____0__25892));
  hi1s1 _______509018(.DIN (___0____26093), .Q (_____9__25891));
  nor2s1 _______509019(.DIN1 (___9____25066), .DIN2 (________25448), .Q
       (________25890));
  nnd2s1 _______509020(.DIN1 (_________38743), .DIN2 (________23544),
       .Q (________25889));
  or2s1 _______509021(.DIN1 (____09__26331), .DIN2 (________24854), .Q
       (________25888));
  nnd2s1 _______509022(.DIN1 (________24981), .DIN2 (___9____23197), .Q
       (________25887));
  nor2s1 _______509023(.DIN1 (________25438), .DIN2 (________24815), .Q
       (________25886));
  hi1s1 ______509024(.DIN (________25884), .Q (________25885));
  nor2s1 ______509025(.DIN1 (________22381), .DIN2 (_____0__25729), .Q
       (________25883));
  nnd2s1 _______509026(.DIN1 (______9__37419), .DIN2 (________22506),
       .Q (_____0__25882));
  nnd2s1 ______509027(.DIN1 (______9__37419), .DIN2 (___9__), .Q
       (_____9__25881));
  nnd2s1 _______509028(.DIN1 (______9__37419), .DIN2 (_______22176), .Q
       (________25880));
  nnd2s1 ____0_509029(.DIN1 (___9____25074), .DIN2 (________25878), .Q
       (________25879));
  and2s1 ____0__509030(.DIN1 (___9____25103), .DIN2 (____9____38898),
       .Q (________25877));
  or2s1 ____0_509031(.DIN1 (___90____39040), .DIN2 (________25015), .Q
       (________25876));
  nnd2s1 ____0__509032(.DIN1 (_____9__24990), .DIN2 (________24978), .Q
       (________25875));
  nnd2s1 _______509033(.DIN1 (_________35394), .DIN2 (_________36761),
       .Q (________25874));
  nor2s1 _______509034(.DIN1 (___00___23218), .DIN2 (____9___25026), .Q
       (________25873));
  nnd2s1 _______509035(.DIN1 (____00__24935), .DIN2 (____09__25871), .Q
       (_____0__25872));
  nnd2s1 ______509036(.DIN1 (___9_0__25048), .DIN2 (____9___24360), .Q
       (____0___25870));
  nnd2s1 _______509037(.DIN1 (________24781), .DIN2 (_________33596),
       .Q (____0___25869));
  xor2s1 _______509038(.DIN1 (________24577), .DIN2 (___9_____39461),
       .Q (____0___25868));
  nor2s1 _______509039(.DIN1 (________24824), .DIN2 (________24871), .Q
       (____0___25867));
  nor2s1 _______509040(.DIN1 (_____________________21748), .DIN2
       (________25743), .Q (____0___25866));
  or2s1 _______509041(.DIN1
       (____________________________________________21864), .DIN2
       (____009__38047), .Q (____0___25865));
  nor2s1 ______509042(.DIN1 (_________41345), .DIN2 (________25014), .Q
       (____0___25864));
  xor2s1 _______509043(.DIN1
       (____________________________________________21830), .DIN2
       (__9_____29971), .Q (____0___25863));
  nnd2s1 _____9_509044(.DIN1 (_________41335), .DIN2 (________24966),
       .Q (____00__25862));
  nor2s1 ______509045(.DIN1 (____9___25860), .DIN2 (________25822), .Q
       (____99__25861));
  nnd2s1 _______509046(.DIN1 (____9___24931), .DIN2 (____0___25498), .Q
       (____9___25859));
  nnd2s1 _____509047(.DIN1 (________24850), .DIN2 (________24697), .Q
       (____9___25858));
  nnd2s1 _______509048(.DIN1 (_________38743), .DIN2 (_____0__23359),
       .Q (____9___25857));
  and2s1 _______509049(.DIN1 (_____0__26428), .DIN2 (_________22014),
       .Q (____9___25856));
  nor2s1 _______509050(.DIN1 (_____00__33066), .DIN2 (____9___25854),
       .Q (____9___25855));
  and2s1 _______509051(.DIN1 (_________36955), .DIN2 (______22158), .Q
       (____9___25853));
  nor2s1 _______509052(.DIN1 (________24956), .DIN2 (________25011), .Q
       (____90__25852));
  nor2s1 _____509053(.DIN1 (________25850), .DIN2 (___9____25112), .Q
       (_____9__25851));
  and2s1 _____9_509054(.DIN1 (_____9__28617), .DIN2 (___09), .Q
       (________25849));
  nnd2s1 ______509055(.DIN1 (________24980), .DIN2 (_____0___37283), .Q
       (________25848));
  nnd2s1 _______509056(.DIN1 (____0___24942), .DIN2 (________22566), .Q
       (________25847));
  or2s1 _______509057(.DIN1 (___0_____40438), .DIN2 (_____9__25795), .Q
       (________25846));
  or2s1 _______509058(.DIN1
       (______________________________________0_______21889), .DIN2
       (_____9__28617), .Q (________25845));
  or2s1 _______509059(.DIN1 (___0_9___40455), .DIN2 (_________38743),
       .Q (________25844));
  nor2s1 ______509060(.DIN1 (____9___25955), .DIN2 (________25548), .Q
       (________25843));
  nnd2s1 _____9_509061(.DIN1 (________25739), .DIN2 (________24625), .Q
       (_____0__25842));
  nor2s1 _____0_509062(.DIN1 (________23742), .DIN2 (________24967), .Q
       (_____9__25841));
  and2s1 _______509063(.DIN1 (_________33769), .DIN2 (_________22014),
       .Q (________25840));
  nor2s1 ______509064(.DIN1 (________25838), .DIN2 (_____9__25738), .Q
       (________25839));
  or2s1 _____509065(.DIN1 (____0___23794), .DIN2 (____9___24932), .Q
       (________25837));
  or2s1 _______509066(.DIN1 (________23914), .DIN2 (________25016), .Q
       (________25836));
  and2s1 _______509067(.DIN1 (___0____27013), .DIN2 (________25834), .Q
       (________25835));
  and2s1 _______509068(.DIN1 (________25792), .DIN2 (___0_____40621),
       .Q (________25833));
  nnd2s1 ______509069(.DIN1 (___9____25080), .DIN2 (________25726), .Q
       (_____0__25832));
  nnd2s1 _______509070(.DIN1 (________24874), .DIN2 (________25829), .Q
       (________25830));
  nor2s1 _______509071(.DIN1 (________26440), .DIN2 (___9____25111), .Q
       (________25828));
  nnd2s1 _______509072(.DIN1 (________24809), .DIN2 (inData[10]), .Q
       (________25827));
  nnd2s1 _______509073(.DIN1 (___9_0__25078), .DIN2 (________25825), .Q
       (________25826));
  nor2s1 ______509074(.DIN1 (_____9__25823), .DIN2 (________25822), .Q
       (_____0__25824));
  hi1s1 _______509075(.DIN (________29173), .Q (________25821));
  hi1s1 ______509076(.DIN (________25819), .Q (________25820));
  hi1s1 _______509077(.DIN (________25817), .Q (________25818));
  nor2s1 _______509078(.DIN1 (________25742), .DIN2 (_____0__25815), .Q
       (________25816));
  and2s1 _______509079(.DIN1 (________24979), .DIN2 (________25813), .Q
       (_____9__25814));
  and2s1 ______509080(.DIN1 (________25811), .DIN2 (____9___22641), .Q
       (________25812));
  nnd2s1 _______509081(.DIN1 (________25754), .DIN2 (_____9__25469), .Q
       (________25810));
  nor2s1 _______509082(.DIN1 (____00__23881), .DIN2 (________24946), .Q
       (________25809));
  and2s1 _______509083(.DIN1 (________25807), .DIN2 (________25552), .Q
       (________25808));
  nnd2s1 _______509084(.DIN1 (________25321), .DIN2 (________24948), .Q
       (_____0__25806));
  nnd2s1 _______509085(.DIN1 (___9____25073), .DIN2 (___9____24114), .Q
       (_____9__25805));
  xor2s1 ______509086(.DIN1 (_________38372), .DIN2 (____9_9__38931),
       .Q (________25804));
  nnd2s1 _______509087(.DIN1 (____0___25772), .DIN2 (_____0__23748), .Q
       (________25803));
  or2s1 _____9_509088(.DIN1 (____0____33465), .DIN2 (_____9__26812), .Q
       (________25802));
  nnd2s1 ______509089(.DIN1 (________25800), .DIN2
       (_____________________________________9_______21883), .Q
       (________25801));
  nor2s1 ______509090(.DIN1 (___0____26067), .DIN2 (_____0__25815), .Q
       (________25799));
  nnd2s1 _____0_509091(.DIN1 (____09__25506), .DIN2 (________25797), .Q
       (________25798));
  nor2s1 ______509092(.DIN1 (___0_____40437), .DIN2 (_____9__25795), .Q
       (_____0__25796));
  nor2s1 _______509093(.DIN1
       (______________________________________________21913), .DIN2
       (_____9__25795), .Q (________25794));
  or2s1 _______509094(.DIN1 (___0_____40621), .DIN2 (________25792), .Q
       (________25793));
  nnd2s1 _______509095(.DIN1 (___9____25044), .DIN2 (________24328), .Q
       (________25791));
  nnd2s1 _______509096(.DIN1 (________24918), .DIN2 (inData[26]), .Q
       (________25790));
  nnd2s1 _______509097(.DIN1 (___9____25043), .DIN2 (________25925), .Q
       (________25789));
  or2s1 _______509098(.DIN1 (________25787), .DIN2 (____0___26687), .Q
       (________25788));
  nnd2s1 _______509099(.DIN1 (_____9__25785), .DIN2 (________23110), .Q
       (_____0__25786));
  nor2s1 _______509100(.DIN1 (________25783), .DIN2 (___0____26096), .Q
       (________25784));
  nnd2s1 _______509101(.DIN1 (____0___24943), .DIN2 (_____9__24021), .Q
       (________25782));
  nor2s1 _______509102(.DIN1 (____9____34341), .DIN2 (________24913),
       .Q (________25781));
  nnd2s1 _______509103(.DIN1 (____0___24938), .DIN2 (________24023), .Q
       (________25780));
  nnd2s1 _____509104(.DIN1 (________24951), .DIN2 (___9____25108), .Q
       (________25779));
  nor2s1 _____509105(.DIN1 (___9____25084), .DIN2 (___9____25072), .Q
       (____09__25777));
  nnd2s1 _____0_509106(.DIN1 (________29441), .DIN2 (____0___25775), .Q
       (____0___25776));
  and2s1 _______509107(.DIN1 (________25752), .DIN2 (____0___25774), .Q
       (_____0__26508));
  hi1s1 __90__0(.DIN (____0___25773), .Q (________26270));
  nnd2s1 ______509108(.DIN1 (____0___25772), .DIN2 (________24771), .Q
       (________25941));
  hi1s1 ___9___509109(.DIN (___0090__30632), .Q (___9_0__26920));
  nor2s1 _______509110(.DIN1 (____0___25771), .DIN2 (____0___25770), .Q
       (___90___25960));
  nnd2s1 _______509111(.DIN1 (___9____25075), .DIN2 (________26272), .Q
       (___90___25966));
  nnd2s1 _______509112(.DIN1 (___90___28649), .DIN2 (____0___27398), .Q
       (____9___25956));
  nnd2s1 ______509113(.DIN1 (________24999), .DIN2 (________25825), .Q
       (____09__27489));
  or2s1 _______509114(.DIN1 (____0___25769), .DIN2 (____00__25768), .Q
       (___9____26938));
  hi1s1 __90__509115(.DIN (____99__25767), .Q (_____0__29227));
  or2s1 _______509116(.DIN1 (________25783), .DIN2 (__909___29720), .Q
       (________26561));
  nnd2s1 _______509117(.DIN1 (________28230), .DIN2 (___90___28653), .Q
       (________28094));
  hi1s1 _____9_509118(.DIN (__9__9__29849), .Q (________26475));
  hi1s1 ___9___509119(.DIN (___9____27782), .Q (____9___26402));
  nor2s1 _____9_509120(.DIN1 (___0_____31324), .DIN2 (___09____31451),
       .Q (________26439));
  or2s1 ______509121(.DIN1 (________24923), .DIN2 (____9___25766), .Q
       (_____0__26448));
  or2s1 ______509122(.DIN1 (__9_____30400), .DIN2 (____9___25765), .Q
       (____9___26494));
  nor2s1 _______509123(.DIN1 (________26174), .DIN2 (___9____25071), .Q
       (____0___26144));
  and2s1 ______509124(.DIN1 (____9___25764), .DIN2 (____9___25763), .Q
       (___0_____31258));
  nor2s1 _______509125(.DIN1 (____9___26680), .DIN2 (____9___25762), .Q
       (___0____26070));
  nnd2s1 _____9_509126(.DIN1 (_________38743), .DIN2 (___0_9__22306),
       .Q (________26458));
  or2s1 _______509127(.DIN1 (____9___25761), .DIN2 (_____9___31789), .Q
       (________26423));
  nor2s1 _______509128(.DIN1 (____9___25760), .DIN2 (____9___25759), .Q
       (________26453));
  nor2s1 _______509129(.DIN1 (_________41351), .DIN2 (____9___25580),
       .Q (________26802));
  nnd2s1 _______509130(.DIN1 (____0_9__33489), .DIN2 (___9____25054),
       .Q (________26472));
  nor2s1 _______509131(.DIN1 (________25337), .DIN2 (___9____25109), .Q
       (____09__26417));
  nnd2s1 _______509132(.DIN1 (____9___24929), .DIN2 (____0____37167),
       .Q (________26190));
  nnd2s1 _______509133(.DIN1 (________24961), .DIN2 (____90__25758), .Q
       (____0___26416));
  hi1s1 _______509134(.DIN (___0____27863), .Q (____09__26598));
  nnd2s1 _______509135(.DIN1 (_____9__25757), .DIN2 (________26151), .Q
       (___0____26118));
  nor2s1 _______509136(.DIN1 (________25756), .DIN2 (________24970), .Q
       (___90___25959));
  nnd2s1 _______509137(.DIN1 (____9____33362), .DIN2 (_________33016),
       .Q (___0____26126));
  hi1s1 _______509138(.DIN (________25755), .Q (________26292));
  nnd2s1 _______509139(.DIN1 (________24855), .DIN2 (________26267), .Q
       (________26420));
  nnd2s1 _______509140(.DIN1 (_____0__24965), .DIN2 (_____0__24775), .Q
       (___0____26103));
  nnd2s1 _______509141(.DIN1 (________24858), .DIN2 (________22953), .Q
       (___0_0__26069));
  or2s1 _______509142(.DIN1 (___9____25974), .DIN2 (________24992), .Q
       (_____0__26738));
  nnd2s1 _______509143(.DIN1 (_____9__24477), .DIN2 (________25754), .Q
       (___0____26084));
  nnd2s1 ____9__509144(.DIN1 (___990__25115), .DIN2 (________26267), .Q
       (___0____26086));
  hi1s1 _______509145(.DIN (________25753), .Q (__9_9___29986));
  nnd2s1 _______509146(.DIN1 (________25752), .DIN2 (________25751), .Q
       (___09___27920));
  nnd2s1 _____9_509147(.DIN1 (___9____25113), .DIN2 (________26258), .Q
       (________26435));
  xor2s1 _______509148(.DIN1 (________24332), .DIN2 (________22788), .Q
       (________26360));
  nor2s1 _______509149(.DIN1 (___00___26054), .DIN2 (___9____25069), .Q
       (________26425));
  dffacs1 ______________________________________509150(.CLRB (reset),
       .CLK (clk), .DIN (________24859), .Q (_____________22098));
  nor2s1 ______509151(.DIN1 (________26433), .DIN2 (___9____25045), .Q
       (__9_____29754));
  nor2s1 _______509152(.DIN1 (________25356), .DIN2 (___9____25055), .Q
       (___9____26917));
  nor2s1 ___9___509153(.DIN1 (________24968), .DIN2 (_____9__24774), .Q
       (___0____27873));
  nor2s1 _______509154(.DIN1 (__9_____30335), .DIN2 (___0____25148), .Q
       (________26520));
  nor2s1 _______509155(.DIN1 (____9____35264), .DIN2 (_________35394),
       .Q (________26514));
  dffacs1 _______________________________________________509156(.CLRB
       (reset), .CLK (clk), .DIN (____99__24838), .Q
       (__________________________________________________________________22005));
  nnd2s1 _______509157(.DIN1 (___9_0__25105), .DIN2 (________25750), .Q
       (_____0__27578));
  hi1s1 _______509158(.DIN (_____0__26168), .Q (____9___28922));
  and2s1 _____0_509159(.DIN1 (____0___25772), .DIN2 (________24630), .Q
       (________26764));
  nnd2s1 ______509160(.DIN1 (_____0__24955), .DIN2 (____0___26146), .Q
       (________29043));
  nor2s1 ______509161(.DIN1 (_________41351), .DIN2 (________29354), .Q
       (____0___26506));
  nnd2s1 _______509162(.DIN1 (________25012), .DIN2 (____9___27298), .Q
       (___9____26925));
  nnd2s1 _______509163(.DIN1 (_________38743), .DIN2 (___0____26098),
       .Q (_________38638));
  and2s1 _____509164(.DIN1 (____9___26317), .DIN2 (_____0__25369), .Q
       (________26532));
  nnd2s1 _______509165(.DIN1 (_____90__32080), .DIN2 (___0_____31366),
       .Q (________29409));
  nnd2s1 _____0_509166(.DIN1 (________27505), .DIN2 (____0___25224), .Q
       (________29256));
  nnd2s1 ______509167(.DIN1 (________24949), .DIN2 (________25925), .Q
       (__9__9__30063));
  xor2s1 _______509168(.DIN1 (________24573), .DIN2 (________24668), .Q
       (___0_09__30841));
  nor2s1 ______509169(.DIN1 (______0__41329), .DIN2 (___0_____30798),
       .Q (_____0__26276));
  hi1s1 ___9___509170(.DIN (___9____27773), .Q (____0_0__32518));
  and2s1 _____0_509171(.DIN1 (___0_0__26092), .DIN2 (___00___27828), .Q
       (_____0__29417));
  nnd2s1 _____509172(.DIN1 (____0___25772), .DIN2 (____0___25229), .Q
       (________28612));
  nnd2s1 _______509173(.DIN1 (____0___25772), .DIN2 (________25375), .Q
       (___9____26921));
  nnd2s1 _______509174(.DIN1 (_____9__24866), .DIN2 (________25749), .Q
       (____9___26587));
  nnd2s1 _______509175(.DIN1 (_____0__25748), .DIN2 (____90__25020), .Q
       (________26422));
  nor2s1 _______509176(.DIN1 (_________32311), .DIN2 (____0___25769),
       .Q (________29341));
  nnd2s1 _______509177(.DIN1 (_____9__25747), .DIN2 (____0___26690), .Q
       (________27627));
  nor2s1 _______509178(.DIN1 (________25929), .DIN2 (___9____25096), .Q
       (________27261));
  nor2s1 _____509179(.DIN1 (___0____26087), .DIN2 (________25822), .Q
       (________26442));
  or2s1 _______509180(.DIN1 (____0____33496), .DIN2 (________25746), .Q
       (__9_____29932));
  nor2s1 _______509181(.DIN1 (________25260), .DIN2 (________24960), .Q
       (___0_____30801));
  nor2s1 _______509182(.DIN1 (___9____25974), .DIN2 (___9____25041), .Q
       (__9_____29773));
  nnd2s1 ______509183(.DIN1 (________24962), .DIN2 (___0____26078), .Q
       (________27494));
  nor2s1 _______509184(.DIN1 (________25745), .DIN2 (________24986), .Q
       (_____9__27138));
  or2s1 _______509185(.DIN1 (________25744), .DIN2 (________25743), .Q
       (___0_____30979));
  nor2s1 _______509186(.DIN1 (________25742), .DIN2 (_____0__25001), .Q
       (__909___29721));
  nnd2s1 _______509187(.DIN1 (________25515), .DIN2 (________24998), .Q
       (__9_____30058));
  nnd2s1 _______509188(.DIN1 (________25727), .DIN2 (____9___24449), .Q
       (____0___27926));
  and2s1 _______509189(.DIN1 (_____0__25243), .DIN2 (____0___25774), .Q
       (________28866));
  hi1s1 _______509190(.DIN (________25741), .Q (__9_0___29899));
  nor2s1 _______509191(.DIN1 (________24814), .DIN2 (____90__25948), .Q
       (___0_____31164));
  hi1s1 _______509192(.DIN (_________31749), .Q (________29110));
  nnd2s1 _______509193(.DIN1 (________24911), .DIN2 (________25931), .Q
       (________28484));
  hi1s1 ___9___509194(.DIN (_____0__25938), .Q (_____0___33821));
  nnd2s1 _______509195(.DIN1 (_________38377), .DIN2 (__90_0__29699),
       .Q (______0__37731));
  nor2s1 _____0_509196(.DIN1 (___9____25053), .DIN2 (_____9__25900), .Q
       (____999__33432));
  and2s1 _______509197(.DIN1 (________24806), .DIN2 (________25923), .Q
       (________27220));
  nor2s1 _______509198(.DIN1 (_____0___38616), .DIN2 (________25800),
       .Q (_________38787));
  nnd2s1 _____9_509199(.DIN1 (____9___25579), .DIN2 (________25740), .Q
       (________29533));
  nnd2s1 _____9_509200(.DIN1 (________24953), .DIN2 (________25605), .Q
       (___0_00__30740));
  and2s1 ______509201(.DIN1 (________25739), .DIN2 (___9____25110), .Q
       (__9_9___29991));
  or2s1 _____9_509202(.DIN1 (_________33217), .DIN2 (________25746), .Q
       (___0_____31194));
  nor2s1 ______509203(.DIN1 (___99___25122), .DIN2 (________26666), .Q
       (___0_00__31216));
  or2s1 _____9_509204(.DIN1 (________25831), .DIN2 (_________34644), .Q
       (____9____34338));
  nnd2s1 _______509205(.DIN1 (_____9__26765), .DIN2 (_____9__25738), .Q
       (_________38253));
  and2s1 _______509206(.DIN1 (____09__24944), .DIN2 (____9___26316), .Q
       (____09__28931));
  nor2s1 _______509207(.DIN1 (________25737), .DIN2 (________25736), .Q
       (___0____28822));
  nor2s1 _____0_509208(.DIN1 (___9____25092), .DIN2 (________29088), .Q
       (____9___28198));
  and2s1 ______509209(.DIN1 (___9_0__25058), .DIN2 (____0___25774), .Q
       (___09___27915));
  nor2s1 _______509210(.DIN1 (________25735), .DIN2 (________25734), .Q
       (________26840));
  nor2s1 ____9__509211(.DIN1 (________26309), .DIN2 (___9_0__25038), .Q
       (___9____29608));
  nor2s1 ____9__509212(.DIN1 (_____9__25434), .DIN2 (________25734), .Q
       (_________31906));
  nnd2s1 ____9__509213(.DIN1 (________26430), .DIN2 (________25733), .Q
       (___00____30625));
  nnd2s1 ____9_509214(.DIN1 (____0___25500), .DIN2 (____0___25774), .Q
       (_________31811));
  nnd2s1 ______509215(.DIN1 (________24795), .DIN2 (________25749), .Q
       (________27526));
  nnd2s1 ____9__509216(.DIN1 (________24958), .DIN2 (________25640), .Q
       (_________31725));
  xor2s1 _______509217(.DIN1 (________24513), .DIN2
       (______________22066), .Q (___9____27758));
  nnd2s1 _______509218(.DIN1 (___9____25070), .DIN2 (___9____25984), .Q
       (___9____27766));
  nnd2s1 ____9__509219(.DIN1 (________25732), .DIN2 (________25731), .Q
       (_________33742));
  nnd2s1 _______509220(.DIN1 (________24810), .DIN2 (________25564), .Q
       (___90___28651));
  hi1s1 _____0_509221(.DIN (________25730), .Q (____9___28196));
  nor2s1 _______509222(.DIN1 (________25324), .DIN2 (_____0__25729), .Q
       (_________31827));
  nnd2s1 ______509223(.DIN1 (________24996), .DIN2 (_____9__24793), .Q
       (________29140));
  nor2s1 ____9__509224(.DIN1 (_____9__25728), .DIN2 (________24921), .Q
       (__90____29692));
  nor2s1 ____9__509225(.DIN1 (________27288), .DIN2 (____9___25021), .Q
       (________28441));
  nor2s1 ____9__509226(.DIN1 (____0___26409), .DIN2 (_________41325),
       .Q (__9_____29750));
  nor2s1 ____9__509227(.DIN1 (________25360), .DIN2 (________25734), .Q
       (_________33580));
  dffacs1 ______________________________________509228(.CLRB (reset),
       .CLK (clk), .DIN (____9___25025), .Q (_____________22101));
  nnd2s1 ____9__509229(.DIN1 (________25727), .DIN2 (_____9__24675), .Q
       (_____0__28481));
  nor2s1 ____9__509230(.DIN1 (___9____24088), .DIN2 (___9____25106), .Q
       (_________37834));
  nor2s1 ____9__509231(.DIN1 (________24884), .DIN2 (___9____25076), .Q
       (_________37884));
  and2s1 _____0_509232(.DIN1 (___9____25051), .DIN2 (________25726), .Q
       (_____0___36285));
  nor2s1 ____9__509233(.DIN1 (________25320), .DIN2 (_____0__24974), .Q
       (_____9___37002));
  hi1s1 ____0__509234(.DIN (________25725), .Q (____99__26498));
  or2s1 ___9__509235(.DIN1 (_____0__24420), .DIN2 (________25723), .Q
       (________25724));
  and2s1 _______509236(.DIN1 (____0___29283), .DIN2 (___0_____40594),
       .Q (________25722));
  nor2s1 ____0__509237(.DIN1 (________23571), .DIN2 (_________35394),
       .Q (_____0__25721));
  nnd2s1 _______509238(.DIN1 (___9____25107), .DIN2 (_____0__23511), .Q
       (_____9__25720));
  and2s1 _______509239(.DIN1 (_____9__25785), .DIN2 (___0_____40621),
       .Q (________25719));
  hi1s1 ___9_0_509240(.DIN (________25717), .Q (________25718));
  hi1s1 ___9_0_509241(.DIN (________25715), .Q (________25716));
  hi1s1 ___9___509242(.DIN (_____0__27345), .Q (________25714));
  hi1s1 ___9__509243(.DIN (_________31783), .Q (________25713));
  nnd2s1 _____0_509244(.DIN1 (_____9__25785), .DIN2 (____9___22931), .Q
       (________25712));
  nnd2s1 ___9___509245(.DIN1 (_____9__25613), .DIN2 (________23380), .Q
       (_____0__25711));
  hi1s1 ___9___509246(.DIN (___9____26924), .Q (_____9__25710));
  hi1s1 _______509247(.DIN (________25707), .Q (________25708));
  hi1s1 _______509248(.DIN (___0____26088), .Q (________25705));
  nnd2s1 ______509249(.DIN1 (___9_9__25067), .DIN2 (_________37722), .Q
       (_____0__25704));
  nnd2s1 ______509250(.DIN1 (___9_9__25104), .DIN2 (________25702), .Q
       (_____9__25703));
  nnd2s1 _______509251(.DIN1 (________25700), .DIN2
       (_____________________________________0______21756), .Q
       (________25701));
  hi1s1 _______509252(.DIN (_________33692), .Q (________25699));
  and2s1 _______509253(.DIN1 (_________38377), .DIN2 (_______22183), .Q
       (________25698));
  hi1s1 ______509254(.DIN (_____0___41315), .Q (________25697));
  nnd2s1 _______509255(.DIN1 (________25700), .DIN2 (____9___23129), .Q
       (________25696));
  nnd2s1 _______509256(.DIN1 (________25008), .DIN2 (________24540), .Q
       (_____0__25695));
  hi1s1 _____0_509257(.DIN (_________31762), .Q (________25693));
  nnd2s1 _______509258(.DIN1 (________25700), .DIN2
       (____________________________________________21764), .Q
       (________25692));
  nnd2s1 _____509259(.DIN1 (________25690), .DIN2 (____99__24745), .Q
       (________25691));
  nor2s1 _____0_509260(.DIN1 (____99__25028), .DIN2 (________25663), .Q
       (________25689));
  nnd2s1 _____0_509261(.DIN1 (_____9__24828), .DIN2
       (_____________________________________________21908), .Q
       (_____0__25688));
  nnd2s1 _______509262(.DIN1 (________25647), .DIN2
       (_____________________________________9_______21881), .Q
       (____09__25687));
  nnd2s1 _______509263(.DIN1 (_________34877), .DIN2 (inData[7]), .Q
       (____0___25686));
  nnd2s1 _______509264(.DIN1 (_________34877), .DIN2 (inData[9]), .Q
       (____0___25685));
  nor2s1 ______509265(.DIN1
       (______________________________________0______21887), .DIN2
       (____0___25683), .Q (____0___25684));
  nnd2s1 ______509266(.DIN1 (____0___25683), .DIN2 (___0__9__40440), .Q
       (____0___25682));
  or2s1 _______509267(.DIN1
       (______________________________________0____), .DIN2
       (____0___25683), .Q (____0___25681));
  nor2s1 _______509268(.DIN1 (___0_____40443), .DIN2 (____0___25683),
       .Q (____0___25680));
  nnd2s1 _______509269(.DIN1 (___0_9___40270), .DIN2
       (______________________________________________21975), .Q
       (____0___25679));
  nnd2s1 ______509270(.DIN1 (___0_9___40270), .DIN2
       (______________________________________________21976), .Q
       (____00__25678));
  nnd2s1 ______509271(.DIN1 (___0_9___40270), .DIN2 (____9___25676), .Q
       (____99__25677));
  nor2s1 _______509272(.DIN1 (___0__0__31061), .DIN2 (________26279),
       .Q (____9___25675));
  or2s1 _______509273(.DIN1 (________23330), .DIN2 (________24780), .Q
       (____9___25674));
  nor2s1 _______509274(.DIN1 (___0_____40415), .DIN2 (________25665),
       .Q (____9___25673));
  nnd2s1 _______509275(.DIN1 (____9___25583), .DIN2 (___90___25034), .Q
       (____9___25672));
  nor2s1 _______509276(.DIN1 (________25257), .DIN2 (___9____25052), .Q
       (____9___25671));
  and2s1 _______509277(.DIN1 (______9__37555), .DIN2 (___0_____40623),
       .Q (____9___25670));
  nnd2s1 ______509278(.DIN1 (________25620), .DIN2 (________25458), .Q
       (_____9__25669));
  nnd2s1 _______509279(.DIN1 (______9__37555), .DIN2 (___0_____40622),
       .Q (________25668));
  and2s1 _______509280(.DIN1 (________25006), .DIN2 (___0____24212), .Q
       (________25667));
  nnd2s1 _______509281(.DIN1 (________25665), .DIN2 (________23850), .Q
       (________25666));
  nor2s1 _______509282(.DIN1 (___0____24230), .DIN2 (________25663), .Q
       (________25664));
  nnd2s1 _______509283(.DIN1 (____0___25683), .DIN2 (____9___23496), .Q
       (________25662));
  nor2s1 _______509284(.DIN1 (________25597), .DIN2 (_________37452),
       .Q (________25661));
  nor2s1 _______509285(.DIN1
       (______________________________________________21945), .DIN2
       (___99____39819), .Q (_____0__25660));
  or2s1 _____9_509286(.DIN1 (_____9__25823), .DIN2 (________25653), .Q
       (_____9__25659));
  nnd2s1 _____509287(.DIN1 (________24826), .DIN2 (___9_0__23182), .Q
       (________25658));
  nnd2s1 _____0_509288(.DIN1 (_____9__26765), .DIN2 (_______22217), .Q
       (________25657));
  nor2s1 _______509289(.DIN1 (________24822), .DIN2 (____90__24355), .Q
       (________25656));
  nnd2s1 _______509290(.DIN1 (________25017), .DIN2 (____9___22934), .Q
       (________25655));
  or2s1 _______509291(.DIN1 (___0____25206), .DIN2 (________25653), .Q
       (________25654));
  nor2s1 ___9_0_509292(.DIN1 (____9___23970), .DIN2 (_____0__24794), .Q
       (________25652));
  nor2s1 ___9_9_509293(.DIN1 (________24347), .DIN2 (________24865), .Q
       (_____0__25651));
  nor2s1 ___9_9_509294(.DIN1 (____0___25594), .DIN2 (_____9__25358), .Q
       (_____9__25650));
  nor2s1 ___9_509295(.DIN1 (________24777), .DIN2 (____0_0__34423), .Q
       (________25649));
  nnd2s1 ___9___509296(.DIN1 (________25647), .DIN2 (________22431), .Q
       (________25648));
  or2s1 ___9___509297(.DIN1 (________29249), .DIN2 (_________32001), .Q
       (________25646));
  nor2s1 ___9___509298(.DIN1 (________25644), .DIN2 (________25554), .Q
       (________25645));
  or2s1 ___9___509299(.DIN1 (________28934), .DIN2 (___9____25999), .Q
       (________25643));
  nor2s1 ___9___509300(.DIN1 (____0___25590), .DIN2 (____0___25588), .Q
       (_____0__25642));
  nnd2s1 ___9___509301(.DIN1 (____09__25595), .DIN2 (________25640), .Q
       (________25641));
  nnd2s1 ___9___509302(.DIN1 (________24770), .DIN2 (________25942), .Q
       (________25639));
  nnd2s1 ___9___509303(.DIN1 (________25562), .DIN2 (________26272), .Q
       (________25638));
  nor2s1 ___9___509304(.DIN1 (____0___23508), .DIN2 (____00__24839), .Q
       (________25637));
  or2s1 ___9__509305(.DIN1 (________25574), .DIN2 (________25723), .Q
       (________25636));
  nnd2s1 ___9___509306(.DIN1 (___900__25029), .DIN2 (________25634), .Q
       (________25635));
  nor2s1 ___9___509307(.DIN1 (_____9__25632), .DIN2 (_____9__25622), .Q
       (_____0__25633));
  hi1s1 ___509308(.DIN (________25630), .Q (________25631));
  hi1s1 ___9_509309(.DIN (________25628), .Q (________25629));
  hi1s1 ___9__509310(.DIN (________25626), .Q (________25627));
  hi1s1 ___9___509311(.DIN (_____0__25928), .Q (________25625));
  hi1s1 ___9___509312(.DIN (________26291), .Q (________25624));
  nor2s1 ___9___509313(.DIN1 (________24594), .DIN2 (_____9__25622), .Q
       (_____0__25623));
  and2s1 ___9___509314(.DIN1 (________25620), .DIN2 (________25640), .Q
       (________25621));
  nor2s1 ___9__509315(.DIN1 (___0____26067), .DIN2 (________24994), .Q
       (________25619));
  nor2s1 ___9_0_509316(.DIN1 (________23770), .DIN2 (________24792), .Q
       (________25618));
  hi1s1 ___9___509317(.DIN (_____9___32965), .Q (________25617));
  nnd2s1 ___9_9_509318(.DIN1 (____0___25587), .DIN2 (____9___23965), .Q
       (________25616));
  nor2s1 ___9___509319(.DIN1 (___9_9__25114), .DIN2 (________24776), .Q
       (________25615));
  nnd2s1 ___9___509320(.DIN1 (_____9__25613), .DIN2 (________22903), .Q
       (_____0__25614));
  nnd2s1 ___9__509321(.DIN1 (_____9__25613), .DIN2 (____9_), .Q
       (________25612));
  nnd2s1 ___9___509322(.DIN1 (________25475), .DIN2 (_____0__24601), .Q
       (________25611));
  nnd2s1 ___9___509323(.DIN1 (________24825), .DIN2 (___90___24071), .Q
       (________25610));
  nnd2s1 ___9___509324(.DIN1 (_________34877), .DIN2 (inData[8]), .Q
       (________25609));
  nor2s1 ___9___509325(.DIN1 (________25607), .DIN2 (____0___25591), .Q
       (________25608));
  nnd2s1 ___9__509326(.DIN1 (________24799), .DIN2 (________25605), .Q
       (________25606));
  nor2s1 ___9___509327(.DIN1 (________25644), .DIN2 (________24787), .Q
       (_____0__25604));
  nnd2s1 ___9___509328(.DIN1 (________25665), .DIN2 (_____0__22568), .Q
       (_____9__25603));
  nor2s1 ___9___509329(.DIN1 (____99__25585), .DIN2 (___9____25065), .Q
       (________26290));
  hi1s1 ___9_0_509330(.DIN (_________37614), .Q (_________33729));
  hi1s1 ___9___509331(.DIN (________26240), .Q (____0___26503));
  hi1s1 ___9___509332(.DIN (________25602), .Q (________26444));
  hi1s1 ___9___509333(.DIN (________25601), .Q (________27183));
  nor2s1 _______509334(.DIN1 (________23984), .DIN2 (________25568), .Q
       (___9_9__25996));
  nnd2s1 _______509335(.DIN1 (____9___25584), .DIN2 (________25923), .Q
       (____99__25957));
  nor2s1 ______509336(.DIN1 (________25600), .DIN2 (________25734), .Q
       (___9____25992));
  hi1s1 ___9___509337(.DIN (________29072), .Q (___00____30627));
  hi1s1 ___9___509338(.DIN (________25599), .Q (__9_0___30182));
  hi1s1 ___9___509339(.DIN (________25598), .Q (_________32246));
  nor2s1 ____9__509340(.DIN1 (_________22019), .DIN2 (_________37199),
       .Q (_________37528));
  nnd2s1 ____9__509341(.DIN1 (____0___25683), .DIN2 (___0_____40617),
       .Q (___9____25971));
  dffacs1 ______________________________________________0_509342(.CLRB
       (reset), .CLK (clk), .DIN (____9___24835), .QN
       (__________________________________________0___21959));
  nnd2s1 _____509343(.DIN1 (_________37452), .DIN2 (________25597), .Q
       (________26376));
  nnd2s1 _______509344(.DIN1 (____90__24829), .DIN2 (________23420), .Q
       (________26373));
  or2s1 ______509345(.DIN1 (____0___25592), .DIN2 (_____0__25596), .Q
       (________26337));
  nnd2s1 ___9___509346(.DIN1 (____09__25595), .DIN2 (________25634), .Q
       (___9_0__26004));
  nnd2s1 ___9__509347(.DIN1 (____0___25594), .DIN2 (____0___25593), .Q
       (________26242));
  or2s1 ___9___509348(.DIN1 (____0___25592), .DIN2 (________26760), .Q
       (________26311));
  nor2s1 ___9__509349(.DIN1 (________25735), .DIN2 (____0___25591), .Q
       (________26436));
  nnd2s1 ___9___509350(.DIN1 (_____9__24819), .DIN2 (________24378), .Q
       (_____0__26266));
  nor2s1 ___9__509351(.DIN1 (____0___25590), .DIN2 (________25663), .Q
       (________26274));
  hi1s1 ___9___509352(.DIN (__9_____29921), .Q (________26293));
  or2s1 ___9___509353(.DIN1 (____0___25589), .DIN2 (___9____25999), .Q
       (________26392));
  nor2s1 _____0_509354(.DIN1 (______0__32803), .DIN2 (____0___24941),
       .Q (___0____26076));
  nor2s1 ___9___509355(.DIN1 (________24531), .DIN2 (____0___25588), .Q
       (________26268));
  nnd2s1 ___9___509356(.DIN1 (________24772), .DIN2 (____0___26590), .Q
       (___9____26006));
  nnd2s1 ___9___509357(.DIN1 (____0___25587), .DIN2 (________24291), .Q
       (________26282));
  nnd2s1 ___9___509358(.DIN1 (____0___25316), .DIN2 (___0____25181), .Q
       (_____9__26265));
  nnd2s1 ___9___509359(.DIN1 (____0___25594), .DIN2 (________24896), .Q
       (_____0__26286));
  nor2s1 ___9___509360(.DIN1 (________25572), .DIN2 (_____9__25328), .Q
       (________26445));
  hi1s1 _______509361(.DIN (________25932), .Q (__9_____30285));
  dffacs1 _________________________________________0__9_(.CLRB (reset),
       .CLK (clk), .DIN (____0___24844), .Q (___0_____40577));
  hi1s1 _______509362(.DIN (________27171), .Q (__9_____29866));
  hi1s1 _______509363(.DIN
       (______________________________________________21932), .Q
       (___9__0__39146));
  nor2s1 _____9_509364(.DIN1 (_____9__24306), .DIN2 (____0___25770), .Q
       (___0____26073));
  hi1s1 ___9___509365(.DIN (___09____31487), .Q (________26287));
  dffacs1 ________________________________________________509366(.CLRB
       (reset), .CLK (clk), .DIN (_____0__24803), .Q
       (______________________________________________21964));
  hi1s1 ___9___509367(.DIN (___9_0__28655), .Q (________26271));
  hi1s1 ___9___509368(.DIN (____00__25586), .Q (________26374));
  nor2s1 ___9___509369(.DIN1 (____0___24845), .DIN2 (________28934), .Q
       (________28029));
  dffacs1 _______________________________________________509370(.CLRB
       (reset), .CLK (clk), .DIN (________24872), .Q
       (_____________________________________________21954));
  nnd2s1 ___9___509371(.DIN1 (___9_0___39344), .DIN2 (___0____25187),
       .Q (________25926));
  hi1s1 __90___(.DIN (___0__9__30984), .Q (_____9__26304));
  hi1s1 __90__509372(.DIN (________26335), .Q (________26283));
  nor2s1 ___9___509373(.DIN1 (____99__25585), .DIN2 (________25483), .Q
       (________27190));
  nnd2s1 _____509374(.DIN1 (____9___25584), .DIN2 (________26269), .Q
       (___0____27012));
  nnd2s1 ___9___509375(.DIN1 (________25665), .DIN2 (________25357), .Q
       (________27094));
  nnd2s1 ___9___509376(.DIN1 (________25003), .DIN2 (________27150), .Q
       (________28895));
  nor2s1 ___9___509377(.DIN1 (_____9__24715), .DIN2 (________25561), .Q
       (____0___27571));
  nnd2s1 ___9__509378(.DIN1 (________24779), .DIN2 (___9____23152), .Q
       (________29309));
  nnd2s1 ___9___509379(.DIN1 (____0___25587), .DIN2 (___0____25156), .Q
       (_____9__27185));
  nor2s1 ___9___509380(.DIN1 (________25376), .DIN2 (___90___25033), .Q
       (________26382));
  nor2s1 ____90_509381(.DIN1 (________24711), .DIN2 (_____0__24867), .Q
       (________26297));
  hi1s1 ______509382(.DIN (___9____26011), .Q (____9___28920));
  nnd2s1 _____509383(.DIN1 (____9___25583), .DIN2 (_____0__23891), .Q
       (____9___27564));
  hi1s1 _______509384(.DIN (___0____26116), .Q (_____0___32288));
  dffacs1 ________________________________________________509385(.CLRB
       (reset), .CLK (clk), .DIN (____9___24836), .Q
       (______________________________________________21961));
  nnd2s1 _______509386(.DIN1 (____9___25582), .DIN2 (________27598), .Q
       (____99__26682));
  nnd2s1 _______509387(.DIN1 (_____9__28617), .DIN2 (____9___25581), .Q
       (__9_____29949));
  nnd2s1 ___9___509388(.DIN1 (____0___25587), .DIN2 (___0____25169), .Q
       (________26344));
  nor2s1 _______509389(.DIN1 (____9___25580), .DIN2 (____9___25762), .Q
       (___09___27916));
  nnd2s1 _______509390(.DIN1 (____9___25579), .DIN2 (________27150), .Q
       (___9_0__26911));
  nnd2s1 ___9___509391(.DIN1 (_____9__25565), .DIN2 (________25550), .Q
       (_____0__27167));
  hi1s1 _______509392(.DIN (______9__31884), .Q (__9_____29818));
  hi1s1 ___9___509393(.DIN (____9___25577), .Q (__99_0__30469));
  nor2s1 ___9__509394(.DIN1 (________25560), .DIN2 (____0_0__34423), .Q
       (_____0__27932));
  nnd2s1 ___9__509395(.DIN1 (_________41327), .DIN2 (________25605), .Q
       (___9____26947));
  hi1s1 ___9___509396(.DIN (___0_____31094), .Q (___9_9__27776));
  nor2s1 ____9__509397(.DIN1 (_____0__25596), .DIN2 (___9____25097), .Q
       (___0____26982));
  hi1s1 ___9___509398(.DIN (____90__25576), .Q (________26394));
  hi1s1 ___9_9_509399(.DIN (___00_0__39902), .Q (________26568));
  nnd2s1 ____9__509400(.DIN1 (_____9__25613), .DIN2 (_____9__25575), .Q
       (_____0__26341));
  or2s1 ___9_9_509401(.DIN1 (___0____28779), .DIN2 (_________33106), .Q
       (________28589));
  nnd2s1 ______509402(.DIN1 (____0___24843), .DIN2 (________26601), .Q
       (________26432));
  hi1s1 __90_90(.DIN (___00____30562), .Q (________26303));
  nor2s1 ___9_509403(.DIN1 (________25002), .DIN2 (________25574), .Q
       (____0___27482));
  nnd2s1 ___9_9_509404(.DIN1 (________24813), .DIN2 (____0_0__34423),
       .Q (________26261));
  nor2s1 ___9___509405(.DIN1 (___0____25139), .DIN2 (________25573), .Q
       (_____9__28360));
  hi1s1 ______509406(.DIN (___0____27016), .Q (____0___26782));
  nnd2s1 ___9___509407(.DIN1 (________24997), .DIN2 (____9____34370),
       .Q (_________38172));
  dffacs1 ______________________________________509408(.CLRB (reset),
       .CLK (clk), .DIN (________24805), .Q (_____________22097));
  nor2s1 ___9__509409(.DIN1 (________25572), .DIN2 (________24790), .Q
       (_________33549));
  nor2s1 __90___509410(.DIN1 (________25571), .DIN2 (________24807), .Q
       (________27554));
  hi1s1 ___9___509411(.DIN (________25570), .Q (________28485));
  nnd2s1 ____9_509412(.DIN1 (________24977), .DIN2 (________25569), .Q
       (_____0__26617));
  and2s1 _____0_509413(.DIN1 (____9___25494), .DIN2 (____9___25763), .Q
       (________28074));
  nor2s1 _____9_509414(.DIN1 (____0___26409), .DIN2 (___90___25031), .Q
       (________29053));
  nnd2s1 ___509415(.DIN1 (____0___24846), .DIN2 (________25558), .Q
       (___90___28650));
  nor2s1 ____99_509416(.DIN1 (___09_9__31465), .DIN2 (_____0__28032),
       .Q (_____0__26390));
  nor2s1 ____9__509417(.DIN1 (___0_9__25154), .DIN2 (________25568), .Q
       (___0__0__30872));
  hi1s1 ___9___509418(.DIN (________25567), .Q (___0_90__31108));
  nor2s1 ____9__509419(.DIN1 (________24679), .DIN2 (____09__27128), .Q
       (________27602));
  nnd2s1 ___9_509420(.DIN1 (________24969), .DIN2 (________24722), .Q
       (_____9__26727));
  nor2s1 _____0_509421(.DIN1 (_____0__25566), .DIN2 (___9____25056), .Q
       (___0__9__40098));
  hi1s1 ______509422(.DIN (____0___26234), .Q (________26559));
  nnd2s1 ____9_509423(.DIN1 (_____9__25565), .DIN2 (________24898), .Q
       (_________32239));
  nnd2s1 _____0_509424(.DIN1 (___9____25046), .DIN2 (________24691), .Q
       (_________37893));
  nnd2s1 _______509425(.DIN1 (________24987), .DIN2 (________25740), .Q
       (________29428));
  nnd2s1 _______509426(.DIN1 (____0___24940), .DIN2 (________25564), .Q
       (_____9__27289));
  nnd2s1 ____9_509427(.DIN1 (________26239), .DIN2 (________25563), .Q
       (_________32931));
  nnd2s1 ___9_9_509428(.DIN1 (________25562), .DIN2 (____0___23316), .Q
       (______0__31825));
  nor2s1 ___9_9_509429(.DIN1 (________24797), .DIN2 (________25561), .Q
       (____0___26325));
  nor2s1 ___9_0_509430(.DIN1 (________25560), .DIN2 (________25946), .Q
       (________26632));
  nnd2s1 ___9_0_509431(.DIN1 (________24788), .DIN2 (________25559), .Q
       (_________31831));
  nnd2s1 ___9___509432(.DIN1 (________25557), .DIN2 (________25558), .Q
       (________27468));
  nnd2s1 ___9___509433(.DIN1 (________25557), .DIN2 (________23912), .Q
       (________28596));
  nor2s1 ___9___509434(.DIN1 (____9___24834), .DIN2 (_____0__25556), .Q
       (____0_0__31523));
  or2s1 ___9__509435(.DIN1 (_____9__25555), .DIN2 (________25554), .Q
       (___090___31415));
  nor2s1 ____9__509436(.DIN1 (________25553), .DIN2 (___9____25099), .Q
       (____0___29374));
  nnd2s1 ___9___509437(.DIN1 (_____0__27411), .DIN2 (___0_0__24218), .Q
       (_____9__27176));
  nnd2s1 ___9___509438(.DIN1 (___9____29574), .DIN2 (_____9__25937), .Q
       (__9_0___29724));
  nor2s1 ___9___509439(.DIN1 (________25573), .DIN2 (_____0__25359), .Q
       (________29090));
  and2s1 ___9___509440(.DIN1 (____0___24842), .DIN2 (_________33172),
       .Q (____9____34322));
  nor2s1 ___9_0_509441(.DIN1 (inData[6]), .DIN2 (_________32001), .Q
       (______0__34524));
  nnd2s1 _______509442(.DIN1 (________24959), .DIN2 (___0____26077), .Q
       (________28122));
  and2s1 ___90__509443(.DIN1 (________25552), .DIN2 (________25551), .Q
       (________28454));
  nnd2s1 ___9__509444(.DIN1 (________24796), .DIN2 (________24544), .Q
       (___09_9__31426));
  hi1s1 _______509445(.DIN (___0_____40380), .Q (________26557));
  nor2s1 ____9__509446(.DIN1 (________26280), .DIN2 (____9___25022), .Q
       (________29217));
  nor2s1 _______509447(.DIN1 (________25745), .DIN2 (________24851), .Q
       (____0___29013));
  nnd2s1 ___9___509448(.DIN1 (____0___25594), .DIN2 (________25550), .Q
       (___0_____31391));
  nnd2s1 ___9___509449(.DIN1 (____0___24841), .DIN2 (___9_0___39344),
       .Q (_________32078));
  nor2s1 ___9___509450(.DIN1 (_____0__25339), .DIN2 (____0___25591), .Q
       (_________32755));
  nor2s1 ___90_509451(.DIN1 (_____0__24820), .DIN2 (________25946), .Q
       (____00___33437));
  dffacs1 _________________________________________0____509452(.CLRB
       (reset), .CLK (clk), .DIN (___9____25083), .Q
       (_____________________________________0______21757));
  nor2s1 _____0_509453(.DIN1 (________24916), .DIN2 (________25549), .Q
       (____0____37113));
  hi1s1 _______509454(.DIN (___9_____39206), .Q (_________36928));
  nor2s1 ___9_0_509455(.DIN1 (___9_0__29602), .DIN2 (_________32001),
       .Q (_________31715));
  nnd2s1 _____509456(.DIN1 (________24856), .DIN2 (________25749), .Q
       (________28034));
  nnd2s1 ___90__509457(.DIN1 (____09__25595), .DIN2 (____9___25405), .Q
       (__9_____29873));
  nor2s1 _______509458(.DIN1 (________25548), .DIN2 (___0____25177), .Q
       (____9___27475));
  nor2s1 ___9_9_509459(.DIN1 (___0____26089), .DIN2 (_____9__24784), .Q
       (______9__32852));
  nnd2s1 ___90__509460(.DIN1 (________25547), .DIN2
       (_____________________21682), .Q (____9___26321));
  nnd2s1 ____9__509461(.DIN1 (___9____25098), .DIN2 (____9___27298), .Q
       (__99____30513));
  nor2s1 ___9_9_509462(.DIN1 (_____9__24983), .DIN2 (________25946), .Q
       (_________31942));
  hi1s1 _______509463(.DIN (_____9__25546), .Q (_________36301));
  nor2s1 _____9_509464(.DIN1 (________25539), .DIN2 (________24864), .Q
       (___0_____31073));
  nor2s1 _____9_509465(.DIN1 (_____0__26247), .DIN2 (___9____25101), .Q
       (___099___31496));
  hi1s1 ______509466(.DIN (________25545), .Q (_________31809));
  hi1s1 ___9_9_509467(.DIN (________26254), .Q (___00____39925));
  ib1s1 ___9_0_509468(.DIN (________25544), .Q (____0____32541));
  nor2s1 ______509469(.DIN1 (________25018), .DIN2 (________25574), .Q
       (________25543));
  nor2s1 _______509470(.DIN1 (___0_9__22323), .DIN2 (________25526), .Q
       (________25542));
  nnd2s1 ______509471(.DIN1 (________24534), .DIN2 (________25343), .Q
       (________25541));
  or2s1 ___9__509472(.DIN1 (________23864), .DIN2 (________25539), .Q
       (________25540));
  nnd2s1 _______509473(.DIN1 (_____9__25537), .DIN2 (______22164), .Q
       (_____0__25538));
  xor2s1 _______509474(.DIN1 (________25535), .DIN2 (___99_9__39836),
       .Q (________25536));
  hi1s1 _______509475(.DIN (___0__0__40571), .Q (________25534));
  nnd2s1 ___9___509476(.DIN1 (________24537), .DIN2 (___9____24123), .Q
       (________25533));
  nnd2s1 _______509477(.DIN1 (________24527), .DIN2 (___9____24093), .Q
       (________25532));
  xor2s1 _______509478(.DIN1 (____0____36194), .DIN2 (_____0___38422),
       .Q (________25531));
  nor2s1 ______509479(.DIN1 (_____9__23616), .DIN2 (________24624), .Q
       (________25530));
  nor2s1 _____0_509480(.DIN1
       (_____________________________________________21908), .DIN2
       (____0___25409), .Q (________25529));
  nnd2s1 _______509481(.DIN1 (________25523), .DIN2 (________25751), .Q
       (_____0__25528));
  nor2s1 ___9___509482(.DIN1 (_____0__22413), .DIN2 (________25526), .Q
       (_____9__25527));
  nnd2s1 _____9_509483(.DIN1 (________25523), .DIN2 (________26259), .Q
       (________25524));
  xor2s1 _______509484(.DIN1 (___0_____40045), .DIN2 (______9__34088),
       .Q (________25522));
  nor2s1 ___9___509485(.DIN1 (___990), .DIN2 (_____9__24505), .Q
       (________25521));
  nnd2s1 ___9__509486(.DIN1 (_________36480), .DIN2 (________22992), .Q
       (_____0__25520));
  and2s1 ___9__509487(.DIN1 (_________38200), .DIN2 (____99___36174),
       .Q (_____9__25519));
  hi1s1 ___9__509488(.DIN (___0_____31376), .Q (________25518));
  hi1s1 _______509489(.DIN (________28131), .Q (________25517));
  hi1s1 ___9___509490(.DIN (____9___25759), .Q (________25516));
  or2s1 _______509491(.DIN1 (_________22029), .DIN2 (________25513), .Q
       (________25514));
  nnd2s1 ______509492(.DIN1 (______0__38711), .DIN2
       (_____________22085), .Q (________25512));
  nor2s1 _______509493(.DIN1 (________25510), .DIN2 (____90__25300), .Q
       (________25511));
  nnd2s1 ______509494(.DIN1 (_____9__24344), .DIN2 (___0____24204), .Q
       (________25509));
  hi1s1 ______509495(.DIN (____09__25506), .Q (_____0__25507));
  nnd2s1 _______509496(.DIN1 (____9___25308), .DIN2 (________23431), .Q
       (____0___25505));
  and2s1 _______509497(.DIN1 (________24437), .DIN2
       (_________________________________________0___21862), .Q
       (____0___25504));
  nnd2s1 _______509498(.DIN1 (________25344), .DIN2 (____0___25502), .Q
       (____0___25503));
  hi1s1 _______509499(.DIN (____0___25500), .Q (____0___25501));
  and2s1 _______509500(.DIN1 (_____9__24419), .DIN2 (____0___25498), .Q
       (____0___25499));
  hi1s1 _______509501(.DIN (___0_____30789), .Q (____00__25497));
  xor2s1 _______509502(.DIN1 (_________33117), .DIN2 (______9__34088),
       .Q (____99__25496));
  nor2s1 _______509503(.DIN1 (________23331), .DIN2 (_____0__24627), .Q
       (____9___25495));
  nor2s1 _____0_509504(.DIN1 (____09__26331), .DIN2 (____9___24551), .Q
       (____9___25493));
  nnd2s1 _____0_509505(.DIN1 (_____0__25748), .DIN2 (________24863), .Q
       (____9___25492));
  nor2s1 _____9_509506(.DIN1 (___0_____40612), .DIN2 (_________37230),
       .Q (____9___25491));
  nnd2s1 _______509507(.DIN1 (____0___24650), .DIN2 (____90__25489), .Q
       (____9___25490));
  nor2s1 ______509508(.DIN1 (________24821), .DIN2 (_____0__25329), .Q
       (_____9__25488));
  hi1s1 _______509509(.DIN (________28876), .Q (________25487));
  nnd2s1 _____0_509510(.DIN1 (____9___24451), .DIN2 (____0___23047), .Q
       (________25486));
  and2s1 _______509511(.DIN1 (_________37230), .DIN2
       (______________________________________________21922), .Q
       (________25485));
  hi1s1 __90___509512(.DIN (________25483), .Q (________25484));
  nor2s1 _____0_509513(.DIN1 (___9_0__29602), .DIN2 (________24615), .Q
       (________25482));
  nor2s1 _____9_509514(.DIN1 (_____0__23019), .DIN2 (________24435), .Q
       (________25481));
  and2s1 _______509515(.DIN1 (____00__24646), .DIN2 (_____0__25479), .Q
       (________25480));
  nnd2s1 _______509516(.DIN1 (_____9__24535), .DIN2 (___0_0__24228), .Q
       (_____9__25478));
  nor2s1 _______509517(.DIN1 (________24013), .DIN2 (________25466), .Q
       (________25477));
  hi1s1 __90__509518(.DIN (________25475), .Q (________25476));
  nnd2s1 ______509519(.DIN1 (________24528), .DIN2 (________25364), .Q
       (________25474));
  nnd2s1 _______509520(.DIN1 (____9___25402), .DIN2 (___0_____40607),
       .Q (________25473));
  nor2s1 _______509521(.DIN1 (inData[1]), .DIN2 (_____0___35834), .Q
       (________25472));
  nnd2s1 _______509522(.DIN1 (_________32712), .DIN2
       (__________________________________________9___21977), .Q
       (________25471));
  nnd2s1 _______509523(.DIN1 (____9___25306), .DIN2 (_____9__25469), .Q
       (_____0__25470));
  nor2s1 _______509524(.DIN1 (________24734), .DIN2 (_____0__25252), .Q
       (________25468));
  nor2s1 _____0_509525(.DIN1 (___0____25186), .DIN2 (________25377), .Q
       (________25467));
  or2s1 _______509526(.DIN1 (_____9__24894), .DIN2 (____0____33465), .Q
       (________25465));
  nnd2s1 _______509527(.DIN1 (_____0__24592), .DIN2 (inData[4]), .Q
       (________25464));
  nnd2s1 _______509528(.DIN1 (________24603), .DIN2 (___00___23217), .Q
       (________25463));
  nor2s1 _______509529(.DIN1 (____0___23888), .DIN2 (_____0__25461), .Q
       (________25462));
  nnd2s1 _______509530(.DIN1 (___0____25182), .DIN2 (_____9__23682), .Q
       (_____9__25460));
  nnd2s1 _______509531(.DIN1 (________25455), .DIN2 (________25458), .Q
       (________25459));
  nnd2s1 ______509532(.DIN1 (________25366), .DIN2 (___99___26049), .Q
       (________25457));
  nnd2s1 _______509533(.DIN1 (________25455), .DIN2 (___0____26099), .Q
       (________25456));
  hi1s1 __90___509534(.DIN (___9____27809), .Q (________25454));
  nnd2s1 ___9_9_509535(.DIN1 (_____0__24526), .DIN2 (________24993), .Q
       (_____0__25453));
  nnd2s1 ___9___509536(.DIN1 (____0___25415), .DIN2 (________25569), .Q
       (_____9__25452));
  nnd2s1 ___9___509537(.DIN1 (____0___24754), .DIN2 (________24046), .Q
       (________25451));
  hi1s1 __90___509538(.DIN (________25560), .Q (________25450));
  nor2s1 ___9___509539(.DIN1 (________23341), .DIN2 (_____9__24410), .Q
       (________25449));
  nor2s1 ______509540(.DIN1 (___0___22203), .DIN2 (_________37230), .Q
       (________25447));
  nor2s1 ___9___509541(.DIN1 (___0____26087), .DIN2 (________25539), .Q
       (________25446));
  nnd2s1 _______509542(.DIN1 (________24539), .DIN2 (________23802), .Q
       (_____0__25445));
  nor2s1 _______509543(.DIN1 (________23828), .DIN2 (________24541), .Q
       (_____9__25444));
  nnd2s1 _______509544(.DIN1 (_________35448), .DIN2 (___9___22268), .Q
       (________25443));
  nor2s1 _______509545(.DIN1 (________25272), .DIN2 (________24434), .Q
       (________25442));
  or2s1 _______509546(.DIN1 (________25440), .DIN2 (________24394), .Q
       (________25441));
  nor2s1 ______509547(.DIN1 (________25438), .DIN2 (________25346), .Q
       (________25439));
  nnd2s1 _______509548(.DIN1 (________24498), .DIN2 (inData[26]), .Q
       (________25437));
  nor2s1 _______509549(.DIN1 (___9____25060), .DIN2 (____9___24453), .Q
       (________25436));
  nor2s1 ______509550(.DIN1 (_____9__25434), .DIN2 (_____9__24764), .Q
       (_____0__25435));
  nnd2s1 ______509551(.DIN1 (________24628), .DIN2 (________23357), .Q
       (________25433));
  xnr2s1 ____0__509552(.DIN1 (___0_0___40569), .DIN2 (___0_9___40556),
       .Q (________25432));
  nnd2s1 ____509553(.DIN1 (_________35448), .DIN2 (________22406), .Q
       (________25431));
  nor2s1 _______509554(.DIN1 (_____00__34847), .DIN2 (_____0__24566),
       .Q (________25430));
  or2s1 ______509555(.DIN1 (___0__9__40412), .DIN2 (_________35448), .Q
       (________25429));
  nnd2s1 _____509556(.DIN1 (_____0__25748), .DIN2 (________24518), .Q
       (________25428));
  nnd2s1 _____9_509557(.DIN1 (___0____24211), .DIN2 (________24402), .Q
       (________25427));
  or2s1 _____0_509558(.DIN1 (_________36402), .DIN2 (_________35448),
       .Q (________25426));
  xor2s1 _______509559(.DIN1 (_________34601), .DIN2 (___900___38985),
       .Q (_____0__25425));
  nor2s1 ______509560(.DIN1 (________22588), .DIN2 (_________37230), .Q
       (_____9__25424));
  nor2s1 _______509561(.DIN1 (________24671), .DIN2 (________24629), .Q
       (________25423));
  nnd2s1 _____0_509562(.DIN1 (____00__25407), .DIN2 (___0____24183), .Q
       (________25422));
  hi1s1 _______509563(.DIN (___9_____39667), .Q (________25421));
  nnd2s1 _____509564(.DIN1 (________25322), .DIN2 (________22974), .Q
       (________25420));
  nor2s1 _____9_509565(.DIN1 (____9___24643), .DIN2 (________24733), .Q
       (________25419));
  nor2s1 _____9_509566(.DIN1 (_____0__25417), .DIN2 (_____0__25271), .Q
       (________25418));
  nnd2s1 _____9_509567(.DIN1 (____0___25415), .DIN2 (________24033), .Q
       (____09__25416));
  nor2s1 _____509568(.DIN1 (________26307), .DIN2 (____9___24639), .Q
       (____0___25414));
  nor2s1 _____0_509569(.DIN1 (____0___25412), .DIN2 (____0___25411), .Q
       (____0___25413));
  nor2s1 _____0_509570(.DIN1
       (______________________________________0___9_), .DIN2
       (____0___25409), .Q (____0___25410));
  or2s1 ______509571(.DIN1
       (______________________________________0_______21894), .DIN2
       (____00__25407), .Q (____0___25408));
  nnd2s1 _______509572(.DIN1 (____9___25405), .DIN2 (____9___25404), .Q
       (____99__25406));
  nnd2s1 _______509573(.DIN1 (____9___25402), .DIN2
       (______________________________________0__0_), .Q
       (____9___25403));
  nnd2s1 _______509574(.DIN1 (_________32712), .DIN2 (___0_____40602),
       .Q (____9___25401));
  nnd2s1 _______509575(.DIN1 (_________32712), .DIN2 (______9__22030),
       .Q (____9___25400));
  nnd2s1 _______509576(.DIN1 (________24674), .DIN2 (________26429), .Q
       (____9___25399));
  nor2s1 _______509577(.DIN1 (_______22239), .DIN2 (_________32712), .Q
       (____90__25398));
  nor2s1 _______509578(.DIN1 (____90__24636), .DIN2 (___0_9__24256), .Q
       (_____9__25397));
  nor2s1 ______509579(.DIN1 (___99___26045), .DIN2 (_________41331), .Q
       (________25396));
  nnd2s1 _______509580(.DIN1 (________25394), .DIN2 (________24442), .Q
       (________25395));
  nnd2s1 _______509581(.DIN1 (________24512), .DIN2 (inData[4]), .Q
       (________25393));
  nor2s1 _______509582(.DIN1 (________25391), .DIN2 (_____0__24430), .Q
       (________25392));
  nor2s1 _______509583(.DIN1 (_____________________21736), .DIN2
       (________24397), .Q (________25390));
  nnd2s1 ______509584(.DIN1 (____9___24638), .DIN2 (inData[0]), .Q
       (_____0__25389));
  nor2s1 _______509585(.DIN1 (___9____24110), .DIN2 (____9___25402), .Q
       (_____9__25388));
  nor2s1 _______509586(.DIN1 (_____22114), .DIN2 (____0_9__38073), .Q
       (________25387));
  nnd2s1 ______509587(.DIN1 (________24520), .DIN2 (___9____24082), .Q
       (________25386));
  nnd2s1 ____0__509588(.DIN1 (_________35448), .DIN2 (________22822),
       .Q (________25385));
  and2s1 _______509589(.DIN1 (________24342), .DIN2 (________26171), .Q
       (________25384));
  nnd2s1 _____9_509590(.DIN1 (________25365), .DIN2 (_____0__24478), .Q
       (________25383));
  nor2s1 _____9_509591(.DIN1 (________24673), .DIN2 (________25285), .Q
       (________25382));
  nnd2s1 _____9_509592(.DIN1 (________28318), .DIN2 (_____9___22051),
       .Q (________25381));
  nor2s1 _______509593(.DIN1 (________25574), .DIN2 (________24405), .Q
       (________26454));
  hi1s1 _______509594(.DIN (___0_0___31031), .Q (___0_0__26082));
  nor2s1 _____0_509595(.DIN1 (______0__35694), .DIN2 (________24606),
       .Q (________25725));
  nor2s1 _______509596(.DIN1 (_____9__24695), .DIN2 (________25334), .Q
       (___0_9__26091));
  nnd2s1 __9009_(.DIN1 (___0____25173), .DIN2 (________25380), .Q
       (________25935));
  hi1s1 _______509597(.DIN (___0____26062), .Q (________26449));
  hi1s1 ___9___509598(.DIN (_____0__25379), .Q (________26424));
  nor2s1 ___90__509599(.DIN1 (________24412), .DIN2 (____9____38909),
       .Q (_____9__25546));
  nor2s1 ___90_509600(.DIN1 (___0_0__25203), .DIN2 (____9___24927), .Q
       (________25741));
  nor2s1 ____9_509601(.DIN1 (_____9__25378), .DIN2 (________25377), .Q
       (________25753));
  nor2s1 ____9__509602(.DIN1 (________25376), .DIN2 (____09__24655), .Q
       (________25755));
  nor2s1 ____9__509603(.DIN1 (_________37321), .DIN2 (_________38200),
       .Q (________25903));
  and2s1 _______509604(.DIN1 (_____0__24585), .DIN2 (________25375), .Q
       (___0____26085));
  hi1s1 ___9__509605(.DIN (________25374), .Q (___0_9__26081));
  and2s1 ___9___509606(.DIN1 (_________38573), .DIN2 (_________32918),
       .Q (___99___26043));
  nnd2s1 _______509607(.DIN1 (__9__0__30206), .DIN2 (________28519), .Q
       (________26799));
  nnd2s1 ___9___509608(.DIN1 (________25363), .DIN2 (________25373), .Q
       (___0_9__26111));
  hi1s1 ______509609(.DIN (________25372), .Q (______0__32823));
  or2s1 ___9___509610(.DIN1 (________25371), .DIN2 (________24508), .Q
       (________26163));
  nnd2s1 _______509611(.DIN1 (________25370), .DIN2 (_____0__25369), .Q
       (________25819));
  nnd2s1 _______509612(.DIN1 (_________38200), .DIN2 (_________37321),
       .Q (________26346));
  nor2s1 ______509613(.DIN1 (____99__25585), .DIN2 (________24427), .Q
       (___9____25994));
  nnd2s1 _______509614(.DIN1 (________25353), .DIN2 (_____9__25368), .Q
       (___9____25982));
  nnd2s1 _______509615(.DIN1 (________25367), .DIN2 (___99___25123), .Q
       (________25706));
  nnd2s1 _______509616(.DIN1 (________25367), .DIN2 (_____9__25348), .Q
       (___0____26124));
  nnd2s1 ______509617(.DIN1 (________24510), .DIN2 (___000__25125), .Q
       (_____9__27056));
  nor2s1 ______509618(.DIN1 (________24604), .DIN2 (___99___25120), .Q
       (________25707));
  nnd2s1 _______509619(.DIN1 (________25366), .DIN2 (________24769), .Q
       (___0_9__26101));
  nnd2s1 __90___509620(.DIN1 (___0____25199), .DIN2 (________25332), .Q
       (___90___25964));
  nnd2s1 _______509621(.DIN1 (___99___25121), .DIN2 (________23764), .Q
       (________25709));
  nnd2s1 _______509622(.DIN1 (________25365), .DIN2 (________25364), .Q
       (________25884));
  dffacs1 ______________________________________________9_509623(.CLRB
       (reset), .CLK (clk), .DIN (_____9__24617), .QN
       (__________________________________________9___21966));
  nnd2s1 _______509624(.DIN1 (________25323), .DIN2 (_____0__24506), .Q
       (___0____26119));
  nnd2s1 _______509625(.DIN1 (________25363), .DIN2 (________25362), .Q
       (___0____26079));
  nor2s1 _______509626(.DIN1 (___0____26078), .DIN2 (________24542), .Q
       (________28151));
  hi1s1 _______509627(.DIN (________25361), .Q (________26716));
  xor2s1 _____509628(.DIN1 (___0____22293), .DIN2 (_________36858), .Q
       (________26188));
  hi1s1 _______509629(.DIN (________28870), .Q (____0____33485));
  nor2s1 ____9__509630(.DIN1 (________25360), .DIN2 (_____9__25338), .Q
       (___0_0__26999));
  hi1s1 __90___509631(.DIN (_____0__25359), .Q (____90__29272));
  hi1s1 ___9__509632(.DIN (______9__31765), .Q (________26734));
  nnd2s1 ___9_9_509633(.DIN1 (_____9__25358), .DIN2 (________25550), .Q
       (___9____27782));
  nor2s1 ___9___509634(.DIN1 (________25357), .DIN2 (_________32712),
       .Q (___9____26023));
  or2s1 _______509635(.DIN1 (_____________________21709), .DIN2
       (________24543), .Q (_____0__27687));
  hi1s1 _______509636(.DIN (__9__0__29946), .Q (___0_____30684));
  nor2s1 ___9_9_509637(.DIN1 (________25356), .DIN2 (________24503), .Q
       (_____0__27345));
  nor2s1 _____9_509638(.DIN1 (________23061), .DIN2 (____0___25771), .Q
       (____0___26231));
  nor2s1 _____9_509639(.DIN1 (___0_0__25155), .DIN2 (________24582), .Q
       (___0_0__26122));
  nor2s1 ____90_509640(.DIN1 (________25336), .DIN2 (________25347), .Q
       (____9___26773));
  nnd2s1 ____90_509641(.DIN1 (________25363), .DIN2 (________25355), .Q
       (_____99__33716));
  nor2s1 ____509642(.DIN1 (________25354), .DIN2 (______0__37872), .Q
       (____0____37139));
  nnd2s1 ____9_509643(.DIN1 (________25366), .DIN2 (____0___26415), .Q
       (________26173));
  nnd2s1 ____9__509644(.DIN1 (________25353), .DIN2 (________25352), .Q
       (___0____26088));
  nor2s1 _______509645(.DIN1 (________26657), .DIN2 (____0___24751), .Q
       (__9_____29737));
  nor2s1 ____9_509646(.DIN1 (________25391), .DIN2 (________25377), .Q
       (________27939));
  nnd2s1 __90___509647(.DIN1 (___0____25160), .DIN2 (___0_9__25164), .Q
       (____9___28917));
  hi1s1 _______509648(.DIN (___90___28653), .Q (___0____26114));
  nor2s1 ____9__509649(.DIN1 (________25351), .DIN2 (________24759), .Q
       (_________32696));
  nnd2s1 ____9_509650(.DIN1 (________25350), .DIN2 (_____0__25349), .Q
       (________27058));
  nnd2s1 ____9__509651(.DIN1 (___0____25179), .DIN2 (____9___24063), .Q
       (__9_____29771));
  nnd2s1 ____9_509652(.DIN1 (________24608), .DIN2 (_____9__25348), .Q
       (________26603));
  nor2s1 ____9__509653(.DIN1 (________24599), .DIN2 (________25347), .Q
       (___0_0__26102));
  nor2s1 ____9__509654(.DIN1 (________24517), .DIN2 (________24446), .Q
       (________26740));
  nor2s1 ____9__509655(.DIN1 (________24632), .DIN2 (________25346), .Q
       (__9__9__29751));
  nor2s1 ____509656(.DIN1 (________25345), .DIN2 (________24660), .Q
       (________25932));
  nor2s1 ___90__509657(.DIN1 (________25335), .DIN2 (________25326), .Q
       (___9____26011));
  nnd2s1 ___90__509658(.DIN1 (____90__24448), .DIN2 (________24602), .Q
       (___0____27016));
  nnd2s1 ___90__509659(.DIN1 (________25344), .DIN2 (________25343), .Q
       (___0____26116));
  hi1s1 ___9___509660(.DIN (________28583), .Q (________29210));
  hi1s1 ___9___509661(.DIN (________25342), .Q (________26726));
  nor2s1 ____90_509662(.DIN1 (_____9__26294), .DIN2 (___0____25158), .Q
       (__9__9__29849));
  hi1s1 ______509663(.DIN (_________38743), .Q (___0____26097));
  hi1s1 ______509664(.DIN (________25341), .Q (________26434));
  hi1s1 _______509665(.DIN (_________33769), .Q (_________32104));
  nnd2s1 ____9__509666(.DIN1 (________25340), .DIN2 (___0_____30958),
       .Q (__9_____30054));
  nnd2s1 ____9__509667(.DIN1 (________24621), .DIN2 (________23535), .Q
       (___0_9__28814));
  nor2s1 _______509668(.DIN1 (________25553), .DIN2 (________24524), .Q
       (_____0__29037));
  nor2s1 ____9_509669(.DIN1 (_____0__25339), .DIN2 (_____9__25338), .Q
       (__99____30463));
  nor2s1 ____9__509670(.DIN1 (________25600), .DIN2 (________25325), .Q
       (___0_____30882));
  nor2s1 ____9__509671(.DIN1 (________25337), .DIN2 (____0___24651), .Q
       (____0___26236));
  nor2s1 ____9__509672(.DIN1 (________25336), .DIN2 (___0____25142), .Q
       (___90___28652));
  nor2s1 ____99_509673(.DIN1 (________25335), .DIN2 (________25330), .Q
       (___0____26117));
  nor2s1 ____99_509674(.DIN1 (________25572), .DIN2 (_____0__24383), .Q
       (___0____28754));
  dffacs1 ______________________________________509675(.CLRB (reset),
       .CLK (clk), .DIN (____0___24561), .Q (_____________22100));
  nor2s1 ___900_509676(.DIN1 (________24634), .DIN2 (________26604), .Q
       (_____0__28148));
  nor2s1 ___900_509677(.DIN1 (________25600), .DIN2 (___0____25147), .Q
       (__9__9__30419));
  and2s1 ___900_509678(.DIN1 (___999__25124), .DIN2 (_____9__25348), .Q
       (________28070));
  nor2s1 ___900_509679(.DIN1 (___0____25137), .DIN2 (________25334), .Q
       (___09___27917));
  nnd2s1 ___900_509680(.DIN1 (________25513), .DIN2 (____99__27741), .Q
       (__90_9__29708));
  nnd2s1 ___900_509681(.DIN1 (____9___24550), .DIN2 (___0____25146), .Q
       (________26523));
  or2s1 ___90__509682(.DIN1 (________25333), .DIN2 (__9__0__29841), .Q
       (___0_____31242));
  nor2s1 ______509683(.DIN1 (____0___26409), .DIN2 (____0___24654), .Q
       (___9_0__26940));
  nnd2s1 __90___509684(.DIN1 (___0____25138), .DIN2 (________25332), .Q
       (___00____30562));
  nnd2s1 ___9__509685(.DIN1 (________24593), .DIN2 (___00___25130), .Q
       (___09____31487));
  nnd2s1 _____0_509686(.DIN1 (________24682), .DIN2 (________25331), .Q
       (________28399));
  dffacs1 ________________________________________________509687(.CLRB
       (reset), .CLK (clk), .DIN (____9___24554), .Q
       (______________________________________________21932));
  nor2s1 ___90__509688(.DIN1 (________25327), .DIN2 (________25330), .Q
       (_____0__26168));
  nnd2s1 __90___509689(.DIN1 (___0____25190), .DIN2 (________25380), .Q
       (__99__));
  nor2s1 ___90__509690(.DIN1 (___0____26089), .DIN2 (_____0__25329), .Q
       (______9__31884));
  hi1s1 _______509691(.DIN (____09__25318), .Q (____99___37096));
  nnd2s1 ___90__509692(.DIN1 (________24390), .DIN2 (________26258), .Q
       (_________31749));
  nor2s1 ___9_9_509693(.DIN1 (________25371), .DIN2 (____9___24356), .Q
       (________28063));
  hi1s1 __90___509694(.DIN (_____9__25328), .Q (________25945));
  nnd2s1 _______509695(.DIN1 (____0___24647), .DIN2 (____90__25758), .Q
       (________28952));
  nor2s1 _______509696(.DIN1 (___0____26120), .DIN2 (_________37230),
       .Q (_________37837));
  nnd2s1 ____9__509697(.DIN1 (________24404), .DIN2 (___0____25157), .Q
       (___0____28811));
  or2s1 ____9__509698(.DIN1 (________25735), .DIN2 (_____9__25338), .Q
       (__99____30506));
  dffacs1 ______________________________________509699(.CLRB (reset),
       .CLK (clk), .DIN (____99__24555), .Q (_____________22102));
  nor2s1 ____9__509700(.DIN1 (________25929), .DIN2 (_____0__24610), .Q
       (____0___27576));
  nor2s1 ___90__509701(.DIN1 (________25327), .DIN2 (________25326), .Q
       (________29170));
  nnd2s1 ___90__509702(.DIN1 (____0___24368), .DIN2 (________23450), .Q
       (_________33692));
  nor2s1 ___90__509703(.DIN1 (________25735), .DIN2 (________25325), .Q
       (____0____31591));
  nor2s1 ____9_509704(.DIN1 (________25324), .DIN2 (___0____25208), .Q
       (_________31762));
  nor2s1 ___90__509705(.DIN1 (___0____25152), .DIN2 (____0___24562), .Q
       (________29173));
  nnd2s1 ___90__509706(.DIN1 (________25323), .DIN2 (________24581), .Q
       (____9___29007));
  nnd2s1 ___90__509707(.DIN1 (___00___25133), .DIN2 (________25944), .Q
       (_________32114));
  nor2s1 ___90__509708(.DIN1 (________23905), .DIN2 (________24670), .Q
       (____9____37036));
  nor2s1 ___90__509709(.DIN1 (____0___24463), .DIN2 (________24611), .Q
       (______0__35711));
  nor2s1 ___9_0_509710(.DIN1 (___9____25079), .DIN2 (________24443), .Q
       (____0____38091));
  nor2s1 ___9___509711(.DIN1 (___0____25168), .DIN2 (________24758), .Q
       (____0___28479));
  hi1s1 ___9_509712(.DIN (_________35394), .Q (____0___26141));
  hi1s1 ___9_9_509713(.DIN (_____9__25795), .Q (________26249));
  nnd2s1 ___90__509714(.DIN1 (________25322), .DIN2 (________23546), .Q
       (___0_____40380));
  nor2s1 ___90__509715(.DIN1 (________25929), .DIN2 (________24578), .Q
       (___0____27863));
  nor2s1 ___90_509716(.DIN1 (___00___25126), .DIN2 (________25347), .Q
       (___0_____31198));
  hi1s1 _______509717(.DIN (_____9__28617), .Q (__9_9___29888));
  hi1s1 _______509718(.DIN (_________38377), .Q (___0_____30688));
  hi1s1 ___9_9_509719(.DIN (________25321), .Q (_________34916));
  nor2s1 ___90_509720(.DIN1 (________25320), .DIN2 (____9___24456), .Q
       (___9_____39312));
  nnd2s1 ___90__509721(.DIN1 (________24416), .DIN2 (_____0__25319), .Q
       (____0___26234));
  nor2s1 ____9__509722(.DIN1 (____9___25023), .DIN2 (________24570), .Q
       (_________35523));
  nnd2s1 ___909_509723(.DIN1 (_____9__24400), .DIN2 (___9____23195), .Q
       (___9_____39582));
  nb1s1 ______509724(.DIN (____09__25318), .Q (_________38435));
  hi1s1 __90___509725(.DIN (____0___25316), .Q (____0___25317));
  nnd2s1 ___9___509726(.DIN1 (____9____37998), .DIN2 (________22487),
       .Q (____0___25315));
  nnd2s1 ___9___509727(.DIN1 (________25267), .DIN2 (________27288), .Q
       (____0___25314));
  nor2s1 ___9___509728(.DIN1 (_______22211), .DIN2 (___9_90__39245), .Q
       (____0___25313));
  nor2s1 ___9___509729(.DIN1 (________25756), .DIN2 (________24374), .Q
       (____0___25312));
  nnd2s1 ___9___509730(.DIN1 (___0_9__25184), .DIN2 (___0____25198), .Q
       (____0___25311));
  nor2s1 ___9___509731(.DIN1 (________22676), .DIN2 (______0__37872),
       .Q (____00__25310));
  nnd2s1 ___9__509732(.DIN1 (____9___25308), .DIN2 (________26259), .Q
       (____99__25309));
  and2s1 ___9___509733(.DIN1 (____9___25306), .DIN2 (________26267), .Q
       (____9___25307));
  nor2s1 ___9___509734(.DIN1 (________25756), .DIN2 (________25259), .Q
       (____9___25305));
  nor2s1 ___9___509735(.DIN1 (________22776), .DIN2 (___9_90__39245),
       .Q (____9___25304));
  nnd2s1 ___9__509736(.DIN1 (________24587), .DIN2 (________25605), .Q
       (____9___25303));
  nor2s1 ___9___509737(.DIN1 (___9____24156), .DIN2 (________24377), .Q
       (____9___25302));
  nor2s1 ___9___509738(.DIN1 (___900__25958), .DIN2 (____90__25300), .Q
       (____9___25301));
  nnd2s1 ___9___509739(.DIN1 (________24662), .DIN2 (________24341), .Q
       (________25299));
  nor2s1 ___9___509740(.DIN1 (________24616), .DIN2 (_____0__24042), .Q
       (________25298));
  nnd2s1 ___9_9_509741(.DIN1 (___0_0__25175), .DIN2 (________25270), .Q
       (________25297));
  and2s1 ___9_9_509742(.DIN1 (________24424), .DIN2 (________25569), .Q
       (________25296));
  nor2s1 ___9_509743(.DIN1 (________25294), .DIN2 (___0_0__25185), .Q
       (________25295));
  nor2s1 ___9_509744(.DIN1 (________24324), .DIN2 (_____9__24857), .Q
       (________25293));
  nnd2s1 ___9_0_509745(.DIN1 (________24491), .DIN2 (____9___22738), .Q
       (________25292));
  and2s1 ___9___509746(.DIN1 (________24391), .DIN2 (________25797), .Q
       (_____0__25291));
  nor2s1 ___9___509747(.DIN1 (________26421), .DIN2 (____0___24367), .Q
       (_____9__25290));
  nnd2s1 ___9___509748(.DIN1 (________25283), .DIN2 (________24302), .Q
       (________25289));
  nnd2s1 ___9___509749(.DIN1 (____0___24559), .DIN2 (___9_0__24139), .Q
       (________25288));
  nor2s1 ___9__509750(.DIN1 (___9_9__25047), .DIN2 (___09___25219), .Q
       (________25287));
  nor2s1 ___9___509751(.DIN1 (________25574), .DIN2 (________25285), .Q
       (________25286));
  nnd2s1 ___9___509752(.DIN1 (________25283), .DIN2 (________25282), .Q
       (________25284));
  nor2s1 ___9__509753(.DIN1 (_____9__25280), .DIN2 (____9___24450), .Q
       (_____0__25281));
  nor2s1 ___9___509754(.DIN1 (________24532), .DIN2 (________25278), .Q
       (________25279));
  nor2s1 ___9___509755(.DIN1 (___0____26083), .DIN2 (____99__24363), .Q
       (________25277));
  nnd2s1 ___9__509756(.DIN1 (________24379), .DIN2 (___9____25085), .Q
       (________25276));
  and2s1 ___9___509757(.DIN1 (_________38573), .DIN2
       (______________________________________________________________________________________0__22096),
       .Q (________25275));
  nnd2s1 ___9___509758(.DIN1 (________24678), .DIN2 (___00___25131), .Q
       (________25274));
  or2s1 ___9___509759(.DIN1 (________25272), .DIN2 (_____0__25271), .Q
       (________25273));
  nnd2s1 ___9___509760(.DIN1 (________24421), .DIN2 (________22855), .Q
       (________25269));
  nnd2s1 ___9___509761(.DIN1 (________25267), .DIN2 (____0___26410), .Q
       (________25268));
  and2s1 ___9__509762(.DIN1 (_____9__24575), .DIN2 (____9___24644), .Q
       (________25266));
  nor2s1 ___9_9_509763(.DIN1 (___0____26080), .DIN2 (___0____25180), .Q
       (________25265));
  nor2s1 ___9_509764(.DIN1 (________24388), .DIN2 (________24860), .Q
       (________25264));
  nor2s1 ___9_0_509765(.DIN1 (________25607), .DIN2 (___0____25178), .Q
       (________25263));
  nor2s1 ___9_0_509766(.DIN1 (____9___25402), .DIN2 (___0____24180), .Q
       (_____0__25262));
  nor2s1 ___9_0_509767(.DIN1 (________25260), .DIN2 (________25259), .Q
       (_____9__25261));
  nor2s1 ___9_0_509768(.DIN1 (____9___24362), .DIN2 (________25257), .Q
       (________25258));
  nnd2s1 ___9___509769(.DIN1 (________24352), .DIN2 (____9___26316), .Q
       (________25256));
  nor2s1 _______509770(.DIN1 (________24337), .DIN2 (________24045), .Q
       (________25255));
  nor2s1 _____0_509771(.DIN1 (_________41333), .DIN2 (____9___24552),
       .Q (________25254));
  nor2s1 _______509772(.DIN1 (____9___25955), .DIN2 (_____0__25252), .Q
       (________25253));
  nnd2s1 _______509773(.DIN1 (________24409), .DIN2 (clk), .Q
       (_____9__25251));
  or2s1 ____509774(.DIN1 (___9__9__39659), .DIN2 (________24406), .Q
       (________25250));
  xor2s1 ___9___509775(.DIN1 (________25248), .DIN2 (_________37687),
       .Q (________25249));
  xor2s1 ___9___509776(.DIN1
       (_____________________________________________21765), .DIN2
       (_____9___37654), .Q (________25247));
  nnd2s1 ___9___509777(.DIN1 (________24816), .DIN2 (________26429), .Q
       (________25245));
  hi1s1 ___9_0_509778(.DIN (_____0__25243), .Q (________25244));
  hi1s1 ___9___509779(.DIN (___0_____31366), .Q (________25242));
  nnd2s1 _______509780(.DIN1 (________24538), .DIN2 (_______22284), .Q
       (________25241));
  hi1s1 ___9___509781(.DIN (______0__33736), .Q (________25240));
  hi1s1 ___9___509782(.DIN (____9____32436), .Q (________25239));
  hi1s1 ___9__509783(.DIN (________25834), .Q (________25238));
  nor2s1 ______509784(.DIN1 (________23582), .DIN2 (________24633), .Q
       (________25237));
  hi1s1 ___9___509785(.DIN (_____0__29262), .Q (________25236));
  nor2s1 ___9___509786(.DIN1 (___0_0__23225), .DIN2 (________25526), .Q
       (________25235));
  nor2s1 ___9_9_509787(.DIN1 (___99___25118), .DIN2 (_____0__24812), .Q
       (________25234));
  hi1s1 ___9__509788(.DIN (___0_____31268), .Q (________25233));
  nnd2s1 ___9___509789(.DIN1 (________24349), .DIN2 (_____9___37752),
       .Q (________25232));
  nnd2s1 ___9___509790(.DIN1 (______0__38711), .DIN2 (___0_9__23243),
       .Q (_____0__25231));
  nor2s1 ___9___509791(.DIN1 (___99___26045), .DIN2 (________24396), .Q
       (____09__25230));
  nor2s1 ___9___509792(.DIN1 (____9___25860), .DIN2 (________25285), .Q
       (____0___25228));
  nor2s1 ___9___509793(.DIN1 (________24693), .DIN2 (____9___24357), .Q
       (____0___25227));
  nor2s1 ___9___509794(.DIN1 (________26440), .DIN2 (____0___24753), .Q
       (____0___25226));
  hi1s1 ___9_509795(.DIN (____0___25224), .Q (____0___25225));
  hi1s1 ___9___509796(.DIN (___9____27820), .Q (____0___25223));
  nor2s1 ___9___509797(.DIN1 (___0____26080), .DIN2 (____09__24372), .Q
       (____00__25222));
  nnd2s1 ___9___509798(.DIN1 (________24626), .DIN2 (____0___25502), .Q
       (___099__25221));
  nor2s1 ___9___509799(.DIN1 (___0____26083), .DIN2 (___09___25219), .Q
       (___09___25220));
  nnd2s1 _____0_509800(.DIN1 (________24672), .DIN2 (______22153), .Q
       (___09___25218));
  nnd2s1 ___9___509801(.DIN1 (_________38262), .DIN2 (____0___24371),
       .Q (___09___25217));
  nor2s1 ___9_9_509802(.DIN1 (________22579), .DIN2 (___9_90__39245),
       .Q (___09___25216));
  nnd2s1 ___9___509803(.DIN1 (________24422), .DIN2 (___9_9__25977), .Q
       (___09___25215));
  or2s1 ___9_9_509804(.DIN1 (___9____25981), .DIN2 (___090__25213), .Q
       (___09___25214));
  hi1s1 __90___509805(.DIN (________26300), .Q (___0_9__25212));
  nor2s1 ___9___509806(.DIN1 (___0____25210), .DIN2 (________24657), .Q
       (___0____25211));
  nor2s1 _______509807(.DIN1 (________22381), .DIN2 (___0____25208), .Q
       (___0____25209));
  or2s1 __90___509808(.DIN1 (___0____25206), .DIN2 (________25574), .Q
       (___0____25207));
  or2s1 __90_0_(.DIN1 (___0____25204), .DIN2 (___0_0__25203), .Q
       (___0____25205));
  or2s1 __90___509809(.DIN1 (________24586), .DIN2 (___0_0__25203), .Q
       (___0_9__25202));
  or2s1 __90___509810(.DIN1 (___00___25132), .DIN2 (___0_0__25203), .Q
       (___0____25201));
  nnd2s1 __90___509811(.DIN1 (___0____25199), .DIN2 (___0____25198), .Q
       (___0____25200));
  and2s1 ___9__509812(.DIN1 (____9___25306), .DIN2 (________25829), .Q
       (___0____25197));
  hi1s1 __90___509813(.DIN (______0__41329), .Q (___0____25196));
  and2s1 ___9___509814(.DIN1 (________25523), .DIN2 (____0___25774), .Q
       (___0____25195));
  nnd2s1 ___9_9_509815(.DIN1 (________24414), .DIN2 (________24343), .Q
       (___0_0__25194));
  xnr2s1 _____9_509816(.DIN1 (___0_0___40565), .DIN2 (___9_____39332),
       .Q (___0_9__25193));
  hi1s1 ___9___509817(.DIN (____9___25583), .Q (___0____25192));
  nnd2s1 ___9___509818(.DIN1 (___0____25190), .DIN2 (____90__23962), .Q
       (___0____25191));
  hi1s1 ___9___509819(.DIN (_____9___32184), .Q (___0____25189));
  hi1s1 ___9___509820(.DIN (___0____25187), .Q (___0____25188));
  nor2s1 ___9___509821(.DIN1 (___0____25186), .DIN2 (___0_0__25185), .Q
       (_____0__25778));
  nnd2s1 ___9___509822(.DIN1 (___0_9__25184), .DIN2 (________25332), .Q
       (____9___25951));
  nnd2s1 ___9___509823(.DIN1 (____9___24359), .DIN2 (________25355), .Q
       (___0____26110));
  nnd2s1 ___9___509824(.DIN1 (___0____25183), .DIN2 (____99__23971), .Q
       (___9____26037));
  nnd2s1 _______509825(.DIN1 (___0____25182), .DIN2 (________23957), .Q
       (________25817));
  nnd2s1 _______509826(.DIN1 (___0____25166), .DIN2 (___0____25181), .Q
       (___9____25976));
  nnd2s1 ____9_509827(.DIN1 (________24620), .DIN2 (________26259), .Q
       (________25730));
  nnd2s1 ___9__509828(.DIN1 (________25523), .DIN2 (____0___23040), .Q
       (________25940));
  nor2s1 _______509829(.DIN1 (_____9__24325), .DIN2 (____00__24458), .Q
       (____9___25950));
  nor2s1 ___9___509830(.DIN1 (________25744), .DIN2 (________24613), .Q
       (________26441));
  nor2s1 ___9__509831(.DIN1 (___0_9__24187), .DIN2 (___0____25180), .Q
       (___0_9__27008));
  hi1s1 ___9___509832(.DIN (________25653), .Q (___9____26002));
  hi1s1 ___9___509833(.DIN (________27638), .Q (___90___25965));
  and2s1 ___9___509834(.DIN1 (___0____25179), .DIN2 (____0___24748), .Q
       (___9_0__25968));
  nor2s1 ___9___509835(.DIN1 (________25391), .DIN2 (___0_0__25185), .Q
       (________25628));
  nor2s1 ___9___509836(.DIN1 (_____0__25339), .DIN2 (___0____25178), .Q
       (________25626));
  nor2s1 _______509837(.DIN1 (________24757), .DIN2 (___0____25208), .Q
       (___0____26090));
  nor2s1 ___9___509838(.DIN1 (________23920), .DIN2 (___0____25177), .Q
       (________25924));
  nnd2s1 ___9___509839(.DIN1 (____0___24370), .DIN2 (___00___25129), .Q
       (________25570));
  hi1s1 ___9___509840(.DIN (_________33570), .Q (___0_____31186));
  nnd2s1 ___9__509841(.DIN1 (___00___25128), .DIN2 (________25373), .Q
       (________25694));
  nor2s1 ___9_9_509842(.DIN1 (________25391), .DIN2 (____0___25411), .Q
       (____00__25586));
  hi1s1 ___9___509843(.DIN (_____0___34487), .Q (________26733));
  hi1s1 ___9__509844(.DIN (____0___29202), .Q (___909__25967));
  and2s1 __90___509845(.DIN1 (___0____25170), .DIN2 (___0____25198), .Q
       (________26284));
  nnd2s1 ___9___509846(.DIN1 (___0____25140), .DIN2 (___0____25176), .Q
       (________25598));
  nnd2s1 ___9___509847(.DIN1 (_____0__24440), .DIN2 (________25375), .Q
       (________25599));
  nnd2s1 ___9___509848(.DIN1 (___0_0__25175), .DIN2 (________25549), .Q
       (________25567));
  hi1s1 ___9___509849(.DIN (___9____28657), .Q (________25939));
  hi1s1 __90__9(.DIN (___0_9__25174), .Q (________26264));
  nnd2s1 __9009_509850(.DIN1 (___0____25173), .DIN2 (___0____25172), .Q
       (________26281));
  hi1s1 __90__509851(.DIN (__9_0___30000), .Q (________25936));
  hi1s1 __90___509852(.DIN (___0____26978), .Q (____9___25954));
  nnd2s1 ___9___509853(.DIN1 (___0_9__25184), .DIN2 (___0____25171), .Q
       (________25601));
  hi1s1 __90_9_(.DIN (_________38576), .Q (___9_0__25988));
  nnd2s1 ___9__509854(.DIN1 (________24773), .DIN2 (________25559), .Q
       (________25715));
  or2s1 ___9___509855(.DIN1 (________24922), .DIN2 (___0____25167), .Q
       (___0____26107));
  nnd2s1 ___9___509856(.DIN1 (____0___24560), .DIN2 (________25944), .Q
       (________25602));
  nnd2s1 ___9__509857(.DIN1 (___90____39051), .DIN2 (_________41337),
       .Q (____90__25576));
  nnd2s1 __90___509858(.DIN1 (___0____25170), .DIN2 (___0____25169), .Q
       (___90___25962));
  nor2s1 ___9_9_509859(.DIN1 (___0____25168), .DIN2 (___0____25167), .Q
       (____9___25577));
  nnd2s1 ___9__509860(.DIN1 (___0____25166), .DIN2 (________24782), .Q
       (________25630));
  nnd2s1 ___9___509861(.DIN1 (___0_0__25165), .DIN2 (____0___26690), .Q
       (________26795));
  nnd2s1 ___9___509862(.DIN1 (___0____25179), .DIN2 (________24720), .Q
       (____0___26147));
  nnd2s1 ___9___509863(.DIN1 (___0____25179), .DIN2 (________23998), .Q
       (___9____25972));
  nnd2s1 __90___509864(.DIN1 (___0____25170), .DIN2 (___0_9__25164), .Q
       (___9____25973));
  nnd2s1 __90___509865(.DIN1 (___0____25162), .DIN2 (________25332), .Q
       (___9____26922));
  nor2s1 ___9___509866(.DIN1 (___0____25163), .DIN2 (________24376), .Q
       (________25717));
  and2s1 __90___509867(.DIN1 (___0____25149), .DIN2 (________25332), .Q
       (____9___25952));
  nor2s1 __90___509868(.DIN1 (____0___23317), .DIN2 (___0_0__25203), .Q
       (____99__25767));
  nnd2s1 __90_0_509869(.DIN1 (___0____25162), .DIN2 (___0____25159), .Q
       (________25943));
  nnd2s1 __90___509870(.DIN1 (________24340), .DIN2 (___9____23169), .Q
       (____0___25773));
  nnd2s1 ___9___509871(.DIN1 (____9___24548), .DIN2 (___0____25161), .Q
       (___0____26104));
  nnd2s1 __90___509872(.DIN1 (___0____25160), .DIN2 (___0____25169), .Q
       (________28162));
  or2s1 ____9__509873(.DIN1 (________25929), .DIN2 (_____0__24676), .Q
       (________25545));
  nnd2s1 _____9_509874(.DIN1 (________24413), .DIN2 (___0____25181), .Q
       (___0____26093));
  nor2s1 _______509875(.DIN1 (_______22228), .DIN2 (________24669), .Q
       (_____9__26210));
  nor2s1 ___9___509876(.DIN1 (___0____25143), .DIN2 (___0____25167), .Q
       (___0_0__26112));
  nor2s1 ____9__509877(.DIN1 (_____9__25434), .DIN2 (_____9__25338), .Q
       (________27665));
  nnd2s1 ____9_509878(.DIN1 (________24667), .DIN2 (________25362), .Q
       (___0____26094));
  nnd2s1 __90___509879(.DIN1 (___0____25160), .DIN2 (___0____25159), .Q
       (___9____25979));
  nnd2s1 ___9_9_509880(.DIN1 (____99__24645), .DIN2 (_____0__26418), .Q
       (_____0__25928));
  nor2s1 ___9_0_509881(.DIN1 (____9___24742), .DIN2 (________25325), .Q
       (____0___27214));
  nnd2s1 ___9___509882(.DIN1 (_____9__25358), .DIN2 (_____0__24905), .Q
       (________26742));
  nor2s1 _______509883(.DIN1 (___0____25158), .DIN2 (____9____34365),
       .Q (___9____29597));
  and2s1 ___9_9_509884(.DIN1 (___00___25127), .DIN2 (___0____25157), .Q
       (___9____26942));
  nnd2s1 __90___509885(.DIN1 (________24677), .DIN2 (___0____25156), .Q
       (___9____25969));
  nor2s1 ___9_0_509886(.DIN1 (___0_0__25155), .DIN2 (________24399), .Q
       (___0____26113));
  nor2s1 ___9___509887(.DIN1 (________25371), .DIN2 (________24350), .Q
       (_____9__25947));
  nnd2s1 __90_00(.DIN1 (___0____25160), .DIN2 (___0____25198), .Q
       (________26335));
  nnd2s1 __90___509888(.DIN1 (___0____25170), .DIN2 (________25332), .Q
       (___0____26095));
  nor2s1 ___9_9_509889(.DIN1 (_________32918), .DIN2 (_________38573),
       .Q (____9___26222));
  nnd2s1 ___9_0_509890(.DIN1 (________24595), .DIN2 (________26272), .Q
       (________27339));
  nor2s1 ___9_509891(.DIN1 (___0_9__25154), .DIN2 (____00__24364), .Q
       (________29336));
  or2s1 ___9___509892(.DIN1 (___0____25153), .DIN2 (________29249), .Q
       (__9__0__30093));
  nor2s1 ___9__509893(.DIN1 (________24698), .DIN2 (________24530), .Q
       (_____0__27270));
  nor2s1 ___9__509894(.DIN1 (___0____25152), .DIN2 (________24339), .Q
       (________27378));
  nor2s1 ___9___509895(.DIN1 (________24886), .DIN2 (_____0__24336), .Q
       (________26291));
  hi1s1 ___9___509896(.DIN (___0____25151), .Q (________29231));
  hi1s1 ___9___509897(.DIN (___0____25150), .Q (___0_____31140));
  nnd2s1 __90___509898(.DIN1 (___0____25149), .DIN2 (___0____25156), .Q
       (____9___25953));
  nor2s1 ___9___509899(.DIN1 (___0_9__25154), .DIN2 (_____9__24354), .Q
       (____9___29544));
  hi1s1 ___9___509900(.DIN (___0____25148), .Q (___0_____30912));
  or2s1 ___9__509901(.DIN1 (___0____25186), .DIN2 (___0____25147), .Q
       (____0___26593));
  nnd2s1 ___9___509902(.DIN1 (________24425), .DIN2 (___0____25146), .Q
       (___0____26061));
  hi1s1 ___9__509903(.DIN (___0_0__25145), .Q (___0__9__30671));
  nor2s1 ___9___509904(.DIN1 (____0___25412), .DIN2 (___0_0__25185), .Q
       (___9____26927));
  dffacs1 _____________________________________________0_509905(.CLRB
       (reset), .CLK (clk), .DIN (____0___24652), .Q
       (_________________________________________0___21952));
  hi1s1 ___9___509906(.DIN (___0____26123), .Q (____9____32446));
  nor2s1 ___9___509907(.DIN1 (_____0__23009), .DIN2 (________24403), .Q
       (________27169));
  nnd2s1 ___9___509908(.DIN1 (_____0__24401), .DIN2 (________25549), .Q
       (________25544));
  nnd2s1 ___9___509909(.DIN1 (_____9__25537), .DIN2 (___0_9__25144), .Q
       (___90___25961));
  nor2s1 ___9__509910(.DIN1 (____09__24565), .DIN2 (_____0__25556), .Q
       (________26614));
  nor2s1 ___9___509911(.DIN1 (________24908), .DIN2 (________24380), .Q
       (________26296));
  nnd2s1 ___9_9_509912(.DIN1 (________24572), .DIN2 (________25355), .Q
       (_____0__25938));
  nnd2s1 ___9___509913(.DIN1 (________24631), .DIN2 (____0___23602), .Q
       (________25934));
  nor2s1 ___9__509914(.DIN1 (____0___24365), .DIN2 (________25946), .Q
       (___0__0__31080));
  hi1s1 __90___509915(.DIN (______9__37555), .Q (______0__37345));
  and2s1 ___9___509916(.DIN1 (___0____25179), .DIN2 (_____0__24895), .Q
       (_____0__29534));
  nnd2s1 ___9___509917(.DIN1 (____9___24549), .DIN2 (___0____25146), .Q
       (__90____29672));
  nor2s1 ___9___509918(.DIN1 (___0____25143), .DIN2 (___0____25142), .Q
       (________29072));
  hi1s1 ___9___509919(.DIN (___0____25141), .Q (____0___27035));
  nnd2s1 ___9__509920(.DIN1 (___0____25140), .DIN2 (________25373), .Q
       (________28084));
  nnd2s1 ___9__509921(.DIN1 (___90___25032), .DIN2 (________25362), .Q
       (___9____27773));
  hi1s1 __90___509922(.DIN (___0____25139), .Q (________28495));
  nnd2s1 ___9___509923(.DIN1 (________24492), .DIN2 (___0____26078), .Q
       (________27545));
  nnd2s1 __90___509924(.DIN1 (___0____25138), .DIN2 (___0____25171), .Q
       (________29384));
  nnd2s1 __90___509925(.DIN1 (___0____25162), .DIN2 (___0____25171), .Q
       (________28507));
  nnd2s1 ___9_0_509926(.DIN1 (_____0__24345), .DIN2 (____9___23037), .Q
       (________26254));
  nor2s1 ___9___509927(.DIN1 (____0___26409), .DIN2 (____0___24461), .Q
       (___9____27801));
  nor2s1 ___9___509928(.DIN1 (___0____25137), .DIN2 (____9___24553), .Q
       (___9_0__28655));
  nnd2s1 __90___509929(.DIN1 (___0____25138), .DIN2 (___0_9__25164), .Q
       (___0__9__30984));
  nor2s1 _____9_509930(.DIN1 (_____0___31994), .DIN2 (________27181),
       .Q (___0__0__30796));
  nor2s1 ____9_509931(.DIN1 (___0_0__25135), .DIN2 (____9___24744), .Q
       (_________32903));
  hi1s1 __90__509932(.DIN (___009__25134), .Q (____0____31527));
  and2s1 ____9__509933(.DIN1 (___00___25133), .DIN2 (________25362), .Q
       (____0____31589));
  nor2s1 ___9_0_509934(.DIN1 (___00___25132), .DIN2 (____0___24366), .Q
       (___00____30587));
  nnd2s1 ____99_509935(.DIN1 (________24381), .DIN2 (___00___25131), .Q
       (____00__27922));
  nnd2s1 ___9_0_509936(.DIN1 (___0____25179), .DIN2 (________24597), .Q
       (________28533));
  nnd2s1 ___9___509937(.DIN1 (___00___25130), .DIN2 (________24334), .Q
       (________26240));
  nor2s1 ___9___509938(.DIN1 (________25360), .DIN2 (________25325), .Q
       (_________32065));
  nnd2s1 ___9__509939(.DIN1 (________24346), .DIN2 (___00___25129), .Q
       (________28040));
  nnd2s1 ___9___509940(.DIN1 (___00___25128), .DIN2 (____99__26407), .Q
       (__9_____29921));
  hi1s1 ___9___509941(.DIN (____00__25768), .Q (_________33000));
  nnd2s1 ___9___509942(.DIN1 (___00___25127), .DIN2 (___00___25129), .Q
       (____9___26491));
  nor2s1 ___9_0_509943(.DIN1 (___00___25126), .DIN2 (___0____25142), .Q
       (________29068));
  nor2s1 ___9_9_509944(.DIN1 (________24589), .DIN2 (________26604), .Q
       (___9____26924));
  or2s1 ___9_0_509945(.DIN1 (_____9__25378), .DIN2 (____0___24649), .Q
       (_________32260));
  nnd2s1 ___9___509946(.DIN1 (_____9__25358), .DIN2 (____0___25593), .Q
       (___0____27014));
  nnd2s1 ___9___509947(.DIN1 (___99___25117), .DIN2 (___000__25125), .Q
       (_________32811));
  nor2s1 ___90__509948(.DIN1 (________24289), .DIN2 (________25334), .Q
       (________27171));
  dffacs1 ______________________________________509949(.CLRB (reset),
       .CLK (clk), .DIN (________24663), .Q (_____________22099));
  and2s1 ___9_0_509950(.DIN1 (_____9__24600), .DIN2 (___0____25157), .Q
       (________28392));
  nor2s1 ____9__509951(.DIN1 (________24569), .DIN2 (________25946), .Q
       (__9_____30115));
  nnd2s1 ___9___509952(.DIN1 (___999__25124), .DIN2 (___99___25123), .Q
       (___0_____31094));
  nnd2s1 ___9__509953(.DIN1 (___00___25128), .DIN2 (________25362), .Q
       (___0090__30632));
  nor2s1 ____99_509954(.DIN1 (___9____24081), .DIN2 (_____9__24545), .Q
       (_________33609));
  hi1s1 ___9___509955(.DIN (___99___25122), .Q (______9__31632));
  hi1s1 ___9___509956(.DIN (___99____39819), .Q (___9_____39743));
  nnd2s1 ___9___509957(.DIN1 (___00___25130), .DIN2 (___99___25121), .Q
       (___0_____31385));
  or2s1 ___90__509958(.DIN1 (___0_0__25135), .DIN2 (___0_0__25185), .Q
       (___0_____30917));
  or2s1 ___90__509959(.DIN1 (_____9__25378), .DIN2 (____0___24563), .Q
       (____0____31517));
  nor2s1 ___90_509960(.DIN1 (___99___25119), .DIN2 (________25330), .Q
       (____0___27925));
  nor2s1 ___9___509961(.DIN1 (___0____25206), .DIN2 (____90__25300), .Q
       (__9_____29766));
  nor2s1 ___90__509962(.DIN1 (___0____26109), .DIN2 (___99___25120), .Q
       (__99____30485));
  nor2s1 ___90__509963(.DIN1 (___99___25119), .DIN2 (________25326), .Q
       (________29225));
  nnd2s1 ___9___509964(.DIN1 (___00___25128), .DIN2 (___0____25176), .Q
       (_____9___32965));
  hi1s1 ___9_9_509965(.DIN (_________36955), .Q (_________36670));
  nor2s1 ___9___509966(.DIN1 (________25294), .DIN2 (____0___25411), .Q
       (____0____31547));
  nnd2s1 ___9___509967(.DIN1 (___9____25064), .DIN2 (___0____25176), .Q
       (_________34243));
  nnd2s1 ___9___509968(.DIN1 (________24982), .DIN2 (___99___25118), .Q
       (_________31868));
  nnd2s1 ___9_9_509969(.DIN1 (____0___24558), .DIN2 (________23933), .Q
       (__90_9__29688));
  nor2s1 ___9_9_509970(.DIN1 (________24387), .DIN2 (____0_0__34423),
       .Q (_________32142));
  nnd2s1 ___9__509971(.DIN1 (___99___25117), .DIN2 (________25944), .Q
       (____9_0__32391));
  nnd2s1 ___909_509972(.DIN1 (________24441), .DIN2 (________23369), .Q
       (___9_____39206));
  dffacs1 _______________________________________509973(.CLRB (reset),
       .CLK (clk), .DIN (________24423), .Q (___0_9___40452));
  nor2s1 ___9___509974(.DIN1 (____9___24830), .DIN2 (_____0__25329), .Q
       (_________31783));
  hi1s1 __90_509975(.DIN (_____9__25613), .Q (_________38177));
  nor2s1 ___9_9_509976(.DIN1 (____99__25585), .DIN2 (____0___24557), .Q
       (_________34207));
  nnd2s1 ___9_0_509977(.DIN1 (________24385), .DIN2 (___9_____39548),
       .Q (___00_0__39902));
  nnd2s1 ___9___509978(.DIN1 (________24375), .DIN2 (________22655), .Q
       (_________37614));
  nnd2s1 ___9___509979(.DIN1 (________24598), .DIN2 (___99___25119), .Q
       (___00____39929));
  hi1s1 ___9_509980(.DIN (___0____25136), .Q (____9____32424));
  hi1s1 ___9_0_509981(.DIN (___99___25116), .Q (____9_9__32410));
  nor2s1 ______509982(.DIN1 (___9_9__25114), .DIN2 (___9____24137), .Q
       (___990__25115));
  nor2s1 _____9_509983(.DIN1 (____00__24267), .DIN2 (________24484), .Q
       (___9____25113));
  nnd2s1 _______509984(.DIN1 (________24947), .DIN2 (________22476), .Q
       (___9____25112));
  nnd2s1 ___9_509985(.DIN1 (_____9__25000), .DIN2 (___9____25110), .Q
       (___9____25111));
  nnd2s1 ______509986(.DIN1 (___9____25108), .DIN2 (____9___22732), .Q
       (___9____25109));
  nor2s1 _______509987(.DIN1 (_____0__23377), .DIN2 (________23996), .Q
       (___9____25107));
  nnd2s1 _______509988(.DIN1 (_____0__24876), .DIN2 (________24020), .Q
       (___9____25106));
  and2s1 ___9_0_509989(.DIN1 (____0___24270), .DIN2 (_____0__26418), .Q
       (___9_0__25105));
  nor2s1 ______509990(.DIN1 (_____9__23718), .DIN2 (___0_0__24208), .Q
       (___9_9__25104));
  or2s1 _______509991(.DIN1 (___9____25102), .DIN2 (___0____24194), .Q
       (___9____25103));
  nnd2s1 _____9_509992(.DIN1 (________24005), .DIN2 (____0___26146), .Q
       (___9____25101));
  or2s1 _______509993(.DIN1 (___0_____40497), .DIN2 (____9____38001),
       .Q (___9____25100));
  nnd2s1 ______509994(.DIN1 (________23954), .DIN2 (________25751), .Q
       (___9____25099));
  nor2s1 _______509995(.DIN1 (________24995), .DIN2 (___9____24152), .Q
       (___9____25098));
  hi1s1 __90___509996(.DIN (________29208), .Q (___9____25097));
  nnd2s1 ___9_0_509997(.DIN1 (________24299), .DIN2 (___9_0__25095), .Q
       (___9____25096));
  nnd2s1 ___9_9_509998(.DIN1 (___9____25093), .DIN2 (_____0__23329), .Q
       (___9_9__25094));
  nor2s1 ___9___509999(.DIN1 (___0____25152), .DIN2 (___9____24115), .Q
       (___9____25092));
  hi1s1 __90___510000(.DIN (___9____27790), .Q (___9____25090));
  nor2s1 ___9___510001(.DIN1 (_________36761), .DIN2 (___0_____40650),
       .Q (___9____25089));
  hi1s1 _______510002(.DIN (________29112), .Q (___9____25088));
  or2s1 _______510003(.DIN1 (________22480), .DIN2 (________25394), .Q
       (___9_0__25087));
  nnd2s1 _____0_510004(.DIN1 (___0____24192), .DIN2 (___9____25085), .Q
       (___9____25086));
  and2s1 _____9_510005(.DIN1 (__9_____30046), .DIN2 (___0_____40445),
       .Q (___9____25084));
  and2s1 ___9___510006(.DIN1 (______0__34855), .DIN2
       (_________________________________________________________________________________________22095),
       .Q (___9____25083));
  nor2s1 _______510007(.DIN1 (_______22285), .DIN2 (___9____25081), .Q
       (___9____25082));
  nor2s1 _______510008(.DIN1 (___9____25079), .DIN2 (___0____24190), .Q
       (___9____25080));
  nor2s1 ______510009(.DIN1 (________25272), .DIN2 (________24873), .Q
       (___9_0__25078));
  nor2s1 ___9__510010(.DIN1 (________25438), .DIN2 (___9_0__24129), .Q
       (___9_9__25077));
  nnd2s1 _______510011(.DIN1 (___0____24213), .DIN2 (________23485), .Q
       (___9____25076));
  nor2s1 ___9___510012(.DIN1 (________25742), .DIN2 (___9____24116), .Q
       (___9____25075));
  nor2s1 ___9___510013(.DIN1 (________23772), .DIN2 (________23940), .Q
       (___9____25074));
  or2s1 ___9_510014(.DIN1 (_____0___32287), .DIN2 (______0__35050), .Q
       (___9____25073));
  nor2s1 _______510015(.DIN1
       (__________________________________________0___21981), .DIN2
       (__9_____30046), .Q (___9____25072));
  nnd2s1 ______510016(.DIN1 (________24024), .DIN2 (___00___25131), .Q
       (___9____25071));
  nor2s1 ___9_0_510017(.DIN1 (________26307), .DIN2 (___09___24259), .Q
       (___9____25070));
  or2s1 _______510018(.DIN1 (___9_0__25068), .DIN2 (___9____24124), .Q
       (___9____25069));
  nor2s1 _______510019(.DIN1 (________23898), .DIN2 (___0____24199), .Q
       (___9_9__25067));
  nnd2s1 _______510020(.DIN1 (___9____24141), .DIN2 (____99__23880), .Q
       (___9____25066));
  hi1s1 __90___510021(.DIN (___9____25064), .Q (___9____25065));
  nor2s1 ______510022(.DIN1 (_______22223), .DIN2 (___0____24246), .Q
       (___9____25063));
  nnd2s1 ___9_0_510023(.DIN1 (________24018), .DIN2 (___000__25125), .Q
       (___9____25062));
  nor2s1 ___9_0_510024(.DIN1 (___9____25060), .DIN2 (________24035), .Q
       (___9____25061));
  nor2s1 ___9_0_510025(.DIN1 (___0____22345), .DIN2 (____9____35258),
       .Q (___9____25059));
  nor2s1 ___9_0_510026(.DIN1 (___9_9__25057), .DIN2 (___9_0__24100), .Q
       (___9_0__25058));
  nnd2s1 ___9_9_510027(.DIN1 (___9_9__24138), .DIN2 (____0___23045), .Q
       (___9____25056));
  nnd2s1 ___9__510028(.DIN1 (________24920), .DIN2 (___0____26099), .Q
       (___9____25055));
  hi1s1 ___9___510029(.DIN (___9____25053), .Q (___9____25054));
  nnd2s1 ___990_510030(.DIN1 (________25282), .DIN2 (________25749), .Q
       (___9____25052));
  nor2s1 ___9___510031(.DIN1 (________24881), .DIN2 (___0_0__24198), .Q
       (___9____25051));
  nnd2s1 ___9__510032(.DIN1 (____9____38001), .DIN2 (_________32159),
       .Q (___9____25050));
  nnd2s1 ___9___510033(.DIN1 (__9_____30046), .DIN2 (________22964), .Q
       (___9____25049));
  nor2s1 _____510034(.DIN1 (___9_9__25047), .DIN2 (________24906), .Q
       (___9_0__25048));
  nor2s1 ___9___510035(.DIN1 (____9___23786), .DIN2 (___9____24130), .Q
       (___9____25046));
  nnd2s1 ___9___510036(.DIN1 (________24596), .DIN2 (___9_9__26020), .Q
       (___9____25045));
  and2s1 _______510037(.DIN1 (___00___24175), .DIN2 (________26269), .Q
       (___9____25044));
  nor2s1 _____9_510038(.DIN1 (________24976), .DIN2 (________24852), .Q
       (___9____25043));
  or2s1 ___9___510039(.DIN1 (___0__0__40581), .DIN2 (____9____38001),
       .Q (___9____25042));
  or2s1 ___9___510040(.DIN1 (________25257), .DIN2 (___0____24225), .Q
       (___9____25041));
  nnd2s1 ___9___510041(.DIN1 (___9____25039), .DIN2 (____0___23409), .Q
       (___9____25040));
  nnd2s1 ___9__510042(.DIN1 (___9____24147), .DIN2 (____0___26146), .Q
       (___9_0__25038));
  nnd2s1 ___9___510043(.DIN1 (___90___25035), .DIN2 (___0_0__22307), .Q
       (___909__25037));
  nnd2s1 ___9___510044(.DIN1 (___90___25035), .DIN2 (___0____22312), .Q
       (___90___25036));
  hi1s1 __90___510045(.DIN (___90___25032), .Q (___90___25033));
  nnd2s1 ___9___510046(.DIN1 (___0____24242), .DIN2 (___90___25030), .Q
       (___90___25031));
  nor2s1 __90__510047(.DIN1 (____99__25028), .DIN2 (_____9__24954), .Q
       (___900__25029));
  or2s1 _______510048(.DIN1 (___0__0__40591), .DIN2 (_____9___36005),
       .Q (____9___25027));
  nnd2s1 ______510049(.DIN1 (___0____24223), .DIN2 (____09__22948), .Q
       (____9___25026));
  nnd2s1 _______510050(.DIN1 (___00___24171), .DIN2 (________23547), .Q
       (____9___25025));
  nor2s1 _______510051(.DIN1 (________24052), .DIN2 (___0____23295), .Q
       (____9___25024));
  nnd2s1 ______510052(.DIN1 (________24281), .DIN2 (________24523), .Q
       (____9___25022));
  nnd2s1 ______510053(.DIN1 (___9____24113), .DIN2 (________25923), .Q
       (____9___25021));
  nor2s1 _______510054(.DIN1 (_____9__25019), .DIN2 (________25018), .Q
       (____90__25020));
  nnd2s1 __90_510055(.DIN1 (___0____24234), .DIN2 (_____9__24635), .Q
       (________25017));
  nnd2s1 _______510056(.DIN1 (____9___24739), .DIN2 (___0____23283), .Q
       (________25016));
  nor2s1 _____510057(.DIN1 (________22612), .DIN2 (___0____24214), .Q
       (________25015));
  nor2s1 _______510058(.DIN1 (________23070), .DIN2 (________25013), .Q
       (________25014));
  nor2s1 _______510059(.DIN1 (____99__25028), .DIN2 (___0____24249), .Q
       (________25012));
  nor2s1 _______510060(.DIN1
       (______________________________________________21982), .DIN2
       (__9_____30046), .Q (________25011));
  nor2s1 ______510061(.DIN1 (_____9__22730), .DIN2 (____99__24934), .Q
       (_____0__25010));
  or2s1 _______510062(.DIN1 (_____00__34847), .DIN2 (___0____24196), .Q
       (_____9__25009));
  nor2s1 _______510063(.DIN1 (_____9__23529), .DIN2 (___9____24107), .Q
       (________25008));
  nnd2s1 _______510064(.DIN1 (___0____24226), .DIN2 (________23388), .Q
       (________25007));
  nor2s1 __9000_(.DIN1 (________23549), .DIN2 (________23943), .Q
       (________25006));
  nnd2s1 _______510065(.DIN1 (________25004), .DIN2 (inData[2]), .Q
       (________25005));
  nor2s1 __90_9_510066(.DIN1 (________23654), .DIN2 (____99__25028), .Q
       (________25003));
  or2s1 __90___510067(.DIN1 (____9___25860), .DIN2 (___0_0__24178), .Q
       (________25002));
  nnd2s1 ___9__510068(.DIN1 (_____9__25000), .DIN2 (____0___25229), .Q
       (_____0__25001));
  and2s1 ___9___510069(.DIN1 (________24998), .DIN2 (____90__25758), .Q
       (________24999));
  hi1s1 __90_9_510070(.DIN (____0_9__38073), .Q (________24997));
  nor2s1 ___9___510071(.DIN1 (________24995), .DIN2 (___9____24133), .Q
       (________24996));
  nnd2s1 __90__510072(.DIN1 (________24284), .DIN2 (________24993), .Q
       (________24994));
  or2s1 ___9___510073(.DIN1 (___9_9__25114), .DIN2 (___9____24098), .Q
       (________24992));
  nor2s1 ___9___510074(.DIN1 (____9___27298), .DIN2 (________24043), .Q
       (_____0__24991));
  nor2s1 _____0_510075(.DIN1 (________23456), .DIN2 (________24989), .Q
       (_____9__24990));
  nor2s1 ___9_0_510076(.DIN1 (____9___22444), .DIN2 (____9____35258),
       .Q (________24988));
  nor2s1 ___9__510077(.DIN1 (________25278), .DIN2 (___0____24231), .Q
       (________24987));
  or2s1 ___9__510078(.DIN1 (___9_9__25114), .DIN2 (___9____24122), .Q
       (________24986));
  or2s1 ___9_9_510079(.DIN1 (________24984), .DIN2 (_________36858), .Q
       (________24985));
  hi1s1 __90___510080(.DIN (________24982), .Q (_____9__24983));
  nor2s1 ___9___510081(.DIN1 (________22673), .DIN2 (________24870), .Q
       (________24981));
  nnd2s1 ___9___510082(.DIN1 (___00___24173), .DIN2 (____0___22648), .Q
       (________24980));
  nnd2s1 _____510083(.DIN1 (___0_9__24207), .DIN2 (________24978), .Q
       (________24979));
  nor2s1 _____9_510084(.DIN1 (________24976), .DIN2 (________24952), .Q
       (________24977));
  nor2s1 ___9__510085(.DIN1 (___0___22275), .DIN2 (________25004), .Q
       (________24975));
  nnd2s1 _____510086(.DIN1 (________24878), .DIN2 (____9___24455), .Q
       (_____0__24974));
  nor2s1 ___9___510087(.DIN1 (________26530), .DIN2 (___9____24132), .Q
       (_____9__24973));
  nnd2s1 ___9___510088(.DIN1 (_____9__24001), .DIN2 (inData[18]), .Q
       (________24972));
  nor2s1 _______510089(.DIN1 (_____9__23834), .DIN2 (________25004), .Q
       (________24971));
  nnd2s1 _______510090(.DIN1 (___9____24097), .DIN2 (________24488), .Q
       (________24970));
  nor2s1 __90__510091(.DIN1 (________24968), .DIN2 (________24353), .Q
       (________24969));
  nor2s1 _____9_510092(.DIN1 (________24475), .DIN2 (________24019), .Q
       (________24967));
  nnd2s1 _____9_510093(.DIN1 (___9_9__24099), .DIN2 (_________32918),
       .Q (________24966));
  nor2s1 _____0_510094(.DIN1 (___0____24224), .DIN2 (_____9__24964), .Q
       (_____0__24965));
  or2s1 _______510095(.DIN1
       (______________________________________0______21886), .DIN2
       (__9_____30046), .Q (________24963));
  nor2s1 _______510096(.DIN1 (___9____24126), .DIN2 (________25278), .Q
       (________24962));
  nor2s1 _______510097(.DIN1 (________23092), .DIN2 (________24014), .Q
       (________24961));
  nnd2s1 _______510098(.DIN1 (_____0__25479), .DIN2 (___0____24255), .Q
       (________24960));
  nor2s1 _______510099(.DIN1 (________26280), .DIN2 (____0___24939), .Q
       (________24959));
  nor2s1 _______510100(.DIN1 (_____0__25417), .DIN2 (_____0__24696), .Q
       (________24958));
  nor2s1 _______510101(.DIN1 (________22917), .DIN2 (____9____35258),
       .Q (________24957));
  and2s1 ______510102(.DIN1 (__9_____30046), .DIN2 (________22895), .Q
       (________24956));
  nor2s1 _______510103(.DIN1 (____0___24272), .DIN2 (_____9__24954), .Q
       (_____0__24955));
  nor2s1 _______510104(.DIN1 (________24853), .DIN2 (________24952), .Q
       (________24953));
  and2s1 _______510105(.DIN1 (___9_0__24109), .DIN2 (________23528), .Q
       (________24951));
  nnd2s1 _______510106(.DIN1 (________24009), .DIN2 (________23542), .Q
       (________24950));
  nor2s1 _______510107(.DIN1 (________25742), .DIN2 (________24417), .Q
       (________24949));
  nnd2s1 _______510108(.DIN1 (________24947), .DIN2 (________24514), .Q
       (________24948));
  nnd2s1 _______510109(.DIN1 (____0___23975), .DIN2 (________23623), .Q
       (________24946));
  nnd2s1 _______510110(.DIN1 (_________41345), .DIN2
       (_____________________________________9_______21881), .Q
       (_____0__24945));
  and2s1 _______510111(.DIN1 (____0___24268), .DIN2 (___90___25030), .Q
       (____09__24944));
  nnd2s1 _______510112(.DIN1 (______9__37314), .DIN2 (inData[26]), .Q
       (____0___24943));
  nnd2s1 _______510113(.DIN1 (________24015), .DIN2 (________23556), .Q
       (____0___24942));
  nnd2s1 _____510114(.DIN1 (_____9__23961), .DIN2 (________23932), .Q
       (____0___24941));
  nor2s1 _____9_510115(.DIN1 (____9___25860), .DIN2 (____0___24939), .Q
       (____0___24940));
  or2s1 _____9_510116(.DIN1 (___0____22299), .DIN2 (___9____25081), .Q
       (____0___24938));
  nor2s1 _____9_510117(.DIN1 (_____0__22403), .DIN2 (___9____25081), .Q
       (____0___24937));
  nnd2s1 _____0_510118(.DIN1 (___0____24206), .DIN2 (___9____24153), .Q
       (____0___24936));
  nor2s1 _____0_510119(.DIN1 (________24661), .DIN2 (____99__24934), .Q
       (____00__24935));
  or2s1 _____0_510120(.DIN1 (__99_9__30508), .DIN2 (___9_9__24128), .Q
       (____9___24933));
  nor2s1 _____0_510121(.DIN1 (________22398), .DIN2 (____9_9__37052),
       .Q (____9___24932));
  nor2s1 ______510122(.DIN1 (________24418), .DIN2 (____00__23972), .Q
       (____9___24931));
  nnd2s1 _______510123(.DIN1 (___0____24209), .DIN2 (________22955), .Q
       (____9___24930));
  nor2s1 _______510124(.DIN1 (____9___24928), .DIN2 (____9___24927), .Q
       (____9___24929));
  nor2s1 _______510125(.DIN1
       (_____________________________________9_______21878), .DIN2
       (____9_9__37052), .Q (____9___24926));
  nor2s1 __90___510126(.DIN1 (___0____23240), .DIN2 (________23899), .Q
       (____90__24925));
  nor2s1 _______510127(.DIN1 (_____0__22919), .DIN2 (___0_9__24227), .Q
       (_____9__24924));
  nor2s1 _______510128(.DIN1 (________24922), .DIN2 (________24900), .Q
       (________24923));
  nnd2s1 _______510129(.DIN1 (________24920), .DIN2 (________25458), .Q
       (________24921));
  and2s1 ______510130(.DIN1 (_____9__24051), .DIN2 (________23736), .Q
       (________24919));
  nnd2s1 _______510131(.DIN1 (___00___24174), .DIN2 (_____0__23068), .Q
       (________24918));
  nor2s1 _______510132(.DIN1 (_______22232), .DIN2 (________25004), .Q
       (________24917));
  or2s1 _______510133(.DIN1 (____9___25023), .DIN2 (________24050), .Q
       (________24916));
  nnd2s1 ______510134(.DIN1 (_________41345), .DIN2
       (_____________________________________9_______21882), .Q
       (_____0__24915));
  nnd2s1 _______510135(.DIN1 (________24054), .DIN2 (____9___23970), .Q
       (_____9__24914));
  and2s1 _______510136(.DIN1 (________24912), .DIN2 (___00___22288), .Q
       (________24913));
  nor2s1 _______510137(.DIN1 (____0___25590), .DIN2 (___0____24185), .Q
       (________24911));
  hi1s1 __90___510138(.DIN (______0__31903), .Q (___0____27870));
  nor2s1 __900__(.DIN1 (____0___24840), .DIN2 (________24968), .Q
       (___0____25187));
  hi1s1 __90__510139(.DIN (_____0__26599), .Q (________25647));
  nor2s1 _______510140(.DIN1 (________24910), .DIN2 (____0___24939), .Q
       (________25752));
  hi1s1 __90___510141(.DIN (________27313), .Q (____0___25589));
  nor2s1 ___9___510142(.DIN1 (________25257), .DIN2 (_____9__24964), .Q
       (____9___25584));
  nnd2s1 ___9___510143(.DIN1 (___9____24135), .DIN2
       (_____________________21682), .Q (_____0__25729));
  hi1s1 __90___510144(.DIN (_____0__25271), .Q (________25620));
  nnd2s1 ___9___510145(.DIN1 (________24899), .DIN2 (________24909), .Q
       (_____0__25379));
  hi1s1 ___9__510146(.DIN (___0____26115), .Q (________26181));
  nor2s1 __90___510147(.DIN1 (____0___29012), .DIN2 (________24908), .Q
       (____0___25316));
  nor2s1 ___9___510148(.DIN1 (________24568), .DIN2 (________24701), .Q
       (___99___25116));
  nnd2s1 ___9___510149(.DIN1 (_____9__24335), .DIN2 (________24704), .Q
       (___0____25150));
  nnd2s1 __90__510150(.DIN1 (________24789), .DIN2 (________24723), .Q
       (________25483));
  nor2s1 ___9___510151(.DIN1 (________25324), .DIN2 (________24756), .Q
       (___99___25122));
  or2s1 ___909_510152(.DIN1 (________23490), .DIN2 (________24680), .Q
       (____09__25318));
  hi1s1 _______510153(.DIN (________24907), .Q (____9___25760));
  hi1s1 ______510154(.DIN (_____9__28100), .Q (____9___25765));
  nor2s1 ___9___510155(.DIN1 (________25360), .DIN2 (________24892), .Q
       (___0_0__25145));
  hi1s1 _______510156(.DIN (_________34154), .Q (________27161));
  nnd2s1 ____9__510157(.DIN1 (_____9__24904), .DIN2 (________25355), .Q
       (________25372));
  nor2s1 ___9_9_510158(.DIN1 (____0___29012), .DIN2 (________24482), .Q
       (___0____25151));
  nor2s1 _______510159(.DIN1 (___9_9__25057), .DIN2 (________24761), .Q
       (____0___25500));
  nnd2s1 _______510160(.DIN1 (________24903), .DIN2 (_____0__24726), .Q
       (________25731));
  nnd2s1 ______510161(.DIN1 (________24887), .DIN2 (___00___25129), .Q
       (_____9__25747));
  nor2s1 _______510162(.DIN1 (________24906), .DIN2 (________23714), .Q
       (____9___25579));
  nnd2s1 _______510163(.DIN1 (________24891), .DIN2 (_____0__24905), .Q
       (________25732));
  nor2s1 _______510164(.DIN1 (________24480), .DIN2 (_____0__26528), .Q
       (________25807));
  nor2s1 ______510165(.DIN1 (_____________________21742), .DIN2
       (____9___23967), .Q (____09__25506));
  nor2s1 _______510166(.DIN1 (________26440), .DIN2 (___0____24210), .Q
       (________25739));
  and2s1 _______510167(.DIN1 (_____9__24904), .DIN2 (________25944), .Q
       (_____0__25901));
  nor2s1 ____9__510168(.DIN1 (_______22278), .DIN2 (___0____24236), .Q
       (________25811));
  nnd2s1 ____9__510169(.DIN1 (________24903), .DIN2 (________24909), .Q
       (_____0__27177));
  nnd2s1 ____90_510170(.DIN1 (________24027), .DIN2 (________24713), .Q
       (___0____26098));
  nnd2s1 _____9_510171(.DIN1 (________25551), .DIN2 (________24902), .Q
       (____0___26687));
  nnd2s1 ____9__510172(.DIN1 (___0_9__24237), .DIN2 (________24490), .Q
       (____9___25764));
  nor2s1 ____9__510173(.DIN1 (________24901), .DIN2 (________24900), .Q
       (_____9__26447));
  nnd2s1 ____9__510174(.DIN1 (___9____24091), .DIN2 (________25559), .Q
       (________28876));
  nor2s1 ____9_510175(.DIN1 (___0____24239), .DIN2 (____0___24750), .Q
       (________28057));
  nnd2s1 ____9__510176(.DIN1 (________24899), .DIN2 (________24898), .Q
       (_____9__25757));
  and2s1 ____9__510177(.DIN1 (____9___23969), .DIN2 (_____9__25348), .Q
       (___0____26096));
  dffacs1 _________________________________________0_____510178(.CLRB
       (reset), .CLK (clk), .DIN (___9_9__24148), .QN
       (_____________________________________0_______21758));
  nnd2s1 __90___510179(.DIN1 (______0__32803), .DIN2 (________24298),
       .Q (_____0___33165));
  hi1s1 ___9___510180(.DIN (_____0__26295), .Q (________28850));
  nnd2s1 ___9___510181(.DIN1 (___99___24160), .DIN2 (_____0__24905), .Q
       (_____0__26832));
  nnd2s1 ____90_510182(.DIN1 (________24890), .DIN2 (___0____25146), .Q
       (_____0__27039));
  hi1s1 __90___510183(.DIN (________24897), .Q (___00___27828));
  nnd2s1 __90___510184(.DIN1 (_____0__25748), .DIN2 (___009__24177), .Q
       (________25723));
  nnd2s1 ___9__510185(.DIN1 (________24717), .DIN2 (________24896), .Q
       (___0____26123));
  hi1s1 __90_9_510186(.DIN (_____9__25358), .Q (____0___25591));
  hi1s1 __90_0_510187(.DIN (_________38871), .Q (___90_0__39025));
  nor2s1 ___9___510188(.DIN1 (___9____24125), .DIN2 (____0_0__34423),
       .Q (________26637));
  hi1s1 ___9__510189(.DIN (________25340), .Q (__9_0___29726));
  nor2s1 ___9___510190(.DIN1 (________24476), .DIN2 (________24694), .Q
       (____9___25580));
  nnd2s1 ____9__510191(.DIN1 (________24903), .DIN2 (________25550), .Q
       (________26151));
  nnd2s1 ___9___510192(.DIN1 (____0___24749), .DIN2 (_____0__24895), .Q
       (________25834));
  and2s1 ___9_510193(.DIN1 (_____0__24755), .DIN2 (________25944), .Q
       (_________33217));
  and2s1 ___9___510194(.DIN1 (___9____24104), .DIN2 (___00___25129), .Q
       (________29088));
  nnd2s1 ___9___510195(.DIN1 (____09__23981), .DIN2 (________25362), .Q
       (__9_____30239));
  nor2s1 ___900_510196(.DIN1 (_____9__24894), .DIN2 (________24893), .Q
       (________29441));
  nnd2s1 ___90__510197(.DIN1 (________24889), .DIN2 (___99___25118), .Q
       (___0_____30789));
  nor2s1 ___90__510198(.DIN1 (________25735), .DIN2 (________24712), .Q
       (__9_____30335));
  nor2s1 ___9___510199(.DIN1 (________25600), .DIN2 (________24892), .Q
       (___09____31451));
  nnd2s1 ___9___510200(.DIN1 (_____0__24885), .DIN2 (____9___24833), .Q
       (__9__0__30234));
  and2s1 ___9___510201(.DIN1 (_____0__24716), .DIN2 (___0____25176), .Q
       (__99____30487));
  nnd2s1 ___9___510202(.DIN1 (________24729), .DIN2 (_____9__23757), .Q
       (___90___28649));
  nor2s1 ___90__510203(.DIN1 (___0____24240), .DIN2 (_____9__25434), .Q
       (___0_____30821));
  nnd2s1 ____9__510204(.DIN1 (________24891), .DIN2 (________24896), .Q
       (______9__32019));
  nor2s1 ____9_510205(.DIN1 (___0____25186), .DIN2 (____9___24743), .Q
       (___0_____31129));
  nnd2s1 ___90__510206(.DIN1 (________24890), .DIN2 (________25362), .Q
       (________28870));
  nnd2s1 ___9___510207(.DIN1 (________24709), .DIN2 (________25944), .Q
       (_________33570));
  nnd2s1 ___900_510208(.DIN1 (___9_0___39344), .DIN2 (________24889),
       .Q (________26239));
  hi1s1 ___9___510209(.DIN (___0____25178), .Q (____0___25594));
  hi1s1 ___9___510210(.DIN (________24888), .Q (___9____29571));
  nnd2s1 ___90__510211(.DIN1 (________24887), .DIN2 (___0____25157), .Q
       (___90___28653));
  nor2s1 __90___510212(.DIN1 (____9___24738), .DIN2 (________24778), .Q
       (___9____29606));
  nor2s1 __90__510213(.DIN1 (________24322), .DIN2 (________24719), .Q
       (________27638));
  dffacs1 _________________________________________0___9_(.CLRB
       (reset), .CLK (clk), .DIN (___09___24262), .Q (___0__0__40571));
  nor2s1 ___9___510214(.DIN1 (________24886), .DIN2 (_____0__24765), .Q
       (________26333));
  nnd2s1 ___9___510215(.DIN1 (___9____24143), .DIN2 (___0____25181), .Q
       (______9__33575));
  hi1s1 _______510216(.DIN (_________37230), .Q (______9__37419));
  nnd2s1 ___9___510217(.DIN1 (_____0__24885), .DIN2 (________24767), .Q
       (___0_____31366));
  nor2s1 ___90__510218(.DIN1 (________23906), .DIN2 (____9____38001),
       .Q (____0____38052));
  nnd2s1 ___90_510219(.DIN1 (________24721), .DIN2 (_____9__25348), .Q
       (________27694));
  nor2s1 ___90__510220(.DIN1 (___0____24184), .DIN2 (________25553), .Q
       (________28131));
  hi1s1 ___9___510221(.DIN (________25513), .Q (___0_9___40270));
  nor2s1 ___90__510222(.DIN1 (________23717), .DIN2 (________24006), .Q
       (_____9__28617));
  hi1s1 ___9___510223(.DIN (_________41335), .Q (_________34877));
  hi1s1 ___9___510224(.DIN (______0__41339), .Q (_________37199));
  nor2s1 ___90__510225(.DIN1 (________24884), .DIN2 (___0_0__24238), .Q
       (_____9___38512));
  nnd2s1 ___90__510226(.DIN1 (________24684), .DIN2 (________23608), .Q
       (_________32140));
  nnd2s1 ___510227(.DIN1 (____0___24271), .DIN2 (________23360), .Q
       (_________38860));
  hi1s1 __90___510228(.DIN (_________36480), .Q (_________37452));
  nor2s1 ___90__510229(.DIN1 (_________34145), .DIN2 (___0____24193),
       .Q (_____0___34932));
  nnd2s1 ___90__510230(.DIN1 (____0___24274), .DIN2 (________24883), .Q
       (_________38271));
  nor2s1 __90___510231(.DIN1 (________24882), .DIN2 (___9____25093), .Q
       (_________38576));
  nnd2s1 ___90_510232(.DIN1 (_____9__24041), .DIN2 (________24280), .Q
       (___9_____39554));
  nnd2s1 ___90__510233(.DIN1 (________24030), .DIN2 (____99__23406), .Q
       (___9_____39542));
  nnd2s1 ___90__510234(.DIN1 (___99___24161), .DIN2 (________23719), .Q
       (___009___39979));
  nor2s1 ___90__510235(.DIN1 (_____0__24411), .DIN2 (________24881), .Q
       (_________36512));
  nnd2s1 ___909_510236(.DIN1 (________24880), .DIN2 (____0___23411), .Q
       (_________38377));
  hi1s1 __90___510237(.DIN (________24879), .Q (_________32001));
  nnd2s1 ___90__510238(.DIN1 (________24878), .DIN2 (___9____23190), .Q
       (_____09__35744));
  nor2s1 ___9___510239(.DIN1 (________24877), .DIN2 (___0____24182), .Q
       (_________35394));
  nnd2s1 ___90_510240(.DIN1 (___0____24241), .DIN2 (_____0__24876), .Q
       (_________38743));
  nor2s1 _______510241(.DIN1 (___9____24112), .DIN2 (________24873), .Q
       (________24874));
  nor2s1 ___9_0_510242(.DIN1 (___0__9__40430), .DIN2 (___0__0__39993),
       .Q (________24872));
  or2s1 ______510243(.DIN1 (_____9__23557), .DIN2 (________24870), .Q
       (________24871));
  or2s1 _______510244(.DIN1 (________25850), .DIN2 (___0____24202), .Q
       (________24869));
  nnd2s1 __90___510245(.DIN1 (________24817), .DIN2 (inData[8]), .Q
       (________24868));
  hi1s1 __90__510246(.DIN (________25323), .Q (_____0__24867));
  and2s1 _____9_510247(.DIN1 (___9____24121), .DIN2 (________25829), .Q
       (_____9__24866));
  nnd2s1 ___9___510248(.DIN1 (________23941), .DIN2 (_____0__23387), .Q
       (________24865));
  hi1s1 ___9_0_510249(.DIN (________24863), .Q (________24864));
  or2s1 ___9___510250(.DIN1 (________24861), .DIN2 (________24860), .Q
       (________24862));
  nor2s1 ___9_9_510251(.DIN1
       (_____________________________________________21969), .DIN2
       (___99_0__39817), .Q (________24859));
  nor2s1 ___9___510252(.DIN1 (________24877), .DIN2 (___999__24167), .Q
       (________24858));
  nor2s1 ___9_9_510253(.DIN1 (________25272), .DIN2 (____0___23976), .Q
       (________24856));
  nor2s1 ___9___510254(.DIN1 (________23860), .DIN2 (_____9__24964), .Q
       (________24855));
  or2s1 ___9__510255(.DIN1 (________24853), .DIN2 (________24852), .Q
       (________24854));
  nnd2s1 ___9___510256(.DIN1 (________23988), .DIN2 (________25829), .Q
       (________24851));
  nor2s1 ___9___510257(.DIN1 (___9____23145), .DIN2 (___09___24264), .Q
       (________24850));
  hi1s1 ___9__510258(.DIN (____09__24848), .Q (_____0__24849));
  hi1s1 ___9__510259(.DIN (___090__25213), .Q (____0___24847));
  hi1s1 ___9___510260(.DIN (________25347), .Q (____0___24846));
  hi1s1 ___9___510261(.DIN (___9_0__27795), .Q (____0___24845));
  nnd2s1 ___9___510262(.DIN1 (______0__34855), .DIN2
       (_________________________________________________________________________________________22094),
       .Q (____0___24844));
  and2s1 ___9___510263(.DIN1 (________23997), .DIN2 (________25942), .Q
       (____0___24843));
  hi1s1 __90___510264(.DIN (_________31958), .Q (____0___24842));
  nor2s1 ___9___510265(.DIN1 (____0___24840), .DIN2 (____0___29012), .Q
       (____0___24841));
  nor2s1 ___9___510266(.DIN1 (_________________9___21685), .DIN2
       (________23945), .Q (____00__24839));
  or2s1 ___9_9_510267(.DIN1 (_________22024), .DIN2 (___99_0__39817),
       .Q (____99__24838));
  nnd2s1 ___9_0_510268(.DIN1 (___0__0__39993), .DIN2 (___0_____40437),
       .Q (____9___24837));
  nor2s1 ___9_0_510269(.DIN1 (______9__22026), .DIN2 (___0__0__39993),
       .Q (____9___24836));
  nor2s1 ___9_0_510270(.DIN1 (________26698), .DIN2 (___0__0__39993),
       .Q (____9___24835));
  nnd2s1 ___9___510271(.DIN1 (____9___24833), .DIN2 (________24766), .Q
       (____9___24834));
  nnd2s1 ___9___510272(.DIN1 (______0__32803), .DIN2 (___9__22165), .Q
       (____9___24832));
  nnd2s1 ___9___510273(.DIN1 (____9___24830), .DIN2 (________23958), .Q
       (____9___24831));
  hi1s1 ___9___510274(.DIN (________25377), .Q (____90__24829));
  hi1s1 ___9__510275(.DIN (____00__25407), .Q (_____9__24828));
  nnd2s1 ___9_9_510276(.DIN1 (______0__32803), .DIN2 (________22490),
       .Q (________24827));
  nnd2s1 ___99_510277(.DIN1 (________23937), .DIN2 (_____9__23444), .Q
       (________24826));
  nor2s1 ___99_510278(.DIN1 (________24824), .DIN2 (___0____24216), .Q
       (________24825));
  nor2s1 __900__510279(.DIN1 (________24821), .DIN2 (________24320), .Q
       (________24822));
  or2s1 __900__510280(.DIN1 (________24968), .DIN2 (________24567), .Q
       (_____0__24820));
  or2s1 __900__510281(.DIN1 (________25571), .DIN2 (_____9__24315), .Q
       (_____9__24819));
  nnd2s1 ___9___510282(.DIN1 (________24817), .DIN2
       (____________________________________________21867), .Q
       (________24818));
  or2s1 ___9__510283(.DIN1 (____9___24928), .DIN2 (________24007), .Q
       (________24815));
  hi1s1 __90___510284(.DIN (_____0__24812), .Q (________24813));
  nnd2s1 _____510285(.DIN1 (________24317), .DIN2
       (______________________________________0_______21894), .Q
       (_____9__24811));
  nor2s1 ___9_510286(.DIN1 (_____9__25823), .DIN2 (________23993), .Q
       (________24810));
  nor2s1 ___9__510287(.DIN1 (___0____22298), .DIN2 (________24808), .Q
       (________24809));
  hi1s1 __9____(.DIN (___0____25190), .Q (________24807));
  nor2s1 ___9___510288(.DIN1 (___9_9__25047), .DIN2 (________24483), .Q
       (________24806));
  and2s1 ___9_0_510289(.DIN1 (________23899), .DIN2 (___0__9__40420),
       .Q (________24805));
  nor2s1 ___9_0_510290(.DIN1 (___0_____40425), .DIN2 (___0__0__39993),
       .Q (_____0__24803));
  hi1s1 __90___510291(.DIN (________24801), .Q (_____9__24802));
  nor2s1 __90___510292(.DIN1 (________22985), .DIN2 (________23899), .Q
       (________24800));
  nor2s1 __90___510293(.DIN1 (________24786), .DIN2 (________24047), .Q
       (________24799));
  or2s1 __90___510294(.DIN1 (________24797), .DIN2 (_____9__24685), .Q
       (________24798));
  nor2s1 __90___510295(.DIN1 (________23709), .DIN2 (________24688), .Q
       (________24796));
  and2s1 ___9_510296(.DIN1 (________24920), .DIN2 (___9____23159), .Q
       (________24795));
  nor2s1 __90_0_510297(.DIN1 (_____9__24793), .DIN2 (________26611), .Q
       (_____0__24794));
  or2s1 __90___510298(.DIN1 (________24791), .DIN2 (________24785), .Q
       (________24792));
  nnd2s1 __90___510299(.DIN1 (________24789), .DIN2 (________24699), .Q
       (________24790));
  and2s1 __90___510300(.DIN1 (________24783), .DIN2 (___90___25034), .Q
       (________24788));
  or2s1 __90___510301(.DIN1 (________24786), .DIN2 (________24785), .Q
       (________24787));
  nnd2s1 __90_9_510302(.DIN1 (________24783), .DIN2 (________24782), .Q
       (_____9__24784));
  nor2s1 _______510303(.DIN1 (_____0___33534), .DIN2 (________24763),
       .Q (________24781));
  nor2s1 __90_0_510304(.DIN1 (________22622), .DIN2 (_____9__24793), .Q
       (________24780));
  nor2s1 __90___510305(.DIN1 (___09___23306), .DIN2 (________24778), .Q
       (________24779));
  or2s1 __90___510306(.DIN1 (_________37722), .DIN2 (____0___29012), .Q
       (________24777));
  nnd2s1 __90__510307(.DIN1 (________25282), .DIN2 (_____0__24775), .Q
       (________24776));
  hi1s1 __90___510308(.DIN (________24773), .Q (_____9__24774));
  and2s1 __90___510309(.DIN1 (________24771), .DIN2 (________25942), .Q
       (________24772));
  and2s1 __90___510310(.DIN1 (________24769), .DIN2 (________24768), .Q
       (________24770));
  nor2s1 _____9_510311(.DIN1 (____99__25028), .DIN2 (________24025), .Q
       (________25361));
  nnd2s1 __900_0(.DIN1 (________24767), .DIN2 (________24766), .Q
       (________25568));
  nor2s1 __90___510312(.DIN1 (____99__25585), .DIN2 (________24692), .Q
       (___009__25134));
  nor2s1 ___9___510313(.DIN1 (________23908), .DIN2 (_____0__24765), .Q
       (___9____25980));
  nnd2s1 _______510314(.DIN1 (_____9__24429), .DIN2 (_____0__24905), .Q
       (________26814));
  nnd2s1 _______510315(.DIN1 (___0____24200), .DIN2
       (____0________________21720), .Q (________25548));
  nor2s1 __90___510316(.DIN1 (________24285), .DIN2 (________24730), .Q
       (_____0__25359));
  hi1s1 ___9___510317(.DIN (_____9__24764), .Q (________25547));
  nor2s1 _______510318(.DIN1 (________25850), .DIN2 (________24763), .Q
       (________25525));
  hi1s1 ___9___510319(.DIN (_____0__25461), .Q (________27421));
  nor2s1 ___9__510320(.DIN1 (________23069), .DIN2 (_________41345), .Q
       (________25792));
  nor2s1 ___9___510321(.DIN1 (________24762), .DIN2 (________24761), .Q
       (________25727));
  nnd2s1 ___9___510322(.DIN1 (_____0__24002), .DIN2 (________24760), .Q
       (____0___25224));
  nnd2s1 ___9___510323(.DIN1 (________24529), .DIN2 (___9____25110), .Q
       (________25743));
  hi1s1 __90___510324(.DIN (________24759), .Q (________29439));
  hi1s1 __90___510325(.DIN (________24758), .Q (________25557));
  nor2s1 ___9___510326(.DIN1 (________24757), .DIN2 (________24756), .Q
       (________25374));
  nnd2s1 ___9___510327(.DIN1 (____9___24741), .DIN2 (___0____25157), .Q
       (____9___25494));
  nnd2s1 ___9___510328(.DIN1 (_____0__24755), .DIN2 (___0____25146), .Q
       (________25246));
  nor2s1 __90_0_510329(.DIN1 (____9___23970), .DIN2 (_____9__24793), .Q
       (________25475));
  nor2s1 ___9___510330(.DIN1 (____0________________21716), .DIN2
       (___0____24181), .Q (________25515));
  hi1s1 __90___510331(.DIN (____0___24754), .Q (_____9__25622));
  hi1s1 __90___510332(.DIN (____0___24753), .Q (________25562));
  hi1s1 __90___510333(.DIN (____0___24752), .Q (____0___25592));
  nnd2s1 ___9___510334(.DIN1 (___00___25130), .DIN2 (________23985), .Q
       (_____0__26371));
  hi1s1 __90___510335(.DIN (___0_9__25184), .Q (________25561));
  nnd2s1 __90__510336(.DIN1 (________24789), .DIN2 (____90__24736), .Q
       (_____9__25328));
  nor2s1 __90__510337(.DIN1 (________25345), .DIN2 (_____0__23952), .Q
       (___0_9__25174));
  nnd2s1 __90__510338(.DIN1 (________23955), .DIN2 (____9___24452), .Q
       (________25554));
  hi1s1 ___9__510339(.DIN (____0___24751), .Q (__90____29649));
  or2s1 ___9__510340(.DIN1 (________25371), .DIN2 (_____9__24011), .Q
       (____9___25582));
  nor2s1 ___9___510341(.DIN1 (___990__24158), .DIN2 (____0___24750), .Q
       (___9____25970));
  nor2s1 ___9___510342(.DIN1 (___0____25186), .DIN2 (_____9__24735), .Q
       (___0____25148));
  hi1s1 ___9___510343(.DIN (_________33016), .Q (________26605));
  nnd2s1 ___9___510344(.DIN1 (____0___24749), .DIN2 (____0___24748), .Q
       (___0_9__26121));
  nor2s1 ___9___510345(.DIN1 (________26280), .DIN2 (_____0__23992), .Q
       (___0____25141));
  nor2s1 ___9___510346(.DIN1 (____0___23977), .DIN2 (________24732), .Q
       (________25736));
  nnd2s1 ___9___510347(.DIN1 (_____0__24686), .DIN2 (________23091), .Q
       (___0____26105));
  nor2s1 __90___510348(.DIN1 (____0___24747), .DIN2 (____9___24737), .Q
       (________26306));
  nnd2s1 __90___510349(.DIN1 (___9____24150), .DIN2 (____00__24746), .Q
       (_____0__26438));
  nnd2s1 __90_9_510350(.DIN1 (_____9__24793), .DIN2 (____99__24745), .Q
       (____0___25588));
  hi1s1 ___9___510351(.DIN (____9___24744), .Q (_____9__25565));
  nor2s1 ____9_510352(.DIN1 (________25600), .DIN2 (____9___24743), .Q
       (________25341));
  nor2s1 ___9___510353(.DIN1 (_____0__25339), .DIN2 (________24892), .Q
       (____9___25761));
  nor2s1 ___9___510354(.DIN1 (____9___24742), .DIN2 (________24728), .Q
       (_____9__26437));
  nor2s1 ___9___510355(.DIN1 (____0________________21716), .DIN2
       (___000__24168), .Q (________25754));
  nnd2s1 ___9_510356(.DIN1 (____9___24741), .DIN2 (___00___25129), .Q
       (________25342));
  nor2s1 ___9___510357(.DIN1 (________23844), .DIN2 (________24761), .Q
       (_____0__25243));
  nor2s1 __90___510358(.DIN1 (________24731), .DIN2 (_____0__24032), .Q
       (___0____25139));
  hi1s1 __90___510359(.DIN (____9___24740), .Q (________28152));
  nnd2s1 ___9_510360(.DIN1 (____9___24739), .DIN2 (_____0__23929), .Q
       (________25321));
  hi1s1 __90___510361(.DIN (________26755), .Q (___9____26010));
  nnd2s1 __90__510362(.DIN1 (____9___26406), .DIN2 (___0_9__23272), .Q
       (________25448));
  or2s1 __90_9_510363(.DIN1 (____9___24738), .DIN2 (____9___24737), .Q
       (___90___25963));
  nor2s1 ___9___510364(.DIN1 (________27043), .DIN2 (___9_____39332),
       .Q (________25898));
  nor2s1 ___9_510365(.DIN1 (_________34145), .DIN2 (________23987), .Q
       (_____9__25738));
  nor2s1 ___9___510366(.DIN1 (________25294), .DIN2 (________24892), .Q
       (____0___29202));
  nnd2s1 ___9_0_510367(.DIN1 (________24724), .DIN2 (____90__24736), .Q
       (____9___25854));
  nnd2s1 ___9_0_510368(.DIN1 (___9_9__24118), .DIN2 (________25355), .Q
       (________26430));
  nor2s1 ___9___510369(.DIN1 (________25360), .DIN2 (_____9__24735), .Q
       (____0___25769));
  or2s1 __90___510370(.DIN1 (____0___24747), .DIN2 (________24288), .Q
       (___0____27013));
  nor2s1 __90___510371(.DIN1 (________24734), .DIN2 (____99__25028), .Q
       (________25690));
  nor2s1 __90___510372(.DIN1 (____99__25028), .DIN2 (________24733), .Q
       (____09__25595));
  or2s1 __90___510373(.DIN1 (____9___24738), .DIN2 (________23956), .Q
       (_____9__25937));
  nnd2s1 __90___510374(.DIN1 (________24386), .DIN2 (________24767), .Q
       (________25560));
  nor2s1 ___9_0_510375(.DIN1 (________23805), .DIN2 (________24732), .Q
       (____9___25762));
  nor2s1 __90__510376(.DIN1 (____0___24747), .DIN2 (________24778), .Q
       (________25573));
  nor2s1 __90_9_510377(.DIN1 (________24731), .DIN2 (________24714), .Q
       (__9_0___30000));
  nor2s1 __90___510378(.DIN1 (____0___24747), .DIN2 (________24730), .Q
       (________26279));
  nnd2s1 _____9_510379(.DIN1 (___9____24151), .DIN2 (________26431), .Q
       (_____0__25815));
  nor2s1 ____90_510380(.DIN1 (________23335), .DIN2 (________24040), .Q
       (________25831));
  hi1s1 __90_0_510381(.DIN (______9__35584), .Q (_________35526));
  nnd2s1 ___9___510382(.DIN1 (________24729), .DIN2 (________24474), .Q
       (____90__27382));
  nor2s1 ___9___510383(.DIN1 (________23866), .DIN2 (________24728), .Q
       (____9____32436));
  nor2s1 ___9__510384(.DIN1 (________24727), .DIN2 (___9____24094), .Q
       (________28500));
  nor2s1 ___9__510385(.DIN1 (________24727), .DIN2 (_____9__24725), .Q
       (____90__25948));
  nnd2s1 ___9___510386(.DIN1 (____0___24648), .DIN2 (_____0__24726), .Q
       (_____9__26737));
  nor2s1 ____9_510387(.DIN1 (___0____23266), .DIN2 (________24728), .Q
       (_____0__26428));
  nor2s1 ___9__510388(.DIN1 (____99__25585), .DIN2 (_____9__24725), .Q
       (_____0__29262));
  and2s1 ___9_0_510389(.DIN1 (________24724), .DIN2 (________24723), .Q
       (_____9__26812));
  nnd2s1 ___9___510390(.DIN1 (____9_9__37052), .DIN2 (________25946),
       .Q (______0__36932));
  nor2s1 __90___510391(.DIN1 (________24821), .DIN2 (________24908), .Q
       (____9___25583));
  nnd2s1 ___9__510392(.DIN1 (_____0__24885), .DIN2 (____00__24746), .Q
       (___9____26915));
  nnd2s1 ___9_0_510393(.DIN1 (________24722), .DIN2 (________23983), .Q
       (___0_0__26092));
  nor2s1 ___9_510394(.DIN1 (________24010), .DIN2 (________24732), .Q
       (____9___25759));
  nor2s1 ___9___510395(.DIN1 (________25294), .DIN2 (_____9__24735), .Q
       (________26666));
  and2s1 ___9__510396(.DIN1 (________24721), .DIN2 (___99___25123), .Q
       (________25783));
  nnd2s1 ____9__510397(.DIN1 (________24891), .DIN2 (________25550), .Q
       (_____0__26758));
  nnd2s1 ___9___510398(.DIN1 (________24899), .DIN2 (_____0__24726), .Q
       (___0_____31376));
  nnd2s1 __90___510399(.DIN1 (_____0__25748), .DIN2 (___90___24074), .Q
       (________25653));
  nnd2s1 ___9_9_510400(.DIN1 (____0___24749), .DIN2 (________24720), .Q
       (________27505));
  nor2s1 __90___510401(.DIN1 (________24731), .DIN2 (________24702), .Q
       (________26289));
  nor2s1 __90___510402(.DIN1 (________24797), .DIN2 (________24719), .Q
       (___0____26100));
  nnd2s1 __90___510403(.DIN1 (________24718), .DIN2 (______22154), .Q
       (________25552));
  dffacs1 _______________________________________________510404(.CLRB
       (reset), .CLK (clk), .DIN (________23942), .QN
       (__________________________________________________________________21992));
  nor2s1 __90___510405(.DIN1 (________26576), .DIN2 (________24719), .Q
       (_____0__28032));
  nnd2s1 __90___510406(.DIN1 (________27150), .DIN2 (____99__24745), .Q
       (________25663));
  nnd2s1 ____9__510407(.DIN1 (________24717), .DIN2 (____0___25593), .Q
       (__9_____29981));
  and2s1 ___9___510408(.DIN1 (___0_____40650), .DIN2 (________27043),
       .Q (________25897));
  nor2s1 ____9__510409(.DIN1 (_____0__24706), .DIN2 (___0____24254), .Q
       (_____9__25900));
  hi1s1 ___9__510410(.DIN (_________34576), .Q (_________33170));
  nnd2s1 ____9__510411(.DIN1 (___9_9__24157), .DIN2 (________23989), .Q
       (________25822));
  nnd2s1 ____9__510412(.DIN1 (_____0__24716), .DIN2 (____99__26407), .Q
       (___0____26062));
  nor2s1 __90_09(.DIN1 (_____9__24715), .DIN2 (________24714), .Q
       (___0____26978));
  nor2s1 ___9___510413(.DIN1 (________25607), .DIN2 (_____9__24735), .Q
       (____00__25768));
  nnd2s1 ___9___510414(.DIN1 (____0___23978), .DIN2 (_____9__25348), .Q
       (___0____26106));
  nor2s1 ___9___510415(.DIN1 (___0_9__25144), .DIN2 (_____9___36005),
       .Q (_________35705));
  or2s1 ___9__510416(.DIN1 (____0___23700), .DIN2 (_____0__26528), .Q
       (____0___25770));
  nor2s1 ____9__510417(.DIN1 (________25360), .DIN2 (____9___24743), .Q
       (___0_0___31031));
  nnd2s1 ___9___510418(.DIN1 (____0___23979), .DIN2 (________24771), .Q
       (______9__31765));
  nnd2s1 ___9_510419(.DIN1 (________24707), .DIN2 (________25558), .Q
       (___9____28657));
  nnd2s1 ___9___510420(.DIN1 (___9____24145), .DIN2 (________24760), .Q
       (________28583));
  hi1s1 ___9_510421(.DIN (_____9___37851), .Q (_____9___34189));
  nnd2s1 ____9__510422(.DIN1 (___0____24222), .DIN2 (________24713), .Q
       (________25800));
  nor2s1 ____9__510423(.DIN1 (________25787), .DIN2 (________23995), .Q
       (____9___26317));
  nor2s1 ___90__510424(.DIN1 (_____0__25339), .DIN2 (________24712), .Q
       (__9__0__29946));
  dffacs1 _________________________________________0___0_510425(.CLRB
       (reset), .CLK (clk), .DIN (________23986), .QN
       (_____________________________________0___0___21760));
  nor2s1 ___9___510426(.DIN1 (________23662), .DIN2 (___99___24166), .Q
       (___0____25136));
  nor2s1 __90___510427(.DIN1 (____9___24738), .DIN2 (________24708), .Q
       (___9____27809));
  nor2s1 ___90_510428(.DIN1 (________24711), .DIN2 (________24732), .Q
       (________27355));
  nor2s1 ____9__510429(.DIN1 (________24785), .DIN2 (____9___24927), .Q
       (___0_____31381));
  nor2s1 ___9_510430(.DIN1 (___99), .DIN2 (________24681), .Q
       (_____9__25795));
  nnd2s1 __90_9_510431(.DIN1 (_____9__23951), .DIN2 (________24767), .Q
       (____0____31554));
  nor2s1 __90___510432(.DIN1 (________24797), .DIN2 (____9___24737), .Q
       (________26300));
  nnd2s1 ____510433(.DIN1 (___9_0__24119), .DIN2 (________24710), .Q
       (__9__9__30319));
  nnd2s1 ____9__510434(.DIN1 (___99___24164), .DIN2
       (_____________________21682), .Q (________25734));
  nnd2s1 ___9_0_510435(.DIN1 (________24709), .DIN2 (____99__26407), .Q
       (____9____33353));
  nor2s1 __90__510436(.DIN1 (________24883), .DIN2 (________24708), .Q
       (________28934));
  or2s1 __90_9_510437(.DIN1 (________26576), .DIN2 (________24730), .Q
       (___9____29574));
  nor2s1 __90___510438(.DIN1 (_____________________21736), .DIN2
       (________24821), .Q (____09__27128));
  nnd2s1 __90_0_510439(.DIN1 (___09___24258), .DIN2 (___000__25125), .Q
       (_____90__33327));
  nnd2s1 ____9__510440(.DIN1 (_________38833), .DIN2 (________24912),
       .Q (____009__38047));
  nnd2s1 ___9___510441(.DIN1 (________24707), .DIN2 (________24690), .Q
       (_____9__27996));
  nor2s1 ___90__510442(.DIN1 (_____0__24706), .DIN2 (___09___24260), .Q
       (_________33769));
  nor2s1 ____9__510443(.DIN1 (_____9__24705), .DIN2 (___9____24140), .Q
       (________27040));
  nnd2s1 ___9___510444(.DIN1 (_____0__24885), .DIN2 (________24704), .Q
       (___0_____31084));
  nor2s1 __90_0_510445(.DIN1 (________24703), .DIN2 (____9___23964), .Q
       (____0___25587));
  nor2s1 __90___510446(.DIN1 (________24700), .DIN2 (________24702), .Q
       (___0__0__31061));
  nnd2s1 __90_9_510447(.DIN1 (________24767), .DIN2 (______22154), .Q
       (_____0__27411));
  nnd2s1 ___9___510448(.DIN1 (__9_____30046), .DIN2 (___0____24179), .Q
       (________26826));
  nor2s1 ____9__510449(.DIN1 (________25371), .DIN2 (___0____24221), .Q
       (___0_____30798));
  nor2s1 __90___510450(.DIN1 (________24883), .DIN2 (________24719), .Q
       (__9__0__29916));
  nor2s1 ____9__510451(.DIN1 (___0____25137), .DIN2 (________24900), .Q
       (________29354));
  nor2s1 ___9___510452(.DIN1 (________25735), .DIN2 (________24689), .Q
       (___0_____31324));
  nor2s1 __90___510453(.DIN1 (_____________________21736), .DIN2
       (________24968), .Q (____0___27484));
  nnd2s1 ___9___510454(.DIN1 (________24729), .DIN2 (________24607), .Q
       (____0___27398));
  nor2s1 ___9___510455(.DIN1 (________24658), .DIN2 (________24687), .Q
       (___0_____31268));
  nor2s1 ____99_510456(.DIN1 (_________41345), .DIN2 (________25013),
       .Q (_____9__25785));
  nor2s1 ____9__510457(.DIN1 (________24886), .DIN2 (________24701), .Q
       (________28310));
  nor2s1 ____9__510458(.DIN1 (_________35663), .DIN2 (________24808),
       .Q (________25700));
  nor2s1 __90___510459(.DIN1 (_____9__24715), .DIN2 (________24000), .Q
       (___9____25999));
  hi1s1 ___9___510460(.DIN (_________32712), .Q (________25665));
  nor2s1 __90_0_510461(.DIN1 (________24700), .DIN2 (________24714), .Q
       (____00__27300));
  hi1s1 _______510462(.DIN (____0_0__38084), .Q (_________37202));
  nnd2s1 ___9___510463(.DIN1 (________24709), .DIN2 (________25373), .Q
       (______0__33736));
  nnd2s1 ___90__510464(.DIN1 (________24724), .DIN2 (________24699), .Q
       (____9____33362));
  nor2s1 ___90_510465(.DIN1 (________24698), .DIN2 (___0_0__24188), .Q
       (_________31673));
  nnd2s1 ___9__510466(.DIN1 (___9____24155), .DIN2 (________24697), .Q
       (__9_99__29992));
  nor2s1 ___90__510467(.DIN1 (________23831), .DIN2 (_____0__24696), .Q
       (________27724));
  nor2s1 ___9___510468(.DIN1 (_____9__24695), .DIN2 (________24694), .Q
       (___9____27774));
  hi1s1 __90___510469(.DIN (______0__37872), .Q (_____9__26765));
  nor2s1 __90___510470(.DIN1 (________24693), .DIN2 (________24692), .Q
       (_________33106));
  nor2s1 __90___510471(.DIN1 (________23950), .DIN2 (___00___25126), .Q
       (_________32305));
  and2s1 ___90__510472(.DIN1 (________24426), .DIN2 (________25944), .Q
       (____0____33496));
  nor2s1 ___9___510473(.DIN1 (___0____25186), .DIN2 (________24892), .Q
       (_____9___31789));
  or2s1 ___9__510474(.DIN1 (________24691), .DIN2 (________24016), .Q
       (______0__31921));
  hi1s1 __90_0_510475(.DIN (___9__9__39569), .Q (___9_____39539));
  nor2s1 ___9___510476(.DIN1 (___99___26045), .DIN2 (___0____24205), .Q
       (_________32071));
  nnd2s1 __90___510477(.DIN1 (___9_0__24149), .DIN2 (________24690), .Q
       (________29066));
  nor2s1 ___90__510478(.DIN1 (________26433), .DIN2 (________24952), .Q
       (____0___25772));
  nnd2s1 __90___510479(.DIN1 (___0____24215), .DIN2 (____9___24062), .Q
       (_____9__25613));
  nnd2s1 ___9___510480(.DIN1 (___0_9__24247), .DIN2 (___000__25125), .Q
       (_____0___34487));
  nor2s1 ___90_510481(.DIN1 (________25600), .DIN2 (________24689), .Q
       (_________32311));
  nor2s1 __90___510482(.DIN1 (_____9__24715), .DIN2 (________24702), .Q
       (___9____27820));
  nor2s1 __90___510483(.DIN1 (_____0__24666), .DIN2 (________24688), .Q
       (_____9___32184));
  nor2s1 ___9___510484(.DIN1 (____0___24564), .DIN2 (________24687), .Q
       (___0_____31345));
  hi1s1 __90_9_510485(.DIN (________26545), .Q (_________32613));
  nnd2s1 ___9_0_510486(.DIN1 (_____0__24686), .DIN2 (___9_____39548),
       .Q (_________36955));
  nnd2s1 ___9_510487(.DIN1 (________24028), .DIN2 (________23901), .Q
       (___9_0___39166));
  nor2s1 __90__510488(.DIN1 (____9___24065), .DIN2 (_____9__24685), .Q
       (____0___29283));
  nnd2s1 ___9___510489(.DIN1 (_____0__24022), .DIN2 (____0___23414), .Q
       (_________35435));
  nnd2s1 ___90__510490(.DIN1 (________24684), .DIN2 (________25559), .Q
       (_____90__32080));
  nor2s1 ___90__510491(.DIN1 (___0____23248), .DIN2 (________24038), .Q
       (___9_____39231));
  hi1s1 ___9__510492(.DIN (________24683), .Q (_________38214));
  hi1s1 __90_0_510493(.DIN (___9_90__39245), .Q (____0___25683));
  nor2s1 __90_0_510494(.DIN1 (________23333), .DIN2 (______0__32803),
       .Q (___99____39819));
  hi1s1 ___9_9_510495(.DIN (________24682), .Q (_________35186));
  nor2s1 ___90_510496(.DIN1 (________23661), .DIN2 (________24681), .Q
       (___9_____39667));
  nor2s1 ___90__510497(.DIN1 (________24278), .DIN2 (________24680), .Q
       (_________34644));
  nor2s1 ___9__510498(.DIN1 (____0___24464), .DIN2 (___09___24261), .Q
       (_________38680));
  nor2s1 __90___510499(.DIN1 (________23903), .DIN2 (_____0__23939), .Q
       (______9__37555));
  nor2s1 __90__510500(.DIN1 (________24282), .DIN2 (________25345), .Q
       (________24679));
  and2s1 __90_9_510501(.DIN1 (____90__23683), .DIN2 (________26618), .Q
       (________24678));
  hi1s1 __90_9_510502(.DIN (________24702), .Q (________24677));
  nnd2s1 _______510503(.DIN1 (________24619), .DIN2 (_____9__24675), .Q
       (_____0__24676));
  nor2s1 __9000_510504(.DIN1 (____9___23874), .DIN2 (________24673), .Q
       (________24674));
  nor2s1 _______510505(.DIN1 (____9___24742), .DIN2 (___99___24163), .Q
       (________24672));
  nor2s1 ___99__510506(.DIN1 (_____9___33157), .DIN2 (____9___23780),
       .Q (________24671));
  nnd2s1 ___9___510507(.DIN1 (____0___24462), .DIN2 (________22897), .Q
       (________24670));
  nor2s1 _____0_510508(.DIN1 (____0___22456), .DIN2 (________24668), .Q
       (________24669));
  nor2s1 ___99__510509(.DIN1 (___9_0__24080), .DIN2 (_____0__24666), .Q
       (________24667));
  nor2s1 _______510510(.DIN1 (________23824), .DIN2 (___9_____39746),
       .Q (_____9__24665));
  nnd2s1 _______510511(.DIN1 (________23853), .DIN2 (inData[26]), .Q
       (________24664));
  and2s1 ___990_510512(.DIN1 (___0_90__40168), .DIN2
       (_____________________________________________21970), .Q
       (________24663));
  nor2s1 ___99__510513(.DIN1 (___0____23278), .DIN2 (________24661), .Q
       (________24662));
  or2s1 __90___510514(.DIN1 (________24659), .DIN2 (________24658), .Q
       (________24660));
  or2s1 __90___510515(.DIN1 (________23391), .DIN2 (________24533), .Q
       (________24657));
  nnd2s1 ______510516(.DIN1 (________23803), .DIN2 (inData[16]), .Q
       (_____0__24656));
  nnd2s1 ___99__510517(.DIN1 (____9___23784), .DIN2 (____9___24358), .Q
       (____09__24655));
  nnd2s1 _____0_510518(.DIN1 (_____9__23944), .DIN2 (_____0__24618), .Q
       (____0___24654));
  nnd2s1 ___99__510519(.DIN1 (________24622), .DIN2 (________22881), .Q
       (____0___24653));
  and2s1 ___99__510520(.DIN1 (___0_90__40168), .DIN2
       (_________________________________________0___21939), .Q
       (____0___24652));
  nnd2s1 ___99__510521(.DIN1 (________23849), .DIN2 (_____9__23463), .Q
       (____0___24651));
  nor2s1 ___9___510522(.DIN1 (________23609), .DIN2 (________24673), .Q
       (____0___24650));
  hi1s1 __90___510523(.DIN (____0___24648), .Q (____0___24649));
  and2s1 _______510524(.DIN1 (_____9__23625), .DIN2 (________25640), .Q
       (____0___24647));
  and2s1 __900__510525(.DIN1 (___9____24096), .DIN2 (____9___24642), .Q
       (____00__24646));
  and2s1 ___99__510526(.DIN1 (____9___24644), .DIN2 (____0___24269), .Q
       (____99__24645));
  nnd2s1 ___99__510527(.DIN1 (____9___24642), .DIN2 (_____9__24296), .Q
       (____9___24643));
  or2s1 ___9__510528(.DIN1 (______22129), .DIN2 (____9___24640), .Q
       (____9___24641));
  or2s1 ___99__510529(.DIN1 (_____0__24536), .DIN2 (___9_9__25057), .Q
       (____9___24639));
  nor2s1 ___9___510530(.DIN1 (____9___24637), .DIN2 (_____0__25349), .Q
       (____9___24638));
  nor2s1 __90_0_510531(.DIN1 (_____9__24635), .DIN2 (___0____24233), .Q
       (____90__24636));
  nnd2s1 ___9___510532(.DIN1 (________23904), .DIN2 (________24502), .Q
       (________24634));
  and2s1 _______510533(.DIN1 (____0___23887), .DIN2
       (_________________0___21687), .Q (________24633));
  and2s1 ___99__510534(.DIN1 (________24395), .DIN2 (________24630), .Q
       (________24631));
  nor2s1 ___9__510535(.DIN1
       (____________________________________________21867), .DIN2
       (___9_9__24089), .Q (________24629));
  nor2s1 ___99_510536(.DIN1 (________23650), .DIN2 (________23320), .Q
       (________24628));
  or2s1 ___99__510537(.DIN1 (________23652), .DIN2 (________23863), .Q
       (_____0__24627));
  and2s1 ___99__510538(.DIN1 (________24630), .DIN2 (________24625), .Q
       (________24626));
  nnd2s1 ___99_510539(.DIN1 (________23740), .DIN2 (___90___23139), .Q
       (________24624));
  nnd2s1 ___99_510540(.DIN1 (________24622), .DIN2 (________22907), .Q
       (________24623));
  nor2s1 ___9_9_510541(.DIN1 (_____0__24706), .DIN2 (________24479), .Q
       (________24621));
  and2s1 _____9_510542(.DIN1 (________24619), .DIN2 (_____0__24618), .Q
       (________24620));
  and2s1 ___9___510543(.DIN1 (___0_90__40168), .DIN2
       (__________________________________________9___21951), .Q
       (_____9__24617));
  nor2s1 ___9___510544(.DIN1 (inData[0]), .DIN2 (____9____34315), .Q
       (________24616));
  nnd2s1 ___99__510545(.DIN1 (________24614), .DIN2
       (______________22111), .Q (________24615));
  or2s1 __90___510546(.DIN1 (___00___25132), .DIN2 (________23808), .Q
       (________24613));
  nnd2s1 _____0_510547(.DIN1 (________24614), .DIN2 (___90___23136), .Q
       (________24612));
  nnd2s1 ___99__510548(.DIN1 (___99___25119), .DIN2 (________23731), .Q
       (________24611));
  nnd2s1 _____0_510549(.DIN1 (________24619), .DIN2 (____9___24644), .Q
       (_____0__24610));
  and2s1 ___510550(.DIN1 (________24607), .DIN2 (________23523), .Q
       (________24608));
  nnd2s1 ___9__510551(.DIN1 (_____0___37283), .DIN2 (___9_9__24108), .Q
       (________24606));
  nor2s1 __90__510552(.DIN1 (________24604), .DIN2 (________24481), .Q
       (________24605));
  or2s1 ___99__510553(.DIN1 (________24602), .DIN2 (________23822), .Q
       (________24603));
  nnd2s1 __90_0_510554(.DIN1 (____9___23684), .DIN2
       (____0_________________21725), .Q (_____0__24601));
  nor2s1 ___9___510555(.DIN1 (________24338), .DIN2 (________24599), .Q
       (_____9__24600));
  nor2s1 ___99__510556(.DIN1 (________24597), .DIN2 (________24283), .Q
       (________24598));
  nor2s1 __90___510557(.DIN1 (________24594), .DIN2 (____9___24547), .Q
       (________24595));
  nor2s1 __90___510558(.DIN1 (___0____26089), .DIN2 (_____0__25556), .Q
       (________24593));
  nor2s1 __90___510559(.DIN1 (___0____22296), .DIN2 (________24408), .Q
       (_____0__24592));
  nnd2s1 ______510560(.DIN1 (________23798), .DIN2 (inData[0]), .Q
       (________24591));
  nnd2s1 __90__510561(.DIN1 (_________33843), .DIN2 (_____9___33157),
       .Q (________24590));
  nnd2s1 ___9_9_510562(.DIN1 (____9___25404), .DIN2 (_____9__23861), .Q
       (________24589));
  nor2s1 ___9_510563(.DIN1 (________24055), .DIN2 (________24436), .Q
       (________24588));
  nor2s1 __90___510564(.DIN1 (________24586), .DIN2 (_____9__23673), .Q
       (________24587));
  hi1s1 ___9__510565(.DIN (________24952), .Q (_____0__24585));
  hi1s1 ___9___510566(.DIN (_____9__28081), .Q (_____9__24584));
  nor2s1 __90___510567(.DIN1 (________22783), .DIN2 (_________33843),
       .Q (________24583));
  nnd2s1 ___9___510568(.DIN1 (________24507), .DIN2 (________24581), .Q
       (________24582));
  nnd2s1 ___9___510569(.DIN1 (____9____34315), .DIN2 (___0____22305),
       .Q (________24580));
  nor2s1 __90___510570(.DIN1 (________23120), .DIN2 (_________33843),
       .Q (________24579));
  nnd2s1 ___9___510571(.DIN1 (____0___24460), .DIN2 (_____0__24618), .Q
       (________24578));
  or2s1 __90___510572(.DIN1 (________23115), .DIN2 (_____0__24576), .Q
       (________24577));
  nor2s1 __90___510573(.DIN1 (________24762), .DIN2 (________24389), .Q
       (_____9__24575));
  or2s1 ___9_510574(.DIN1 (___0_____40579), .DIN2 (_________34796), .Q
       (________24574));
  xor2s1 ___9__510575(.DIN1 (____90__23493), .DIN2 (______9__31640), .Q
       (________24573));
  and2s1 __90_9_510576(.DIN1 (____00__24556), .DIN2 (____90__24736), .Q
       (________24572));
  xnr2s1 ___9___510577(.DIN1 (___0_9___40556), .DIN2 (_________38675),
       .Q (________24571));
  nnd2s1 ___9_0_510578(.DIN1 (_____0__23816), .DIN2 (________23079), .Q
       (________24570));
  or2s1 ___9___510579(.DIN1 (________24568), .DIN2 (________24567), .Q
       (________24569));
  nnd2s1 ___9___510580(.DIN1 (________25331), .DIN2 (_____9__22596), .Q
       (_____0__24566));
  or2s1 __90___510581(.DIN1 (____0___24564), .DIN2 (________25345), .Q
       (____09__24565));
  hi1s1 ___9___510582(.DIN (________24903), .Q (____0___24563));
  nnd2s1 ___9__510583(.DIN1 (____09__24467), .DIN2 (________24398), .Q
       (____0___24562));
  nnd2s1 ___9___510584(.DIN1 (____0___23883), .DIN2 (___0____23296), .Q
       (____0___24561));
  hi1s1 __90___510585(.DIN (_____9__24725), .Q (____0___24560));
  nor2s1 __90___510586(.DIN1 (_____9__24705), .DIN2 (_____9__24439), .Q
       (____0___24559));
  hi1s1 __90___510587(.DIN (________24694), .Q (____0___24558));
  nnd2s1 __90___510588(.DIN1 (____00__24556), .DIN2 (________24699), .Q
       (____0___24557));
  nnd2s1 _______510589(.DIN1 (_____0__23530), .DIN2 (________23675), .Q
       (____99__24555));
  nnd2s1 ___9__510590(.DIN1 (________23550), .DIN2 (________23846), .Q
       (____9___24554));
  hi1s1 __90___510591(.DIN (________24707), .Q (____9___24553));
  nnd2s1 __90__510592(.DIN1 (________23632), .DIN2 (________23367), .Q
       (____9___24552));
  nnd2s1 ___9___510593(.DIN1 (________23771), .DIN2 (________25508), .Q
       (____9___24551));
  nor2s1 ___9___510594(.DIN1 (_____9__24486), .DIN2 (________24509), .Q
       (____9___24550));
  nor2s1 __90__510595(.DIN1 (________23637), .DIN2 (________24504), .Q
       (____9___24549));
  nor2s1 ___9___510596(.DIN1 (________23894), .DIN2 (____9___24547), .Q
       (____9___24548));
  nor2s1 __90___510597(.DIN1 (________22756), .DIN2 (_________34796),
       .Q (____90__24546));
  nnd2s1 ___9__510598(.DIN1 (_____9__23710), .DIN2 (________24544), .Q
       (_____9__24545));
  nnd2s1 _______510599(.DIN1 (________23848), .DIN2 (___00___25129), .Q
       (________24543));
  or2s1 _______510600(.DIN1 (________26470), .DIN2 (________23869), .Q
       (________24542));
  nnd2s1 _____9_510601(.DIN1 (________23622), .DIN2 (________22875), .Q
       (________24541));
  nor2s1 _______510602(.DIN1 (________23352), .DIN2 (________23809), .Q
       (________24540));
  nnd2s1 _______510603(.DIN1 (____00__23692), .DIN2
       (_____________________21691), .Q (________24539));
  nnd2s1 _____510604(.DIN1 (________23804), .DIN2 (_________22038), .Q
       (________24538));
  nor2s1 ___9___510605(.DIN1 (________25510), .DIN2 (_____0__24536), .Q
       (________24537));
  or2s1 ___9___510606(.DIN1 (_____________________21688), .DIN2
       (________23936), .Q (_____9__24535));
  nor2s1 ___9___510607(.DIN1 (________24533), .DIN2 (________24329), .Q
       (________24534));
  or2s1 __90_0_510608(.DIN1 (___9____24085), .DIN2 (________24531), .Q
       (________24532));
  hi1s1 __90___510609(.DIN (________24529), .Q (________24530));
  nor2s1 ___9___510610(.DIN1 (_____0__24393), .DIN2 (________24673), .Q
       (________24528));
  nor2s1 ___9___510611(.DIN1 (________23458), .DIN2 (_____9__23825), .Q
       (________24527));
  nor2s1 ___9___510612(.DIN1 (_____9__24525), .DIN2 (________24438), .Q
       (_____0__24526));
  nnd2s1 ___9___510613(.DIN1 (____9___26316), .DIN2 (________24523), .Q
       (________24524));
  nor2s1 ___9___510614(.DIN1 (________22926), .DIN2 (_________34796),
       .Q (________24522));
  and2s1 ___9___510615(.DIN1 (________23854), .DIN2 (_____9___37656),
       .Q (________24521));
  and2s1 ___9___510616(.DIN1 (________24519), .DIN2 (________23570), .Q
       (________24520));
  nor2s1 ___9___510617(.DIN1 (________24517), .DIN2 (________23865), .Q
       (________24518));
  nnd2s1 ___9900(.DIN1 (____9___23781), .DIN2 (___0_9__24217), .Q
       (_____0__24516));
  xor2s1 ___9___510618(.DIN1 (________24514), .DIN2 (_________34647),
       .Q (_____9__24515));
  xor2s1 ___9___510619(.DIN1 (____________), .DIN2 (___0____24235), .Q
       (________24513));
  nnd2s1 ___9___510620(.DIN1 (____9___23686), .DIN2 (________24511), .Q
       (________24512));
  nor2s1 ___9___510621(.DIN1 (________23926), .DIN2 (________24509), .Q
       (________24510));
  nnd2s1 __90___510622(.DIN1 (________24507), .DIN2 (_____0__24506), .Q
       (________24508));
  or2s1 __90___510623(.DIN1 (_____9__23635), .DIN2 (________24504), .Q
       (_____9__24505));
  nnd2s1 ___9___510624(.DIN1 (____9___25404), .DIN2 (________24502), .Q
       (________24503));
  nnd2s1 ___9___510625(.DIN1 (________24500), .DIN2 (____0_), .Q
       (________24501));
  nor2s1 ___9__510626(.DIN1 (___0_____40443), .DIN2 (_____0__24497), .Q
       (________24499));
  nor2s1 ___9___510627(.DIN1 (___0__0__40619), .DIN2 (_____0__24497),
       .Q (________24498));
  nor2s1 ___9___510628(.DIN1 (_________33206), .DIN2 (_________33843),
       .Q (_____9__24496));
  nnd2s1 ___9__510629(.DIN1 (________24500), .DIN2 (________24494), .Q
       (________24495));
  nnd2s1 ___9_510630(.DIN1 (____99__23691), .DIN2 (inData[2]), .Q
       (________24493));
  nor2s1 ___99__510631(.DIN1 (_____0__23711), .DIN2 (___9_9__25114), .Q
       (________24492));
  nnd2s1 ___9_9_510632(.DIN1 (_____9__23727), .DIN2
       (____0________________21717), .Q (________24491));
  nor2s1 _______510633(.DIN1 (____9___25578), .DIN2 (________24473), .Q
       (___9____25091));
  nnd2s1 ____90_510634(.DIN1 (________23647), .DIN2 (________24490), .Q
       (________24907));
  hi1s1 __90___510635(.DIN (________24489), .Q (________25370));
  nnd2s1 __900_9(.DIN1 (________23893), .DIN2 (________24488), .Q
       (________25259));
  nnd2s1 __900__510636(.DIN1 (____99__24457), .DIN2 (_____0__24487), .Q
       (___99___25120));
  hi1s1 ___9___510637(.DIN (_____0__24696), .Q (________25455));
  nnd2s1 __90___510638(.DIN1 (________24472), .DIN2 (________25558), .Q
       (________24888));
  or2s1 __90___510639(.DIN1 (______22154), .DIN2 (________25345), .Q
       (________25350));
  nnd2s1 __90__510640(.DIN1 (_____0__25556), .DIN2 (_____0__23086), .Q
       (_____0__24812));
  nnd2s1 __90___510641(.DIN1 (________23949), .DIN2 (________24507), .Q
       (___0_0__25165));
  nor2s1 __90_9_510642(.DIN1 (_____9__24486), .DIN2 (________24485), .Q
       (___9____25064));
  nnd2s1 __900__510643(.DIN1 (____9___24642), .DIN2 (________24433), .Q
       (_____0__25252));
  nor2s1 __90_0_510644(.DIN1 (________24470), .DIN2 (________24485), .Q
       (___0____25140));
  hi1s1 __90_9_510645(.DIN (________29181), .Q (_____0__26305));
  nor2s1 __900__510646(.DIN1 (________23935), .DIN2 (________24293), .Q
       (___0____25158));
  hi1s1 __90___510647(.DIN (________24484), .Q (________25365));
  hi1s1 __90___510648(.DIN (________24483), .Q (________25283));
  nor2s1 __900__510649(.DIN1 (________24348), .DIN2 (________24471), .Q
       (________25933));
  nor2s1 ___9__510650(.DIN1 (___00___26054), .DIN2 (_____0__23835), .Q
       (________24863));
  nor2s1 ___9__510651(.DIN1 (___9____25983), .DIN2 (________24482), .Q
       (____0___24751));
  nor2s1 __90___510652(.DIN1 (_____________________21682), .DIN2
       (________23679), .Q (___0_0__25175));
  nnd2s1 ___9__510653(.DIN1 (___9_0__24090), .DIN2 (___00___25130), .Q
       (___0____26108));
  nor2s1 __90___510654(.DIN1 (___0____26089), .DIN2 (________24481), .Q
       (________26805));
  nor2s1 __90_9_510655(.DIN1 (____0___24465), .DIN2 (_____9__24695), .Q
       (____9___25766));
  nnd2s1 __90___510656(.DIN1 (_____0__24287), .DIN2 (______22153), .Q
       (____9___24744));
  nor2s1 __900__510657(.DIN1 (_____0__23626), .DIN2 (________24480), .Q
       (_____0__25369));
  nor2s1 __900__510658(.DIN1 (________24300), .DIN2 (________24479), .Q
       (___00___25133));
  nnd2s1 __900__510659(.DIN1 (________24697), .DIN2 (_____0__24478), .Q
       (________24804));
  nor2s1 __90__510660(.DIN1 (_____0__24706), .DIN2 (________23641), .Q
       (________25333));
  hi1s1 __90___510661(.DIN (_____9__24477), .Q (___0____25177));
  nor2s1 __9009_510662(.DIN1 (___900__24070), .DIN2 (________24305), .Q
       (________25351));
  nor2s1 __90_0_510663(.DIN1 (________24476), .DIN2 (________24312), .Q
       (___999__25124));
  nor2s1 __900__510664(.DIN1 (________23651), .DIN2 (________24318), .Q
       (________25813));
  nnd2s1 __90__510665(.DIN1 (________23706), .DIN2
       (_____________________21681), .Q (_____9__24764));
  hi1s1 __90___510666(.DIN (___0_9___31401), .Q (____0___25775));
  hi1s1 __90_99(.DIN (____9_9__37052), .Q (________25526));
  nnd2s1 __90___510667(.DIN1 (________23619), .DIN2 (________24475), .Q
       (________25326));
  nnd2s1 ___9___510668(.DIN1 (_____9__23806), .DIN2 (_____9__25348), .Q
       (_____0__26295));
  nnd2s1 ___9___510669(.DIN1 (_____9__23851), .DIN2 (___0____25176), .Q
       (________25733));
  nnd2s1 __90___510670(.DIN1 (________24474), .DIN2 (________24313), .Q
       (___0____25167));
  nor2s1 ___9___510671(.DIN1 (________23820), .DIN2 (________24908), .Q
       (________26657));
  dffacs1 ________________________________________________510672(.CLRB
       (reset), .CLK (clk), .DIN (________23621), .Q
       (______________________________________________21956));
  nor2s1 ___9___510673(.DIN1 (________24604), .DIN2 (________24473), .Q
       (___0_____31088));
  hi1s1 __90_0_510674(.DIN (_____9___36005), .Q (_____9__25537));
  nnd2s1 __90___510675(.DIN1 (________23743), .DIN2 (________24475), .Q
       (________25330));
  nnd2s1 ____9_510676(.DIN1 (________24303), .DIN2 (________25373), .Q
       (____0_9__33489));
  nor2s1 ____9_510677(.DIN1 (_____0__24706), .DIN2 (________23630), .Q
       (_____9__26294));
  hi1s1 ___9___510678(.DIN (__9_____30046), .Q (____9___25402));
  nnd2s1 __90__510679(.DIN1 (________24469), .DIN2 (____0___23697), .Q
       (____0___25411));
  nnd2s1 ___90__510680(.DIN1 (________23707), .DIN2 (_____9__23900), .Q
       (____0_0__38084));
  nnd2s1 ___90__510681(.DIN1 (_____0__24468), .DIN2 (________23921), .Q
       (_____9__28100));
  nnd2s1 __90___510682(.DIN1 (________24472), .DIN2 (____9___23500), .Q
       (________27598));
  nor2s1 ___9__510683(.DIN1 (________23870), .DIN2 (________24908), .Q
       (________27181));
  hi1s1 __9____510684(.DIN (________24730), .Q (___0____25160));
  nnd2s1 __90___510685(.DIN1 (________24290), .DIN2 (____0___24466), .Q
       (_____9__27646));
  nor2s1 __90__510686(.DIN1 (________23813), .DIN2 (______9__33955), .Q
       (______0__34259));
  nor2s1 __90___510687(.DIN1 (________24471), .DIN2 (________24886), .Q
       (_____0___31994));
  nor2s1 __90___510688(.DIN1 (________24470), .DIN2 (________24504), .Q
       (___00___25128));
  nor2s1 __90_9_510689(.DIN1 (________24330), .DIN2 (_____0__23646), .Q
       (__909___29720));
  nnd2s1 __90___510690(.DIN1 (________24469), .DIN2
       (_____________________21679), .Q (________25377));
  nnd2s1 __90___510691(.DIN1 (____0___23791), .DIN2
       (_____________________21682), .Q (________25325));
  hi1s1 ___9___510692(.DIN (_________38833), .Q (____9____34341));
  nor2s1 __90__510693(.DIN1 (____0___23042), .DIN2 (________23644), .Q
       (___0_9__25184));
  nor2s1 __90___510694(.DIN1 (________26576), .DIN2 (________24321), .Q
       (______0__31903));
  nnd2s1 __90_0_510695(.DIN1 (________23722), .DIN2 (_____0__23728), .Q
       (________25513));
  and2s1 ___90__510696(.DIN1 (_____0__24468), .DIN2 (____09__24467), .Q
       (__9_____30400));
  nor2s1 ___9___510697(.DIN1 (________23814), .DIN2 (________24908), .Q
       (_________32056));
  nnd2s1 ___90__510698(.DIN1 (_____0__24468), .DIN2 (___0____24219), .Q
       (________29112));
  nor2s1 __90___510699(.DIN1 (____0___24369), .DIN2 (_____9__24447), .Q
       (____9___27389));
  hi1s1 __90_9_510700(.DIN (___0_9__27017), .Q (___0_____30695));
  nnd2s1 __90___510701(.DIN1 (________24310), .DIN2 (____0___24466), .Q
       (___9_0__27795));
  nnd2s1 __90___510702(.DIN1 (_____0__24297), .DIN2 (___0____25159), .Q
       (___0_____30958));
  and2s1 ___90__510703(.DIN1 (___0____24253), .DIN2 (________25944), .Q
       (____9____34365));
  nnd2s1 __90___510704(.DIN1 (___0_9__24197), .DIN2 (____99__23787), .Q
       (___9__9__39569));
  hi1s1 __90___510705(.DIN (____9____38001), .Q (____9____37998));
  nor2s1 __90___510706(.DIN1 (___0____25168), .DIN2 (____0___24465), .Q
       (___0_____31274));
  nor2s1 __90__510707(.DIN1 (____0___24464), .DIN2 (________23659), .Q
       (______9__35584));
  nor2s1 __90_9_510708(.DIN1 (________24475), .DIN2 (________23627), .Q
       (___0____25179));
  nnd2s1 ___90__510709(.DIN1 (_____0__24468), .DIN2 (________23752), .Q
       (________28230));
  hi1s1 __90__510710(.DIN (_____0___38616), .Q (______0__38711));
  nnd2s1 ___9___510711(.DIN1 (________23620), .DIN2 (____0___23041), .Q
       (_____9___37851));
  hi1s1 __90_510712(.DIN (________25004), .Q (_____0___35834));
  nnd2s1 __90___510713(.DIN1 (_________38385), .DIN2 (________23827),
       .Q (_________38573));
  nnd2s1 ___909_510714(.DIN1 (_____0__23768), .DIN2 (___9____24087), .Q
       (_________37230));
  nor2s1 ___9___510715(.DIN1 (____0___24463), .DIN2 (________23829), .Q
       (_________35968));
  nnd2s1 __90___510716(.DIN1 (____0___24462), .DIN2 (________24517), .Q
       (_________38200));
  or2s1 ___9_0_510717(.DIN1 (______0__35694), .DIN2 (_____9___35559),
       .Q (_________35448));
  nnd2s1 __90__510718(.DIN1 (____0___24460), .DIN2 (________26258), .Q
       (____0___24461));
  or2s1 ___99__510719(.DIN1 (____0_0__38093), .DIN2 (_____9__23777), .Q
       (____0___24459));
  nnd2s1 ___99__510720(.DIN1 (____99__24457), .DIN2 (________23734), .Q
       (____00__24458));
  nnd2s1 ___99__510721(.DIN1 (____9___23877), .DIN2 (____9___24455), .Q
       (____9___24456));
  nnd2s1 ___999_510722(.DIN1 (________23823), .DIN2 (________23475), .Q
       (____9___24454));
  nnd2s1 ___999_510723(.DIN1 (________23895), .DIN2 (____9___24452), .Q
       (____9___24453));
  nor2s1 ___999_510724(.DIN1 (________23628), .DIN2 (___9_9__23208), .Q
       (____9___24451));
  nnd2s1 ___999_510725(.DIN1 (________23561), .DIN2 (____9___24449), .Q
       (____9___24450));
  nor2s1 ___510726(.DIN1 (________23847), .DIN2 (_____9__24447), .Q
       (____90__24448));
  nnd2s1 __9000_510727(.DIN1 (________25920), .DIN2 (____0___23790), .Q
       (________24446));
  or2s1 __9000_510728(.DIN1 (___9_0__29602), .DIN2 (____0___23885), .Q
       (________24445));
  and2s1 __900__510729(.DIN1 (________24902), .DIN2 (________23466), .Q
       (________24444));
  nnd2s1 __900_510730(.DIN1 (_____0__23843), .DIN2 (________22925), .Q
       (________24443));
  nnd2s1 __900_510731(.DIN1 (____9____34315), .DIN2
       (_____________________________________9_______21884), .Q
       (________24442));
  nor2s1 __900__510732(.DIN1 (________23634), .DIN2 (_____0__23702), .Q
       (________24441));
  nor2s1 __900__510733(.DIN1 (_____9__24439), .DIN2 (________24438), .Q
       (_____0__24440));
  nnd2s1 __900__510734(.DIN1 (________24436), .DIN2 (________23733), .Q
       (________24437));
  nnd2s1 __900_510735(.DIN1 (____9___24644), .DIN2 (________25364), .Q
       (________24435));
  nnd2s1 __900__510736(.DIN1 (________24327), .DIN2 (________24433), .Q
       (________24434));
  nnd2s1 ___9_9_510737(.DIN1 (___99____39861), .DIN2 (________24431),
       .Q (________24432));
  hi1s1 ___9___510738(.DIN (_____9__24429), .Q (_____0__24430));
  xor2s1 __90___510739(.DIN1 (___0__0__40511), .DIN2 (___9_____39372),
       .Q (________24428));
  hi1s1 ___9___510740(.DIN (________24426), .Q (________24427));
  nor2s1 ___990_510741(.DIN1 (_____9__24382), .DIN2 (________24509), .Q
       (________24425));
  nor2s1 __90_9_510742(.DIN1 (________24786), .DIN2 (________24698), .Q
       (________24424));
  nnd2s1 ___99__510743(.DIN1 (_____0__23807), .DIN2 (________23355), .Q
       (________24423));
  nor2s1 __90___510744(.DIN1 (________23016), .DIN2 (________24533), .Q
       (________24422));
  nor2s1 ___9___510745(.DIN1 (_____0__24420), .DIN2 (_____9__24392), .Q
       (________24421));
  nor2s1 ___9___510746(.DIN1 (________24418), .DIN2 (____9___23875), .Q
       (_____9__24419));
  nor2s1 __90__510747(.DIN1 (________24415), .DIN2 (________23830), .Q
       (________24416));
  nor2s1 ___99__510748(.DIN1 (________23730), .DIN2 (________23512), .Q
       (________24414));
  nor2s1 ___99__510749(.DIN1 (________24886), .DIN2 (________24658), .Q
       (________24413));
  or2s1 __9000_510750(.DIN1 (________23732), .DIN2 (_____0__24411), .Q
       (________24412));
  nnd2s1 __90___510751(.DIN1 (________23769), .DIN2 (________23653), .Q
       (_____9__24410));
  nor2s1 ___990_510752(.DIN1 (___0__0__40599), .DIN2 (________24408),
       .Q (________24409));
  nnd2s1 ___9___510753(.DIN1 (________23859), .DIN2 (inData[26]), .Q
       (________24407));
  nor2s1 _______510754(.DIN1 (____0________________21714), .DIN2
       (____0___23886), .Q (________24406));
  nnd2s1 ___9__510755(.DIN1 (____9___26316), .DIN2 (________23810), .Q
       (________24405));
  nor2s1 ___99__510756(.DIN1 (________24323), .DIN2 (________24599), .Q
       (________24404));
  nnd2s1 ___9__510757(.DIN1 (_____0__23666), .DIN2 (____9___24361), .Q
       (________24403));
  nnd2s1 ___9___510758(.DIN1 (________24500), .DIN2 (________23815), .Q
       (________24402));
  hi1s1 __90_9_510759(.DIN (________24892), .Q (_____0__24401));
  nor2s1 __90___510760(.DIN1 (________22902), .DIN2 (____0___23698), .Q
       (_____9__24400));
  nnd2s1 __90___510761(.DIN1 (________24474), .DIN2 (________24398), .Q
       (________24399));
  and2s1 __90___510762(.DIN1 (____0___26594), .DIN2 (________25345), .Q
       (________24397));
  nnd2s1 __90___510763(.DIN1 (________24395), .DIN2 (________25375), .Q
       (________24396));
  or2s1 ___99__510764(.DIN1 (_____0__24393), .DIN2 (_____9__24392), .Q
       (________24394));
  and2s1 __90__510765(.DIN1 (________24314), .DIN2 (________23911), .Q
       (________24391));
  nor2s1 __90___510766(.DIN1 (________24389), .DIN2 (___0____25206), .Q
       (________24390));
  nnd2s1 __90___510767(.DIN1 (___0____23282), .DIN2 (________23680), .Q
       (________24388));
  nnd2s1 __90___510768(.DIN1 (________24386), .DIN2 (________24704), .Q
       (________24387));
  nor2s1 __90___510769(.DIN1 (________23477), .DIN2 (________24384), .Q
       (________24385));
  or2s1 __90___510770(.DIN1 (_____9__24382), .DIN2 (________24504), .Q
       (_____0__24383));
  nor2s1 __90___510771(.DIN1 (_____9__25632), .DIN2 (_____9__23655), .Q
       (________24381));
  or2s1 __90___510772(.DIN1 (____0___26594), .DIN2 (_____0__25556), .Q
       (________24380));
  nnd2s1 __90__510773(.DIN1 (________24292), .DIN2 (________22952), .Q
       (________24379));
  nnd2s1 __90___510774(.DIN1 (________24301), .DIN2 (___0____25169), .Q
       (________24378));
  nnd2s1 __90___510775(.DIN1 (________25920), .DIN2 (________24351), .Q
       (________24377));
  or2s1 __90___510776(.DIN1 (____9___24928), .DIN2 (________23948), .Q
       (________24376));
  nnd2s1 __90__510777(.DIN1 (________23663), .DIN2 (________23754), .Q
       (________24375));
  nnd2s1 __90_9_510778(.DIN1 (____9___25404), .DIN2 (___0_0__23291), .Q
       (________24374));
  nnd2s1 ___9__510779(.DIN1 (________23657), .DIN2 (inData[4]), .Q
       (_____0__24373));
  or2s1 __90_0_510780(.DIN1 (________24791), .DIN2 (____9___24547), .Q
       (____09__24372));
  nor2s1 __90_0_510781(.DIN1 (________23545), .DIN2 (________23723), .Q
       (____0___24371));
  nor2s1 __90___510782(.DIN1 (____0___24369), .DIN2 (_____9__24695), .Q
       (____0___24370));
  nor2s1 __90__510783(.DIN1 (____9___24068), .DIN2 (____0___25412), .Q
       (____0___24368));
  or2s1 __90___510784(.DIN1 (________24594), .DIN2 (________24533), .Q
       (____0___24367));
  or2s1 __90___510785(.DIN1 (___0____25163), .DIN2 (_____0__23674), .Q
       (____0___24366));
  or2s1 __90___510786(.DIN1 (________25345), .DIN2 (________24311), .Q
       (____0___24365));
  or2s1 __90___510787(.DIN1 (____0___24564), .DIN2 (________24886), .Q
       (____00__24364));
  nnd2s1 __90___510788(.DIN1 (____9___25404), .DIN2 (_____0__24775), .Q
       (____99__24363));
  nnd2s1 __90___510789(.DIN1 (____9___24361), .DIN2 (____9___24360), .Q
       (____9___24362));
  and2s1 __90_9_510790(.DIN1 (________23896), .DIN2 (____9___24358), .Q
       (____9___24359));
  or2s1 __90_0_510791(.DIN1 (________24319), .DIN2 (________24504), .Q
       (____9___24357));
  nnd2s1 __90_0_510792(.DIN1 (________25558), .DIN2 (________24607), .Q
       (____9___24356));
  nor2s1 __90_0_510793(.DIN1 (___9____25983), .DIN2 (________24481), .Q
       (____90__24355));
  or2s1 __90___510794(.DIN1 (___9____25983), .DIN2 (________24353), .Q
       (_____9__24354));
  and2s1 __90___510795(.DIN1 (____0___24460), .DIN2 (________24351), .Q
       (________24352));
  nnd2s1 __90___510796(.DIN1 (___0____24220), .DIN2 (____09__24467), .Q
       (________24350));
  nor2s1 __90___510797(.DIN1 (____9___23034), .DIN2 (________24348), .Q
       (________24349));
  nnd2s1 __90__510798(.DIN1 (____0___23793), .DIN2 (___0____23242), .Q
       (________24347));
  nor2s1 __90___510799(.DIN1 (________24476), .DIN2 (____0___24369), .Q
       (________24346));
  nor2s1 __90___510800(.DIN1 (________23096), .DIN2 (________24384), .Q
       (_____0__24345));
  nor2s1 ___99__510801(.DIN1 (________23365), .DIN2 (________23818), .Q
       (_____9__24344));
  nor2s1 ___9___510802(.DIN1 (________22825), .DIN2 (________23708), .Q
       (________24343));
  and2s1 ___9___510803(.DIN1 (________23856), .DIN2 (________24341), .Q
       (________24342));
  nor2s1 __9__9_(.DIN1 (_____9__22858), .DIN2 (________24295), .Q
       (________24340));
  or2s1 __90___510804(.DIN1 (________24338), .DIN2 (___00___25126), .Q
       (________24339));
  nor2s1 ___9___510805(.DIN1 (_________36883), .DIN2 (________24436),
       .Q (________24337));
  hi1s1 __90__510806(.DIN (_____9__24335), .Q (_____0__24336));
  nor2s1 __90___510807(.DIN1 (________24659), .DIN2 (___0____26109), .Q
       (________24334));
  xor2s1 ___9___510808(.DIN1
       (__________________________________________________________________21988),
       .DIN2 (_________34647), .Q (________24333));
  xor2s1 ___9___510809(.DIN1 (________23514), .DIN2
       (_____________22097), .Q (________24332));
  nnd2s1 ___9_9_510810(.DIN1 (___99____39861), .DIN2 (___0_____40616),
       .Q (________24331));
  nor2s1 __90___510811(.DIN1 (___0____25168), .DIN2 (________24330), .Q
       (________25737));
  nnd2s1 ___9_0_510812(.DIN1 (_____9___35467), .DIN2 (________23799),
       .Q (________24682));
  or2s1 __90___510813(.DIN1 (___00___25132), .DIN2 (________24698), .Q
       (___0____25180));
  nor2s1 __900__510814(.DIN1 (_____9__24525), .DIN2 (________24329), .Q
       (________25344));
  nor2s1 __90___510815(.DIN1 (___9____25060), .DIN2 (________24329), .Q
       (___0____25182));
  nnd2s1 __90_0_510816(.DIN1 (______0__37673), .DIN2 (________23712),
       .Q (________24683));
  nnd2s1 __90_510817(.DIN1 (________24328), .DIN2 (________24327), .Q
       (________25466));
  nor2s1 __90_0_510818(.DIN1 (________25257), .DIN2 (_____9__24954), .Q
       (____9___25405));
  nor2s1 __90__510819(.DIN1 (________24017), .DIN2 (_____0__24326), .Q
       (___99___25117));
  nor2s1 __900_510820(.DIN1 (________24348), .DIN2 (________24658), .Q
       (___0____25166));
  nor2s1 __900__510821(.DIN1 (_____9__24325), .DIN2 (________23735), .Q
       (________25353));
  nor2s1 __90099(.DIN1 (________24324), .DIN2 (________23897), .Q
       (________24816));
  nor2s1 __900_510822(.DIN1 (________24323), .DIN2 (___00___25126), .Q
       (________25367));
  dffacs1 _______________________________________________510823(.CLRB
       (reset), .CLK (clk), .DIN (________23720), .Q
       (_____________________________________________21925));
  nor2s1 __90___510824(.DIN1 (________24322), .DIN2 (________24321), .Q
       (___0____25153));
  nor2s1 __90___510825(.DIN1 (____0___26594), .DIN2 (________24481), .Q
       (________24801));
  or2s1 __90_510826(.DIN1 (____0___26594), .DIN2 (________24320), .Q
       (________25563));
  nor2s1 __90_0_510827(.DIN1 (________24319), .DIN2 (________24485), .Q
       (___90___25032));
  nnd2s1 __90_0_510828(.DIN1 (________25920), .DIN2 (____9___24061), .Q
       (_____9__24857));
  nor2s1 __90_0_510829(.DIN1 (________23811), .DIN2 (________24318), .Q
       (___0____25183));
  nnd2s1 __90_0_510830(.DIN1 (________24294), .DIN2 (_____9__25348), .Q
       (________24823));
  nor2s1 __90___510831(.DIN1 (________24604), .DIN2 (________24320), .Q
       (____9___24740));
  nnd2s1 __900_510832(.DIN1 (____0___23889), .DIN2 (___00___25131), .Q
       (________25346));
  nor2s1 __90__510833(.DIN1 (_____0__24706), .DIN2 (________23649), .Q
       (________24759));
  nor2s1 __90___510834(.DIN1 (________24308), .DIN2 (___0____26089), .Q
       (___99___25121));
  hi1s1 ___9___510835(.DIN (________24317), .Q (____0___25409));
  or2s1 __90_510836(.DIN1 (_____0__24316), .DIN2 (________24531), .Q
       (___09___25219));
  nnd2s1 __90___510837(.DIN1 (_____9__23938), .DIN2 (_____0__24876), .Q
       (________26260));
  nor2s1 __90___510838(.DIN1 (________26426), .DIN2 (________24698), .Q
       (____0___24754));
  hi1s1 __9____510839(.DIN (_____9__24685), .Q (___0____25199));
  hi1s1 __9____510840(.DIN (_____9__24315), .Q (___0____25173));
  nnd2s1 __90___510841(.DIN1 (________24314), .DIN2 (________24768), .Q
       (____0___24753));
  nor2s1 __900_510842(.DIN1 (_____0__23919), .DIN2 (________24309), .Q
       (___9____25053));
  nnd2s1 __90___510843(.DIN1 (________24607), .DIN2 (________24313), .Q
       (________24758));
  nor2s1 __90090(.DIN1 (___9____23196), .DIN2 (________24312), .Q
       (___00___25127));
  nor2s1 __9009_510844(.DIN1 (____0___23312), .DIN2 (________24614), .Q
       (________25322));
  nor2s1 __90__510845(.DIN1 (____0_______________), .DIN2
       (_____9__23645), .Q (________25267));
  nor2s1 __90_0_510846(.DIN1 (________24311), .DIN2 (____9___24830), .Q
       (________24982));
  nnd2s1 __90___510847(.DIN1 (________24310), .DIN2 (_____0__23339), .Q
       (____0___24752));
  nor2s1 __9009_510848(.DIN1 (___909__24079), .DIN2 (________24309), .Q
       (________24814));
  nor2s1 __90___510849(.DIN1 (_____9__23586), .DIN2 (________24976), .Q
       (____0___25415));
  nor2s1 __90_0_510850(.DIN1 (_____0__24326), .DIN2 (________24309), .Q
       (____09__24848));
  nor2s1 __90_0_510851(.DIN1 (___0____26109), .DIN2 (________24481), .Q
       (________24897));
  nor2s1 __90___510852(.DIN1 (________24308), .DIN2 (________24353), .Q
       (________24773));
  or2s1 __90_0_510853(.DIN1 (________23705), .DIN2 (________24757), .Q
       (___0____25147));
  hi1s1 __90_0_510854(.DIN (________24714), .Q (___0____25149));
  nor2s1 __900__510855(.DIN1 (________23759), .DIN2 (________23704), .Q
       (____9___25308));
  or2s1 __90___510856(.DIN1 (_____0__24307), .DIN2 (_____9__24306), .Q
       (____0___25771));
  nor2s1 __90___510857(.DIN1 (________24693), .DIN2 (________24305), .Q
       (________26739));
  nnd2s1 __90__510858(.DIN1 (____99__24457), .DIN2 (________24304), .Q
       (_____0__25329));
  and2s1 ____510859(.DIN1 (________24303), .DIN2 (________25944), .Q
       (________25746));
  hi1s1 __90_0_510860(.DIN (_________35806), .Q (__9_____29971));
  nor2s1 __90___510861(.DIN1 (____0___26590), .DIN2 (________23639), .Q
       (________25366));
  hi1s1 __90___510862(.DIN (________27150), .Q (________25745));
  hi1s1 __90___510863(.DIN (_____9___37654), .Q (_________34907));
  nor2s1 __90___510864(.DIN1 (________24901), .DIN2 (____0___24465), .Q
       (___090__25213));
  nor2s1 __90___510865(.DIN1 (____9___23689), .DIN2 (________24722), .Q
       (_____0__26599));
  nnd2s1 __90__510866(.DIN1 (____09__24467), .DIN2 (___90___24073), .Q
       (________25334));
  nnd2s1 __90___510867(.DIN1 (________23668), .DIN2 (___00___25129), .Q
       (____9___25763));
  nnd2s1 __90_9_510868(.DIN1 (____90__25758), .DIN2 (________24302), .Q
       (_____0__25271));
  nor2s1 __90__510869(.DIN1 (_____________________21736), .DIN2
       (___0____26089), .Q (_____0__25461));
  and2s1 __90__510870(.DIN1 (________24301), .DIN2 (___0____25156), .Q
       (________26760));
  nor2s1 __90___510871(.DIN1 (________24922), .DIN2 (________24330), .Q
       (____9___26680));
  nnd2s1 ___9___510872(.DIN1 (________24722), .DIN2 (____9___23785), .Q
       (___9____25975));
  nor2s1 __90__510873(.DIN1 (________24300), .DIN2 (_____0__23636), .Q
       (________25363));
  nor2s1 __90___510874(.DIN1 (________25371), .DIN2 (___00___25126), .Q
       (________25323));
  nnd2s1 __90___510875(.DIN1 (_____0__24506), .DIN2 (________24313), .Q
       (___0____25142));
  hi1s1 __90__510876(.DIN (________24299), .Q (________25539));
  nor2s1 __90__510877(.DIN1 (________23946), .DIN2 (_____9__24447), .Q
       (___0____26115));
  hi1s1 __9____510878(.DIN (________24778), .Q (___0____25162));
  hi1s1 __9____510879(.DIN (____9___24737), .Q (___0____25138));
  nor2s1 __90___510880(.DIN1 (________24298), .DIN2 (___99____39861),
       .Q (_________32956));
  or2s1 __90___510881(.DIN1 (________26576), .DIN2 (________23671), .Q
       (________24879));
  nnd2s1 __90___510882(.DIN1 (____9____34315), .DIN2 (________22481),
       .Q (___9_____39283));
  or2s1 __90___510883(.DIN1 (______________________21698), .DIN2
       (________23841), .Q (________25285));
  nnd2s1 __90_9_510884(.DIN1 (_____0__24297), .DIN2 (___0_9__25164), .Q
       (________25340));
  and2s1 __90___510885(.DIN1 (________24327), .DIN2 (_____9__24296), .Q
       (____9___25306));
  nnd2s1 ____9__510886(.DIN1 (________23868), .DIN2
       (_____________________21682), .Q (___0____25208));
  nor2s1 __9____510887(.DIN1 (________24700), .DIN2 (________24295), .Q
       (___0____25190));
  nnd2s1 __90__510888(.DIN1 (________24294), .DIN2 (___99___25123), .Q
       (____9___26862));
  nor2s1 __90___510889(.DIN1 (________24504), .DIN2 (________24293), .Q
       (___9____27790));
  nnd2s1 __90___510890(.DIN1 (________24875), .DIN2 (____9___24449), .Q
       (____90__25300));
  nnd2s1 __90_510891(.DIN1 (________23819), .DIN2
       (_____________________21679), .Q (___0____25178));
  nnd2s1 __90___510892(.DIN1 (________24292), .DIN2 (___0_____40616),
       .Q (____00__25407));
  nnd2s1 __90___510893(.DIN1 (________24301), .DIN2 (________24291), .Q
       (________26755));
  xor2s1 __90__510894(.DIN1 (_____0___34938), .DIN2 (________22537), .Q
       (________26545));
  or2s1 ___510895(.DIN1 (___0____26109), .DIN2 (________24473), .Q
       (___0__0__30787));
  nor2s1 __90___510896(.DIN1 (________24727), .DIN2 (________23638), .Q
       (___0____28779));
  nnd2s1 __90_0_510897(.DIN1 (____09__23796), .DIN2 (___0____25176), .Q
       (_________33172));
  nnd2s1 __90___510898(.DIN1 (_____9__24031), .DIN2 (____0___24466), .Q
       (________27313));
  nnd2s1 __90___510899(.DIN1 (_____0__24297), .DIN2 (___0____25171), .Q
       (________28519));
  nnd2s1 __90_0_510900(.DIN1 (________24290), .DIN2 (___0____25171), .Q
       (____9___29190));
  nnd2s1 __90_9_510901(.DIN1 (___9____24086), .DIN2 (___9____24083), .Q
       (_________34576));
  nor2s1 __90_510902(.DIN1 (________24289), .DIN2 (_____9__24286), .Q
       (___9____27771));
  hi1s1 __9____510903(.DIN (________24288), .Q (___0____25170));
  nnd2s1 __90___510904(.DIN1 (________24581), .DIN2 (________24313), .Q
       (________25347));
  hi1s1 __9____510905(.DIN (_____9__24793), .Q (___9____25974));
  nor2s1 __90_0_510906(.DIN1 (___9_0__25068), .DIN2 (________24389), .Q
       (________25523));
  nnd2s1 __90___510907(.DIN1 (_____0__24287), .DIN2
       (_____________________21682), .Q (_____9__25338));
  nor2s1 __90___510908(.DIN1 (________24922), .DIN2 (_____9__24286), .Q
       (________28318));
  nnd2s1 __90___510909(.DIN1 (________24472), .DIN2 (________24690), .Q
       (____9___29463));
  nor2s1 __90__510910(.DIN1 (____99__25585), .DIN2 (________24305), .Q
       (____0____33465));
  or2s1 __90_9_510911(.DIN1 (_____________________21679), .DIN2
       (________23725), .Q (___0_0__25185));
  nor2s1 __90___510912(.DIN1 (______22153), .DIN2 (________23633), .Q
       (_____9__25358));
  nnd2s1 ___90_510913(.DIN1 (________24303), .DIN2 (___000__25125), .Q
       (_________34154));
  or2s1 __90___510914(.DIN1 (________25376), .DIN2 (________24305), .Q
       (_____0___33721));
  nor2s1 __90_510915(.DIN1 (________24285), .DIN2 (________23716), .Q
       (________29249));
  hi1s1 __9____510916(.DIN (________24284), .Q (___0_0__25203));
  nnd2s1 __90___510917(.DIN1 (________24301), .DIN2 (________25332), .Q
       (________29208));
  nnd2s1 __90_9_510918(.DIN1 (_____0__23738), .DIN2 (________25355), .Q
       (_________33016));
  nor2s1 __90___510919(.DIN1 (________24727), .DIN2 (___090__24257), .Q
       (_________31958));
  nor2s1 __90___510920(.DIN1 (________24883), .DIN2 (________23631), .Q
       (___09_9__31465));
  nor2s1 __90_510921(.DIN1 (________23062), .DIN2 (________24283), .Q
       (___9_____39784));
  nor2s1 __90___510922(.DIN1 (________24282), .DIN2 (________24886), .Q
       (________28860));
  nnd2s1 __90__510923(.DIN1 (___9_____39384), .DIN2 (______0__38256),
       .Q (_________36480));
  hi1s1 __9____510924(.DIN (________24281), .Q (________25574));
  nor2s1 __90__510925(.DIN1 (________24720), .DIN2 (________23833), .Q
       (_________38372));
  nnd2s1 __90___510926(.DIN1 (________23857), .DIN2 (______0__37673),
       .Q (_____9___36360));
  nor2s1 __90___510927(.DIN1 (________22824), .DIN2 (________23713), .Q
       (___9__9__39125));
  nnd2s1 __90___510928(.DIN1 (________23855), .DIN2 (________22765), .Q
       (_________38871));
  nor2s1 __90___510929(.DIN1 (________23370), .DIN2 (________23681), .Q
       (_____9___36721));
  nor2s1 __90___510930(.DIN1 (_____9__23453), .DIN2 (________23729), .Q
       (___9_90__39245));
  nor2s1 __90_0_510931(.DIN1 (________23721), .DIN2 (________24279), .Q
       (_________32712));
  nor2s1 __90___510932(.DIN1 (____9___23036), .DIN2 (________23858), .Q
       (___9_0___39619));
  nor2s1 __90__510933(.DIN1 (________24278), .DIN2 (_____0__24277), .Q
       (______0__37872));
  nnd2s1 __90___510934(.DIN1 (_____0__24277), .DIN2 (________23678), .Q
       (____0_9__38073));
  nnd2s1 ___9__510935(.DIN1 (________23471), .DIN2 (________24475), .Q
       (____09__24276));
  nor2s1 __900__510936(.DIN1 (____9___23878), .DIN2 (____9___23499), .Q
       (____0___24275));
  nor2s1 __900__510937(.DIN1 (___09___23307), .DIN2 (________23741), .Q
       (____0___24274));
  nor2s1 ___99__510938(.DIN1 (________26530), .DIN2 (________23344), .Q
       (____0___24273));
  nnd2s1 ___9___510939(.DIN1 (___9____24120), .DIN2 (________24433), .Q
       (____0___24272));
  nor2s1 __900__510940(.DIN1 (_____0__22781), .DIN2 (________23551), .Q
       (____0___24271));
  and2s1 __900__510941(.DIN1 (_____9__24675), .DIN2 (____0___24269), .Q
       (____0___24270));
  nor2s1 __900__510942(.DIN1 (____00__24267), .DIN2 (________25440), .Q
       (____0___24268));
  nor2s1 __900__510943(.DIN1 (________23534), .DIN2 (___09___24265), .Q
       (___099__24266));
  nnd2s1 ___99_510944(.DIN1 (___09___24263), .DIN2 (____0___23789), .Q
       (___09___24264));
  nnd2s1 __90___510945(.DIN1 (_________38262), .DIN2 (_________37320),
       .Q (___09___24262));
  nnd2s1 __900_510946(.DIN1 (___0____24189), .DIN2 (________25726), .Q
       (___09___24261));
  nnd2s1 __900__510947(.DIN1 (___9____24117), .DIN2 (____0___23603), .Q
       (___09___24260));
  nnd2s1 __900__510948(.DIN1 (___09___24263), .DIN2 (___00___24176), .Q
       (___09___24259));
  hi1s1 __9____510949(.DIN (___090__24257), .Q (___09___24258));
  nnd2s1 __900__510950(.DIN1 (____9___23398), .DIN2 (________23342), .Q
       (___0_9__24256));
  nor2s1 __900__510951(.DIN1 (___9_9__25047), .DIN2 (___9____24111), .Q
       (___0____24255));
  hi1s1 ___9___510952(.DIN (___0____24253), .Q (___0____24254));
  nnd2s1 __900_510953(.DIN1 (___0____24251), .DIN2 (___0____24250), .Q
       (___0____24252));
  nnd2s1 __9000_510954(.DIN1 (___9____24136), .DIN2 (_____9__25469), .Q
       (___0____24249));
  nor2s1 ___99__510955(.DIN1 (_____9__24382), .DIN2 (___90___24077), .Q
       (___0_9__24247));
  nor2s1 ___999_510956(.DIN1 (____0__22215), .DIN2 (___0____24251), .Q
       (___0____24246));
  nnd2s1 ___999_510957(.DIN1 (________23562), .DIN2
       (_________________9___21749), .Q (___0____24245));
  nor2s1 ___510958(.DIN1 (_____________________21691), .DIN2
       (_____0__23483), .Q (___0____24244));
  and2s1 ___99__510959(.DIN1 (___9____24131), .DIN2 (______22159), .Q
       (___0____24243));
  nor2s1 ___99__510960(.DIN1 (____00__24267), .DIN2 (________23750), .Q
       (___0____24242));
  nor2s1 ___9___510961(.DIN1 (________23007), .DIN2 (________24058), .Q
       (___0____24241));
  or2s1 ___99__510962(.DIN1 (___99___24159), .DIN2 (___0____24239), .Q
       (___0____24240));
  nnd2s1 ___99__510963(.DIN1 (________23902), .DIN2 (________23050), .Q
       (___0_0__24238));
  nor2s1 ___99_510964(.DIN1 (________24711), .DIN2 (________25336), .Q
       (___0_9__24237));
  nor2s1 ___99__510965(.DIN1 (___0____22336), .DIN2 (___0____24235), .Q
       (___0____24236));
  hi1s1 __90___510966(.DIN (___0____24233), .Q (___0____24234));
  nor2s1 ___99__510967(.DIN1 (_____9__23338), .DIN2 (_____9__23567), .Q
       (___0____24232));
  or2s1 ___99__510968(.DIN1 (___0____24230), .DIN2 (________25257), .Q
       (___0____24231));
  nnd2s1 ___99__510969(.DIN1 (________23487), .DIN2 (_____9__22988), .Q
       (___0____24229));
  nnd2s1 ___9___510970(.DIN1 (________23378), .DIN2
       (_____________________21691), .Q (___0_0__24228));
  nor2s1 ___99_510971(.DIN1 (_____________________21669), .DIN2
       (________23484), .Q (___0_9__24227));
  nor2s1 ___99_510972(.DIN1 (_____0__22597), .DIN2 (________23489), .Q
       (___0____24226));
  or2s1 ___99__510973(.DIN1 (___0____24224), .DIN2 (____0___25590), .Q
       (___0____24225));
  nnd2s1 __90___510974(.DIN1 (________23536), .DIN2 (________23364), .Q
       (___0____24223));
  nor2s1 ___99_510975(.DIN1 (________22517), .DIN2 (________24026), .Q
       (___0____24222));
  nnd2s1 ___9___510976(.DIN1 (___0____24220), .DIN2 (___0____24219), .Q
       (___0____24221));
  nnd2s1 __9____510977(.DIN1 (____9___24067), .DIN2 (___0_9__24217), .Q
       (___0_0__24218));
  nnd2s1 __90__510978(.DIN1 (___0_9__23290), .DIN2 (___0____23277), .Q
       (___0____24216));
  hi1s1 __90_9_510979(.DIN (_____0__24277), .Q (___0____24215));
  nnd2s1 ___99__510980(.DIN1 (________23543), .DIN2 (inData[18]), .Q
       (___0____24214));
  nor2s1 ___9___510981(.DIN1 (________22779), .DIN2 (___09___23308), .Q
       (___0____24213));
  nor2s1 ___99__510982(.DIN1 (________23459), .DIN2 (_____0__23548), .Q
       (___0____24212));
  nnd2s1 __90___510983(.DIN1 (______9__33955), .DIN2
       (______________22067), .Q (___0____24211));
  nnd2s1 ___99__510984(.DIN1 (________23925), .DIN2 (___9_9__25977), .Q
       (___0____24210));
  and2s1 ___9___510985(.DIN1 (____0___23980), .DIN2 (________23089), .Q
       (___0____24209));
  nnd2s1 __90___510986(.DIN1 (____9___23403), .DIN2 (___0____23279), .Q
       (___0_0__24208));
  nnd2s1 ___99__510987(.DIN1 (___0____24206), .DIN2 (________23345), .Q
       (___0_9__24207));
  nnd2s1 __90___510988(.DIN1 (____00__23788), .DIN2 (____0___23315), .Q
       (___0____24205));
  nor2s1 ___9___510989(.DIN1 (____9___22739), .DIN2 (________23585), .Q
       (___0____24204));
  nor2s1 ___99__510990(.DIN1 (inData[24]), .DIN2 (___9_____39183), .Q
       (___0____24203));
  nnd2s1 ___99__510991(.DIN1 (___0____24201), .DIN2
       (_____________________________________0______21755), .Q
       (___0____24202));
  nor2s1 ___9___510992(.DIN1 (________23424), .DIN2 (___9____24146), .Q
       (___0____24200));
  and2s1 _______510993(.DIN1 (_____9___37656), .DIN2 (________23395),
       .Q (___0____24199));
  nnd2s1 ___99__510994(.DIN1 (___0_9__24197), .DIN2 (_____0__22949), .Q
       (___0_0__24198));
  or2s1 ___9_9_510995(.DIN1
       (______________________________________0______21886), .DIN2
       (___0____24195), .Q (___0____24196));
  nnd2s1 ___99_510996(.DIN1 (___9____24127), .DIN2 (___90__22262), .Q
       (___0____24194));
  nnd2s1 ___99_510997(.DIN1 (_____0__23521), .DIN2 (___9____24084), .Q
       (___0____24193));
  or2s1 ___9_9_510998(.DIN1
       (______________________________________0_______21894), .DIN2
       (___0____24191), .Q (___0____24192));
  nor2s1 ___99__510999(.DIN1 (_____9__23842), .DIN2 (___0____24189), .Q
       (___0____24190));
  or2s1 ___9___511000(.DIN1 (___0_9__24187), .DIN2 (___0____25204), .Q
       (___0_0__24188));
  nnd2s1 ___9__511001(.DIN1 (___0____23285), .DIN2 (inData[2]), .Q
       (___0____24186));
  nnd2s1 ___99__511002(.DIN1 (____99__24745), .DIN2 (________24488), .Q
       (___0____24185));
  nnd2s1 ___9___511003(.DIN1 (________23468), .DIN2 (________26259), .Q
       (___0____24184));
  or2s1 ___990_511004(.DIN1 (________24431), .DIN2 (___0____24191), .Q
       (___0____24183));
  or2s1 ___990_511005(.DIN1 (________25337), .DIN2 (____90__23397), .Q
       (___0____24182));
  nnd2s1 ___9___511006(.DIN1 (_____9__24296), .DIN2 (________23428), .Q
       (___0____24181));
  or2s1 __90___511007(.DIN1 (________23054), .DIN2 (___0____24179), .Q
       (___0____24180));
  nnd2s1 __9____511008(.DIN1 (___009__24177), .DIN2 (___00___24176), .Q
       (___0_0__24178));
  nor2s1 ___9__511009(.DIN1 (_____0__23436), .DIN2 (_____0__24012), .Q
       (___00___24175));
  nnd2s1 ___9___511010(.DIN1 (___09___24265), .DIN2 (______22145), .Q
       (___00___24174));
  nor2s1 ___9_9_511011(.DIN1 (_____0__22899), .DIN2 (________23332), .Q
       (___00___24173));
  or2s1 ___9___511012(.DIN1 (___9____25102), .DIN2 (_____0__23540), .Q
       (___00___24172));
  or2s1 ___9___511013(.DIN1 (__99_9__30508), .DIN2 (____09__23318), .Q
       (___00___24171));
  nnd2s1 __90___511014(.DIN1 (___00___24169), .DIN2 (____09), .Q
       (___00___24170));
  nnd2s1 ___9_511015(.DIN1 (________24433), .DIN2 (_____9__23435), .Q
       (___000__24168));
  nnd2s1 ___9___511016(.DIN1 (________23323), .DIN2 (___0____22321), .Q
       (___999__24167));
  or2s1 __90___511017(.DIN1 (___99___24165), .DIN2 (________23390), .Q
       (___99___24166));
  hi1s1 ___9___511018(.DIN (___99___24163), .Q (___99___24164));
  nnd2s1 __90___511019(.DIN1 (___9____24102), .DIN2 (___0____22348), .Q
       (___99___24162));
  nor2s1 ___9___511020(.DIN1 (___9_9__23191), .DIN2 (_____0__23578), .Q
       (___99___24161));
  nor2s1 __90___511021(.DIN1 (___99___24159), .DIN2 (___990__24158), .Q
       (___99___24160));
  nor2s1 __90__511022(.DIN1 (________24517), .DIN2 (___9____24156), .Q
       (___9_9__24157));
  nor2s1 ___9___511023(.DIN1 (________25510), .DIN2 (_____9__23991), .Q
       (___9____24155));
  nnd2s1 __90_511024(.DIN1 (________23462), .DIN2 (_____0__24876), .Q
       (___9____24154));
  nor2s1 ___9___511025(.DIN1 (___9____23180), .DIN2 (________23569), .Q
       (___9____24153));
  nnd2s1 __90___511026(.DIN1 (____99__24745), .DIN2 (____0___26146), .Q
       (___9____24152));
  nor2s1 __90_511027(.DIN1 (___0____26080), .DIN2 (________23392), .Q
       (___9____24151));
  hi1s1 __9____511028(.DIN (________24481), .Q (___9____24150));
  hi1s1 __9____511029(.DIN (_____9__24286), .Q (___9_0__24149));
  and2s1 __90__511030(.DIN1 (_____9___35467), .DIN2 (_________36556),
       .Q (___9_9__24148));
  nor2s1 __90___511031(.DIN1 (___9____24146), .DIN2 (_____9__25728), .Q
       (___9____24147));
  and2s1 __90__511032(.DIN1 (___9____24144), .DIN2 (_____0__24895), .Q
       (___9____24145));
  nor2s1 __90__511033(.DIN1 (________24604), .DIN2 (_____0__23982), .Q
       (___9____24143));
  nnd2s1 __90___511034(.DIN1 (___00___24169), .DIN2 (___009__23224), .Q
       (___9____24142));
  nor2s1 ___9___511035(.DIN1 (____0___22652), .DIN2 (________23354), .Q
       (___9____24141));
  nnd2s1 ___9__511036(.DIN1 (____90__23587), .DIN2 (___9_0__24139), .Q
       (___9____24140));
  nor2s1 ___9___511037(.DIN1 (________23532), .DIN2 (____0___23310), .Q
       (___9_9__24138));
  nnd2s1 __90___511038(.DIN1 (________25749), .DIN2 (___9____24136), .Q
       (___9____24137));
  and2s1 __90___511039(.DIN1 (_____0__24726), .DIN2 (___9____24134), .Q
       (___9____24135));
  nnd2s1 __90___511040(.DIN1 (___9____24136), .DIN2 (________25829), .Q
       (___9____24133));
  nnd2s1 ___9___511041(.DIN1 (___9____24131), .DIN2 (___0____22350), .Q
       (___9____24132));
  nnd2s1 ___9__511042(.DIN1 (_____0__23558), .DIN2 (________22906), .Q
       (___9____24130));
  nnd2s1 __90___511043(.DIN1 (________24034), .DIN2 (________25343), .Q
       (___9_0__24129));
  nnd2s1 ___9___511044(.DIN1 (___9____24127), .DIN2 (____90__23124), .Q
       (___9_9__24128));
  nnd2s1 ___9___511045(.DIN1 (___9____24095), .DIN2 (________25825), .Q
       (___9____24126));
  nnd2s1 __90_9_511046(.DIN1 (_____9__23928), .DIN2 (________23746), .Q
       (___9____24125));
  nnd2s1 ___9___511047(.DIN1 (________23703), .DIN2 (___9____24123), .Q
       (___9____24124));
  nnd2s1 __90_511048(.DIN1 (_____0__25479), .DIN2 (___9____24136), .Q
       (___9____24122));
  and2s1 __90___511049(.DIN1 (___9____24120), .DIN2 (_____9__24296), .Q
       (___9____24121));
  nor2s1 __900__511050(.DIN1 (___90___24078), .DIN2 (____0___24840), .Q
       (___9_0__24119));
  and2s1 __90_9_511051(.DIN1 (___9____24117), .DIN2 (____90__24736), .Q
       (___9_9__24118));
  nnd2s1 __90___511052(.DIN1 (____9___23966), .DIN2 (____9___24452), .Q
       (___9____24116));
  or2s1 __90___511053(.DIN1 (________24338), .DIN2 (____9___23968), .Q
       (___9____24115));
  or2s1 ___9_0_511054(.DIN1 (_____00__34847), .DIN2 (________23537), .Q
       (___9____24114));
  nor2s1 ___9___511055(.DIN1 (___9____24112), .DIN2 (___9____24111), .Q
       (___9____24113));
  or2s1 ___9___511056(.DIN1
       (_____________________________________________21897), .DIN2
       (___0____24179), .Q (___9____24110));
  or2s1 ___9__511057(.DIN1 (_____________________21746), .DIN2
       (___9_9__24108), .Q (___9_0__24109));
  and2s1 ___9_511058(.DIN1 (_____0__25566), .DIN2
       (_____________________21688), .Q (___9____24107));
  nor2s1 __90___511059(.DIN1 (____9__22246), .DIN2 (___9_____39183), .Q
       (___9____24106));
  nnd2s1 ___9_9_511060(.DIN1 (________23584), .DIN2 (inData[30]), .Q
       (___9____24105));
  nor2s1 __90___511061(.DIN1 (________24338), .DIN2 (________25336), .Q
       (___9____24104));
  nnd2s1 ___9_9_511062(.DIN1 (___9____24102), .DIN2 (________23122), .Q
       (___9____24103));
  nnd2s1 ___9___511063(.DIN1 (________23763), .DIN2
       (__________________________________________9___21951), .Q
       (___9____24101));
  nnd2s1 __90___511064(.DIN1 (____9___23595), .DIN2 (___90___24072), .Q
       (___9_0__24100));
  nnd2s1 __90___511065(.DIN1 (________23321), .DIN2 (_________33686),
       .Q (___9_9__24099));
  nnd2s1 __90__511066(.DIN1 (_____0__25479), .DIN2 (_____0__24775), .Q
       (___9____24098));
  and2s1 __90__511067(.DIN1 (___9____24096), .DIN2 (___9____24095), .Q
       (___9____24097));
  nnd2s1 __90__511068(.DIN1 (___9____24117), .DIN2 (____9___23588), .Q
       (___9____24094));
  nnd2s1 ___9___511069(.DIN1 (________23479), .DIN2 (________24475), .Q
       (___9____24093));
  nnd2s1 ___9___511070(.DIN1 (________23337), .DIN2 (inData[26]), .Q
       (___9____24092));
  nor2s1 ___9___511071(.DIN1 (________24567), .DIN2 (________24713), .Q
       (___9____24091));
  hi1s1 __90___511072(.DIN (___9_0__24090), .Q (________24687));
  hi1s1 __9___9(.DIN (___9_9__24089), .Q (________24817));
  nor2s1 __90_0_511073(.DIN1 (___9____24088), .DIN2 (________23343), .Q
       (______0__35745));
  nor2s1 __90_0_511074(.DIN1 (____99__23596), .DIN2 (___9____24087), .Q
       (________24681));
  hi1s1 __9____511075(.DIN (___9____24086), .Q (________24688));
  nor2s1 __900__511076(.DIN1 (________23923), .DIN2 (___990__24158), .Q
       (_____9__24429));
  or2s1 __900__511077(.DIN1 (___9____24085), .DIN2 (___0____24230), .Q
       (________24906));
  nnd2s1 __90_0_511078(.DIN1 (________23346), .DIN2 (___9____24084), .Q
       (________24680));
  nor2s1 __9009_511079(.DIN1 (____9___23876), .DIN2 (____9___23401), .Q
       (________24878));
  and2s1 __900__511080(.DIN1 (________23761), .DIN2 (________24723), .Q
       (________24890));
  hi1s1 __90__511081(.DIN (________24886), .Q (____9___24833));
  nor2s1 __90_9_511082(.DIN1 (________25376), .DIN2 (____99__24069), .Q
       (________24893));
  nor2s1 __9009_511083(.DIN1 (________23382), .DIN2 (_____0__23049), .Q
       (___9____25108));
  nor2s1 __9____511084(.DIN1 (________22697), .DIN2 (____9___24928), .Q
       (________24284));
  hi1s1 __9___511085(.DIN (________24853), .Q (________24769));
  nnd2s1 __9_0__(.DIN1 (____9___23590), .DIN2 (___9____24083), .Q
       (________24692));
  nnd2s1 __90_9_511086(.DIN1 (___9____24082), .DIN2 (________22821), .Q
       (________24989));
  nor2s1 __90___511087(.DIN1 (___9____24081), .DIN2 (____0___23795), .Q
       (_____9__24894));
  nor2s1 __90___511088(.DIN1 (___9_0__24080), .DIN2 (___909__24079), .Q
       (_____0__24755));
  nor2s1 __90_511089(.DIN1 (_____9__25632), .DIN2 (___0____25204), .Q
       (________24529));
  nnd2s1 __90_0_511090(.DIN1 (___90___24076), .DIN2 (_____9__23909), .Q
       (________24689));
  nor2s1 __90_511091(.DIN1 (___90___24078), .DIN2 (________24567), .Q
       (________24889));
  nor2s1 __90___511092(.DIN1 (________24319), .DIN2 (___90___24077), .Q
       (________24426));
  nor2s1 __90___511093(.DIN1 (____90__24060), .DIN2 (___9____24082), .Q
       (____99__24934));
  nnd2s1 __90___511094(.DIN1 (________24328), .DIN2 (___9____24095), .Q
       (________24483));
  nor2s1 __900__511095(.DIN1 (____00__22939), .DIN2 (________23389), .Q
       (____9___24739));
  nnd2s1 __900__511096(.DIN1 (___90___24075), .DIN2 (___90___24076), .Q
       (________24712));
  nor2s1 __90___511097(.DIN1 (________23340), .DIN2 (________25371), .Q
       (___9____25981));
  nnd2s1 __90___511098(.DIN1 (____9___23687), .DIN2 (________26272), .Q
       (____9___24927));
  nnd2s1 __90___511099(.DIN1 (___9____24117), .DIN2 (________23640), .Q
       (_____9__24725));
  or2s1 __9____511100(.DIN1 (____09__26331), .DIN2 (____9___24928), .Q
       (________24785));
  dffacs1 ________________________________________________511101(.CLRB
       (reset), .CLK (clk), .DIN (___0____23288), .Q
       (______________________________________________21958));
  nnd2s1 __90___511102(.DIN1 (___90___24075), .DIN2 (_____0__23910), .Q
       (____9___24743));
  nnd2s1 __90___511103(.DIN1 (___90___24074), .DIN2 (________23460), .Q
       (____0___24939));
  nnd2s1 __90__511104(.DIN1 (___0____24219), .DIN2 (___90___24073), .Q
       (________24900));
  dffacs1 _________________________________________0_____511105(.CLRB
       (reset), .CLK (clk), .DIN (____9___23402), .Q (___0_0___40569));
  or2s1 __90___511106(.DIN1 (___0_____40582), .DIN2 (___9_____39183),
       .Q (________25394));
  and2s1 __90___511107(.DIN1 (___0____24220), .DIN2 (_____9__25348), .Q
       (________24729));
  nor2s1 __90___511108(.DIN1 (______9__36337), .DIN2 (____0___23505),
       .Q (____0___24749));
  nnd2s1 __90___511109(.DIN1 (___09___24263), .DIN2 (___90___24072), .Q
       (________25018));
  nor2s1 __90___511110(.DIN1 (____0___23311), .DIN2 (________23934), .Q
       (________24880));
  or2s1 __90___511111(.DIN1 (___90___24071), .DIN2 (________23572), .Q
       (___0_9___31214));
  nor2s1 __90__511112(.DIN1 (___900__24070), .DIN2 (____99__24069), .Q
       (_________33553));
  or2s1 __90___511113(.DIN1 (________24797), .DIN2 (____9___24064), .Q
       (__9__0__30206));
  nor2s1 __90__511114(.DIN1 (____9___24068), .DIN2 (________23916), .Q
       (________24903));
  nnd2s1 __9____511115(.DIN1 (____9___23963), .DIN2 (________25380), .Q
       (________24702));
  nnd2s1 __9___0(.DIN1 (____9___24067), .DIN2 (____9___24066), .Q
       (________24821));
  nor2s1 __90___511116(.DIN1 (____9___24065), .DIN2 (____9___24064), .Q
       (___0_0___30746));
  nnd2s1 __9____511117(.DIN1 (________23999), .DIN2 (____9___24063), .Q
       (________24730));
  nnd2s1 __90_9_511118(.DIN1 (________23525), .DIN2 (_____9__25348), .Q
       (____0___26690));
  nnd2s1 __90__511119(.DIN1 (________23670), .DIN2 (____0___24466), .Q
       (________29181));
  nor2s1 __90__511120(.DIN1 (________24476), .DIN2 (____9___23498), .Q
       (_____9__28081));
  nor2s1 __90___511121(.DIN1 (________23457), .DIN2 (___90___25034), .Q
       (________25004));
  nor2s1 __90_9_511122(.DIN1 (________23554), .DIN2 (________23516), .Q
       (______0__34855));
  nnd2s1 __90_0_511123(.DIN1 (________23491), .DIN2 (____9___24062), .Q
       (_________38833));
  hi1s1 __90___511124(.DIN (________26604), .Q (________26611));
  nor2s1 __90___511125(.DIN1 (____9___24061), .DIN2 (________23564), .Q
       (___0_____40323));
  or2s1 __90___511126(.DIN1 (____9___24061), .DIN2 (____0___23313), .Q
       (___99_9__39836));
  nor2s1 __9__9_511127(.DIN1 (____90__24060), .DIN2 (_____9__24059), .Q
       (________27150));
  nor2s1 __90___511128(.DIN1 (________24710), .DIN2 (________24058), .Q
       (_____9___36005));
  and2s1 __90___511129(.DIN1 (________23486), .DIN2 (________24280), .Q
       (___9_____39332));
  nnd2s1 __90___511130(.DIN1 (___0____23294), .DIN2 (_____9__23425), .Q
       (__9_____30046));
  nor2s1 __90___511131(.DIN1 (____0___23412), .DIN2 (____9____38898),
       .Q (____9____38001));
  hi1s1 __9____511132(.DIN (________23899), .Q (___0__0__39993));
  and2s1 _______511133(.DIN1 (_____9___37656), .DIN2 (________23375),
       .Q (________24057));
  nnd2s1 ___99__511134(.DIN1 (________24044), .DIN2 (________24055), .Q
       (________24056));
  nnd2s1 __900__511135(.DIN1 (________27288), .DIN2 (_____0__23473), .Q
       (________24054));
  nnd2s1 ___99__511136(.DIN1 (________24003), .DIN2 (___9___22192), .Q
       (________24053));
  nnd2s1 ___99__511137(.DIN1 (___0_0__23273), .DIN2 (________23326), .Q
       (________24052));
  nnd2s1 __900__511138(.DIN1 (____9___23685), .DIN2 (_____9__23871), .Q
       (_____9__24051));
  nnd2s1 ___9___511139(.DIN1 (________24049), .DIN2 (_____0__23349), .Q
       (________24050));
  nnd2s1 ___99_511140(.DIN1 (________23565), .DIN2 (inData[18]), .Q
       (________24048));
  nnd2s1 __9__99(.DIN1 (________24046), .DIN2 (________23669), .Q
       (________24047));
  and2s1 ___99__511141(.DIN1 (________24044), .DIN2 (_________36883),
       .Q (________24045));
  nnd2s1 ___99__511142(.DIN1 (____9___27649), .DIN2 (________23080), .Q
       (________24043));
  nor2s1 __90___511143(.DIN1 (________22893), .DIN2 (___9_____39183),
       .Q (_____0__24042));
  nor2s1 __900__511144(.DIN1 (________22995), .DIN2 (____0___23408), .Q
       (_____9__24041));
  or2s1 __9000_511145(.DIN1 (________23913), .DIN2 (____9___23405), .Q
       (________24040));
  nor2s1 __9000_511146(.DIN1 (___99____39814), .DIN2 (_____9__23358),
       .Q (________24039));
  nnd2s1 __900_511147(.DIN1 (________24037), .DIN2 (___0____23274), .Q
       (________24038));
  nnd2s1 ___9___511148(.DIN1 (________23381), .DIN2 (clk), .Q
       (________24036));
  nnd2s1 __90___511149(.DIN1 (________24034), .DIN2 (________24033), .Q
       (________24035));
  hi1s1 __90___511150(.DIN (_____9__24031), .Q (_____0__24032));
  nor2s1 __900__511151(.DIN1 (________22951), .DIN2 (________23366), .Q
       (________24030));
  nor2s1 ___9__511152(.DIN1 (inData[29]), .DIN2 (____9____38898), .Q
       (________24029));
  nor2s1 __90__511153(.DIN1 (________22921), .DIN2 (________23361), .Q
       (________24028));
  nor2s1 ___9___511154(.DIN1 (________22966), .DIN2 (________24026), .Q
       (________24027));
  nnd2s1 __90___511155(.DIN1 (________23560), .DIN2 (____0___26146), .Q
       (________24025));
  nor2s1 __90___511156(.DIN1 (____0___22841), .DIN2 (_____9__23577), .Q
       (________24024));
  or2s1 __90___511157(.DIN1 (_________35587), .DIN2 (____9____38898),
       .Q (________24023));
  nor2s1 __90___511158(.DIN1 (___0____23251), .DIN2 (________23488), .Q
       (_____0__24022));
  nnd2s1 __90___511159(.DIN1 (________23334), .DIN2 (inData[22]), .Q
       (_____9__24021));
  nnd2s1 __90___511160(.DIN1 (________23385), .DIN2 (___09___22354), .Q
       (________24020));
  nor2s1 __90___511161(.DIN1 (____0___24466), .DIN2 (___09___23303), .Q
       (________24019));
  nor2s1 __90__511162(.DIN1 (________24017), .DIN2 (___909__24079), .Q
       (________24018));
  or2s1 __90___511163(.DIN1 (___90___24071), .DIN2 (________25324), .Q
       (________24016));
  nnd2s1 __90___511164(.DIN1 (___9_9__24108), .DIN2 (____9___22830), .Q
       (________24015));
  or2s1 __90_9_511165(.DIN1 (________24013), .DIN2 (_____0__24012), .Q
       (________24014));
  or2s1 __90_511166(.DIN1 (________24010), .DIN2 (___0____25168), .Q
       (_____9__24011));
  or2s1 ___9_0_511167(.DIN1 (____0____________0_), .DIN2
       (___0_9__23300), .Q (________24009));
  nor2s1 __90___511168(.DIN1 (___09____40687), .DIN2 (___9_____39746),
       .Q (________24008));
  nnd2s1 __90___511169(.DIN1 (________24034), .DIN2 (_____0__23617), .Q
       (________24007));
  nor2s1 __90___511170(.DIN1 (____0________________21720), .DIN2
       (________23960), .Q (________24006));
  nor2s1 __90__511171(.DIN1 (___9____24146), .DIN2 (____9___25955), .Q
       (________24005));
  nnd2s1 __90___511172(.DIN1 (________24003), .DIN2 (________22370), .Q
       (________24004));
  and2s1 __90___511173(.DIN1 (___9____24144), .DIN2 (________24720), .Q
       (_____0__24002));
  and2s1 __90___511174(.DIN1 (___0____24201), .DIN2 (________22991), .Q
       (_____9__24001));
  nnd2s1 __9____511175(.DIN1 (________23999), .DIN2 (________23998), .Q
       (________24000));
  and2s1 __90___511176(.DIN1 (________24034), .DIN2 (________24993), .Q
       (________23997));
  nor2s1 __90___511177(.DIN1 (________23573), .DIN2 (_____9__23328), .Q
       (________23996));
  nor2s1 __90___511178(.DIN1 (________24282), .DIN2 (___90___24078), .Q
       (________23995));
  nnd2s1 __90___511179(.DIN1 (______9__35170), .DIN2 (___0__0__40413),
       .Q (________23994));
  or2s1 __90_511180(.DIN1 (___9____24156), .DIN2 (_____0__24420), .Q
       (________23993));
  or2s1 __90_9_511181(.DIN1 (________25440), .DIN2 (_____9__23991), .Q
       (_____0__23992));
  and2s1 __90_9_511182(.DIN1 (____9___26316), .DIN2 (________23989), .Q
       (________23990));
  and2s1 __90_9_511183(.DIN1 (___9____24096), .DIN2 (___9____24120), .Q
       (________23988));
  nnd2s1 __90_9_511184(.DIN1 (___0____23293), .DIN2 (____9___24062), .Q
       (________23987));
  and2s1 __90_511185(.DIN1 (_________38262), .DIN2 (_________37412), .Q
       (________23986));
  nor2s1 __90_0_511186(.DIN1 (________23984), .DIN2 (________24604), .Q
       (________23985));
  nor2s1 __90_0_511187(.DIN1 (____9___25578), .DIN2 (_____0__23982), .Q
       (________23983));
  and2s1 __90__511188(.DIN1 (____0___23980), .DIN2 (________23629), .Q
       (____09__23981));
  and2s1 __90___511189(.DIN1 (___0____23287), .DIN2 (________24993), .Q
       (____0___23979));
  nor2s1 __90__511190(.DIN1 (____0___23977), .DIN2 (________25336), .Q
       (____0___23978));
  nnd2s1 __90___511191(.DIN1 (________24328), .DIN2 (___9____24120), .Q
       (____0___23976));
  nnd2s1 __90___511192(.DIN1 (___0____23286), .DIN2 (________23580), .Q
       (____0___23975));
  nor2s1 ___9_511193(.DIN1 (inData[8]), .DIN2 (___9_____39183), .Q
       (____0___23974));
  nnd2s1 __900__511194(.DIN1 (________23465), .DIN2 (inData[16]), .Q
       (____0___23973));
  nnd2s1 ___99__511195(.DIN1 (_____9__24675), .DIN2 (________23765), .Q
       (____00__23972));
  or2s1 __9__0_(.DIN1 (____9___23970), .DIN2 (_____9__24059), .Q
       (____99__23971));
  nor2s1 __900_511196(.DIN1 (________24323), .DIN2 (____9___23968), .Q
       (____9___23969));
  nnd2s1 __90009(.DIN1 (_____0__23607), .DIN2 (____9___23966), .Q
       (____9___23967));
  or2s1 __9____511197(.DIN1 (___0____25156), .DIN2 (___0____25169), .Q
       (____9___23965));
  nnd2s1 __9____511198(.DIN1 (____9___23963), .DIN2 (____90__23962), .Q
       (____9___23964));
  nnd2s1 ___9___511199(.DIN1 (________23960), .DIN2 (________23959), .Q
       (_____9__23961));
  nor2s1 __9___511200(.DIN1 (________23760), .DIN2 (____9___24067), .Q
       (________23958));
  hi1s1 __9____511201(.DIN (________24698), .Q (________23957));
  hi1s1 __9___511202(.DIN (________24290), .Q (________23956));
  hi1s1 __9____511203(.DIN (_____9__24439), .Q (________23955));
  and2s1 ___9__511204(.DIN1 (________23762), .DIN2 (________23953), .Q
       (________23954));
  hi1s1 __9____511205(.DIN (_____9__23951), .Q (_____0__23952));
  hi1s1 __9____511206(.DIN (________23949), .Q (________23950));
  nnd2s1 ___9___511207(.DIN1 (___0____23237), .DIN2 (________23574), .Q
       (________23947));
  nor2s1 __9_0__511208(.DIN1 (____9___23495), .DIN2 (________24824), .Q
       (________23945));
  and2s1 __90___511209(.DIN1 (________25362), .DIN2
       (____0________________21664), .Q (________23943));
  nnd2s1 __90___511210(.DIN1 (___9_9), .DIN2
       (_____________________________________________21908), .Q
       (________23942));
  or2s1 __90___511211(.DIN1 (____0________________21663), .DIN2
       (________25572), .Q (________23941));
  nor2s1 ___99__511212(.DIN1 (____9___23970), .DIN2 (________23579), .Q
       (________23940));
  hi1s1 __90___511213(.DIN (_____9__23938), .Q (_____0__23939));
  hi1s1 __90___511214(.DIN (________23936), .Q (________23937));
  nnd2s1 __900_511215(.DIN1 (________23559), .DIN2 (________23930), .Q
       (________24881));
  nor2s1 __900__511216(.DIN1 (_____9__24486), .DIN2 (________23935), .Q
       (_____0__24716));
  nor2s1 __90___511217(.DIN1 (____0_________________21724), .DIN2
       (___9____24082), .Q (________24860));
  nor2s1 __900__511218(.DIN1 (____9___23589), .DIN2 (________25572), .Q
       (________26198));
  nor2s1 __900__511219(.DIN1 (________22685), .DIN2 (________23934), .Q
       (_____0__24686));
  nor2s1 __90__511220(.DIN1 (________24324), .DIN2 (_____0__24420), .Q
       (________24299));
  and2s1 __900__511221(.DIN1 (________23931), .DIN2 (________23933), .Q
       (____9___24741));
  hi1s1 __90_511222(.DIN (________24353), .Q (________24783));
  and2s1 __900__511223(.DIN1 (________23350), .DIN2 (________23932), .Q
       (____9___25581));
  nor2s1 __900__511224(.DIN1 (________24323), .DIN2 (________25336), .Q
       (________24887));
  nnd2s1 __900__511225(.DIN1 (_____0__23464), .DIN2 (____0___22944), .Q
       (________24609));
  and2s1 __9009_511226(.DIN1 (________23931), .DIN2 (________24690), .Q
       (________24721));
  hi1s1 __90___511227(.DIN (___0____26109), .Q (________24718));
  nor2s1 __90___511228(.DIN1 (___0_____40616), .DIN2 (___0____24191),
       .Q (________24317));
  nor2s1 __900__511229(.DIN1 (____0___24840), .DIN2 (________24713), .Q
       (________24684));
  dffacs1 ________________________________________________511230(.CLRB
       (reset), .CLK (clk), .DIN (____9___23399), .Q
       (______________________________________________21957));
  or2s1 __90_9_511231(.DIN1 (___99___24159), .DIN2 (________25391), .Q
       (____0___24750));
  nor2s1 __90__511232(.DIN1 (________23455), .DIN2 (________24713), .Q
       (_____9__24335));
  nor2s1 __90___511233(.DIN1 (________26433), .DIN2 (________23526), .Q
       (_____9__25000));
  nor2s1 __90__511234(.DIN1 (________26530), .DIN2 (________23812), .Q
       (___90___25035));
  nor2s1 __90___511235(.DIN1 (________23930), .DIN2 (________23924), .Q
       (____0___24648));
  nnd2s1 __900__511236(.DIN1 (________23336), .DIN2 (_____0__23929), .Q
       (________24947));
  nnd2s1 __90__511237(.DIN1 (_____9__23928), .DIN2 (________24710), .Q
       (_____0__24765));
  or2s1 __90___511238(.DIN1 (________23867), .DIN2 (___90___24071), .Q
       (________24756));
  nnd2s1 __9__0_511239(.DIN1 (________23999), .DIN2 (________24597), .Q
       (________24288));
  nnd2s1 __9____511240(.DIN1 (___0____23280), .DIN2 (________23927), .Q
       (________24861));
  nor2s1 __90___511241(.DIN1 (_____9__25728), .DIN2 (____0___23314), .Q
       (_____9__24477));
  or2s1 __9____511242(.DIN1 (________23753), .DIN2 (________25335), .Q
       (________24708));
  nnd2s1 __90__511243(.DIN1 (________25750), .DIN2 (________23953), .Q
       (________24484));
  nor2s1 __900__511244(.DIN1 (________23926), .DIN2 (___90___24077), .Q
       (_____9__24904));
  nnd2s1 __9____511245(.DIN1 (_____0__23758), .DIN2 (___0____25156), .Q
       (_____9__24315));
  nor2s1 __90_511246(.DIN1 (________25272), .DIN2 (_____0__24012), .Q
       (________24998));
  nnd2s1 __900_511247(.DIN1 (________23925), .DIN2 (____0___25229), .Q
       (________24417));
  nor2s1 __9___511248(.DIN1 (___9____23149), .DIN2 (________23581), .Q
       (____00__26408));
  nnd2s1 __90___511249(.DIN1 (________25607), .DIN2 (_____0__25339), .Q
       (________24870));
  nor2s1 __900__511250(.DIN1 (________23917), .DIN2 (________23922), .Q
       (________24717));
  nor2s1 __90___511251(.DIN1 (_____________________21736), .DIN2
       (____0___26594), .Q (________24489));
  nor2s1 __9____511252(.DIN1 (________23989), .DIN2 (________24517), .Q
       (________24281));
  nor2s1 __90___511253(.DIN1 (_____9__23918), .DIN2 (____0___23507), .Q
       (________24763));
  nnd2s1 __90___511254(.DIN1 (_____9__23928), .DIN2 (___99___25118), .Q
       (________24701));
  nor2s1 __90___511255(.DIN1 (___00___25132), .DIN2 (_____9__23472), .Q
       (________24596));
  hi1s1 __9____511256(.DIN (_____0__25349), .Q (___9____25039));
  nor2s1 __90___511257(.DIN1 (___0_0__25155), .DIN2 (________24010), .Q
       (________24707));
  or2s1 __90___511258(.DIN1 (_____________________21736), .DIN2
       (___9____25983), .Q (________25551));
  or2s1 __90___511259(.DIN1 (________24691), .DIN2 (________23924), .Q
       (________24728));
  nor2s1 __90__511260(.DIN1 (________23923), .DIN2 (________23922), .Q
       (________24899));
  hi1s1 __90___511261(.DIN (_____0__24326), .Q (________24789));
  nnd2s1 __90___511262(.DIN1 (____99__23501), .DIN2 (___00___25129), .Q
       (___0_9__27017));
  hi1s1 __90___511263(.DIN (________24976), .Q (________24771));
  nnd2s1 __90__511264(.DIN1 (________23921), .DIN2 (___90___24073), .Q
       (________24694));
  nor2s1 __90___511265(.DIN1 (________23920), .DIN2 (___9_9__25114), .Q
       (________24920));
  hi1s1 __90___511266(.DIN (_________37717), .Q (___9____25093));
  nor2s1 __90___511267(.DIN1 (________25376), .DIN2 (________23480), .Q
       (__9__0__29841));
  nnd2s1 __90___511268(.DIN1 (________24875), .DIN2 (___9_0__25095), .Q
       (________24761));
  nor2s1 __90__511269(.DIN1 (_____0__23919), .DIN2 (________25572), .Q
       (________24724));
  hi1s1 __9____511270(.DIN (____9___24830), .Q (____00__24746));
  nor2s1 __90___511271(.DIN1 (________23613), .DIN2 (___909__24079), .Q
       (________24709));
  nor2s1 __90___511272(.DIN1 (_____9__23918), .DIN2 (_____0__23568), .Q
       (________24808));
  nnd2s1 __90__511273(.DIN1 (________23925), .DIN2 (________26426), .Q
       (________24852));
  nor2s1 __90_0_511274(.DIN1 (____99__25585), .DIN2 (____99__24069), .Q
       (___0_9___31401));
  nnd2s1 __9__9_511275(.DIN1 (________23999), .DIN2 (________24720), .Q
       (_____9__24685));
  hi1s1 __90___511276(.DIN (___9_____39301), .Q (___9_____39688));
  nor2s1 __90___511277(.DIN1 (_____9__23348), .DIN2 (___0____25181), .Q
       (________25013));
  nor2s1 __90__511278(.DIN1 (____9___24738), .DIN2 (____9___24064), .Q
       (_____0__25596));
  nor2s1 __90___511279(.DIN1 (________23917), .DIN2 (________23916), .Q
       (________24891));
  nnd2s1 __90___511280(.DIN1 (________23915), .DIN2 (________24302), .Q
       (________24873));
  nnd2s1 __90___511281(.DIN1 (________23915), .DIN2 (________23624), .Q
       (_____0__24696));
  or2s1 __90__511282(.DIN1 (________23914), .DIN2 (________23913), .Q
       (________24912));
  hi1s1 __90___511283(.DIN (___0_90__40168), .Q (___99_0__39817));
  nnd2s1 __9____511284(.DIN1 (________23999), .DIN2 (____0___24748), .Q
       (________24778));
  nnd2s1 __9____511285(.DIN1 (________23999), .DIN2 (_____0__24895), .Q
       (____9___24737));
  hi1s1 ___9___511286(.DIN (_________36854), .Q (___900___38985));
  and2s1 __90_511287(.DIN1 (________23374), .DIN2 (________24710), .Q
       (_____0__24885));
  nnd2s1 __90___511288(.DIN1 (________23912), .DIN2 (________24490), .Q
       (________24732));
  nnd2s1 __90___511289(.DIN1 (________23925), .DIN2 (________23911), .Q
       (________24952));
  nnd2s1 __9____511290(.DIN1 (____9___23963), .DIN2 (___0____25172), .Q
       (________24714));
  hi1s1 ___9__511291(.DIN (___9_____39123), .Q (___9_____39274));
  nnd2s1 __9____511292(.DIN1 (____9___25023), .DIN2
       (_____________________21684), .Q (____9___26406));
  nnd2s1 __90___511293(.DIN1 (____9____38898), .DIN2 (___9____24127),
       .Q (___9____25081));
  hi1s1 __9___511294(.DIN (________24733), .Q (________25282));
  or2s1 __90_9_511295(.DIN1 (________27288), .DIN2 (____0___25590), .Q
       (_____9__24964));
  nor2s1 __90___511296(.DIN1 (_____________________21736), .DIN2
       (________24604), .Q (_____0__26528));
  or2s1 __9__0_511297(.DIN1 (________23715), .DIN2 (________25335), .Q
       (________24719));
  dffacs1 _________________________________________0__0_(.CLRB (reset),
       .CLK (clk), .DIN (___0____23298), .QN (___0__0__40581));
  nnd2s1 __90___511298(.DIN1 (_____0__23910), .DIN2 (_____9__23909), .Q
       (_____9__24735));
  hi1s1 __90__511299(.DIN (________25553), .Q (___9____25984));
  nnd2s1 __9__0_511300(.DIN1 (____9___24067), .DIN2
       (_____________________21732), .Q (________24968));
  nor2s1 __9__511301(.DIN1 (____09__23416), .DIN2 (___0_0__23281), .Q
       (_____9___37654));
  hi1s1 __9___511302(.DIN (________23908), .Q (________24767));
  nnd2s1 __90___511303(.DIN1 (________23394), .DIN2 (_____9__23909), .Q
       (________24892));
  hi1s1 __90___511304(.DIN (________25559), .Q (____0___29012));
  nor2s1 __9___511305(.DIN1 (____0_________________21724), .DIN2
       (_____9__24059), .Q (_____9__24793));
  hi1s1 __90__511306(.DIN (________23907), .Q (_________37687));
  nor2s1 __90___511307(.DIN1 (________24693), .DIN2 (____99__24069), .Q
       (_____0___34102));
  nnd2s1 __90___511308(.DIN1 (____0___23506), .DIN2 (___99___24165), .Q
       (_________35806));
  hi1s1 __9____511309(.DIN (___9_0__25978), .Q (_____0__25748));
  nor2s1 __90_0_511310(.DIN1 (________23906), .DIN2 (________23745), .Q
       (______9__37314));
  nor2s1 __90___511311(.DIN1 (________22981), .DIN2 (________23470), .Q
       (______0__35050));
  nor2s1 __90___511312(.DIN1 (________23363), .DIN2 (________23905), .Q
       (______9__34088));
  hi1s1 __9____511313(.DIN (________23904), .Q (____99__25028));
  nor2s1 __90___511314(.DIN1 (________23903), .DIN2 (___0____23275), .Q
       (_____0___38616));
  hi1s1 __9____511315(.DIN (___99____39861), .Q (______0__32803));
  nnd2s1 __90___511316(.DIN1 (________23902), .DIN2 (___9____23142), .Q
       (_________38842));
  nnd2s1 __90___511317(.DIN1 (________24713), .DIN2 (________23384), .Q
       (____9_9__37052));
  nnd2s1 __90___511318(.DIN1 (____9___23404), .DIN2 (________23901), .Q
       (_________36858));
  nnd2s1 __90___511319(.DIN1 (___9_9), .DIN2 (_____9__23520), .Q
       (___90____39051));
  nnd2s1 __90___511320(.DIN1 (______0__37673), .DIN2 (____9___23497),
       .Q (___90____39001));
  nor2s1 __90_0_511321(.DIN1 (________22753), .DIN2 (___0____24201), .Q
       (____9____35258));
  dffacs1 __________________511322(.CLRB (reset), .CLK (clk), .DIN
       (_____9__23396), .QN (_______________22076));
  nnd2s1 __90___511323(.DIN1 (________23576), .DIN2 (_____9__23900), .Q
       (_____0___38422));
  nor2s1 __909__(.DIN1 (inData[30]), .DIN2 (_____9___37656), .Q
       (________23898));
  hi1s1 __90___511324(.DIN (___90___24074), .Q (________23897));
  and2s1 __9____511325(.DIN1 (________23766), .DIN2 (_______22249), .Q
       (________23896));
  nor2s1 __909__511326(.DIN1 (________23672), .DIN2 (________23894), .Q
       (________23895));
  hi1s1 __90___511327(.DIN (___9____24111), .Q (________23893));
  nnd2s1 __90_9_511328(.DIN1 (_____0__23891), .DIN2 (________22463), .Q
       (________23892));
  xor2s1 __90___511329(.DIN1 (____0____36215), .DIN2 (____99___36174),
       .Q (____09__23890));
  nor2s1 __909__511330(.DIN1 (___0____23268), .DIN2 (___0_9__24187), .Q
       (____0___23889));
  nor2s1 __90_9_511331(.DIN1 (________24282), .DIN2 (____9___25578), .Q
       (____0___23888));
  nnd2s1 __90__511332(.DIN1 (___0____23245), .DIN2 (________23531), .Q
       (____0___23887));
  nnd2s1 ___99__511333(.DIN1 (___9____23206), .DIN2 (inData[24]), .Q
       (____0___23886));
  nnd2s1 __90___511334(.DIN1 (_____0___36728), .DIN2
       (_____________________________________________21812), .Q
       (____0___23885));
  or2s1 __90___511335(.DIN1
       (____________________________________________21866), .DIN2
       (_____0__23929), .Q (____0___23884));
  or2s1 __90900(.DIN1 (___0_____40419), .DIN2 (____0___23882), .Q
       (____0___23883));
  nor2s1 __900__511336(.DIN1 (______22153), .DIN2 (____99__23880), .Q
       (____00__23881));
  nor2s1 __90___511337(.DIN1 (____9___23878), .DIN2 (___9_9__23200), .Q
       (____9___23879));
  nor2s1 __909__511338(.DIN1 (________22796), .DIN2 (____9___23876), .Q
       (____9___23877));
  or2s1 __90___511339(.DIN1 (____0___23044), .DIN2 (____9___23874), .Q
       (____9___23875));
  or2s1 __900__511340(.DIN1 (___9_0__29602), .DIN2 (___00___23220), .Q
       (____9___23873));
  nnd2s1 __90___511341(.DIN1 (_____0___36728), .DIN2 (_____9__23871),
       .Q (____90__23872));
  nnd2s1 __90___511342(.DIN1 (_____0__23417), .DIN2 (___90___25034), .Q
       (________23870));
  nor2s1 __90_511343(.DIN1 (____0_______________), .DIN2
       (_____9__23057), .Q (________23869));
  nor2s1 __90___511344(.DIN1 (________23867), .DIN2 (________23866), .Q
       (________23868));
  or2s1 __90___511345(.DIN1 (________23864), .DIN2 (_____9__25823), .Q
       (________23865));
  and2s1 __909_9(.DIN1 (________26643), .DIN2
       (____0_________________21726), .Q (________23863));
  nnd2s1 __90___511346(.DIN1 (_________34145), .DIN2 (___00___23216),
       .Q (_____0__23862));
  nor2s1 __90___511347(.DIN1 (________23860), .DIN2 (________24734), .Q
       (_____9__23861));
  nor2s1 __90___511348(.DIN1 (________22990), .DIN2 (____9___23690), .Q
       (________23859));
  nnd2s1 __909__511349(.DIN1 (________23084), .DIN2 (____9___22832), .Q
       (________23858));
  nor2s1 __90___511350(.DIN1 (____9___24063), .DIN2 (____0___24463), .Q
       (________23857));
  nor2s1 __90___511351(.DIN1 (________23074), .DIN2 (___0____23229), .Q
       (________23856));
  nnd2s1 __9__9_511352(.DIN1 (________25320), .DIN2 (________23362), .Q
       (________23855));
  nnd2s1 __90__511353(.DIN1 (___0____23246), .DIN2 (clk), .Q
       (________23854));
  nor2s1 __90___511354(.DIN1 (_____0__23852), .DIN2 (___0____23232), .Q
       (________23853));
  nor2s1 __900__511355(.DIN1 (_____9__24382), .DIN2 (_____9__23767), .Q
       (_____9__23851));
  nnd2s1 ___9_9_511356(.DIN1 (___9____23199), .DIN2 (inData[30]), .Q
       (________23850));
  nnd2s1 __9099_(.DIN1 (________24877), .DIN2 (____09__23048), .Q
       (________23849));
  nor2s1 __90000(.DIN1 (________23847), .DIN2 (_____9__24695), .Q
       (________23848));
  or2s1 __90___511357(.DIN1 (___0_____40436), .DIN2 (________23845), .Q
       (________23846));
  hi1s1 __90___511358(.DIN (________26258), .Q (________23844));
  or2s1 __9_0__511359(.DIN1 (_____9__23842), .DIN2 (________23930), .Q
       (_____0__23843));
  nnd2s1 __9_0__511360(.DIN1 (___90___25030), .DIN2 (________23011), .Q
       (________23841));
  nnd2s1 ___99_511361(.DIN1 (________23085), .DIN2 (inData[18]), .Q
       (________23839));
  nnd2s1 __90___511362(.DIN1 (_____9___38509), .DIN2 (___0____23231),
       .Q (________23838));
  xor2s1 __90___511363(.DIN1
       (____________________________________________21848), .DIN2
       (___99_0__39864), .Q (________23837));
  nor2s1 ___9__511364(.DIN1 (___99____39814), .DIN2 (___0____23230), .Q
       (________23836));
  or2s1 __90___511365(.DIN1 (_____0__26149), .DIN2 (_____9__25823), .Q
       (_____0__23835));
  nor2s1 ___9___511366(.DIN1 (________26530), .DIN2 (________23119), .Q
       (_____9__23834));
  nnd2s1 __9___511367(.DIN1 (________23432), .DIN2 (____0___23600), .Q
       (________23833));
  xnr2s1 __90___511368(.DIN1
       (__________________________________________9___21934), .DIN2
       (_________36349), .Q (________23832));
  nnd2s1 ___99__511369(.DIN1 (_____9__25469), .DIN2 (___9_0__23173), .Q
       (________23831));
  and2s1 __909_511370(.DIN1 (__90_0__29699), .DIN2 (________23100), .Q
       (________23830));
  nnd2s1 __90___511371(.DIN1 (_____0__23105), .DIN2 (_____0__22989), .Q
       (________23829));
  nnd2s1 __9____511372(.DIN1 (___000), .DIN2 (____0___23599), .Q
       (________23827));
  nor2s1 __90___511373(.DIN1 (___9_0__29602), .DIN2 (___0____23241), .Q
       (_____0__23826));
  nor2s1 __9____511374(.DIN1 (________24475), .DIN2 (________24322), .Q
       (_____9__23825));
  nor2s1 __90_0_511375(.DIN1 (____0_0__38093), .DIN2 (_____9__23113),
       .Q (________23824));
  nnd2s1 __9____511376(.DIN1 (___0____25176), .DIN2 (____9___24358), .Q
       (________23823));
  nor2s1 __9_00_(.DIN1 (________23440), .DIN2 (________23755), .Q
       (________23822));
  xor2s1 __90___511377(.DIN1 (______0__38256), .DIN2 (_________38456),
       .Q (________23821));
  or2s1 __90___511378(.DIN1 (________23984), .DIN2 (____9___25578), .Q
       (________23820));
  nor2s1 __9____511379(.DIN1 (________23724), .DIN2 (________23922), .Q
       (________23819));
  and2s1 __90___511380(.DIN1 (___0____25176), .DIN2
       (____0________________21663), .Q (________23818));
  nor2s1 __90__511381(.DIN1 (___0_____40416), .DIN2 (________23845), .Q
       (________23817));
  nnd2s1 __90___511382(.DIN1 (___9____23198), .DIN2 (______22153), .Q
       (_____0__23816));
  nnd2s1 __90___511383(.DIN1 (___9____23193), .DIN2 (inData[28]), .Q
       (________23815));
  or2s1 __90___511384(.DIN1 (___0_9__25154), .DIN2 (____9___25578), .Q
       (________23814));
  hi1s1 __90___511385(.DIN (________23812), .Q (________23813));
  hi1s1 __90_511386(.DIN (___9____24082), .Q (________23811));
  nor2s1 __90___511387(.DIN1 (________24910), .DIN2 (___9____24156), .Q
       (________23810));
  nor2s1 ___990_511388(.DIN1 (________23800), .DIN2 (____0___23046), .Q
       (________23809));
  nnd2s1 __9__0_511389(.DIN1 (________23419), .DIN2 (___9____25110), .Q
       (________23808));
  nnd2s1 __909__511390(.DIN1 (________23845), .DIN2 (________23099), .Q
       (_____0__23807));
  nor2s1 __90__511391(.DIN1 (________23805), .DIN2 (___0____25143), .Q
       (_____9__23806));
  nnd2s1 ___99_511392(.DIN1 (___9____23194), .DIN2 (______9__32360), .Q
       (________23804));
  nor2s1 __90___511393(.DIN1 (_____0__23852), .DIN2 (___90___23135), .Q
       (________23803));
  nnd2s1 __9____511394(.DIN1 (________23801), .DIN2 (________23800), .Q
       (________23802));
  and2s1 __90___511395(.DIN1 (____0___23598), .DIN2 (________22816), .Q
       (________23799));
  nor2s1 __90__511396(.DIN1 (_____9__22908), .DIN2 (_____0__23656), .Q
       (________23798));
  or2s1 __90___511397(.DIN1 (________22374), .DIN2 (________25946), .Q
       (_____0__23797));
  hi1s1 __9____511398(.DIN (____0___23795), .Q (____09__23796));
  nor2s1 __90___511399(.DIN1 (___9____23204), .DIN2 (________25946), .Q
       (____0___23794));
  nnd2s1 __9____511400(.DIN1 (___9____23188), .DIN2 (________23517), .Q
       (____0___23793));
  xor2s1 __90___511401(.DIN1 (___0___22274), .DIN2 (____0____36215), .Q
       (____0___23792));
  nor2s1 __9__0_511402(.DIN1 (________23930), .DIN2 (________23922), .Q
       (____0___23791));
  and2s1 __909_0(.DIN1 (___90___25030), .DIN2 (____0___23789), .Q
       (____0___23790));
  or2s1 __9__9_511403(.DIN1 (____9___23786), .DIN2 (____0___23696), .Q
       (____99__23787));
  nor2s1 __90___511404(.DIN1 (____0___24564), .DIN2 (____9___25578), .Q
       (____9___23785));
  nor2s1 __9____511405(.DIN1 (________22852), .DIN2 (_____9__23737), .Q
       (____9___23784));
  and2s1 __9____511406(.DIN1 (________26643), .DIN2 (____9___23782), .Q
       (____9___23783));
  nnd2s1 __90___511407(.DIN1 (________23433), .DIN2 (___0____23267), .Q
       (____9___23781));
  nnd2s1 __90___511408(.DIN1 (_____0__23891), .DIN2
       (____________________________________________21867), .Q
       (____9___23780));
  xor2s1 __90__511409(.DIN1 (___0_9___40558), .DIN2 (_________38533),
       .Q (____9___23779));
  xor2s1 __90___511410(.DIN1 (___0_____40525), .DIN2 (_____9___35917),
       .Q (____90__23778));
  nnd2s1 __90___511411(.DIN1 (_____0___36728), .DIN2 (____0_0__36258),
       .Q (_____9__23777));
  or2s1 __90___511412(.DIN1 (___0_____40418), .DIN2 (________23845), .Q
       (________23776));
  xor2s1 __90___511413(.DIN1 (____90__22929), .DIN2
       (_________________________________________________________________________________________22090),
       .Q (________23775));
  xor2s1 __90___511414(.DIN1 (________22987), .DIN2 (____0___22746), .Q
       (________23774));
  nor2s1 __90_0_511415(.DIN1 (____0____37167), .DIN2 (___9____23184),
       .Q (________23773));
  nor2s1 __9____511416(.DIN1 (________22536), .DIN2 (________24978), .Q
       (________23772));
  nor2s1 __90_0_511417(.DIN1 (________23770), .DIN2 (________24594), .Q
       (________23771));
  nnd2s1 __9____511418(.DIN1 (___9____26025), .DIN2 (____0___26410), .Q
       (________23769));
  nnd2s1 __90___511419(.DIN1 (___9_9), .DIN2 (___00___23219), .Q
       (_____0__23768));
  nor2s1 __900__511420(.DIN1 (_____9__24486), .DIN2 (_____9__23767), .Q
       (___0____24253));
  xnr2s1 __90___511421(.DIN1 (____9_9__37984), .DIN2 (____0___22647),
       .Q (________24668));
  nnd2s1 __9____511422(.DIN1 (________23766), .DIN2 (____0___22844), .Q
       (________24479));
  nor2s1 __9___511423(.DIN1 (____0___22745), .DIN2 (___99___23211), .Q
       (________24279));
  hi1s1 __90___511424(.DIN (________23765), .Q (_____0__24536));
  and2s1 __9____511425(.DIN1 (___0____23258), .DIN2 (________23667), .Q
       (________24294));
  nnd2s1 __90___511426(.DIN1 (________23764), .DIN2 (_____0__23891), .Q
       (________24482));
  nnd2s1 __9_0__511427(.DIN1 (_____0__23454), .DIN2 (________23073), .Q
       (________24298));
  and2s1 __9_0__511428(.DIN1 (____0___23699), .DIN2 (____0___23601), .Q
       (________24480));
  hi1s1 __90__511429(.DIN (________23763), .Q (________26731));
  hi1s1 __90___511430(.DIN (________23762), .Q (_____9__24392));
  nor2s1 __90__511431(.DIN1 (________24308), .DIN2 (____9___25578), .Q
       (___9_0__24090));
  hi1s1 __9____511432(.DIN (________23761), .Q (_____0__24666));
  hi1s1 __9____511433(.DIN (___00___24169), .Q (________24408));
  nnd2s1 __9____511434(.DIN1 (________23760), .DIN2
       (_____________________21732), .Q (________23908));
  hi1s1 __9___511435(.DIN (______9__35170), .Q (________24622));
  nor2s1 __9_0__511436(.DIN1 (________23860), .DIN2 (___0____24224), .Q
       (________24502));
  nor2s1 __900__511437(.DIN1 (________23759), .DIN2 (____9___23874), .Q
       (_____9__23944));
  hi1s1 __90___511438(.DIN (___9__9__39459), .Q (___9____25085));
  nnd2s1 __900_511439(.DIN1 (___9____23202), .DIN2
       (_____________________21681), .Q (___99___24163));
  nnd2s1 __9_0__511440(.DIN1 (_____0__23929), .DIN2 (________22752), .Q
       (_____9__25575));
  hi1s1 __9___511441(.DIN (___0____24191), .Q (________24292));
  nor2s1 __9_0__511442(.DIN1 (________23056), .DIN2 (________23461), .Q
       (_____9__23938));
  hi1s1 __9__0_511443(.DIN (_____0__23758), .Q (________24295));
  nor2s1 __9__00(.DIN1 (________22684), .DIN2 (________23751), .Q
       (________23907));
  nnd2s1 __9____511444(.DIN1 (_________38164), .DIN2 (___0_0___40567),
       .Q (________24436));
  hi1s1 __90_0_511445(.DIN (____0___23980), .Q (________24485));
  hi1s1 __90_0_511446(.DIN (________23921), .Q (____0___24369));
  nnd2s1 __9____511447(.DIN1 (________24033), .DIN2
       (_____________________21742), .Q (________24329));
  hi1s1 __90___511448(.DIN (___9_0__25068), .Q (____9___24449));
  and2s1 __9___511449(.DIN1 (_____9__23757), .DIN2 (___0____25157), .Q
       (________24472));
  nnd2s1 __9____511450(.DIN1 (_____9__23757), .DIN2 (________24490), .Q
       (________24330));
  hi1s1 __9____511451(.DIN (____0___23977), .Q (_____0__24506));
  nnd2s1 __9___511452(.DIN1 (______9__35039), .DIN2 (________26426), .Q
       (____9___24640));
  hi1s1 __9____511453(.DIN (___90___24078), .Q (________24704));
  hi1s1 __9____511454(.DIN (_____9__25019), .Q (________24697));
  hi1s1 __90__511455(.DIN (____9___23968), .Q (________24507));
  nnd2s1 __9____511456(.DIN1 (____9___23127), .DIN2 (___9_0__24139), .Q
       (____9___24547));
  nor2s1 __9__09(.DIN1 (_____________________21709), .DIN2
       (________23756), .Q (________24474));
  nnd2s1 __9____511457(.DIN1 (___99___25123), .DIN2 (________23933), .Q
       (_____9__24447));
  nor2s1 __9_090(.DIN1 (________24602), .DIN2 (________23756), .Q
       (________24581));
  nnd2s1 __9____511458(.DIN1 (________23755), .DIN2 (________23754), .Q
       (________24599));
  nor2s1 __9____511459(.DIN1 (________23753), .DIN2 (___99___25119), .Q
       (________24290));
  hi1s1 __90_0_511460(.DIN (_____9__23991), .Q (____0___24460));
  nor2s1 __9_09_(.DIN1 (___9_9__23163), .DIN2 (________23098), .Q
       (____99__24457));
  nnd2s1 __9_09_511461(.DIN1 (___90___24073), .DIN2 (________23752), .Q
       (____0___24465));
  nnd2s1 __9____511462(.DIN1 (________23751), .DIN2
       (____0________________21667), .Q (_____0__24326));
  hi1s1 __9___511463(.DIN (______9__33955), .Q (________24500));
  hi1s1 __9____511464(.DIN (________23750), .Q (____9___24644));
  hi1s1 __9____511465(.DIN (________25607), .Q (________25549));
  nor2s1 __9____511466(.DIN1 (________23024), .DIN2 (________23749), .Q
       (________24614));
  hi1s1 __9____511467(.DIN (________24010), .Q (________24607));
  nor2s1 __90___511468(.DIN1 (___0____25152), .DIN2 (________24901), .Q
       (_____0__24468));
  nnd2s1 __9____511469(.DIN1 (________23906), .DIN2 (______22154), .Q
       (________24353));
  nnd2s1 __9____511470(.DIN1 (_____0__23748), .DIN2 (________26601), .Q
       (________24976));
  hi1s1 __9____511471(.DIN (________25923), .Q (________25278));
  hi1s1 __9____511472(.DIN (________24909), .Q (____0___25412));
  hi1s1 __90___511473(.DIN (___9____24146), .Q (____90__25758));
  nnd2s1 __9____511474(.DIN1 (________23059), .DIN2
       (_____________________21690), .Q (___900__25958));
  nor2s1 __9___511475(.DIN1 (________24602), .DIN2 (________23847), .Q
       (____09__24467));
  hi1s1 __9___511476(.DIN (_____9__23747), .Q (________25920));
  nnd2s1 __9____511477(.DIN1 (________23744), .DIN2
       (____0________________21667), .Q (________24504));
  nnd2s1 __90___511478(.DIN1 (___9____23178), .DIN2
       (_____________________21705), .Q (___9_____39123));
  hi1s1 __9___511479(.DIN (________24995), .Q (____9___25404));
  hi1s1 __9___511480(.DIN (___00___25130), .Q (________24908));
  hi1s1 __90___511481(.DIN (___9_____39183), .Q (____9____34315));
  dffacs1 _________________________________________0_____511482(.CLRB
       (reset), .CLK (clk), .DIN (___00___23223), .Q (___0_0___40568));
  hi1s1 __90_0_511483(.DIN (_________34775), .Q (____9____38948));
  hi1s1 __90__511484(.DIN (_________33596), .Q (_________33843));
  nor2s1 __9__9_511485(.DIN1 (____9___24066), .DIN2 (________23664), .Q
       (________25559));
  hi1s1 __90___511486(.DIN (________24722), .Q (_____0__25556));
  hi1s1 __9____511487(.DIN (________25750), .Q (____0___26409));
  nor2s1 __9__9_511488(.DIN1 (_____0__22375), .DIN2 (_____0___36728),
       .Q (_________37717));
  nnd2s1 __9___511489(.DIN1 (____0___23694), .DIN2 (____9___24066), .Q
       (________24886));
  hi1s1 __90___511490(.DIN (________23746), .Q (________25345));
  hi1s1 __9____511491(.DIN (________23745), .Q (_________34796));
  nor2s1 __9__0_511492(.DIN1 (________22980), .DIN2 (___00___23221), .Q
       (_________38876));
  nor2s1 __9____511493(.DIN1 (________22679), .DIN2 (________23744), .Q
       (___0_____40308));
  nor2s1 __909_511494(.DIN1 (________23618), .DIN2 (________24322), .Q
       (________23743));
  and2s1 __90___511495(.DIN1 (________23741), .DIN2 (________23356), .Q
       (________23742));
  or2s1 __90___511496(.DIN1 (____0______________), .DIN2
       (________23090), .Q (________23740));
  nnd2s1 __90__511497(.DIN1 (___9____26025), .DIN2 (________23611), .Q
       (________23739));
  nor2s1 __90_511498(.DIN1 (_____9__23737), .DIN2 (________24470), .Q
       (_____0__23738));
  nnd2s1 __90_511499(.DIN1 (_____0___36728), .DIN2 (____9__22234), .Q
       (________23736));
  nnd2s1 __9090_(.DIN1 (____0___23605), .DIN2 (________23734), .Q
       (________23735));
  nnd2s1 __909__511500(.DIN1 (_________38164), .DIN2 (_________36883),
       .Q (________23733));
  nnd2s1 __909__511501(.DIN1 (___9____23186), .DIN2 (___900), .Q
       (________23732));
  or2s1 __909_511502(.DIN1 (__________________0_), .DIN2
       (___99___23214), .Q (________23731));
  and2s1 __909__511503(.DIN1 (________23741), .DIN2
       (_____________________21671), .Q (________23730));
  nnd2s1 __9__511504(.DIN1 (_____0__23728), .DIN2 (________23063), .Q
       (________23729));
  nnd2s1 __909__511505(.DIN1 (________23749), .DIN2 (________23726), .Q
       (_____9__23727));
  or2s1 __909__511506(.DIN1 (________23724), .DIN2 (___0____24239), .Q
       (________23725));
  nor2s1 __9____511507(.DIN1
       (______________________________________________________________________________________0__22093),
       .DIN2 (_________38164), .Q (________23723));
  nor2s1 __909_511508(.DIN1 (_____9__22800), .DIN2 (________23721), .Q
       (________23722));
  nor2s1 __909__511509(.DIN1 (______), .DIN2 (________23660), .Q
       (________23720));
  nor2s1 __909__511510(.DIN1 (________22972), .DIN2 (________23064), .Q
       (________23719));
  nor2s1 __9099_511511(.DIN1 (____0________________21662), .DIN2
       (___90_), .Q (_____9__23718));
  nor2s1 __9____511512(.DIN1 (________25931), .DIN2 (_________41353),
       .Q (________23717));
  or2s1 __9___511513(.DIN1 (________23614), .DIN2 (________23715), .Q
       (________23716));
  hi1s1 __9____511514(.DIN (________26269), .Q (________23714));
  nor2s1 __9_0__511515(.DIN1 (________23754), .DIN2 (________23088), .Q
       (________23713));
  nor2s1 __9_0__511516(.DIN1 (_____0__23058), .DIN2 (________22799), .Q
       (________23712));
  or2s1 __9_0__511517(.DIN1 (___0____24224), .DIN2 (_____0__24316), .Q
       (_____0__23711));
  nor2s1 __9____511518(.DIN1 (________23709), .DIN2 (___9_0__24080), .Q
       (_____9__23710));
  nor2s1 __9090_511519(.DIN1 (________24475), .DIN2 (________23103), .Q
       (________23708));
  nor2s1 ___99__511520(.DIN1 (________22722), .DIN2 (___099__23309), .Q
       (________23707));
  nor2s1 __909__511521(.DIN1 (___9_0__23201), .DIN2 (___0____24239), .Q
       (________23706));
  hi1s1 __90_9_511522(.DIN (___90___24075), .Q (________23705));
  hi1s1 __90__511523(.DIN (________23703), .Q (________23704));
  and2s1 __9090_511524(.DIN1 (_________38164), .DIN2 (___0_____40494),
       .Q (____09__23701));
  and2s1 __9____511525(.DIN1 (____0___23699), .DIN2 (___0_9__24217), .Q
       (____0___23700));
  nor2s1 __9____511526(.DIN1 (____0___23697), .DIN2 (____0___23696), .Q
       (____0___23698));
  and2s1 __9____511527(.DIN1 (_____9__23067), .DIN2 (____0___23694), .Q
       (____0___23695));
  nnd2s1 __90___511528(.DIN1 (_____9__23918), .DIN2 (________23053), .Q
       (____0___23693));
  nnd2s1 ___999_511529(.DIN1 (________23112), .DIN2 (________23481), .Q
       (____00__23692));
  nor2s1 __9__9_511530(.DIN1 (________22492), .DIN2 (____9___23690), .Q
       (____99__23691));
  nnd2s1 __9__0_511531(.DIN1 (___0____23255), .DIN2 (________24308), .Q
       (____9___23689));
  nor2s1 ___99__511532(.DIN1 (___0_____40622), .DIN2 (________25946),
       .Q (____9___23688));
  hi1s1 __90___511533(.DIN (____9___23685), .Q (____9___23686));
  nor2s1 __9____511534(.DIN1 (___9____23167), .DIN2 (___0_9__23234), .Q
       (____9___23684));
  and2s1 __9__0_511535(.DIN1 (_____9__23682), .DIN2 (________24033), .Q
       (____90__23683));
  nor2s1 __9__0_511536(.DIN1 (_____________________21705), .DIN2
       (___0____25152), .Q (________23681));
  nnd2s1 __9____511537(.DIN1 (___0____23228), .DIN2 (___9____23187), .Q
       (________23680));
  or2s1 __9__511538(.DIN1 (________24691), .DIN2 (________24757), .Q
       (________23679));
  nnd2s1 __9__9_511539(.DIN1 (____0___23604), .DIN2 (____0___26590), .Q
       (________23678));
  xor2s1 __90__511540(.DIN1 (___0__9__40550), .DIN2 (_________36527),
       .Q (________23677));
  nor2s1 ___9___511541(.DIN1 (__99_9__30508), .DIN2 (________23060), .Q
       (________23676));
  nnd2s1 ___9___511542(.DIN1 (________23441), .DIN2 (___0____23233), .Q
       (________23675));
  nnd2s1 __9____511543(.DIN1 (____9___23593), .DIN2 (___0_0__24248), .Q
       (_____0__23674));
  or2s1 __9___511544(.DIN1 (________23672), .DIN2 (___0_9__24187), .Q
       (_____9__23673));
  hi1s1 __9____511545(.DIN (________23670), .Q (________23671));
  and2s1 __9____511546(.DIN1 (________23933), .DIN2 (________23667), .Q
       (________23668));
  nor2s1 __9__9_511547(.DIN1 (_____0__25417), .DIN2 (_____0__24316), .Q
       (_____0__23666));
  nor2s1 __9_00_511548(.DIN1 (________23066), .DIN2 (________23664), .Q
       (_____9__23665));
  nnd2s1 __9____511549(.DIN1 (___0____25152), .DIN2 (________23662), .Q
       (________23663));
  nor2s1 __9____511550(.DIN1 (________23959), .DIN2 (________23660), .Q
       (________23661));
  nor2s1 __9___511551(.DIN1 (_____9__23842), .DIN2 (________24691), .Q
       (________23659));
  nor2s1 __9__0_511552(.DIN1 (________22804), .DIN2 (___99___23209), .Q
       (________23658));
  nor2s1 __9__90(.DIN1 (________22494), .DIN2 (_____0__23656), .Q
       (________23657));
  nnd2s1 __9__9_511553(.DIN1 (_____9__23682), .DIN2 (________24993), .Q
       (_____9__23655));
  or2s1 __9__0_511554(.DIN1 (________25272), .DIN2 (_____0__24316), .Q
       (________23654));
  or2s1 __9__0_511555(.DIN1 (___9____23151), .DIN2 (________24978), .Q
       (________23653));
  and2s1 __9____511556(.DIN1 (________23651), .DIN2
       (____0_________________21725), .Q (________23652));
  and2s1 __9____511557(.DIN1 (________23741), .DIN2 (____0___23504), .Q
       (________23650));
  or2s1 __9____511558(.DIN1 (_____9__23737), .DIN2 (________24017), .Q
       (________23649));
  nnd2s1 __9__511559(.DIN1 (________26450), .DIN2
       (____0_______________), .Q (________23648));
  nor2s1 __900__511560(.DIN1 (________24711), .DIN2 (_____0__23646), .Q
       (________23647));
  or2s1 __9___511561(.DIN1 (________23429), .DIN2 (________23651), .Q
       (_____9__23645));
  or2s1 __9____511562(.DIN1 (________24703), .DIN2 (___0_0__23253), .Q
       (________23644));
  nor2s1 __9____511563(.DIN1 (________22973), .DIN2 (________23642), .Q
       (________23643));
  nnd2s1 __9____511564(.DIN1 (________23640), .DIN2 (________23766), .Q
       (________23641));
  or2s1 __9____511565(.DIN1 (___0____25163), .DIN2 (________24786), .Q
       (________23639));
  or2s1 __9___511566(.DIN1 (_____9__23737), .DIN2 (________23637), .Q
       (________23638));
  or2s1 __9____511567(.DIN1 (_____9__23635), .DIN2 (_____9__23737), .Q
       (_____0__23636));
  nor2s1 __9____511568(.DIN1 (_____0__23445), .DIN2 (___9____23176), .Q
       (________23634));
  or2s1 __9____511569(.DIN1 (________24691), .DIN2 (________23922), .Q
       (________23633));
  nnd2s1 __9__0_511570(.DIN1 (________23664), .DIN2 (______22154), .Q
       (________23632));
  or2s1 __9____511571(.DIN1 (________23715), .DIN2 (___99___25119), .Q
       (________23631));
  nnd2s1 __900__511572(.DIN1 (________23629), .DIN2 (________23448), .Q
       (________23630));
  nor2s1 __9___511573(.DIN1 (____9___23591), .DIN2 (________23078), .Q
       (________23628));
  nnd2s1 __9__9_511574(.DIN1 (___0____25198), .DIN2 (________24760), .Q
       (________23627));
  nor2s1 __9__0_511575(.DIN1 (______22154), .DIN2 (________23664), .Q
       (_____0__23626));
  and2s1 __900__511576(.DIN1 (________25458), .DIN2 (________23624), .Q
       (_____9__23625));
  nnd2s1 __9____511577(.DIN1 (___9____23183), .DIN2 (___0____23276), .Q
       (________23623));
  and2s1 ___99__511578(.DIN1 (___0____23226), .DIN2 (____9___23125), .Q
       (________23622));
  nor2s1 __90___511579(.DIN1 (___0_____40428), .DIN2 (___9_____39575),
       .Q (________23621));
  nor2s1 ___9_9_511580(.DIN1 (________23102), .DIN2 (________23097), .Q
       (________23620));
  nor2s1 __909_511581(.DIN1 (________23618), .DIN2 (________24731), .Q
       (________23619));
  nor2s1 __9_0__511582(.DIN1 (_____0__22721), .DIN2 (________26450), .Q
       (________24519));
  and2s1 __9____511583(.DIN1 (___9_0__24139), .DIN2 (________25343), .Q
       (________24314));
  nor2s1 __9____511584(.DIN1 (________23423), .DIN2 (___9_____39575),
       .Q (________23899));
  nor2s1 __9_0__511585(.DIN1 (________23930), .DIN2 (________23916), .Q
       (_____0__24287));
  and2s1 __9__0_511586(.DIN1 (_____9__26616), .DIN2
       (____0_________________21725), .Q (________24318));
  nor2s1 __9_0_0(.DIN1 (____9___23400), .DIN2 (________23055), .Q
       (____0___24462));
  nor2s1 __9____511587(.DIN1 (________23724), .DIN2 (___990__24158), .Q
       (________24469));
  and2s1 __9____511588(.DIN1 (________23760), .DIN2 (___0_9__24217), .Q
       (_____0__24307));
  nor2s1 __9____511589(.DIN1 (____0________________21716), .DIN2
       (________28994), .Q (________23904));
  nor2s1 __9____511590(.DIN1 (____0___24564), .DIN2 (________24308), .Q
       (_____9__23951));
  xor2s1 __9___511591(.DIN1 (___0_0__22324), .DIN2 (______0__34897), .Q
       (_____0__24576));
  nnd2s1 __9____511592(.DIN1 (_____0__23617), .DIN2 (________24625), .Q
       (________23948));
  nor2s1 __9____511593(.DIN1 (_____9__23616), .DIN2 (________23446), .Q
       (________25702));
  or2s1 __9____511594(.DIN1 (________25327), .DIN2 (________23753), .Q
       (________24321));
  nor2s1 __9_0__511595(.DIN1 (________23109), .DIN2 (________23615), .Q
       (________23936));
  nor2s1 __9____511596(.DIN1 (________24338), .DIN2 (___0____23250), .Q
       (________23949));
  nnd2s1 __9___511597(.DIN1 (________23629), .DIN2 (________25355), .Q
       (________24293));
  nor2s1 __9_0__511598(.DIN1 (________23614), .DIN2 (________23612), .Q
       (________24310));
  nor2s1 __9____511599(.DIN1 (________23613), .DIN2 (________25376), .Q
       (___9____24086));
  nor2s1 __9_0_511600(.DIN1 (________23612), .DIN2 (________25327), .Q
       (_____9__24031));
  and2s1 __9_0__511601(.DIN1 (___9____26025), .DIN2
       (____0_________________21727), .Q (________24661));
  hi1s1 __90_9_511602(.DIN (________23931), .Q (________24312));
  nnd2s1 __9_0__511603(.DIN1 (________26643), .DIN2 (________23611), .Q
       (________25878));
  nnd2s1 __9_0__511604(.DIN1 (______0__37673), .DIN2 (_____0__23114),
       .Q (________24283));
  nor2s1 __9_0_9(.DIN1 (________23610), .DIN2 (________23107), .Q
       (___0____24233));
  nnd2s1 __9_0__511605(.DIN1 (_____0___36728), .DIN2 (___9__22156), .Q
       (________24511));
  nor2s1 __90__511606(.DIN1 (________23609), .DIN2 (___9____24156), .Q
       (________24523));
  nnd2s1 __9_0__511607(.DIN1 (________24782), .DIN2 (________24766), .Q
       (________24471));
  hi1s1 __9____511608(.DIN (________23608), .Q (________24568));
  hi1s1 __90___511609(.DIN (_____0__23607), .Q (________24438));
  hi1s1 __90___511610(.DIN (___909__24079), .Q (____00__24556));
  hi1s1 __90_511611(.DIN (____09__23606), .Q (_____0__24497));
  hi1s1 __90___511612(.DIN (________24328), .Q (________25260));
  nnd2s1 __9____511613(.DIN1 (_____0__23891), .DIN2 (_____9___33157),
       .Q (___9_9__24089));
  nnd2s1 __9____511614(.DIN1 (________23629), .DIN2 (________23766), .Q
       (___090__24257));
  hi1s1 __90___511615(.DIN (___9_9__25114), .Q (____9___24361));
  nnd2s1 __9__9_511616(.DIN1 (___99___23215), .DIN2
       (_____________________21745), .Q (________24853));
  or2s1 __9____511617(.DIN1 (_____________________21732), .DIN2
       (________23664), .Q (________24348));
  and2s1 __9____511618(.DIN1 (_____0__23748), .DIN2 (________26272), .Q
       (________24630));
  nor2s1 __9____511619(.DIN1 (____00__23597), .DIN2 (____9___23690), .Q
       (________24327));
  nnd2s1 __9____511620(.DIN1 (_____9__23757), .DIN2 (________24313), .Q
       (_____9__24286));
  nor2s1 __9____511621(.DIN1 (________23065), .DIN2 (________23664), .Q
       (________25787));
  nor2s1 __90___511622(.DIN1 (________23020), .DIN2 (____9___23874), .Q
       (________24619));
  nnd2s1 __9____511623(.DIN1 (________24304), .DIN2 (____0___23605), .Q
       (________24320));
  nnd2s1 __9__511624(.DIN1 (___9____24084), .DIN2 (____0___23604), .Q
       (_____0__24277));
  nnd2s1 __90___511625(.DIN1 (________23764), .DIN2 (___90___25034), .Q
       (________24473));
  nnd2s1 __9____511626(.DIN1 (___9_____39575), .DIN2
       (____0________________21716), .Q (________24531));
  nnd2s1 __9___511627(.DIN1 (___000__25125), .DIN2 (____0___23603), .Q
       (________24309));
  hi1s1 __9____511628(.DIN (___0____24195), .Q (________24384));
  nnd2s1 __9____511629(.DIN1 (___0_0__23244), .DIN2 (____0___23602), .Q
       (_____9__24439));
  nor2s1 __90__511630(.DIN1 (________23926), .DIN2 (_____9__23767), .Q
       (________24303));
  nnd2s1 __9__0_511631(.DIN1 (____0___23694), .DIN2 (____0___23601), .Q
       (________24902));
  nor2s1 __9_0__511632(.DIN1 (____0___23600), .DIN2 (________23753), .Q
       (_____0__24297));
  nnd2s1 __9_0__511633(.DIN1 (________23751), .DIN2 (____0___23599), .Q
       (________24509));
  nnd2s1 __90___511634(.DIN1 (____0___23598), .DIN2 (____90__23029), .Q
       (________25331));
  nor2s1 __9_0_511635(.DIN1 (____00__23597), .DIN2 (________28994), .Q
       (____9___24642));
  nnd2s1 __9___511636(.DIN1 (____99__23596), .DIN2 (____9___23970), .Q
       (________24733));
  hi1s1 __90_9_511637(.DIN (____9___23595), .Q (________24389));
  nnd2s1 __9____511638(.DIN1 (________23905), .DIN2 (________23989), .Q
       (________24673));
  nnd2s1 __9____511639(.DIN1 (___0____26077), .DIN2 (________25751), .Q
       (___0____25206));
  nor2s1 __9__9_511640(.DIN1 (____09__26331), .DIN2 (_____9__24705), .Q
       (________25375));
  nnd2s1 __9__9_511641(.DIN1 (________26450), .DIN2 (____90__24060), .Q
       (_____9__24954));
  nnd2s1 __9___511642(.DIN1 (____9___23593), .DIN2 (________25605), .Q
       (________24533));
  hi1s1 __90___511643(.DIN (________25360), .Q (____0___25593));
  nnd2s1 __9___511644(.DIN1 (_________36973), .DIN2
       (______________________21698), .Q (___9_0__25978));
  nor2s1 __9__9_511645(.DIN1 (________25571), .DIN2 (___0____23264), .Q
       (________24301));
  nnd2s1 __9__0_511646(.DIN1 (____0___23694), .DIN2 (____9___23592), .Q
       (_____0__25349));
  hi1s1 __90___511647(.DIN (_____9__25434), .Q (_____0__24905));
  nnd2s1 __9____511648(.DIN1 (________23766), .DIN2 (____0___23603), .Q
       (________24305));
  nnd2s1 __9____511649(.DIN1 (________23905), .DIN2
       (_____________________21691), .Q (________25553));
  nnd2s1 __90_9_511650(.DIN1 (____0___23598), .DIN2 (________22900), .Q
       (_____9___35559));
  nnd2s1 __90___511651(.DIN1 (___0____23249), .DIN2 (____9___23591), .Q
       (_________36854));
  nnd2s1 __9___511652(.DIN1 (____0___23694), .DIN2
       (_____________________21732), .Q (____9___24830));
  nnd2s1 __9____511653(.DIN1 (________23906), .DIN2
       (_____________________21736), .Q (________24658));
  nnd2s1 __9__0_511654(.DIN1 (________26450), .DIN2
       (____0_________________21724), .Q (________26604));
  hi1s1 __9____511655(.DIN (____9___23594), .Q (____9____38944));
  nnd2s1 __9____511656(.DIN1 (___9____25110), .DIN2 (___99___26049), .Q
       (________24698));
  nnd2s1 __9____511657(.DIN1 (________23755), .DIN2
       (_____________________21705), .Q (___00___25126));
  and2s1 __90___511658(.DIN1 (____0___23598), .DIN2 (________23515), .Q
       (_____0___37283));
  nnd2s1 __9____511659(.DIN1 (_____0__24487), .DIN2 (____0___23605), .Q
       (________24481));
  nnd2s1 __9____511660(.DIN1 (____0___23699), .DIN2 (____9___24066), .Q
       (___0____26109));
  nnd2s1 __9__511661(.DIN1 (___0____23238), .DIN2 (_____9__23076), .Q
       (___9_____39301));
  nnd2s1 __9____511662(.DIN1 (________23760), .DIN2 (____9___24066), .Q
       (___0____26089));
  nnd2s1 __9____511663(.DIN1 (________24691), .DIN2 (________22975), .Q
       (____9____38909));
  nor2s1 __9____511664(.DIN1 (___0____23227), .DIN2 (________23022), .Q
       (___9_____39384));
  nnd2s1 __9__0_511665(.DIN1 (________23847), .DIN2 (________23756), .Q
       (_____99__37662));
  nnd2s1 __9____511666(.DIN1 (______9__35039), .DIN2
       (_____________________21742), .Q (____0____35361));
  nnd2s1 __9____511667(.DIN1 (_____9__23094), .DIN2
       (____0________________21720), .Q (___99____39861));
  nor2s1 __9____511668(.DIN1 (_____0__23426), .DIN2 (___9_____39575),
       .Q (___0_90__40168));
  hi1s1 __9___511669(.DIN (___9_0__24080), .Q (____9___23590));
  nnd2s1 __909__511670(.DIN1 (____9___23588), .DIN2 (___9____24083), .Q
       (____9___23589));
  nor2s1 __909__511671(.DIN1 (________23894), .DIN2 (_____9__23586), .Q
       (____90__23587));
  nor2s1 __9____511672(.DIN1 (________22866), .DIN2 (___0____26125), .Q
       (________23585));
  nor2s1 __90___511673(.DIN1
       (______________________________________________21903), .DIN2
       (________23583), .Q (________23584));
  and2s1 __9__0_511674(.DIN1 (________23615), .DIN2 (___9____23165), .Q
       (________23582));
  nnd2s1 __9____511675(.DIN1 (________23580), .DIN2 (________22672), .Q
       (________23581));
  and2s1 __9___511676(.DIN1 (________23927), .DIN2
       (____0_________________21725), .Q (________23579));
  nor2s1 __909__511677(.DIN1 (____0___22846), .DIN2 (____9___24455), .Q
       (_____0__23578));
  or2s1 __9____511678(.DIN1 (________24632), .DIN2 (________24586), .Q
       (_____9__23577));
  nor2s1 __909__511679(.DIN1 (____0___22946), .DIN2 (___9_9__23154), .Q
       (________23576));
  nnd2s1 __9___511680(.DIN1 (________23012), .DIN2 (___0_9__24217), .Q
       (________23575));
  or2s1 __9____511681(.DIN1 (___0____23289), .DIN2 (________23573), .Q
       (________23574));
  nnd2s1 __9___511682(.DIN1 (_____0__23910), .DIN2 (___9____24134), .Q
       (________23572));
  xor2s1 __90___511683(.DIN1 (____9___22637), .DIN2 (_______22220), .Q
       (________23571));
  nnd2s1 __909__511684(.DIN1 (________22802), .DIN2 (____9___23970), .Q
       (________23570));
  nor2s1 __9____511685(.DIN1 (____0_________________21725), .DIN2
       (____09__25871), .Q (________23569));
  nnd2s1 __9099_511686(.DIN1 (________22764), .DIN2 (________22595), .Q
       (_____0__23568));
  and2s1 __9____511687(.DIN1 (________23566), .DIN2
       (_____________________21690), .Q (_____9__23567));
  and2s1 __9_0__511688(.DIN1 (_____9__23918), .DIN2 (___0_____40528),
       .Q (________23565));
  nnd2s1 __909__511689(.DIN1 (________23563), .DIN2 (____9___24455), .Q
       (________23564));
  nnd2s1 __909__511690(.DIN1 (________22914), .DIN2 (________22806), .Q
       (________23562));
  nor2s1 __90_9_511691(.DIN1 (___9____23166), .DIN2 (________23759), .Q
       (________23561));
  nor2s1 __9____511692(.DIN1 (________23860), .DIN2 (___9____26019), .Q
       (________23560));
  or2s1 __909__511693(.DIN1 (_____9__23842), .DIN2 (________23867), .Q
       (________23559));
  nnd2s1 __9___511694(.DIN1 (________23447), .DIN2
       (_____________________21678), .Q (_____0__23558));
  nor2s1 __9____511695(.DIN1 (___9___22195), .DIN2 (________23573), .Q
       (_____9__23557));
  or2s1 __909__511696(.DIN1 (________23555), .DIN2 (________23554), .Q
       (________23556));
  nnd2s1 __90__511697(.DIN1 (________23552), .DIN2 (____0___22941), .Q
       (________23553));
  nor2s1 __9090_511698(.DIN1 (________22994), .DIN2 (________24280), .Q
       (________23551));
  nnd2s1 __90___511699(.DIN1 (___9____23153), .DIN2
       (______________22104), .Q (________23550));
  nor2s1 __90__511700(.DIN1 (____0______________), .DIN2
       (___0____26125), .Q (________23549));
  nor2s1 __90___511701(.DIN1 (_____9__24635), .DIN2 (________23106), .Q
       (_____0__23548));
  nnd2s1 __90__511702(.DIN1 (___9_____39746), .DIN2
       (_____________________________________________21973), .Q
       (________23547));
  or2s1 __9____511703(.DIN1 (___9____23147), .DIN2 (____0___23410), .Q
       (________23546));
  nor2s1 __9____511704(.DIN1 (_____0__22529), .DIN2 (_____9___37943),
       .Q (________23545));
  or2s1 ___99__511705(.DIN1 (____0_0__38093), .DIN2 (_____9__22720), .Q
       (________23544));
  nor2s1 __9____511706(.DIN1 (________22677), .DIN2 (________22962), .Q
       (________23543));
  or2s1 __9_00_511707(.DIN1 (________23474), .DIN2 (________23541), .Q
       (________23542));
  nnd2s1 __90___511708(.DIN1 (_____9___38509), .DIN2
       (______________________________________0_______21892), .Q
       (_____0__23540));
  and2s1 __90__511709(.DIN1 (________23538), .DIN2 (___0_____40417), .Q
       (_____9__23539));
  nnd2s1 __90___511710(.DIN1 (_____9__23918), .DIN2
       (____________________________________________21762), .Q
       (________23537));
  or2s1 __9____511711(.DIN1 (________23535), .DIN2 (________23518), .Q
       (________23536));
  nor2s1 __909_511712(.DIN1 (____0____36220), .DIN2 (________23533), .Q
       (________23534));
  nor2s1 __9____511713(.DIN1 (________22408), .DIN2 (________23531), .Q
       (________23532));
  nnd2s1 __90___511714(.DIN1 (___9_____39746), .DIN2
       (_____________________________________________21974), .Q
       (_____0__23530));
  nor2s1 __909__511715(.DIN1 (________22884), .DIN2 (________23531), .Q
       (_____9__23529));
  nnd2s1 __9__511716(.DIN1 (________23437), .DIN2 (________22861), .Q
       (________23528));
  nor2s1 __90__511717(.DIN1 (_____________22101), .DIN2
       (___9_____39746), .Q (________23527));
  or2s1 __9__9_511718(.DIN1 (___99___26045), .DIN2 (________24791), .Q
       (________23526));
  and2s1 __9____511719(.DIN1 (________24690), .DIN2 (________23667), .Q
       (________23525));
  nnd2s1 __9_00_511720(.DIN1 (___9_9___39339), .DIN2 (inData[9]), .Q
       (________23524));
  nor2s1 __9__9_511721(.DIN1 (_____0__22499), .DIN2 (________22961), .Q
       (________23522));
  nor2s1 __9_0__511722(.DIN1 (________23914), .DIN2 (_____0__22671), .Q
       (_____0__23521));
  nor2s1 __9__511723(.DIN1 (________22757), .DIN2 (________22808), .Q
       (_____9__23520));
  and2s1 __9___511724(.DIN1 (________23518), .DIN2 (________23517), .Q
       (________23519));
  nnd2s1 __9_0_511725(.DIN1 (________23515), .DIN2 (________22954), .Q
       (________23516));
  xnr2s1 __9____511726(.DIN1 (__________), .DIN2 (________23513), .Q
       (________23514));
  nor2s1 __909__511727(.DIN1 (_____________________21670), .DIN2
       (____0___23503), .Q (________23512));
  nnd2s1 __9____511728(.DIN1 (____0___23509), .DIN2 (_______22255), .Q
       (_____0__23511));
  nnd2s1 __9____511729(.DIN1 (____0___23413), .DIN2 (____0___23509), .Q
       (____09__23510));
  nor2s1 __9____511730(.DIN1 (_____9__23376), .DIN2 (________23573), .Q
       (____0___23508));
  nnd2s1 __9099_511731(.DIN1 (________23422), .DIN2 (_______22174), .Q
       (____0___23507));
  nor2s1 __9__0_511732(.DIN1 (____0___22651), .DIN2 (____0___22749), .Q
       (____0___23506));
  or2s1 __9____511733(.DIN1 (____0___23504), .DIN2 (____0___23503), .Q
       (____0___23505));
  nnd2s1 __909__511734(.DIN1 (___9_9___39339), .DIN2 (______22119), .Q
       (____00__23502));
  and2s1 __9099_511735(.DIN1 (____9___23500), .DIN2 (________23752), .Q
       (____99__23501));
  nnd2s1 __9_00_511736(.DIN1 (________22767), .DIN2 (________22657), .Q
       (____9___23499));
  or2s1 __909__511737(.DIN1 (________23946), .DIN2 (________23027), .Q
       (____9___23498));
  nor2s1 __90999(.DIN1 (_____9__23104), .DIN2 (________22768), .Q
       (____9___23497));
  nnd2s1 __9_0__511738(.DIN1 (________22814), .DIN2 (inData[8]), .Q
       (____9___23496));
  and2s1 __9___511739(.DIN1 (________23580), .DIN2
       (_____________________21684), .Q (____9___23495));
  nor2s1 __9___511740(.DIN1 (________26530), .DIN2 (________23001), .Q
       (____9___23494));
  xor2s1 __9____511741(.DIN1 (___00____41368), .DIN2 (_____9__23492),
       .Q (____90__23493));
  nor2s1 __9_0__511742(.DIN1 (_______22279), .DIN2 (________23490), .Q
       (________23491));
  nor2s1 __9_0_511743(.DIN1 (___9_9__23181), .DIN2 (________23531), .Q
       (________23489));
  nor2s1 __9____511744(.DIN1 (________23469), .DIN2 (____0___22947), .Q
       (________23488));
  nnd2s1 __9____511745(.DIN1 (________23518), .DIN2 (____9___22933), .Q
       (________23487));
  and2s1 __9_0__511746(.DIN1 (________23901), .DIN2 (________23485), .Q
       (________23486));
  nor2s1 __909__511747(.DIN1 (____0___22557), .DIN2 (____0___22945), .Q
       (________23484));
  and2s1 __9090_511748(.DIN1 (_____9__23482), .DIN2 (________23481), .Q
       (_____0__23483));
  or2s1 __9___511749(.DIN1 (________23017), .DIN2 (________24470), .Q
       (________23480));
  nnd2s1 __9_0__511750(.DIN1 (_____0__22889), .DIN2 (________22813), .Q
       (________23479));
  nnd2s1 __9_0__511751(.DIN1 (________23477), .DIN2 (________23476), .Q
       (________23478));
  nnd2s1 __909__511752(.DIN1 (________23518), .DIN2 (________23474), .Q
       (________23475));
  nor2s1 __909__511753(.DIN1 (___9____23168), .DIN2 (________23442), .Q
       (_____0__23473));
  or2s1 __9____511754(.DIN1 (________25644), .DIN2 (________24632), .Q
       (_____9__23472));
  nnd2s1 __909__511755(.DIN1 (________24797), .DIN2 (________22896), .Q
       (________23471));
  nor2s1 __9____511756(.DIN1 (________23469), .DIN2 (_____0__22969), .Q
       (________23470));
  nor2s1 __909_511757(.DIN1 (_____0__24393), .DIN2 (____00__24267), .Q
       (________23468));
  nor2s1 __90_9_511758(.DIN1 (____9), .DIN2 (_________38249), .Q
       (________23467));
  nnd2s1 __9__0_511759(.DIN1 (________23430), .DIN2 (______22154), .Q
       (________23466));
  and2s1 __90___511760(.DIN1 (___9_9___39339), .DIN2 (___0_____40502),
       .Q (________23465));
  or2s1 __90___511761(.DIN1 (____0________________21664), .DIN2
       (___9____24081), .Q (_____0__23464));
  nor2s1 __909__511762(.DIN1 (____0___22649), .DIN2 (________22916), .Q
       (_____9__23463));
  nor2s1 __9_000(.DIN1 (________22877), .DIN2 (________23461), .Q
       (________23462));
  hi1s1 __90___511763(.DIN (___9____24156), .Q (________23460));
  and2s1 __90___511764(.DIN1 (_____0__22791), .DIN2
       (____0____________0_), .Q (________23459));
  and2s1 __90___511765(.DIN1 (________23434), .DIN2
       (_____________________21670), .Q (________23458));
  nnd2s1 __909__511766(.DIN1 (______0__35181), .DIN2 (________22586),
       .Q (________23457));
  nor2s1 __90___511767(.DIN1 (____0_________________21726), .DIN2
       (_____9__23018), .Q (________23456));
  hi1s1 __9___511768(.DIN (________24700), .Q (________24291));
  hi1s1 __9____511769(.DIN (________23455), .Q (________24386));
  nnd2s1 __9___511770(.DIN1 (_____0__23454), .DIN2 (________25756), .Q
       (________23960));
  nnd2s1 __9_0__511771(.DIN1 (________23347), .DIN2 (_____9__22878), .Q
       (________24026));
  nor2s1 __9___511772(.DIN1 (________23014), .DIN2 (_____9__23453), .Q
       (________25357));
  nor2s1 __9_0__511773(.DIN1 (___0___22201), .DIN2 (________23452), .Q
       (____9___23685));
  nor2s1 __9__0_511774(.DIN1 (________22986), .DIN2 (____0___22748), .Q
       (___0____24235));
  nor2s1 __9_0__511775(.DIN1 (____90__26673), .DIN2 (________23451), .Q
       (_____0__23607));
  nnd2s1 __9_0__511776(.DIN1 (________22787), .DIN2 (____00__23407), .Q
       (________23902));
  nor2s1 __9___511777(.DIN1 (____0___23600), .DIN2 (________23715), .Q
       (________23670));
  nnd2s1 __9____511778(.DIN1 (________23450), .DIN2 (______22153), .Q
       (________23924));
  nor2s1 __9_0__511779(.DIN1 (_____________________21669), .DIN2
       (________22811), .Q (________26199));
  nor2s1 __9_09_511780(.DIN1 (________23449), .DIN2 (___0____23265), .Q
       (________23765));
  nor2s1 __9_0__511781(.DIN1 (_____________________21671), .DIN2
       (____0___23503), .Q (________23840));
  nnd2s1 __9____511782(.DIN1 (________23533), .DIN2 (_________37722),
       .Q (________23745));
  nor2s1 __9_0__511783(.DIN1 (________22880), .DIN2 (___9____23160), .Q
       (________23812));
  nor2s1 __9____511784(.DIN1 (____0________________21667), .DIN2
       (________23418), .Q (________23761));
  hi1s1 __9____511785(.DIN (________23448), .Q (________23935));
  nnd2s1 __9___511786(.DIN1 (________23447), .DIN2 (____0___23697), .Q
       (___0____24189));
  nor2s1 __9_0_511787(.DIN1 (________22421), .DIN2 (________22812), .Q
       (___9____24131));
  nnd2s1 __9_0__511788(.DIN1 (________23443), .DIN2
       (_____________________21682), .Q (________23917));
  hi1s1 __9__0_511789(.DIN (________23446), .Q (________26257));
  nnd2s1 __9___511790(.DIN1 (________26575), .DIN2 (___0____23239), .Q
       (________23828));
  nor2s1 __9_0_511791(.DIN1 (_____0__23445), .DIN2 (___0____23257), .Q
       (________23703));
  nnd2s1 __9____511792(.DIN1 (________23421), .DIN2
       (_____________________21691), .Q (________23750));
  nor2s1 __9_0__511793(.DIN1 (______________________21698), .DIN2
       (______0__38256), .Q (________23762));
  nor2s1 __9_0__511794(.DIN1 (________24475), .DIN2 (________22901), .Q
       (____0___26501));
  nnd2s1 __9_0__511795(.DIN1 (____0___22940), .DIN2 (_____9__23444), .Q
       (________26577));
  nnd2s1 __9____511796(.DIN1 (________23443), .DIN2 (______22153), .Q
       (____9___24068));
  nor2s1 __9_0__511797(.DIN1 (____0___26590), .DIN2 (________22823), .Q
       (________25930));
  hi1s1 __9____511798(.DIN (_____0__26247), .Q (________25634));
  nnd2s1 __9_0_511799(.DIN1 (________23583), .DIN2 (________22867), .Q
       (____99__27741));
  nnd2s1 __9___511800(.DIN1 (________23442), .DIN2
       (____0_______________), .Q (________26171));
  nor2s1 __9____511801(.DIN1 (_____________________21710), .DIN2
       (________22784), .Q (________23931));
  nor2s1 __9____511802(.DIN1 (_______22286), .DIN2 (________22789), .Q
       (___0____24251));
  nnd2s1 __9_0_511803(.DIN1 (________23441), .DIN2 (____00__23597), .Q
       (___9____24111));
  nor2s1 __9__0_511804(.DIN1 (________24602), .DIN2 (________23439), .Q
       (___0____24219));
  nnd2s1 __9____511805(.DIN1 (________23440), .DIN2
       (_____________________21705), .Q (____9___23968));
  nor2s1 __9_0__511806(.DIN1 (________23989), .DIN2 (________23563), .Q
       (___90___24074));
  or2s1 __9_0__511807(.DIN1 (________23715), .DIN2 (________25327), .Q
       (____9___24064));
  nor2s1 __9____511808(.DIN1 (_____________________21709), .DIN2
       (________23439), .Q (________23921));
  nor2s1 __9_099(.DIN1
       (_____________________________________________21841), .DIN2
       (________23533), .Q (___09___24265));
  nnd2s1 __90__511809(.DIN1 (____9___22735), .DIN2 (________23662), .Q
       (_________34775));
  hi1s1 __90_9_511810(.DIN (________24289), .Q (___0____24220));
  and2s1 __9_0__511811(.DIN1 (____9___24061), .DIN2
       (_____________________21691), .Q (_____0__24618));
  nor2s1 __9_0__511812(.DIN1 (___0_0___40567), .DIN2 (_____9___37943),
       .Q (________24044));
  nor2s1 __9____511813(.DIN1 (________26431), .DIN2 (_____9__23586), .Q
       (________24395));
  nnd2s1 __9____511814(.DIN1 (________23427), .DIN2
       (_____________________21709), .Q (____0___23977));
  nor2s1 __9__0_511815(.DIN1 (________23438), .DIN2 (________22923), .Q
       (________24488));
  nnd2s1 __9___511816(.DIN1 (________23437), .DIN2
       (_____________________21745), .Q (___9_9__24108));
  or2s1 __9__0_511817(.DIN1 (____00__23597), .DIN2 (_____0__23436), .Q
       (___0____24230));
  and2s1 __9____511818(.DIN1 (_____9__23435), .DIN2
       (____0________________21716), .Q (________23915));
  nor2s1 __9__0_511819(.DIN1 (_____________________21682), .DIN2
       (________23867), .Q (___90___24075));
  nnd2s1 __9____511820(.DIN1 (____0___24269), .DIN2 (________25564), .Q
       (_____9__23991));
  nnd2s1 __9__0_511821(.DIN1 (________23533), .DIN2 (________22716), .Q
       (___9____24127));
  and2s1 __9____511822(.DIN1 (________23434), .DIN2 (___9____23156), .Q
       (___9____24144));
  nnd2s1 __9____511823(.DIN1 (____9___24061), .DIN2 (________23989), .Q
       (________25440));
  hi1s1 __9____511824(.DIN (________23433), .Q (____9___24067));
  hi1s1 __9____511825(.DIN (________23432), .Q (_____0__24895));
  nnd2s1 __9____511826(.DIN1 (________23431), .DIN2 (________23989), .Q
       (___9_0__25068));
  nnd2s1 __9____511827(.DIN1 (________23002), .DIN2
       (____0_______________), .Q (____9___27649));
  nnd2s1 __9____511828(.DIN1 (________23430), .DIN2 (____9___24066), .Q
       (___90___24078));
  nnd2s1 __9__0_511829(.DIN1 (________25270), .DIN2
       (_____________________21683), .Q (_____9__25378));
  hi1s1 __9____511830(.DIN (____9___24065), .Q (___0_9__25164));
  nor2s1 __9__511831(.DIN1 (____0________________21720), .DIN2
       (___0____23259), .Q (_____9__24296));
  nor2s1 __9___511832(.DIN1 (________26431), .DIN2 (________22967), .Q
       (________23925));
  hi1s1 __9____511833(.DIN (________23429), .Q (_____9__24059));
  nnd2s1 __9____511834(.DIN1 (________23428), .DIN2
       (____0________________21716), .Q (___9____24146));
  nnd2s1 __9___511835(.DIN1 (________23427), .DIN2 (________24602), .Q
       (________24010));
  or2s1 __9____511836(.DIN1 (_____________________21691), .DIN2
       (________23563), .Q (_____0__24420));
  and2s1 __9___511837(.DIN1 (_____0__23426), .DIN2
       (____0________________21716), .Q (___9____24120));
  hi1s1 __9__9_511838(.DIN (________24734), .Q (___0____26099));
  nnd2s1 __9____511839(.DIN1 (___0_9__23262), .DIN2
       (____0________________21667), .Q (___909__24079));
  nor2s1 __9____511840(.DIN1 (________23959), .DIN2 (_____9__23425), .Q
       (____99__24745));
  nor2s1 __9___511841(.DIN1 (____0________________21720), .DIN2
       (________23424), .Q (________25640));
  nor2s1 __9___511842(.DIN1 (________23423), .DIN2 (________23441), .Q
       (___0____24191));
  nnd2s1 __9___511843(.DIN1 (________23422), .DIN2 (________22497), .Q
       (___0____24201));
  nnd2s1 __9____511844(.DIN1 (____0___23415), .DIN2 (___0____23252), .Q
       (_____9__25434));
  nnd2s1 __9____511845(.DIN1 (________22826), .DIN2
       (____0_______________), .Q (___9____24082));
  hi1s1 __9____511846(.DIN (____9___24742), .Q (________25550));
  nnd2s1 __9____511847(.DIN1 (________23421), .DIN2 (________23989), .Q
       (___9_9__25057));
  hi1s1 __9____511848(.DIN (________23420), .Q (________25294));
  hi1s1 __9____511849(.DIN (________23419), .Q (____9___24928));
  nnd2s1 __9__0_511850(.DIN1 (________23418), .DIN2 (________22683), .Q
       (_________38675));
  nnd2s1 __9___511851(.DIN1 (________23440), .DIN2 (________23754), .Q
       (________25336));
  hi1s1 __90___511852(.DIN (_____0__23417), .Q (___9____25983));
  nor2s1 __9____511853(.DIN1 (____9___23970), .DIN2 (_____9__25927), .Q
       (________25923));
  nnd2s1 __9____511854(.DIN1 (________24415), .DIN2 (________23959), .Q
       (________25257));
  nor2s1 __9____511855(.DIN1 (____09__23416), .DIN2 (________22805), .Q
       (_________38395));
  nnd2s1 __9____511856(.DIN1 (________23430), .DIN2
       (_____________________21732), .Q (____0___26594));
  nnd2s1 __9____511857(.DIN1 (____0___23415), .DIN2
       (_____________________21683), .Q (________25391));
  nnd2s1 __9__0_511858(.DIN1 (___0_0__23263), .DIN2 (___9____23164), .Q
       (_________34647));
  nor2s1 __9____511859(.DIN1 (_____9__22760), .DIN2 (________23554), .Q
       (_____9___35467));
  nor2s1 __9___511860(.DIN1 (_____9__22819), .DIN2 (________23427), .Q
       (_________38306));
  nnd2s1 __9____511861(.DIN1 (_____0__23426), .DIN2 (____00__23597), .Q
       (___9_9__25114));
  nnd2s1 __9____511862(.DIN1 (________22982), .DIN2 (____0___23414), .Q
       (______9__35170));
  and2s1 __9___511863(.DIN1 (_____9__23425), .DIN2 (________23726), .Q
       (___90____39040));
  nnd2s1 __9__9_511864(.DIN1 (____0___23413), .DIN2
       (_____________________21683), .Q (________25360));
  nor2s1 __9____511865(.DIN1 (____0___23412), .DIN2 (____0____33482),
       .Q (______9__33955));
  nor2s1 __9____511866(.DIN1 (________22728), .DIN2 (___9____23143), .Q
       (___9_____39183));
  nnd2s1 __9__9_511867(.DIN1 (_________38543), .DIN2 (________22580),
       .Q (_________38262));
  or2s1 __9_0__511868(.DIN1 (____0________________21717), .DIN2
       (____0___23410), .Q (____0___23411));
  xor2s1 __90___511869(.DIN1 (________22658), .DIN2 (___0____22322), .Q
       (____0___23409));
  nor2s1 __909__511870(.DIN1 (____00__23407), .DIN2 (____99__23406), .Q
       (____0___23408));
  nor2s1 __9_00_511871(.DIN1 (___0____23292), .DIN2 (________23451), .Q
       (____9___23405));
  nor2s1 __909__511872(.DIN1 (________22922), .DIN2 (________22807), .Q
       (____9___23404));
  nnd2s1 __9____511873(.DIN1 (________23518), .DIN2 (___99_), .Q
       (____9___23403));
  or2s1 __9____511874(.DIN1 (_______________22077), .DIN2
       (_________38583), .Q (____9___23402));
  and2s1 __909__511875(.DIN1 (____9___23400), .DIN2
       (_____________________21692), .Q (____9___23401));
  and2s1 __909_511876(.DIN1 (______9__38496), .DIN2
       (______________________________________________21945), .Q
       (____9___23399));
  or2s1 __90_9_511877(.DIN1 (____0________________21664), .DIN2
       (________24727), .Q (____9___23398));
  or2s1 __909__511878(.DIN1 (____0___22742), .DIN2 (_____9__22780), .Q
       (____90__23397));
  nnd2s1 __909_511879(.DIN1 (_____9__22968), .DIN2 (________22521), .Q
       (_____9__23396));
  nnd2s1 __90___511880(.DIN1 (________22912), .DIN2 (inData[14]), .Q
       (________23395));
  hi1s1 __9___511881(.DIN (________24757), .Q (________23394));
  nnd2s1 __9____511882(.DIN1 (___9_9___39339), .DIN2 (___0____22309),
       .Q (________23393));
  or2s1 __9___511883(.DIN1 (________23391), .DIN2 (___9____23157), .Q
       (________23392));
  or2s1 __9_0__511884(.DIN1 (____9___22734), .DIN2 (________23946), .Q
       (________23390));
  nor2s1 __909__511885(.DIN1 (____0___26590), .DIN2 (___9____24084), .Q
       (________23389));
  or2s1 __909__511886(.DIN1 (________23989), .DIN2 (________22886), .Q
       (________23388));
  nnd2s1 __90___511887(.DIN1 (________25944), .DIN2
       (____0________________21664), .Q (_____0__23387));
  nnd2s1 ___99_511888(.DIN1 (_____9__22790), .DIN2 (inData[24]), .Q
       (_____9__23386));
  nnd2s1 __909__511889(.DIN1 (________23384), .DIN2 (________23383), .Q
       (________23385));
  nor2s1 __909__511890(.DIN1 (_____________________21744), .DIN2
       (_____0__22761), .Q (________23382));
  xor2s1 __90___511891(.DIN1 (____09__22653), .DIN2 (_______22222), .Q
       (________23381));
  nnd2s1 __90___511892(.DIN1 (_____0__22959), .DIN2 (inData[12]), .Q
       (________23380));
  nor2s1 __90___511893(.DIN1 (_____0__22979), .DIN2 (_________37744),
       .Q (________23379));
  nnd2s1 __90_9_511894(.DIN1 (________23351), .DIN2 (________22817), .Q
       (________23378));
  nor2s1 __9____511895(.DIN1 (_____9__23376), .DIN2 (________23325), .Q
       (_____0__23377));
  nnd2s1 ___9__511896(.DIN1 (________22910), .DIN2 (inData[24]), .Q
       (________23375));
  hi1s1 __90_9_511897(.DIN (________24311), .Q (________23374));
  or2s1 __90___511898(.DIN1 (________23372), .DIN2 (________22920), .Q
       (________23373));
  nnd2s1 ___990_511899(.DIN1 (________22773), .DIN2 (inData[30]), .Q
       (________23371));
  and2s1 __9____511900(.DIN1 (________24313), .DIN2
       (_____________________21705), .Q (________23370));
  or2s1 __9____511901(.DIN1 (______________________21698), .DIN2
       (________23485), .Q (________23369));
  and2s1 __9____511902(.DIN1 (________23327), .DIN2 (________23580), .Q
       (_____0__23368));
  nnd2s1 __90___511903(.DIN1 (___0____23271), .DIN2 (____9___23592), .Q
       (________23367));
  and2s1 __90___511904(.DIN1 (________22882), .DIN2
       (____________________), .Q (________23366));
  and2s1 __9___511905(.DIN1 (________23518), .DIN2 (________23364), .Q
       (________23365));
  nor2s1 __90_9_511906(.DIN1 (________23362), .DIN2 (________22793), .Q
       (________23363));
  nnd2s1 __90_9_511907(.DIN1 (________23360), .DIN2 (________22769), .Q
       (________23361));
  or2s1 __9090_511908(.DIN1 (__99____30501), .DIN2 (________22797), .Q
       (_____0__23359));
  nnd2s1 __909__511909(.DIN1 (________22997), .DIN2 (___0____26120), .Q
       (_____9__23358));
  nnd2s1 __909__511910(.DIN1 (________23434), .DIN2 (________23356), .Q
       (________23357));
  nnd2s1 __909__511911(.DIN1 (________23538), .DIN2 (___0_____40611),
       .Q (________23355));
  and2s1 __9__0_511912(.DIN1 (____0___23413), .DIN2
       (_____________________21682), .Q (________23354));
  nnd2s1 __909_511913(.DIN1 (___9_9___39339), .DIN2 (inData[13]), .Q
       (________23353));
  nor2s1 __909_511914(.DIN1 (_____________________21691), .DIN2
       (________23351), .Q (________23352));
  and2s1 __909__511915(.DIN1 (________22803), .DIN2 (___909), .Q
       (________23350));
  or2s1 __909__511916(.DIN1 (_____________________21682), .DIN2
       (____09__22750), .Q (_____0__23349));
  nnd2s1 __909__511917(.DIN1 (________23347), .DIN2 (___0____23269), .Q
       (_____9__23348));
  nor2s1 __909__511918(.DIN1 (________22915), .DIN2 (________23914), .Q
       (________23346));
  nnd2s1 __909__511919(.DIN1 (________22778), .DIN2 (____9___23970), .Q
       (________23345));
  nnd2s1 __909__511920(.DIN1 (___9_9___39339), .DIN2 (____9___23131),
       .Q (________23344));
  nnd2s1 __909__511921(.DIN1 (________23347), .DIN2 (________22775), .Q
       (________23343));
  nnd2s1 __909__511922(.DIN1 (________22758), .DIN2 (________23517), .Q
       (________23342));
  nor2s1 __9__9_511923(.DIN1 (________22862), .DIN2 (________24341), .Q
       (________23341));
  nnd2s1 __9_0_511924(.DIN1 (________24398), .DIN2 (________23752), .Q
       (________23340));
  hi1s1 __9____511925(.DIN (________24731), .Q (_____0__23339));
  nor2s1 __909__511926(.DIN1 (________23989), .DIN2 (________22785), .Q
       (_____9__23338));
  and2s1 __9_0_511927(.DIN1 (________23423), .DIN2
       (__________________________________________0___21919), .Q
       (________23337));
  nor2s1 __9_0__511928(.DIN1 (____00__23039), .DIN2 (________23335), .Q
       (________23336));
  nor2s1 __9__511929(.DIN1 (___090), .DIN2 (________23533), .Q
       (________23334));
  nnd2s1 __9____511930(.DIN1 (_____9__25927), .DIN2 (________23000), .Q
       (________23333));
  nnd2s1 __9___511931(.DIN1 (________23437), .DIN2 (________22820), .Q
       (________23332));
  nor2s1 __909__511932(.DIN1 (________23330), .DIN2 (________23927), .Q
       (________23331));
  nnd2s1 ___999_511933(.DIN1 (________22911), .DIN2 (inData[26]), .Q
       (_____0__23329));
  nor2s1 __9__9_511934(.DIN1 (________25270), .DIN2 (________23327), .Q
       (_____9__23328));
  or2s1 __9___511935(.DIN1 (__________________0___21686), .DIN2
       (________23325), .Q (________23326));
  nor2s1 __9___511936(.DIN1 (____9___22443), .DIN2 (_________37744), .Q
       (________23324));
  nnd2s1 __909__511937(.DIN1 (________23554), .DIN2 (________23555), .Q
       (________23323));
  nnd2s1 __909__511938(.DIN1 (________22774), .DIN2 (inData[6]), .Q
       (________23322));
  nor2s1 __9___511939(.DIN1 (___9_0__23155), .DIN2 (___90___25034), .Q
       (________23321));
  nor2s1 __9___511940(.DIN1 (________24475), .DIN2 (________24797), .Q
       (________23320));
  nor2s1 __9__9_511941(.DIN1 (___99____39814), .DIN2 (____9___22936),
       .Q (_____0__23319));
  nnd2s1 __909__511942(.DIN1 (________23441), .DIN2
       (_____________22102), .Q (____09__23318));
  nnd2s1 __9____511943(.DIN1 (____0___23316), .DIN2 (____0___23315), .Q
       (____0___23317));
  hi1s1 __90___511944(.DIN (________25829), .Q (____0___23314));
  nnd2s1 __9__511945(.DIN1 (____00__22741), .DIN2 (___9____23170), .Q
       (____0___23313));
  and2s1 __9____511946(.DIN1 (____0___23410), .DIN2 (____0___23311), .Q
       (____0___23312));
  and2s1 __9__9_511947(.DIN1 (________23566), .DIN2 (_____9__23444), .Q
       (____0___23310));
  nor2s1 __9__0_511948(.DIN1 (________22871), .DIN2 (________23901), .Q
       (___09___23308));
  nor2s1 __9____511949(.DIN1 (________22719), .DIN2 (___09___23306), .Q
       (___09___23307));
  nnd2s1 __9____511950(.DIN1 (_________35663), .DIN2 (_________34167),
       .Q (___09___23305));
  nor2s1 __9____511951(.DIN1 (________22664), .DIN2 (________22971), .Q
       (___09___23304));
  nnd2s1 __9___511952(.DIN1 (________26576), .DIN2 (____9___24738), .Q
       (___09___23303));
  xnr2s1 __9____511953(.DIN1 (_________22041), .DIN2 (___090__23301),
       .Q (___09___23302));
  nor2s1 __9____511954(.DIN1 (____9___22733), .DIN2 (___0____23299), .Q
       (___0_9__23300));
  or2s1 __9____511955(.DIN1 (___0____23297), .DIN2 (____0____33482), .Q
       (___0____23298));
  nnd2s1 __9____511956(.DIN1 (________23441), .DIN2 (________22438), .Q
       (___0____23296));
  and2s1 __9__9_511957(.DIN1 (________23327), .DIN2 (________23325), .Q
       (___0____23295));
  nnd2s1 __9____511958(.DIN1 (____9___22736), .DIN2 (___99___23210), .Q
       (___0____23294));
  and2s1 __9__9_511959(.DIN1 (_____0__22801), .DIN2 (___0____23292), .Q
       (___0____23293));
  nor2s1 __9__9_511960(.DIN1 (________24013), .DIN2 (_____0__24316), .Q
       (___0_0__23291));
  or2s1 __9____511961(.DIN1 (___0____23289), .DIN2 (________23325), .Q
       (___0_9__23290));
  and2s1 __909__511962(.DIN1 (______9__38496), .DIN2
       (______________________________________________21946), .Q
       (___0____23288));
  and2s1 __9____511963(.DIN1 (___0_0__24248), .DIN2 (________23911), .Q
       (___0____23287));
  or2s1 __9____511964(.DIN1 (____9___22834), .DIN2 (____0___23413), .Q
       (___0____23286));
  and2s1 __9___511965(.DIN1 (___9_9___39339), .DIN2 (________22482), .Q
       (___0____23285));
  xnr2s1 __90___511966(.DIN1
       (____________________________________________21792), .DIN2
       (_____9___38412), .Q (___0____23284));
  nnd2s1 __909__511967(.DIN1 (____90__22829), .DIN2 (____0___26590), .Q
       (___0____23283));
  nnd2s1 __9____511968(.DIN1 (___0____26064), .DIN2 (____9___23970), .Q
       (___0____23282));
  hi1s1 __9____511969(.DIN (________23756), .Q (___0_0__23281));
  hi1s1 __9____511970(.DIN (________26450), .Q (___0____23280));
  nnd2s1 __9____511971(.DIN1 (___0____23299), .DIN2 (________23517), .Q
       (___0____23279));
  nnd2s1 __9__0_511972(.DIN1 (____0___23509), .DIN2 (___0____23276), .Q
       (___0____23277));
  nor2s1 __9____511973(.DIN1 (_____9__22770), .DIN2 (___90___25034), .Q
       (___0____23275));
  nnd2s1 __9____511974(.DIN1 (____90__22731), .DIN2 (_____9__23900), .Q
       (___0____23274));
  nnd2s1 __9__0_511975(.DIN1 (________25270), .DIN2 (______22153), .Q
       (___0_0__23273));
  nnd2s1 __9__0_511976(.DIN1 (________23580), .DIN2 (____9___22635), .Q
       (___0_9__23272));
  and2s1 __9____511977(.DIN1 (________23430), .DIN2 (____9___23592), .Q
       (_____9__24306));
  hi1s1 __9____511978(.DIN (___0____25171), .Q (________24285));
  nor2s1 __9__511979(.DIN1 (____9___24066), .DIN2 (___0____23271), .Q
       (________23746));
  hi1s1 __9__0_511980(.DIN (___0____23270), .Q (________24046));
  hi1s1 __9____511981(.DIN (____9_9__38931), .Q (_________32987));
  nnd2s1 __9_0__511982(.DIN1 (________22718), .DIN2 (______22153), .Q
       (________23923));
  nnd2s1 __9____511983(.DIN1 (________22905), .DIN2 (___0____23269), .Q
       (________24058));
  nnd2s1 __9_09_511984(.DIN1 (_____0__23436), .DIN2 (________22856), .Q
       (____09__23606));
  hi1s1 __90_511985(.DIN (___0____25143), .Q (________23912));
  nor2s1 __9_0__511986(.DIN1 (___0____23268), .DIN2 (___0____26067), .Q
       (____9___23687));
  hi1s1 __9____511987(.DIN (________24324), .Q (___00___24176));
  nor2s1 __9____511988(.DIN1 (____9___24066), .DIN2 (___0____23267), .Q
       (________23608));
  nor2s1 __9____511989(.DIN1 (__________________0___21750), .DIN2
       (________22794), .Q (________24278));
  hi1s1 __90_0_511990(.DIN (________23764), .Q (_____0__23982));
  nor2s1 __9__0_511991(.DIN1 (_____________________21669), .DIN2
       (______0__34897), .Q (_____0__23758));
  nnd2s1 __9_0__511992(.DIN1 (___0____23236), .DIN2 (________23573), .Q
       (________24049));
  and2s1 __9____511993(.DIN1 (_____9__23918), .DIN2 (inData[22]), .Q
       (___9____24102));
  and2s1 __9____511994(.DIN1 (_________38543), .DIN2 (________22894),
       .Q (___00___26056));
  hi1s1 __9____511995(.DIN (________24594), .Q (____9___23966));
  nnd2s1 __9____511996(.DIN1 (________24699), .DIN2 (___0____23260), .Q
       (____0___23795));
  and2s1 __9_0__511997(.DIN1 (________23451), .DIN2
       (______________________21753), .Q (________23913));
  nnd2s1 __9_0_511998(.DIN1 (_____0__24411), .DIN2
       (_____________________21681), .Q (___0_9__24197));
  nor2s1 __9____511999(.DIN1 (___9____23177), .DIN2 (_____9__25555), .Q
       (____00__23788));
  hi1s1 __90___512000(.DIN (___0____23266), .Q (________24898));
  nor2s1 __9_0__512001(.DIN1 (___0____22318), .DIN2 (________22983), .Q
       (________24003));
  nnd2s1 __9_09_512002(.DIN1 (________23932), .DIN2
       (____0________________21720), .Q (________23763));
  nnd2s1 __9____512003(.DIN1 (_____9__25927), .DIN2 (________23959), .Q
       (___9____24087));
  and2s1 __9____512004(.DIN1 (____0___23410), .DIN2 (_____0__23095), .Q
       (________23934));
  nor2s1 __9____512005(.DIN1 (______________________21699), .DIN2
       (___0____23265), .Q (____9___23595));
  nnd2s1 __9____512006(.DIN1 (____90__25489), .DIN2 (________23989), .Q
       (_____9__23747));
  or2s1 __9_0__512007(.DIN1 (____0_________________21725), .DIN2
       (_____9__22898), .Q (_____0__24012));
  nnd2s1 __9____512008(.DIN1 (_____0__22751), .DIN2 (______22153), .Q
       (___99___24159));
  nor2s1 __9___512009(.DIN1 (____0________________21716), .DIN2
       (______9__38496), .Q (___9____24095));
  hi1s1 __9____512010(.DIN (___0____23264), .Q (____9___23963));
  nnd2s1 __9____512011(.DIN1 (________24351), .DIN2
       (_____________________21691), .Q (_____9__25019));
  nor2s1 __9____512012(.DIN1 (____0___23599), .DIN2 (___0_0__23263), .Q
       (____0___23980));
  and2s1 __9____512013(.DIN1 (___9____24134), .DIN2 (______22153), .Q
       (_____9__23909));
  nnd2s1 __9____512014(.DIN1 (___0____23261), .DIN2 (________22585), .Q
       (____9___23594));
  hi1s1 __90___512015(.DIN (________25735), .Q (________24896));
  nor2s1 __9____512016(.DIN1 (____0________________21720), .DIN2
       (_____0__25319), .Q (___9____24096));
  hi1s1 __9____512017(.DIN (____0____38106), .Q (_____0___34938));
  nnd2s1 __9____512018(.DIN1 (________23423), .DIN2 (____00__23597), .Q
       (________24995));
  nnd2s1 __9___512019(.DIN1 (________24415), .DIN2
       (____0________________21716), .Q (___0____24195));
  nnd2s1 __9_0__512020(.DIN1 (___0_9__23262), .DIN2 (____0___23599), .Q
       (___90___24077));
  nor2s1 __9__0_512021(.DIN1 (_____0__23445), .DIN2 (___0____23261), .Q
       (_____0__24478));
  nnd2s1 __9____512022(.DIN1 (____0___22744), .DIN2 (________22965), .Q
       (___0_9__25144));
  nor2s1 __9____512023(.DIN1 (____0___23311), .DIN2 (_____9___38509),
       .Q (___0____24179));
  nor2s1 __9_09_512024(.DIN1 (_____________________21689), .DIN2
       (________23108), .Q (_____0__25566));
  nor2s1 __9____512025(.DIN1 (___0____23256), .DIN2 (_____9__23482), .Q
       (________25750));
  nnd2s1 __9__512026(.DIN1 (___0____23260), .DIN2 (____0___23603), .Q
       (____99__24069));
  hi1s1 __9____512027(.DIN (________23866), .Q (_____0__24726));
  nor2s1 __9__0_512028(.DIN1 (________23959), .DIN2 (___0____23259), .Q
       (________24433));
  nnd2s1 __9__9_512029(.DIN1 (________23023), .DIN2 (________25605), .Q
       (_____9__24525));
  nor2s1 __9__0_512030(.DIN1 (___0____25163), .DIN2 (___0____26067), .Q
       (________24034));
  hi1s1 __90___512031(.DIN (_____0__23919), .Q (___9____24117));
  nor2s1 __9____512032(.DIN1 (________23989), .DIN2 (___0____23254), .Q
       (_____9__24675));
  nor2s1 __9_99_(.DIN1 (________22627), .DIN2 (________23325), .Q
       (____9___25023));
  hi1s1 __9___512033(.DIN (___0____23258), .Q (________24476));
  hi1s1 __9____512034(.DIN (___9____24085), .Q (_____0__24775));
  nor2s1 __9____512035(.DIN1 (______________________21698), .DIN2
       (___0____23257), .Q (________24875));
  nnd2s1 __9____512036(.DIN1 (________25270), .DIN2 (________23580), .Q
       (___90___24071));
  nor2s1 __9____512037(.DIN1 (___0____23256), .DIN2 (________22763), .Q
       (___09___24263));
  nor2s1 __9__9_512038(.DIN1 (_____________________21736), .DIN2
       (_________37722), .Q (_____9__23928));
  nor2s1 __9____512039(.DIN1 (_____________________21683), .DIN2
       (________22883), .Q (________24909));
  nnd2s1 __9____512040(.DIN1 (____9___22937), .DIN2 (________23021), .Q
       (________24323));
  nor2s1 __9__512041(.DIN1 (____0________________21714), .DIN2
       (___9__9__39659), .Q (___00___24169));
  hi1s1 __9__9_512042(.DIN (____0___24463), .Q (________25335));
  hi1s1 __9__0_512043(.DIN (___0____26083), .Q (________26267));
  hi1s1 __9__0_512044(.DIN (________25320), .Q (________24517));
  nor2s1 __9___512045(.DIN1 (____0________________21720), .DIN2
       (_____9__23425), .Q (___9____24136));
  nor2s1 __9___512046(.DIN1 (____9___23970), .DIN2 (_____0__23454), .Q
       (_____0__25479));
  hi1s1 __9____512047(.DIN (___0____23255), .Q (________24710));
  hi1s1 __9___512048(.DIN (_____9__24715), .Q (___0____25169));
  nnd2s1 __9____512049(.DIN1 (________23441), .DIN2
       (____0________________21716), .Q (____0___25590));
  or2s1 __9____512050(.DIN1 (_____________________21742), .DIN2
       (___0____23268), .Q (___0____25204));
  hi1s1 __90__512051(.DIN (_____0__23646), .Q (________25558));
  nor2s1 __9__9_512052(.DIN1 (________22727), .DIN2 (_____0__24876), .Q
       (________24722));
  nor2s1 __9____512053(.DIN1 (________23959), .DIN2 (_____0__25319), .Q
       (________24328));
  hi1s1 __9____512054(.DIN (____99__26407), .Q (________25572));
  nor2s1 __9____512055(.DIN1 (_____________________21691), .DIN2
       (___0____23254), .Q (________26258));
  nnd2s1 __9____512056(.DIN1 (________23461), .DIN2 (________23734), .Q
       (________24713));
  hi1s1 __9____512057(.DIN (___0_0__23253), .Q (________23999));
  nnd2s1 __9__0_512058(.DIN1 (________22777), .DIN2 (________22692), .Q
       (____9_0__38941));
  hi1s1 __90___512059(.DIN (____0_0__34423), .Q (___9_0___39344));
  nor2s1 __9____512060(.DIN1 (_____________________21736), .DIN2
       (________23533), .Q (___00___25130));
  nor2s1 __9____512061(.DIN1 (____0_______________), .DIN2
       (_____9__25927), .Q (________26269));
  nnd2s1 __9____512062(.DIN1 (____0___23413), .DIN2 (___0____23252), .Q
       (________25607));
  nor2s1 __9____512063(.DIN1 (_____________________21689), .DIN2
       (________23351), .Q (____9___26316));
  nnd2s1 __9____512064(.DIN1 (________22729), .DIN2 (________22864), .Q
       (___9__9__39459));
  or2s1 __9___512065(.DIN1 (_____________________21732), .DIN2
       (___0____23271), .Q (________24604));
  hi1s1 __9____512066(.DIN (_____0___35660), .Q (___9_____39372));
  nor2s1 __9__0_512067(.DIN1 (___0____23251), .DIN2 (________22755), .Q
       (_________33596));
  hi1s1 __9____512068(.DIN (________24693), .Q (________25362));
  nnd2s1 __9____512069(.DIN1 (________23533), .DIN2 (____0___22550), .Q
       (____9____38898));
  hi1s1 __9____512070(.DIN (___0____23250), .Q (_____9__25348));
  nor2s1 __9099_512071(.DIN1 (___0____23248), .DIN2 (___0____23247), .Q
       (___0____23249));
  xor2s1 __9____512072(.DIN1 (_______________22077), .DIN2
       (___90___23134), .Q (___0____23246));
  or2s1 __909_512073(.DIN1 (_____________________21691), .DIN2
       (________23481), .Q (___0____23245));
  and2s1 __9___512074(.DIN1 (____0___25502), .DIN2 (________24768), .Q
       (___0_0__23244));
  nnd2s1 __9____512075(.DIN1 (________22656), .DIN2 (inData[26]), .Q
       (___0_9__23243));
  nnd2s1 __9____512076(.DIN1 (________23535), .DIN2 (________23364), .Q
       (___0____23242));
  xnr2s1 __9____512077(.DIN1 (________22493), .DIN2 (___0_____40596),
       .Q (___0____23241));
  nor2s1 __9____512078(.DIN1 (___9_0__29602), .DIN2 (________22569), .Q
       (___0____23240));
  dffacs1 _____________0_(.CLRB (reset), .CLK (clk), .DIN
       (________22537), .Q (outData[0]));
  or2s1 __9____512079(.DIN1 (___99___23213), .DIN2 (________23101), .Q
       (___0____23238));
  nnd2s1 __909__512080(.DIN1 (___0____23236), .DIN2
       (_____________________21682), .Q (___0____23237));
  nor2s1 __9____512081(.DIN1 (________23071), .DIN2 (________23093), .Q
       (___0_0__23235));
  nor2s1 __9____512082(.DIN1 (____90__24060), .DIN2 (____0___26410), .Q
       (___0_9__23234));
  xor2s1 __90___512083(.DIN1 (___0____22338), .DIN2 (_______22216), .Q
       (___0____23233));
  xor2s1 __9____512084(.DIN1 (________22372), .DIN2
       (_____________________________________________21842), .Q
       (___0____23232));
  xor2s1 __9____512085(.DIN1
       (______________________________________0___0_), .DIN2
       (___0____22308), .Q (___0____23231));
  nnd2s1 __9_009(.DIN1 (________22573), .DIN2
       (____0_____________0___21723), .Q (___0____23230));
  and2s1 __9___512086(.DIN1 (___0____23228), .DIN2
       (____0_________________21727), .Q (___0____23229));
  and2s1 __9____512087(.DIN1 (___9_9__23172), .DIN2
       (______________________21700), .Q (___0____23227));
  nnd2s1 __9_00_512088(.DIN1 (________22572), .DIN2 (_____9__24635), .Q
       (___0____23226));
  xor2s1 __9____512089(.DIN1 (_____________22079), .DIN2
       (___9____23203), .Q (___0_0__23225));
  xor2s1 __9____512090(.DIN1
       (______________________________________________21922), .DIN2
       (________22475), .Q (___009__23224));
  nnd2s1 __9____512091(.DIN1 (_____9___38319), .DIN2 (____9___22639),
       .Q (___00___23223));
  xor2s1 __9____512092(.DIN1
       (_____________________________________________21766), .DIN2
       (________22425), .Q (___00___23222));
  nor2s1 __9____512093(.DIN1 (____0___22363), .DIN2 (________23662), .Q
       (___00___23221));
  nnd2s1 __90___512094(.DIN1 (________23552), .DIN2 (____0____36220),
       .Q (___00___23220));
  or2s1 __90__512095(.DIN1 (____0________________21721), .DIN2
       (____0___22646), .Q (___00___23219));
  and2s1 __9___512096(.DIN1 (________23517), .DIN2
       (____0________________21664), .Q (___00___23218));
  nnd2s1 __90990(.DIN1 (___0____23247), .DIN2 (____9___23032), .Q
       (___00___23217));
  xor2s1 __9___512097(.DIN1
       (____________________________________________21830), .DIN2
       (________22429), .Q (___00___23216));
  nnd2s1 __9____512098(.DIN1 (____0___22845), .DIN2 (___999), .Q
       (___000));
  nor2s1 __9____512099(.DIN1 (________25744), .DIN2 (________26433), .Q
       (___99___23215));
  nor2s1 __9____512100(.DIN1 (________22865), .DIN2 (___99___23213), .Q
       (___99___23214));
  nnd2s1 __9___512101(.DIN1 (________22603), .DIN2
       (______________22067), .Q (___99___23212));
  nor2s1 __9____512102(.DIN1 (____9___22638), .DIN2 (___99___23210), .Q
       (___99___23211));
  nor2s1 __9____512103(.DIN1 (___99_), .DIN2 (___990), .Q
       (___99___23209));
  and2s1 __9_0__512104(.DIN1 (___9____23207), .DIN2
       (_____________________21709), .Q (___9_9__23208));
  xnr2s1 __9____512105(.DIN1
       (_________________________________________9___21943), .DIN2
       (___0____22315), .Q (___9____23206));
  xor2s1 __9____512106(.DIN1
       (_________________________________________________________________22000),
       .DIN2 (________22766), .Q (___9____23205));
  xnr2s1 __9____512107(.DIN1
       (_____________________________________9_______21878), .DIN2
       (___9____23203), .Q (___9____23204));
  nor2s1 __9__9_512108(.DIN1 (___9_0__23201), .DIN2 (________23916), .Q
       (___9____23202));
  xnr2s1 __9__9_512109(.DIN1 (________22960), .DIN2 (_________22039),
       .Q (___9_9__23200));
  xor2s1 __9__9_512110(.DIN1 (___0_____40449), .DIN2 (________22460),
       .Q (___9____23199));
  nnd2s1 __9____512111(.DIN1 (___9____23197), .DIN2 (_____9__22604), .Q
       (___9____23198));
  hi1s1 __9___512112(.DIN (________23523), .Q (___9____23196));
  nnd2s1 __9____512113(.DIN1 (____0___24464), .DIN2 (____0___23697), .Q
       (___9____23195));
  nor2s1 __9____512114(.DIN1 (_________32611), .DIN2 (____9___22642),
       .Q (___9____23194));
  xor2s1 __9__0_512115(.DIN1 (_________22045), .DIN2 (___9_0__23192),
       .Q (___9____23193));
  nor2s1 __9____512116(.DIN1 (_____________________21695), .DIN2
       (___9____23190), .Q (___9_9__23191));
  nnd2s1 __9__0_512117(.DIN1 (________23552), .DIN2 (________22464), .Q
       (___9____23189));
  hi1s1 __9___512118(.DIN (___0____26125), .Q (___9____23188));
  nnd2s1 __9__512119(.DIN1 (________23081), .DIN2 (________23611), .Q
       (___9____23187));
  nnd2s1 __9____512120(.DIN1 (____0___24464), .DIN2 (________22924), .Q
       (___9____23186));
  xnr2s1 __9____512121(.DIN1
       (______________________________________________21905), .DIN2
       (___90___23137), .Q (___9____23185));
  xnr2s1 __9____512122(.DIN1 (___0_0___40568), .DIN2 (________22913),
       .Q (___9____23184));
  hi1s1 __9_90_(.DIN (________23573), .Q (___9____23183));
  nnd2s1 __9__9_512123(.DIN1 (___9____23148), .DIN2 (___9_9__23181), .Q
       (___9_0__23182));
  nor2s1 __9____512124(.DIN1 (________23330), .DIN2 (____9___26581), .Q
       (___9____23180));
  nnd2s1 __90909(.DIN1 (________22670), .DIN2 (inData[22]), .Q
       (___9____23179));
  nnd2s1 __9____512125(.DIN1 (____9___22836), .DIN2 (________23662), .Q
       (___9____23178));
  nnd2s1 __9__512126(.DIN1 (___00___26054), .DIN2
       (____________________), .Q (___9____23176));
  nnd2s1 __9___512127(.DIN1 (___9____23161), .DIN2 (______22154), .Q
       (________23455));
  nor2s1 __9_0_512128(.DIN1 (___0____23236), .DIN2 (___9____23175), .Q
       (____99__23880));
  nnd2s1 __9___512129(.DIN1 (___9____23174), .DIN2 (________22610), .Q
       (____0____35302));
  nnd2s1 __9_0_512130(.DIN1 (________22686), .DIN2 (____9___23591), .Q
       (___099__23309));
  hi1s1 __9____512131(.DIN (________23418), .Q (________23744));
  nnd2s1 __9_90_512132(.DIN1 (___9____23162), .DIN2 (________24475), .Q
       (________23612));
  nnd2s1 __9__512133(.DIN1 (________25740), .DIN2
       (____0_______________), .Q (___0____24206));
  or2s1 __9_9__(.DIN1 (____0________________21717), .DIN2
       (___99___23210), .Q (_____0__23728));
  hi1s1 __9___512134(.DIN (___9____26019), .Q (________23624));
  or2s1 __9_0__512135(.DIN1 (_____________________21709), .DIN2
       (___99___24165), .Q (________24037));
  nnd2s1 __9____512136(.DIN1 (___99___23213), .DIN2 (____90__23962), .Q
       (________23432));
  hi1s1 __9____512137(.DIN (___9_0__23173), .Q (___9____24112));
  and2s1 __9_9__512138(.DIN1 (___9_9__23172), .DIN2 (________22872), .Q
       (____0___23789));
  hi1s1 __9__0_512139(.DIN (___9_____39746), .Q (____0___23882));
  nor2s1 __9____512140(.DIN1 (____0_________________21725), .DIN2
       (____9___26581), .Q (________23429));
  nnd2s1 __9_0__512141(.DIN1 (________23087), .DIN2
       (_____________________21704), .Q (___0____23250));
  hi1s1 __9____512142(.DIN (_____9__25555), .Q (____9___23593));
  nnd2s1 __9___512143(.DIN1 (___9____23171), .DIN2 (________22582), .Q
       (________25535));
  nor2s1 __9__0_512144(.DIN1 (________26174), .DIN2 (________26433), .Q
       (________23419));
  nor2s1 __9____512145(.DIN1 (___0____23252), .DIN2 (___9____23197), .Q
       (________23420));
  nor2s1 __9____512146(.DIN1 (____0___23599), .DIN2 (_____9__22680), .Q
       (________23448));
  hi1s1 __9____512147(.DIN (________23447), .Q (____0___23696));
  nnd2s1 __9__0_512148(.DIN1 (________24760), .DIN2 (________24475), .Q
       (___0_0__23253));
  nnd2s1 __9___512149(.DIN1 (___9_____39627), .DIN2
       (_____________________21669), .Q (___0____23264));
  nor2s1 __9_90_512150(.DIN1 (________23026), .DIN2 (___9____23170), .Q
       (____9___23876));
  nnd2s1 __9_09_512151(.DIN1 (________23327), .DIN2
       (_____________________21683), .Q (___0____23266));
  nnd2s1 __9__0_512152(.DIN1 (________25942), .DIN2 (________25508), .Q
       (___0____23270));
  nnd2s1 __9_0_512153(.DIN1 (________22607), .DIN2
       (_____________________21735), .Q (________23433));
  hi1s1 __9____512154(.DIN (_____0__23454), .Q (____99__23596));
  nnd2s1 __9____512155(.DIN1 (___9____23169), .DIN2 (___9____23158), .Q
       (____9___24065));
  nnd2s1 __9___512156(.DIN1 (_____9___36725), .DIN2 (_____99__36913),
       .Q (_____0___35660));
  nnd2s1 __9____512157(.DIN1 (________23669), .DIN2 (________26272), .Q
       (________23672));
  nnd2s1 __9___512158(.DIN1 (___9____23175), .DIN2
       (_____________________21684), .Q (________23866));
  hi1s1 __9__512159(.DIN (________23423), .Q (____9___23690));
  and2s1 __9_9__512160(.DIN1 (____0___22554), .DIN2 (___9____23168), .Q
       (________26470));
  hi1s1 __9__9_512161(.DIN (________24398), .Q (___0____25137));
  hi1s1 __9____512162(.DIN (________24659), .Q (________24782));
  nnd2s1 __9____512163(.DIN1 (___9____23207), .DIN2
       (_____________________21705), .Q (_____0__23646));
  hi1s1 __9____512164(.DIN (________23640), .Q (________24017));
  and2s1 __9____512165(.DIN1 (___0____23228), .DIN2 (___9____23167), .Q
       (________23651));
  nnd2s1 __9_0__512166(.DIN1 (____9___23035), .DIN2 (____0___23599), .Q
       (_____9__23767));
  or2s1 __9____512167(.DIN1 (_____________________21683), .DIN2
       (___9____23197), .Q (___0_0__25135));
  nor2s1 __9_09_512168(.DIN1 (________23449), .DIN2 (___9____23166), .Q
       (________25364));
  nor2s1 __9__0_512169(.DIN1 (____9___23031), .DIN2 (________25744), .Q
       (_____9__23682));
  or2s1 __9____512170(.DIN1 (___999), .DIN2 (____0___22942), .Q
       (________24319));
  and2s1 __9____512171(.DIN1 (_____9__22700), .DIN2 (________25352), .Q
       (________24304));
  nnd2s1 __9____512172(.DIN1 (___9____23165), .DIN2 (____9___22835), .Q
       (________24762));
  hi1s1 __9____512173(.DIN (___9____23164), .Q (________23751));
  hi1s1 __9__9_512174(.DIN (________23422), .Q (_____9___35464));
  nor2s1 __9____512175(.DIN1 (_____________________21736), .DIN2
       (_____0__22879), .Q (________23764));
  nnd2s1 __9____512176(.DIN1 (____0___23602), .DIN2 (________25508), .Q
       (___0_9__24187));
  nnd2s1 __9_99_512177(.DIN1 (________23025), .DIN2
       (_____________________21678), .Q (___0____24239));
  and2s1 __9_9__512178(.DIN1 (________22584), .DIN2
       (_____________________21735), .Q (________23760));
  hi1s1 __9____512179(.DIN (___9_9), .Q (________23660));
  nor2s1 __9_99_512180(.DIN1 (___9_9__23163), .DIN2 (_____0__23852), .Q
       (________23906));
  or2s1 __9____512181(.DIN1 (____0_______________), .DIN2
       (____0___26410), .Q (________24978));
  nor2s1 __9____512182(.DIN1 (____0___26410), .DIN2 (________22621), .Q
       (_____9__26616));
  hi1s1 __9____512183(.DIN (____0___24466), .Q (________24322));
  hi1s1 __9__0_512184(.DIN (_________34145), .Q (_____0__23929));
  nnd2s1 __9_99_512185(.DIN1 (___9____23162), .DIN2
       (_____________________21669), .Q (________23753));
  hi1s1 __9__512186(.DIN (____9___23500), .Q (________24922));
  nor2s1 __9____512187(.DIN1 (____0_______________), .DIN2
       (_____9__23008), .Q (________25458));
  or2s1 __9_512188(.DIN1 (_________________9___21711), .DIN2
       (____99__22643), .Q (________23847));
  or2s1 __9__9_512189(.DIN1 (____0_________________21724), .DIN2
       (___9_0), .Q (_____9__25728));
  or2s1 __9___512190(.DIN1 (_____________________21705), .DIN2
       (___99___24165), .Q (________24901));
  nor2s1 __9____512191(.DIN1 (____0_______________), .DIN2
       (___9____23146), .Q (_____9__25469));
  hi1s1 __9____512192(.DIN (___90___24076), .Q (________25324));
  hi1s1 __9____512193(.DIN (________25564), .Q (________26307));
  nnd2s1 __9__512194(.DIN1 (___9____23161), .DIN2
       (_____________________21736), .Q (____0___24840));
  nnd2s1 __9____512195(.DIN1 (___9____23160), .DIN2
       (_____________________21736), .Q (________24567));
  hi1s1 __9____512196(.DIN (___9____23159), .Q (_____0__25417));
  and2s1 __9____512197(.DIN1 (___9____23158), .DIN2 (________24475), .Q
       (________23741));
  hi1s1 __9____512198(.DIN (___9____23157), .Q (___9_0__24139));
  and2s1 __9____512199(.DIN1 (___9____23156), .DIN2 (___9____23158), .Q
       (___0____25198));
  nnd2s1 __9____512200(.DIN1 (___9____23169), .DIN2 (_____0__22810), .Q
       (_____9__24715));
  and2s1 __9____512201(.DIN1 (________22798), .DIN2 (___99___23213), .Q
       (________24720));
  hi1s1 __9____512202(.DIN (________23450), .Q (________23922));
  nnd2s1 __9____512203(.DIN1 (_____9__23028), .DIN2 (___9____23158), .Q
       (________24731));
  hi1s1 __9____512204(.DIN (___9_0__23155), .Q (________24308));
  nnd2s1 __9____512205(.DIN1 (___9_9__23154), .DIN2
       (_____________________21705), .Q (___0____25168));
  nnd2s1 __9_0__512206(.DIN1 (________25931), .DIN2 (____9___23030), .Q
       (___0____26083));
  hi1s1 __9___512207(.DIN (___9____23153), .Q (________28994));
  nor2s1 __9____512208(.DIN1 (___0____25163), .DIN2 (________25644), .Q
       (___9____25110));
  hi1s1 __9__0_512209(.DIN (________23538), .Q (________23845));
  nnd2s1 __9___512210(.DIN1 (___9____23169), .DIN2 (___9____23152), .Q
       (____0___24747));
  or2s1 __9____512211(.DIN1 (________23754), .DIN2 (___99___24165), .Q
       (_____9__24695));
  nnd2s1 __9____512212(.DIN1 (____99__23133), .DIN2 (____0___23697), .Q
       (________23930));
  nor2s1 __9_0__512213(.DIN1 (________22704), .DIN2 (_____0__23077), .Q
       (________23933));
  and2s1 __9____512214(.DIN1 (___0____23228), .DIN2 (___9____23151), .Q
       (________26643));
  or2s1 __9__9_512215(.DIN1 (___9____23150), .DIN2 (________24013), .Q
       (________25272));
  nnd2s1 __9___512216(.DIN1 (________23010), .DIN2
       (_____________________21683), .Q (___0____25186));
  hi1s1 __9____512217(.DIN (___99___25123), .Q (___0____25152));
  nnd2s1 __9____512218(.DIN1 (___9____23175), .DIN2 (___9____23149), .Q
       (_____0__25339));
  nnd2s1 __9____512219(.DIN1 (___9____23148), .DIN2 (___9____23165), .Q
       (___0____26087));
  and2s1 __9____512220(.DIN1 (________25337), .DIN2
       (_____________________21744), .Q (______0__35694));
  nnd2s1 __9___512221(.DIN1 (________23111), .DIN2
       (_____________________21690), .Q (_____9__25823));
  or2s1 __9__9_512222(.DIN1 (___9____23147), .DIN2 (___99___23210), .Q
       (___9_____39548));
  nor2s1 __9__0_512223(.DIN1 (____99__22548), .DIN2 (________22674), .Q
       (_________35084));
  nor2s1 __9____512224(.DIN1 (____9___23970), .DIN2 (___9____23146), .Q
       (________25829));
  nor2s1 __9____512225(.DIN1 (____90__24060), .DIN2 (___9_0), .Q
       (________25749));
  nnd2s1 __9__0_512226(.DIN1 (________24768), .DIN2 (___0____25161), .Q
       (___00___25132));
  hi1s1 __9___512227(.DIN (________23452), .Q (_____0___36728));
  nor2s1 __9____512228(.DIN1 (____0_________________21725), .DIN2
       (____0___26410), .Q (________26450));
  hi1s1 __9____512229(.DIN (________25376), .Q (________25355));
  nnd2s1 __9__512230(.DIN1 (___9____23148), .DIN2 (____0___25498), .Q
       (________26280));
  nnd2s1 __9__9_512231(.DIN1 (___0____23236), .DIN2 (___0____23252), .Q
       (________25735));
  nor2s1 __9___512232(.DIN1 (___9____23145), .DIN2 (___00___26054), .Q
       (___0____26077));
  or2s1 __9____512233(.DIN1 (_____________________21732), .DIN2
       (___9____23144), .Q (____9___25578));
  nnd2s1 __9____512234(.DIN1 (___9____23143), .DIN2
       (_____________________21730), .Q (____0_0__34423));
  nor2s1 __9_512235(.DIN1 (_______22213), .DIN2 (________23083), .Q
       (____9_9__38931));
  hi1s1 __9____512236(.DIN (________24727), .Q (___0____25176));
  xor2s1 __9____512237(.DIN1 (___9____23140), .DIN2 (______9__36337),
       .Q (___9____23141));
  xor2s1 __9____512238(.DIN1 (_________22023), .DIN2 (________22996),
       .Q (___9__));
  nnd2s1 __9____512239(.DIN1 (____9___24358), .DIN2 (________23517), .Q
       (___90___23139));
  xor2s1 __9___512240(.DIN1 (_________22019), .DIN2 (___90___23137), .Q
       (___90___23138));
  xor2s1 __90___512241(.DIN1 (_____0__22459), .DIN2 (_____9__22468), .Q
       (___90___23136));
  xnr2s1 __9____512242(.DIN1 (_________22044), .DIN2 (___90___23134),
       .Q (___90___23135));
  nnd2s1 __9____512243(.DIN1 (________23535), .DIN2 (________23474), .Q
       (___90_));
  nnd2s1 __9____512244(.DIN1 (____99__23133), .DIN2
       (_____________________21678), .Q (___900));
  xor2s1 __9____512245(.DIN1 (____9___23131), .DIN2 (____0____36245),
       .Q (____9___23132));
  xnr2s1 __9____512246(.DIN1 (________22970), .DIN2
       (____________________________________________21804), .Q
       (____9___23130));
  xor2s1 __90__512247(.DIN1 (________22484), .DIN2 (___0____22329), .Q
       (____9___23129));
  xor2s1 __9____512248(.DIN1
       (______________________________________________21903), .DIN2
       (______9__36337), .Q (____9___23128));
  hi1s1 __9__9_512249(.DIN (___0____26067), .Q (____9___23127));
  nnd2s1 __909__512250(.DIN1 (________22682), .DIN2 (____0___22552), .Q
       (____9___23126));
  or2s1 __9____512251(.DIN1 (____0________________21664), .DIN2
       (___99_), .Q (____9___23125));
  xnr2s1 __9___512252(.DIN1
       (_____________________________________________21875), .DIN2
       (_____9__23123), .Q (____90__23124));
  xor2s1 __90__512253(.DIN1 (________22405), .DIN2 (___00_), .Q
       (________23122));
  xor2s1 __9____512254(.DIN1 (___0_____40411), .DIN2 (____9___22935),
       .Q (________23121));
  xor2s1 __9____512255(.DIN1 (_________22046), .DIN2 (________22782),
       .Q (________23120));
  xor2s1 __90___512256(.DIN1 (_____0__22469), .DIN2 (___0___22198), .Q
       (________23119));
  xor2s1 __9____512257(.DIN1
       (______________________________________________21982), .DIN2
       (________23117), .Q (________23118));
  and2s1 __9____512258(.DIN1 (___9_____39627), .DIN2 (________23115),
       .Q (________23116));
  or2s1 __9__9_512259(.DIN1 (__________________0_), .DIN2
       (________23075), .Q (_____0__23114));
  xor2s1 __9____512260(.DIN1 (_____________22099), .DIN2
       (________22608), .Q (_____9__23113));
  nor2s1 __9090_512261(.DIN1 (________22526), .DIN2 (________23111), .Q
       (________23112));
  xor2s1 __9____512262(.DIN1 (_____________22083), .DIN2
       (___0____22342), .Q (________23110));
  hi1s1 __9____512263(.DIN (________23108), .Q (________23109));
  hi1s1 __9___512264(.DIN (________23106), .Q (________23107));
  nor2s1 __9_0__512265(.DIN1 (_____9__23104), .DIN2 (________22688), .Q
       (_____0__23105));
  nnd2s1 __9____512266(.DIN1 (___9____23158), .DIN2 (________23356), .Q
       (________23103));
  nor2s1 __9__9_512267(.DIN1 (_____________________21674), .DIN2
       (________23101), .Q (________23102));
  nnd2s1 __9____512268(.DIN1 (________23726), .DIN2
       (____0________________21717), .Q (________23100));
  nnd2s1 __9____512269(.DIN1 (________22570), .DIN2
       (______________22103), .Q (________23099));
  or2s1 __9___512270(.DIN1 (__________________0___21738), .DIN2
       (____9___23033), .Q (________23098));
  and2s1 __909__512271(.DIN1 (________22571), .DIN2
       (_____________________21674), .Q (________23097));
  nor2s1 __9____512272(.DIN1 (_____0__23095), .DIN2 (___99___23210), .Q
       (________23096));
  nnd2s1 __9____512273(.DIN1 (________23093), .DIN2 (________23092), .Q
       (_____9__23094));
  or2s1 __9__512274(.DIN1 (_____0__23095), .DIN2 (________23726), .Q
       (________23091));
  nor2s1 __9____512275(.DIN1 (________23089), .DIN2 (________23535), .Q
       (________23090));
  or2s1 __9___512276(.DIN1 (_____________________21704), .DIN2
       (________23087), .Q (________23088));
  nor2s1 __9____512277(.DIN1 (________22483), .DIN2 (_____0__23852), .Q
       (________23085));
  nnd2s1 __9__0_512278(.DIN1 (________23083), .DIN2 (____0___23599), .Q
       (________23084));
  nor2s1 __9____512279(.DIN1 (________23081), .DIN2 (________23080), .Q
       (________23082));
  nnd2s1 __9__9_512280(.DIN1 (________23327), .DIN2
       (_____________________21682), .Q (________23079));
  and2s1 __9____512281(.DIN1 (_____0__23077), .DIN2 (____99__22838), .Q
       (________23078));
  or2s1 __9____512282(.DIN1 (_________________9_), .DIN2
       (________23075), .Q (_____9__23076));
  nor2s1 __9____512283(.DIN1 (________23330), .DIN2 (________23081), .Q
       (________23074));
  nnd2s1 __9___512284(.DIN1 (________23072), .DIN2 (________23071), .Q
       (________23073));
  and2s1 __909__512285(.DIN1 (________23069), .DIN2 (____9___22930), .Q
       (________23070));
  nnd2s1 __9____512286(.DIN1 (________23552), .DIN2 (_______22207), .Q
       (_____0__23068));
  nnd2s1 __9____512287(.DIN1 (________23066), .DIN2 (________23065), .Q
       (_____9__23067));
  nor2s1 __9__0_512288(.DIN1 (________22715), .DIN2 (___9____23170), .Q
       (________23064));
  nnd2s1 __9____512289(.DIN1 (________23726), .DIN2 (____0___23311), .Q
       (________23063));
  nor2s1 __9__9_512290(.DIN1 (_____________________21675), .DIN2
       (________23101), .Q (________23062));
  nor2s1 __9____512291(.DIN1 (___9____23144), .DIN2 (________23065), .Q
       (________23061));
  xor2s1 __90__512292(.DIN1 (________22516), .DIN2 (_______22229), .Q
       (________23060));
  and2s1 __9____512293(.DIN1 (___9____23165), .DIN2
       (_________________0___21687), .Q (________23059));
  and2s1 __9____512294(.DIN1 (___99___23213), .DIN2
       (__________________0_), .Q (_____0__23058));
  and2s1 __9____512295(.DIN1 (___9_0), .DIN2 (________23081), .Q
       (_____9__23057));
  and2s1 __9___512296(.DIN1 (________25352), .DIN2 (_____9__24325), .Q
       (________23056));
  nor2s1 __9___512297(.DIN1 (________22461), .DIN2 (___9____23170), .Q
       (________23055));
  xor2s1 __9____512298(.DIN1 (______9__22017), .DIN2 (________22963),
       .Q (________23054));
  xor2s1 __9____512299(.DIN1
       (____________________________________________21774), .DIN2
       (________23052), .Q (________23053));
  xor2s1 __9____512300(.DIN1 (_________22039), .DIN2 (___9_____39461),
       .Q (________23051));
  or2s1 __9__9_512301(.DIN1 (________22950), .DIN2 (___00___26054), .Q
       (________23050));
  nor2s1 __9__512302(.DIN1 (____09__23048), .DIN2 (________23515), .Q
       (_____0__23049));
  nnd2s1 __9_00_512303(.DIN1 (___9_9__23154), .DIN2 (________24602), .Q
       (____0___23047));
  and2s1 __9_0__512304(.DIN1 (____0___23045), .DIN2 (____0___22843), .Q
       (____0___23046));
  hi1s1 __9____512305(.DIN (____0___23316), .Q (________23770));
  hi1s1 __9__0_512306(.DIN (_________35663), .Q (________26525));
  hi1s1 __9____512307(.DIN (________24723), .Q (________23613));
  hi1s1 __9_512308(.DIN (____0___23044), .Q (___009__24177));
  xor2s1 __9____512309(.DIN1 (___0____22332), .DIN2 (___9_9___39790),
       .Q (____0___28839));
  hi1s1 __9____512310(.DIN (_____9__23482), .Q (________23801));
  hi1s1 __9___512311(.DIN (________23629), .Q (________23637));
  nnd2s1 __9____512312(.DIN1 (____0___23043), .DIN2 (________22565), .Q
       (_________34684));
  or2s1 __9____512313(.DIN1 (____0___23042), .DIN2 (________23075), .Q
       (________23614));
  hi1s1 __9__512314(.DIN (____0___23041), .Q (________23998));
  hi1s1 __9____512315(.DIN (____0___23040), .Q (________23609));
  hi1s1 __9____512316(.DIN (________24586), .Q (_____0__23617));
  nor2s1 __9_9__512317(.DIN1 (____0________________21718), .DIN2
       (________23726), .Q (________23721));
  hi1s1 __9____512318(.DIN (________24910), .Q (___90___24072));
  hi1s1 __9____512319(.DIN (________23477), .Q (_____0__23656));
  and2s1 __9_9__512320(.DIN1 (________23535), .DIN2
       (____0____________0_), .Q (________23610));
  nor2s1 __9____512321(.DIN1 (____0_________________21724), .DIN2
       (____0___26410), .Q (___0____23278));
  nor2s1 __9____512322(.DIN1 (____9___24066), .DIN2 (___9____23144), .Q
       (_____0__23417));
  nor2s1 __9__512323(.DIN1 (________24300), .DIN2 (___99_), .Q
       (________23446));
  nor2s1 __9____512324(.DIN1 (_____0__23077), .DIN2 (____9___22837), .Q
       (___0____23258));
  hi1s1 __9__0_512325(.DIN (____00__23039), .Q (____0___23604));
  nor2s1 __9____512326(.DIN1 (____99__23038), .DIN2 (________22593), .Q
       (________26209));
  nor2s1 __9____512327(.DIN1 (____9___23037), .DIN2 (___99___23210), .Q
       (________23642));
  nnd2s1 __9____512328(.DIN1 (________23006), .DIN2 (________25352), .Q
       (___0____23255));
  hi1s1 __9__0_512329(.DIN (________24883), .Q (___0____25159));
  hi1s1 __9____512330(.DIN (_____9___35917), .Q (___9_____39319));
  hi1s1 __9____512331(.DIN (___0____23267), .Q (____0___23699));
  nnd2s1 __9____512332(.DIN1 (________23535), .DIN2 (____9___23036), .Q
       (________23926));
  nnd2s1 __9____512333(.DIN1 (____0___23311), .DIN2 (________23015), .Q
       (___9____24085));
  nnd2s1 __9____512334(.DIN1 (___9_9__23154), .DIN2 (________23754), .Q
       (________24289));
  nnd2s1 __9____512335(.DIN1 (____9___23035), .DIN2
       (____0________________21667), .Q (_____0__23919));
  nnd2s1 __9____512336(.DIN1 (___9____23160), .DIN2 (______22154), .Q
       (________24311));
  nor2s1 __9____512337(.DIN1 (________23075), .DIN2 (________23101), .Q
       (____0___24748));
  nor2s1 __9_9__512338(.DIN1 (____9___23034), .DIN2 (____9___23033), .Q
       (____0___23605));
  nor2s1 __9_9__512339(.DIN1 (____9___23032), .DIN2 (_____0__23077), .Q
       (________23755));
  nor2s1 __9_9__512340(.DIN1 (________22689), .DIN2 (____9___23033), .Q
       (________24766));
  nor2s1 __9____512341(.DIN1 (___9____26912), .DIN2 (____9___23031), .Q
       (_____0__23748));
  or2s1 __9_9__512342(.DIN1 (____0________________21718), .DIN2
       (___99___23210), .Q (________23749));
  nnd2s1 __9_9__512343(.DIN1 (_____0__22999), .DIN2 (____9___23030), .Q
       (___0____24224));
  nnd2s1 __9___512344(.DIN1 (____9___24358), .DIN2 (________23083), .Q
       (___9_0__24080));
  hi1s1 __9____512345(.DIN (____90__23029), .Q (________24877));
  nnd2s1 __9____512346(.DIN1 (_____9__23028), .DIN2 (____0___22650), .Q
       (________24700));
  hi1s1 __9___512347(.DIN (________23027), .Q (___90___24073));
  hi1s1 __9____512348(.DIN (____0___23315), .Q (________24786));
  hi1s1 __9____512349(.DIN (___0____25181), .Q (___0_9__25154));
  hi1s1 __9____512350(.DIN (________23805), .Q (_____9__23757));
  nnd2s1 __9____512351(.DIN1 (_____9__22587), .DIN2 (________26431), .Q
       (____0___23598));
  nnd2s1 __9____512352(.DIN1 (________23327), .DIN2 (___0____23252), .Q
       (____9___24742));
  nor2s1 __9_00_512353(.DIN1 (________23026), .DIN2 (___9____23190), .Q
       (________23905));
  hi1s1 __9____512354(.DIN (________25825), .Q (________26309));
  nnd2s1 __9____512355(.DIN1 (________23025), .DIN2 (_____9__23842), .Q
       (___990__24158));
  hi1s1 __9____512356(.DIN (______0__38256), .Q (_________36973));
  nor2s1 __9_0__512357(.DIN1 (_____________________21693), .DIN2
       (___9____23190), .Q (________25320));
  nnd2s1 __9_00_512358(.DIN1 (___99___23210), .DIN2 (________23024), .Q
       (__90_0__29699));
  hi1s1 __9____512359(.DIN (________23023), .Q (_____9__24705));
  nnd2s1 __9__0_512360(.DIN1 (________23022), .DIN2 (_____0__23445), .Q
       (____9___23874));
  or2s1 __9____512361(.DIN1 (________23075), .DIN2 (________22860), .Q
       (________25571));
  hi1s1 __9___512362(.DIN (___00___25131), .Q (________25742));
  nnd2s1 __9_0__512363(.DIN1 (____9___23030), .DIN2 (________23072), .Q
       (________24734));
  nnd2s1 __9____512364(.DIN1 (___9____23207), .DIN2 (________23754), .Q
       (___0____25143));
  nnd2s1 __9_0__512365(.DIN1 (________23013), .DIN2 (________23021), .Q
       (________23756));
  or2s1 __9____512366(.DIN1 (________24300), .DIN2 (___999), .Q
       (_____9__24382));
  hi1s1 __9____512367(.DIN (___0____25210), .Q (________24033));
  hi1s1 __9____512368(.DIN (_________35680), .Q (______9__35039));
  nor2s1 __9_0__512369(.DIN1 (________22854), .DIN2 (________23101), .Q
       (____0___24463));
  nnd2s1 __9_0__512370(.DIN1 (___9_9__23172), .DIN2 (________22696), .Q
       (________24324));
  hi1s1 __9____512371(.DIN (________23020), .Q (_____0__26418));
  hi1s1 __9____512372(.DIN (_____0__23019), .Q (___90___25030));
  nnd2s1 __9____512373(.DIN1 (___9____23148), .DIN2 (________22885), .Q
       (____9___25860));
  hi1s1 __9__9_512374(.DIN (___0____23260), .Q (_____9__23737));
  nnd2s1 __9____512375(.DIN1 (________23517), .DIN2
       (____0________________21662), .Q (________24693));
  hi1s1 __9___512376(.DIN (_____9__23018), .Q (___9____26025));
  hi1s1 __9____512377(.DIN (_________33686), .Q (_____0__23891));
  hi1s1 __9____512378(.DIN (________23017), .Q (________23766));
  hi1s1 __9____512379(.DIN (________23016), .Q (________24993));
  nnd2s1 __9____512380(.DIN1 (____9___22640), .DIN2
       (_____________________21744), .Q (________24594));
  nnd2s1 __9____512381(.DIN1 (____0___22556), .DIN2 (___9____23151), .Q
       (____9___25955));
  nnd2s1 __9___512382(.DIN1 (___00____41368), .DIN2 (_____9__23842), .Q
       (________24757));
  and2s1 __9_0__512383(.DIN1 (________22668), .DIN2
       (_____________________21735), .Q (____0___23694));
  nnd2s1 __9__512384(.DIN1 (________23015), .DIN2 (________23014), .Q
       (_____0__26247));
  nor2s1 __9____512385(.DIN1 (________23013), .DIN2 (________22818), .Q
       (____0____38106));
  hi1s1 __9__512386(.DIN (________23012), .Q (________23664));
  or2s1 __9____512387(.DIN1 (________24703), .DIN2 (________23101), .Q
       (___99___25119));
  hi1s1 __9__0_512388(.DIN (____90__25489), .Q (________25929));
  nnd2s1 __9___512389(.DIN1 (________23011), .DIN2
       (______________________21698), .Q (___9____24156));
  nor2s1 __9_0_512390(.DIN1 (____0________________21662), .DIN2
       (___99_), .Q (____99__26407));
  hi1s1 __9____512391(.DIN (___0____25146), .Q (_____0__24706));
  hi1s1 __9___512392(.DIN (_____9__25280), .Q (____0___25774));
  hi1s1 __9____512393(.DIN (________23864), .Q (________26429));
  hi1s1 __9___512394(.DIN (________25356), .Q (____9___27298));
  nnd2s1 __9__0_512395(.DIN1 (____99__23133), .DIN2
       (_____________________21679), .Q (________24691));
  nnd2s1 __9____512396(.DIN1 (________23010), .DIN2 (___0____23252), .Q
       (________25600));
  hi1s1 __9____512397(.DIN (______9__38496), .Q (___9_____39575));
  hi1s1 __9____512398(.DIN (___9____24081), .Q (___000__25125));
  hi1s1 __9____512399(.DIN (_____9___37943), .Q (_________38164));
  nor2s1 __9____512400(.DIN1 (_____9__22918), .DIN2 (________22574), .Q
       (___0____25171));
  hi1s1 __9____512401(.DIN (_____0__23009), .Q (___0____26078));
  nor2s1 __9____512402(.DIN1 (____9___23970), .DIN2 (_____9__23008), .Q
       (____0___26146));
  hi1s1 __9____512403(.DIN (________25373), .Q (____99__25585));
  or2s1 __9_0__512404(.DIN1 (_____________________21703), .DIN2
       (________23662), .Q (________25371));
  nnd2s1 __9_0__512405(.DIN1 (_____0__23852), .DIN2 (_____9__22690), .Q
       (_____9___37656));
  nnd2s1 __9__9_512406(.DIN1 (___9____23143), .DIN2 (________23734), .Q
       (________25946));
  and2s1 __9__512407(.DIN1 (________23006), .DIN2
       (_________________0___21728), .Q (________23007));
  or2s1 __9_9__512408(.DIN1 (________23004), .DIN2 (________23003), .Q
       (________23005));
  nor2s1 __9____512409(.DIN1 (____90__24060), .DIN2 (________23438), .Q
       (________23002));
  or2s1 __9___512410(.DIN1 (________22414), .DIN2 (________23117), .Q
       (________23001));
  nnd2s1 __9____512411(.DIN1 (_____0__22999), .DIN2 (________23959), .Q
       (________23000));
  nor2s1 __9___512412(.DIN1 (_____0__22393), .DIN2 (____9___23591), .Q
       (_____9__22998));
  nor2s1 __9____512413(.DIN1 (________22471), .DIN2 (________22996), .Q
       (________22997));
  and2s1 __9___512414(.DIN1 (________24884), .DIN2 (________22994), .Q
       (________22995));
  xor2s1 __9__0_512415(.DIN1 (___0___22199), .DIN2
       (_______________________________________________________________9),
       .Q (________22993));
  nor2s1 __9__9_512416(.DIN1 (_______22257), .DIN2 (________25597), .Q
       (________22992));
  xnr2s1 __9__0_512417(.DIN1 (___00), .DIN2 (___0__0__40511), .Q
       (________22991));
  xor2s1 __9___512418(.DIN1 (______), .DIN2 (________22984), .Q
       (________22990));
  nnd2s1 __9____512419(.DIN1 (____90__23962), .DIN2 (________24703), .Q
       (_____0__22989));
  or2s1 __9____512420(.DIN1 (____0___22943), .DIN2 (________22379), .Q
       (_____9__22988));
  or2s1 __9_90_512421(.DIN1 (________22986), .DIN2 (____0___22747), .Q
       (________22987));
  xor2s1 __9____512422(.DIN1
       (______________________________________________21911), .DIN2
       (________22984), .Q (________22985));
  nor2s1 __9____512423(.DIN1
       (_______________________________________________________________0__22010),
       .DIN2 (____0___22452), .Q (________22983));
  nnd2s1 __9__0_512424(.DIN1 (________22981), .DIN2
       (_____________________21742), .Q (________22982));
  nor2s1 __9___512425(.DIN1 (________23754), .DIN2 (___00___22289), .Q
       (________22980));
  nor2s1 __9__9_512426(.DIN1 (___99____39814), .DIN2 (___0____22327),
       .Q (_____0__22979));
  nnd2s1 __9____512427(.DIN1 (________22977), .DIN2 (________22437), .Q
       (_____9__22978));
  nor2s1 __9__0_512428(.DIN1 (_____________________21731), .DIN2
       (____00__22839), .Q (________22976));
  nnd2s1 __9____512429(.DIN1 (____9___23786), .DIN2 (____0___22457), .Q
       (________22975));
  nnd2s1 __9____512430(.DIN1 (________22973), .DIN2 (____9___23037), .Q
       (________22974));
  nor2s1 __9____512431(.DIN1 (________23362), .DIN2 (________22795), .Q
       (________22972));
  nor2s1 __9____512432(.DIN1
       (____________________________________________21804), .DIN2
       (________22970), .Q (________22971));
  and2s1 __9__0_512433(.DIN1 (____0___23414), .DIN2
       (_________________0___21740), .Q (_____0__22969));
  nnd2s1 __9____512434(.DIN1 (________22977), .DIN2
       (_____________________________________________21815), .Q
       (_____9__22968));
  nnd2s1 __9__0_512435(.DIN1 (________25942), .DIN2 (________26618), .Q
       (________22967));
  nor2s1 __9__0_512436(.DIN1 (___9____24088), .DIN2 (________22965), .Q
       (________22966));
  or2s1 __9____512437(.DIN1 (___0____22352), .DIN2 (________22963), .Q
       (________22964));
  nor2s1 __9____512438(.DIN1 (____0________________21716), .DIN2
       (_____0__23095), .Q (________22962));
  or2s1 __9____512439(.DIN1 (________22407), .DIN2 (________22960), .Q
       (________22961));
  xnr2s1 __9____512440(.DIN1
       (____________________________________________21772), .DIN2
       (___00__22196), .Q (_____0__22959));
  nnd2s1 __9____512441(.DIN1 (________24882), .DIN2 (___0_____40505),
       .Q (_____9__22958));
  nor2s1 __9__0_512442(.DIN1 (___9____25102), .DIN2 (___0____22326), .Q
       (________22957));
  and2s1 __9____512443(.DIN1 (________22955), .DIN2
       (____0________________21663), .Q (________22956));
  or2s1 __9____512444(.DIN1 (_____________________21746), .DIN2
       (________22953), .Q (________22954));
  xnr2s1 __9____512445(.DIN1
       (______________________________________0_______21891), .DIN2
       (_______22243), .Q (________22952));
  nor2s1 __9____512446(.DIN1 (________22994), .DIN2 (________22950), .Q
       (________22951));
  or2s1 __9___512447(.DIN1 (_____________________21678), .DIN2
       (___9_0__23201), .Q (_____0__22949));
  nnd2s1 __9____512448(.DIN1 (____9___22932), .DIN2 (_____9__22868), .Q
       (____09__22948));
  nor2s1 __9____512449(.DIN1 (________26426), .DIN2 (________22981), .Q
       (____0___22947));
  nor2s1 __9___512450(.DIN1 (_____________________21706), .DIN2
       (____9___23591), .Q (____0___22946));
  and2s1 __9____512451(.DIN1 (___9____23152), .DIN2
       (_____________________21670), .Q (____0___22945));
  or2s1 __9____512452(.DIN1 (____0___22943), .DIN2 (____0___22942), .Q
       (____0___22944));
  xnr2s1 __9____512453(.DIN1 (___9___22193), .DIN2
       (____________________________________________21834), .Q
       (____0___22941));
  and2s1 __9__9_512454(.DIN1 (________23800), .DIN2 (________22386), .Q
       (____0___22940));
  nor2s1 __9____512455(.DIN1 (_____9__22828), .DIN2 (____9___24062), .Q
       (____00__22939));
  nnd2s1 __90_9_512456(.DIN1 (________22373), .DIN2 (inData[24]), .Q
       (____99__22938));
  and2s1 __9___512457(.DIN1 (________22702), .DIN2
       (__________________0___21712), .Q (____9___22937));
  or2s1 __9____512458(.DIN1 (________22411), .DIN2 (____9___22935), .Q
       (____9___22936));
  nnd2s1 __9__9_512459(.DIN1 (____9___22933), .DIN2 (____9___22932), .Q
       (____9___22934));
  xor2s1 __9____512460(.DIN1 (____9___22930), .DIN2 (____9___22544), .Q
       (____9___22931));
  xor2s1 __9____512461(.DIN1 (___________________), .DIN2
       (_________33117), .Q (____90__22929));
  or2s1 __9____512462(.DIN1 (______0___22057), .DIN2 (________22927),
       .Q (_____9__22928));
  nor2s1 __9__9_512463(.DIN1 (___9____25102), .DIN2 (__9____22287), .Q
       (________22926));
  nnd2s1 __9____512464(.DIN1 (____9___23786), .DIN2 (________22924), .Q
       (________22925));
  nnd2s1 __9___512465(.DIN1 (________24302), .DIN2 (____9___24360), .Q
       (________22923));
  and2s1 __9__0_512466(.DIN1 (________22921), .DIN2
       (____________________), .Q (________22922));
  xor2s1 __9____512467(.DIN1 (______22161), .DIN2 (___0_____40537), .Q
       (________22920));
  nor2s1 __9__512468(.DIN1 (_____________________21672), .DIN2
       (_____9__22918), .Q (_____0__22919));
  nor2s1 __9__512469(.DIN1 (____00), .DIN2 (____0___22455), .Q
       (________22917));
  nor2s1 __9____512470(.DIN1 (________23555), .DIN2 (________22953), .Q
       (________22916));
  nor2s1 __9____512471(.DIN1 (____0___26590), .DIN2 (___0____23292), .Q
       (________22915));
  nnd2s1 __9____512472(.DIN1 (________22913), .DIN2 (___0_0___40568),
       .Q (________22914));
  xor2s1 __9___512473(.DIN1 (_____0__22909), .DIN2
       (_____________________________________________21843), .Q
       (________22912));
  nor2s1 __9____512474(.DIN1 (_____________________21747), .DIN2
       (________22465), .Q (________22911));
  xor2s1 __9___512475(.DIN1
       (______________________________________________________________________________________0__22093),
       .DIN2 (_____0__22909), .Q (________22910));
  xor2s1 __9____512476(.DIN1
       (__________________________________________________________________21994),
       .DIN2 (_____0__22771), .Q (_____9__22908));
  nnd2s1 __9____512477(.DIN1 (________23469), .DIN2 (______22131), .Q
       (________22907));
  or2s1 __9____512478(.DIN1 (___9_0__23201), .DIN2 (________22708), .Q
       (________22906));
  hi1s1 __9____512479(.DIN (___9____23143), .Q (________22905));
  nor2s1 __9____512480(.DIN1 (________22887), .DIN2 (_____9__23900), .Q
       (________22904));
  xor2s1 __9____512481(.DIN1 (________22675), .DIN2 (__________22063),
       .Q (________22903));
  nor2s1 __9__0_512482(.DIN1 (_____________________21678), .DIN2
       (_____0__22849), .Q (________22902));
  or2s1 __9____512483(.DIN1 (_____________________21672), .DIN2
       (____0___23504), .Q (________22901));
  or2s1 __9____512484(.DIN1 (_____0__22899), .DIN2 (________22850), .Q
       (________22900));
  nnd2s1 __9____512485(.DIN1 (____0___22847), .DIN2 (____90__24060), .Q
       (_____9__22898));
  or2s1 __9____512486(.DIN1 (_____________________21695), .DIN2
       (________22462), .Q (________22897));
  or2s1 __9____512487(.DIN1 (_____________________21673), .DIN2
       (____0___23504), .Q (________22896));
  nnd2s1 __9____512488(.DIN1 (___0____22319), .DIN2 (inData[12]), .Q
       (________22895));
  nnd2s1 __9___512489(.DIN1 (________24882), .DIN2
       (_____________________21747), .Q (________22894));
  nor2s1 __9___512490(.DIN1 (____9___23878), .DIN2 (________22435), .Q
       (________22893));
  nor2s1 __9_9__512491(.DIN1 (________22891), .DIN2 (________22890), .Q
       (________22892));
  or2s1 __9____512492(.DIN1 (___09___23306), .DIN2 (___9____23152), .Q
       (_____0__22889));
  and2s1 __9____512493(.DIN1 (________22887), .DIN2
       (_____________________21706), .Q (_____9__22888));
  nnd2s1 __9____512494(.DIN1 (________22885), .DIN2 (________22884), .Q
       (________22886));
  or2s1 __9____512495(.DIN1 (__________________0___21686), .DIN2
       (___0____23289), .Q (________22883));
  or2s1 __9____512496(.DIN1 (__________________0___21697), .DIN2
       (________22921), .Q (________22882));
  nnd2s1 __9____512497(.DIN1 (________23469), .DIN2 (______22128), .Q
       (________22881));
  hi1s1 __9____512498(.DIN (_____0__22879), .Q (________22880));
  hi1s1 __9____512499(.DIN (________22877), .Q (_____9__22878));
  nor2s1 __9_0__512500(.DIN1 (____0________________21714), .DIN2
       (________22876), .Q (___9____23153));
  or2s1 __9___512501(.DIN1 (____0________________21662), .DIN2
       (________22875), .Q (________23541));
  and2s1 __9____512502(.DIN1 (____0___22842), .DIN2
       (__________________0___21750), .Q (________23490));
  nor2s1 __9____512503(.DIN1 (________22874), .DIN2 (________22873), .Q
       (_________33859));
  nnd2s1 __9____512504(.DIN1 (____0___25502), .DIN2
       (_____________________21744), .Q (________23016));
  nnd2s1 __9_9__512505(.DIN1 (________22872), .DIN2 (____9___22545), .Q
       (___0____23265));
  nnd2s1 __9_9__512506(.DIN1 (________22871), .DIN2 (_____0__23445), .Q
       (________23360));
  nor2s1 __9_909(.DIN1 (_____9__24325), .DIN2 (____9___22445), .Q
       (________23383));
  nor2s1 __9_9__512507(.DIN1 (________22870), .DIN2 (_____0__22869), .Q
       (________29123));
  nor2s1 __9_9_9(.DIN1 (________22391), .DIN2 (___9____23147), .Q
       (___9_0__23173));
  nnd2s1 __9____512508(.DIN1 (___9____24088), .DIN2 (________22965), .Q
       (_____0__23086));
  nnd2s1 __9__512509(.DIN1 (____9___24358), .DIN2 (_____9__22868), .Q
       (________23106));
  nor2s1 __9____512510(.DIN1 (____0___22743), .DIN2 (________22851), .Q
       (___9_0__23155));
  nor2s1 __9___512511(.DIN1 (________22867), .DIN2 (____0__22247), .Q
       (_____9__23453));
  nnd2s1 __9_9__512512(.DIN1 (____9___26583), .DIN2
       (____________________), .Q (___9____23142));
  nor2s1 __9____512513(.DIN1 (________22866), .DIN2 (____0___22942), .Q
       (_____9__23616));
  nor2s1 __9_9__512514(.DIN1 (_______22256), .DIN2 (________26419), .Q
       (____0___23040));
  nnd2s1 __9____512515(.DIN1 (____90__23962), .DIN2 (________22865), .Q
       (____0___23041));
  nnd2s1 __9____512516(.DIN1 (________25569), .DIN2 (_______22248), .Q
       (___9____23157));
  nnd2s1 __9_9__512517(.DIN1 (________22863), .DIN2
       (____0_____________0_), .Q (___9____23164));
  nnd2s1 __9_0__512518(.DIN1 (________22871), .DIN2 (________22714), .Q
       (_____0__23019));
  nor2s1 __9_90_512519(.DIN1 (________22857), .DIN2 (________22864), .Q
       (________23428));
  nnd2s1 __9_90_512520(.DIN1 (________23800), .DIN2 (________22884), .Q
       (________23108));
  nnd2s1 __9____512521(.DIN1 (________22625), .DIN2 (________22863), .Q
       (________23017));
  nnd2s1 __9_0__512522(.DIN1 (________22616), .DIN2
       (_____________________21703), .Q (________23027));
  nnd2s1 __9__512523(.DIN1 (________22862), .DIN2
       (____0_______________), .Q (_____9__23018));
  nor2s1 __9____512524(.DIN1 (___9____23149), .DIN2 (________22693), .Q
       (____0___23415));
  nnd2s1 __9_9_512525(.DIN1 (________23014), .DIN2 (________22705), .Q
       (___0____23259));
  and2s1 __9_9__512526(.DIN1 (________24544), .DIN2
       (____0_____________0_), .Q (___0_9__23262));
  nor2s1 __9__9_512527(.DIN1 (____0________________21714), .DIN2
       (________22864), .Q (_____9__23435));
  hi1s1 __9____512528(.DIN (________23022), .Q (___0____23261));
  nnd2s1 __9__9_512529(.DIN1 (________23071), .DIN2
       (____0_____________0___21723), .Q (___909));
  nnd2s1 __9____512530(.DIN1 (________22861), .DIN2
       (_____________________21744), .Q (____90__23029));
  nnd2s1 __9_9_512531(.DIN1 (________22762), .DIN2 (___0____23256), .Q
       (________23351));
  nor2s1 __9_9__512532(.DIN1 (________23989), .DIN2 (________24418), .Q
       (________23615));
  nor2s1 __9____512533(.DIN1 (____0___23042), .DIN2 (_____0__22859), .Q
       (____9___24063));
  nor2s1 __9__9_512534(.DIN1 (________23391), .DIN2 (________22619), .Q
       (____0___23315));
  nnd2s1 __9_9__512535(.DIN1 (____9___22833), .DIN2 (________23014), .Q
       (________23920));
  nor2s1 __9____512536(.DIN1 (________25644), .DIN2 (________26440), .Q
       (____0___23316));
  nnd2s1 __9__9_512537(.DIN1 (________24625), .DIN2 (___0____25161), .Q
       (_____9__23586));
  nor2s1 __9__9_512538(.DIN1 (________22860), .DIN2 (_____0__22859), .Q
       (________24597));
  nnd2s1 __9_0__512539(.DIN1 (________23469), .DIN2
       (_____________________21741), .Q (________23422));
  or2s1 __9____512540(.DIN1 (________24475), .DIN2 (_____9__22858), .Q
       (____0___23503));
  or2s1 __9____512541(.DIN1 (________24300), .DIN2 (____0___22943), .Q
       (________26575));
  nor2s1 __9_9__512542(.DIN1 (________22857), .DIN2 (________22856), .Q
       (_____0__23426));
  nor2s1 __9__9_512543(.DIN1 (____09__26331), .DIN2 (________26421), .Q
       (____9___24452));
  nor2s1 __9____512544(.DIN1 (________22867), .DIN2 (____9___23037), .Q
       (________23477));
  nnd2s1 __9____512545(.DIN1 (________22871), .DIN2 (________22855), .Q
       (________23864));
  nor2s1 __9_9_0(.DIN1 (________22854), .DIN2 (____0___23042), .Q
       (___0____25172));
  nor2s1 __9____512546(.DIN1 (_____________________21745), .DIN2
       (________22853), .Q (________25797));
  nor2s1 __9___512547(.DIN1 (________22852), .DIN2 (___990), .Q
       (________23640));
  nor2s1 __9_9__512548(.DIN1 (_____9__24325), .DIN2 (________22851), .Q
       (________23461));
  nor2s1 __9_0__512549(.DIN1 (____0___22365), .DIN2 (________23709), .Q
       (___0____23260));
  nnd2s1 __9__9_512550(.DIN1 (________25569), .DIN2
       (_____________________21744), .Q (___0____25210));
  nnd2s1 __9____512551(.DIN1 (________22850), .DIN2 (________22953), .Q
       (________23437));
  nnd2s1 __9____512552(.DIN1 (_____0__22849), .DIN2 (____09__22848), .Q
       (________23447));
  nnd2s1 __9_9__512553(.DIN1 (____9___22831), .DIN2 (________22857), .Q
       (_____0__23436));
  or2s1 __9_9__512554(.DIN1 (_____________________21735), .DIN2
       (________22667), .Q (___0____23271));
  nnd2s1 __9____512555(.DIN1 (___9____24123), .DIN2 (____0___22840), .Q
       (________24910));
  or2s1 __9____512556(.DIN1 (_____________________21679), .DIN2
       (____09__22848), .Q (________23867));
  nnd2s1 __9_0__512557(.DIN1 (________25931), .DIN2 (_______22252), .Q
       (_____0__23454));
  nnd2s1 __9____512558(.DIN1 (____0___22847), .DIN2
       (____0_________________21725), .Q (________23927));
  nnd2s1 __9_00_512559(.DIN1 (___0_9__22353), .DIN2
       (_____________________21691), .Q (________23531));
  nnd2s1 __9____512560(.DIN1 (________23006), .DIN2 (___9____24088), .Q
       (________23984));
  nnd2s1 __9____512561(.DIN1 (________22867), .DIN2 (__9___22168), .Q
       (____0___23410));
  nnd2s1 __9____512562(.DIN1 (____9___24358), .DIN2 (____9___23036), .Q
       (_____9__24486));
  or2s1 __9_9__512563(.DIN1 (_____________________21747), .DIN2
       (________24882), .Q (_________38543));
  nor2s1 __9____512564(.DIN1 (___9____26912), .DIN2 (________22850), .Q
       (________23554));
  nnd2s1 __9_0__512565(.DIN1 (________22792), .DIN2 (____0___22846), .Q
       (________23563));
  nnd2s1 __9____512566(.DIN1 (____0___25502), .DIN2 (________26431), .Q
       (________24586));
  nor2s1 __9____512567(.DIN1 (____0___22845), .DIN2 (____0___22942), .Q
       (________24723));
  nnd2s1 __9____512568(.DIN1 (____9___24358), .DIN2 (____0___22844), .Q
       (________24470));
  hi1s1 __9__9_512569(.DIN (___0_0__25155), .Q (________24490));
  nnd2s1 __9____512570(.DIN1 (________22871), .DIN2 (___9____24123), .Q
       (_____0__24393));
  nor2s1 __9__0_512571(.DIN1 (_____0__26149), .DIN2 (________22786), .Q
       (________25564));
  nor2s1 __9_0_512572(.DIN1 (____0___22843), .DIN2 (________24418), .Q
       (____90__25489));
  nnd2s1 __9_999(.DIN1 (____0___22842), .DIN2 (________26217), .Q
       (___9____24084));
  nnd2s1 __9____512573(.DIN1 (________23669), .DIN2 (___99___26049), .Q
       (_____9__25555));
  nor2s1 __9____512574(.DIN1 (____0___22841), .DIN2 (___0____26080), .Q
       (___0_0__24248));
  nor2s1 __9_00_512575(.DIN1 (________22854), .DIN2 (________22860), .Q
       (________25380));
  or2s1 __9____512576(.DIN1 (__________________0___21750), .DIN2
       (___0____23292), .Q (____9____34370));
  nor2s1 __9___512577(.DIN1 (________22617), .DIN2 (________22965), .Q
       (___99___25118));
  nnd2s1 __9____512578(.DIN1 (________23364), .DIN2 (_____9__24635), .Q
       (___9____24081));
  or2s1 __9____512579(.DIN1 (________22950), .DIN2 (____0___22840), .Q
       (________23901));
  nor2s1 __9_0_512580(.DIN1 (________22628), .DIN2 (________22707), .Q
       (________23914));
  nor2s1 __9___512581(.DIN1 (____0___22845), .DIN2 (___990), .Q
       (____90__24736));
  nor2s1 __9___512582(.DIN1 (________24418), .DIN2 (____9___22540), .Q
       (________25751));
  nor2s1 __9____512583(.DIN1 (_____________________21742), .DIN2
       (________25644), .Q (___00___25131));
  hi1s1 __9____512584(.DIN (_________38591), .Q (_________36291));
  nor2s1 __9____512585(.DIN1 (________22632), .DIN2 (___9____23147), .Q
       (________25825));
  nor2s1 __9_0__512586(.DIN1 (_____________________21735), .DIN2
       (________22583), .Q (________23430));
  nnd2s1 __9_0__512587(.DIN1 (____9___24358), .DIN2 (_____9__24635), .Q
       (___0____26125));
  or2s1 __9_0__512588(.DIN1 (_________________0___21728), .DIN2
       (________22965), .Q (_____0__24876));
  nor2s1 __9_0_512589(.DIN1 (_____________________21694), .DIN2
       (________22706), .Q (____9___24061));
  nnd2s1 __9____512590(.DIN1 (____00__22839), .DIN2 (________23006), .Q
       (_________33686));
  nor2s1 __9____512591(.DIN1 (____99__22838), .DIN2 (____9___22837), .Q
       (________24690));
  nnd2s1 __9____512592(.DIN1 (______22153), .DIN2 (___0____23252), .Q
       (________23325));
  nor2s1 __9___512593(.DIN1 (_____9__23635), .DIN2 (____0___22942), .Q
       (________23629));
  or2s1 __9____512594(.DIN1 (___09___23306), .DIN2 (_____9__22858), .Q
       (____9___24738));
  hi1s1 __9__9_512595(.DIN (____9___22836), .Q (________24313));
  nor2s1 __9___512596(.DIN1 (________22385), .DIN2 (_____9__22918), .Q
       (___0____25156));
  and2s1 __9__9_512597(.DIN1 (________22973), .DIN2 (_____0__23095), .Q
       (_____9___38509));
  nnd2s1 __9____512598(.DIN1 (______22153), .DIN2
       (_____________________21683), .Q (________23573));
  nor2s1 __9____512599(.DIN1 (________22857), .DIN2 (________22876), .Q
       (________23441));
  and2s1 __9___512600(.DIN1 (___0____23251), .DIN2
       (_____________________21742), .Q (_____9__23918));
  and2s1 __9____512601(.DIN1 (____9___22835), .DIN2 (____0___25498), .Q
       (________26259));
  and2s1 __9__9_512602(.DIN1 (____9___22834), .DIN2
       (_____________________21684), .Q (________25270));
  nor2s1 __9_0__512603(.DIN1 (_____________________21704), .DIN2
       (________22631), .Q (___99___25123));
  and2s1 __9____512604(.DIN1 (________23372), .DIN2
       (_________________9___21749), .Q (____0____38117));
  nor2s1 __9_0__512605(.DIN1 (____0____________0_), .DIN2
       (____0___22943), .Q (___0____25146));
  nor2s1 __9____512606(.DIN1 (________23384), .DIN2 (________22965), .Q
       (___0____25181));
  nnd2s1 __9_0__512607(.DIN1 (_____0__23095), .DIN2 (____9___22833), .Q
       (_____0__24316));
  nor2s1 __9___512608(.DIN1 (_________________9___21749), .DIN2
       (________22703), .Q (_____9___37943));
  nor2s1 __9_0__512609(.DIN1 (_____________________21704), .DIN2
       (_______22282), .Q (___0____25157));
  or2s1 __9_0__512610(.DIN1 (____0________________21665), .DIN2
       (____9___22832), .Q (_________38385));
  or2s1 __9____512611(.DIN1 (________22419), .DIN2 (________24544), .Q
       (___99_0__39864));
  nnd2s1 __9____512612(.DIN1 (________23364), .DIN2
       (____0________________21662), .Q (________25376));
  nor2s1 __9____512613(.DIN1 (_________38301), .DIN2 (________22666),
       .Q (_________38456));
  or2s1 __9__0_512614(.DIN1 (_____9__22918), .DIN2 (_____9__22858), .Q
       (________24797));
  hi1s1 __9___512615(.DIN (________23552), .Q (________23533));
  nnd2s1 __9___512616(.DIN1 (________22876), .DIN2 (________22864), .Q
       (_________37744));
  and2s1 __9____512617(.DIN1 (_____9___38319), .DIN2 (________23372),
       .Q (_________38249));
  nnd2s1 __9_09_512618(.DIN1 (____9___22831), .DIN2
       (____0________________21714), .Q (______9__38496));
  or2s1 __9____512619(.DIN1 (_____9___37752), .DIN2 (____9___23034), .Q
       (_________37722));
  nnd2s1 __9____512620(.DIN1 (________22850), .DIN2 (___9____26912), .Q
       (____9___22830));
  and2s1 __9____512621(.DIN1 (_____9__22828), .DIN2
       (______________________21751), .Q (____90__22829));
  nnd2s1 __9____512622(.DIN1 (________24882), .DIN2 (___0__9__40550),
       .Q (________22827));
  nor2s1 __9____512623(.DIN1 (___9____23151), .DIN2 (________23438), .Q
       (________22826));
  nor2s1 __9____512624(.DIN1 (________22510), .DIN2
       (_____________________21669), .Q (________22825));
  nor2s1 __9___512625(.DIN1 (________22514), .DIN2
       (_____________________21705), .Q (________22824));
  nor2s1 __9___512626(.DIN1 (________26217), .DIN2 (___0____23292), .Q
       (________22823));
  xor2s1 __9____512627(.DIN1 (_______22185), .DIN2 (_________33591), .Q
       (________22822));
  nnd2s1 __9____512628(.DIN1 (___9____23168), .DIN2 (____9___23970), .Q
       (________22821));
  nnd2s1 __9____512629(.DIN1 (________22953), .DIN2 (________23555), .Q
       (________22820));
  and2s1 __9____512630(.DIN1 (________22818), .DIN2
       (_________________9___21711), .Q (_____9__22819));
  nnd2s1 __9____512631(.DIN1 (________22885), .DIN2 (___0____23256), .Q
       (________22817));
  nnd2s1 __9____512632(.DIN1 (________22861), .DIN2
       (_____________________21743), .Q (________22816));
  nnd2s1 __9____512633(.DIN1 (___0____22341), .DIN2 (inData[10]), .Q
       (________22815));
  nnd2s1 __9____512634(.DIN1 (___9___22264), .DIN2
       (__________________________________________________________________21986),
       .Q (________22814));
  or2s1 __9____512635(.DIN1 (_____________________21670), .DIN2
       (_____9__22858), .Q (________22813));
  nor2s1 __9___512636(.DIN1 (____0___28017), .DIN2 (___9___22265), .Q
       (________22812));
  nnd2s1 __9____512637(.DIN1 (_____0__22810), .DIN2 (________23356), .Q
       (________22811));
  xor2s1 __9____512638(.DIN1
       (__________________________________________________________________21988),
       .DIN2 (_______22209), .Q (________22809));
  nor2s1 __9__0_512639(.DIN1 (____0____________9___21722), .DIN2
       (_____0__22701), .Q (________22808));
  and2s1 __9__512640(.DIN1 (____9___26583), .DIN2
       (______________________21698), .Q (________22807));
  nnd2s1 __9____512641(.DIN1 (________22501), .DIN2 (_____9__22392), .Q
       (________22806));
  nor2s1 __9____512642(.DIN1 (_________________9___21711), .DIN2
       (________22818), .Q (________22805));
  and2s1 __9____512643(.DIN1 (____9___22932), .DIN2
       (____0______________), .Q (________22804));
  nnd2s1 __9__0_512644(.DIN1 (___90____38993), .DIN2 (________23959),
       .Q (________22803));
  nor2s1 __9__0_512645(.DIN1 (________22400), .DIN2 (________22862), .Q
       (________22802));
  nnd2s1 __9____512646(.DIN1 (____0___22842), .DIN2
       (______________________21751), .Q (_____0__22801));
  nor2s1 __9__0_512647(.DIN1 (________22867), .DIN2 (___9____23147), .Q
       (_____9__22800));
  and2s1 __9____512648(.DIN1 (________22798), .DIN2
       (_____________________21674), .Q (________22799));
  nor2s1 __9____512649(.DIN1 (________22502), .DIN2 (________22505), .Q
       (________22797));
  nor2s1 __9__9_512650(.DIN1 (_____________________21695), .DIN2
       (________22795), .Q (________22796));
  nor2s1 __9____512651(.DIN1 (___0____22330), .DIN2 (____0___22842), .Q
       (________22794));
  nor2s1 __9____512652(.DIN1 (________22416), .DIN2 (________22792), .Q
       (________22793));
  or2s1 __9____512653(.DIN1 (___0___22202), .DIN2 (________23089), .Q
       (_____0__22791));
  xor2s1 __9__0_512654(.DIN1 (___0_____40588), .DIN2 (______22162), .Q
       (_____9__22790));
  nor2s1 __9____512655(.DIN1 (_______22283), .DIN2 (________22788), .Q
       (________22789));
  nnd2s1 __9___512656(.DIN1 (________22786), .DIN2 (________26419), .Q
       (________22787));
  nnd2s1 __9__0_512657(.DIN1 (____9___22835), .DIN2 (_____9__23444), .Q
       (________22785));
  nnd2s1 __9____512658(.DIN1 (________22699), .DIN2
       (__________________0___21712), .Q (________22784));
  nor2s1 __9____512659(.DIN1 (_____0__22433), .DIN2 (________22782), .Q
       (________22783));
  and2s1 __9____512660(.DIN1 (________24884), .DIN2 (____9___26583), .Q
       (_____0__22781));
  nor2s1 __9____512661(.DIN1 (________23555), .DIN2 (________22850), .Q
       (_____9__22780));
  and2s1 __9__0_512662(.DIN1 (________22871), .DIN2 (________22950), .Q
       (________22779));
  nor2s1 __9____512663(.DIN1 (____0_________________21725), .DIN2
       (___9____23167), .Q (________22778));
  nnd2s1 __9____512664(.DIN1 (____9___23036), .DIN2 (____0___23599), .Q
       (________22777));
  nor2s1 __9__9_512665(.DIN1 (___99____39814), .DIN2 (___0_0__22334),
       .Q (________22776));
  nnd2s1 __9____512666(.DIN1 (____00__22839), .DIN2 (_____9__24325), .Q
       (________22775));
  nor2s1 __9____512667(.DIN1 (___0_____40495), .DIN2 (________23372),
       .Q (________22774));
  xor2s1 __9____512668(.DIN1 (________22772), .DIN2 (_____0__22771), .Q
       (________22773));
  and2s1 __9____512669(.DIN1 (________22965), .DIN2 (________22851), .Q
       (_____9__22770));
  nnd2s1 __9__9_512670(.DIN1 (________24884), .DIN2
       (__________________0___21697), .Q (________22769));
  and2s1 __9___512671(.DIN1 (________22798), .DIN2 (________24703), .Q
       (________22768));
  or2s1 __9____512672(.DIN1 (___), .DIN2 (________22766), .Q
       (________22767));
  nnd2s1 __9____512673(.DIN1 (________22620), .DIN2 (________22792), .Q
       (________22765));
  nnd2s1 __9___512674(.DIN1 (________23469), .DIN2 (________22754), .Q
       (________22764));
  nnd2s1 __9____512675(.DIN1 (________22762), .DIN2 (_____9__23444), .Q
       (________22763));
  hi1s1 __9____512676(.DIN (_____9__22760), .Q (_____0__22761));
  xor2s1 __9____512677(.DIN1 (________22599), .DIN2 (______0___22055),
       .Q (________22759));
  nnd2s1 __9____512678(.DIN1 (____0___22942), .DIN2 (____0___22454), .Q
       (________22758));
  nor2s1 __9___512679(.DIN1 (________23959), .DIN2 (________23092), .Q
       (________22757));
  nor2s1 __9____512680(.DIN1 (____9___23878), .DIN2 (________22430), .Q
       (________22756));
  nor2s1 __9____512681(.DIN1 (________22754), .DIN2 (________22753), .Q
       (________22755));
  nnd2s1 __9___512682(.DIN1 (____0___22842), .DIN2 (____0___26590), .Q
       (________22752));
  nor2s1 __9____512683(.DIN1 (_____________________21679), .DIN2
       (________22717), .Q (_____0__22751));
  nor2s1 __9____512684(.DIN1 (___0__), .DIN2 (___0____23276), .Q
       (____09__22750));
  nor2s1 __9____512685(.DIN1 (_____9__22538), .DIN2 (____9___23591), .Q
       (____0___22749));
  nor2s1 __9___512686(.DIN1 (____0___22747), .DIN2 (____0___22746), .Q
       (____0___22748));
  nor2s1 __9__9_512687(.DIN1 (_____0__23095), .DIN2 (_____0__22614), .Q
       (____0___22745));
  nnd2s1 __9__512688(.DIN1 (____00__22839), .DIN2 (____0___22743), .Q
       (____0___22744));
  nor2s1 __9____512689(.DIN1 (___9____26912), .DIN2 (________22953), .Q
       (____0___22742));
  nor2s1 __9____512690(.DIN1 (________22792), .DIN2 (____9___22541), .Q
       (____00__22741));
  nnd2s1 __9____512691(.DIN1 (________22977), .DIN2 (____99___36174),
       .Q (____99__22740));
  nor2s1 __9___512692(.DIN1 (________22615), .DIN2 (____0___22942), .Q
       (____9___22739));
  or2s1 __9____512693(.DIN1 (____0________________21717), .DIN2
       (________22867), .Q (____9___22738));
  nor2s1 __9____512694(.DIN1 (_____9__22422), .DIN2 (_________38838),
       .Q (____9___22737));
  or2s1 __9____512695(.DIN1 (_____0__23095), .DIN2 (________22973), .Q
       (____9___22736));
  xnr2s1 __9____512696(.DIN1 (_________________0___21702), .DIN2
       (____9___22734), .Q (____9___22735));
  nor2s1 __9____512697(.DIN1 (____0________________21662), .DIN2
       (____0___22942), .Q (____9___22733));
  or2s1 __9____512698(.DIN1 (_____________________21745), .DIN2
       (________22953), .Q (____9___22732));
  nnd2s1 __9____512699(.DIN1 (_______22253), .DIN2 (____9___23591), .Q
       (____90__22731));
  nor2s1 __9__0_512700(.DIN1 (_____0__22711), .DIN2 (________23080), .Q
       (_____9__22730));
  nnd2s1 __9____512701(.DIN1 (________22856), .DIN2 (________22857), .Q
       (________22729));
  nor2s1 __9____512702(.DIN1 (________22727), .DIN2 (________22965), .Q
       (________22728));
  or2s1 __9_9_512703(.DIN1 (________22725), .DIN2 (________22724), .Q
       (________22726));
  xnr2s1 __9___512704(.DIN1 (_____0__22681), .DIN2
       (__________________________________________0_), .Q
       (________22723));
  and2s1 __9____512705(.DIN1 (________22887), .DIN2
       (_____________________21708), .Q (________22722));
  nor2s1 __9____512706(.DIN1 (____0_______________), .DIN2
       (____0___22362), .Q (_____0__22721));
  and2s1 __9099_512707(.DIN1 (___9____26034), .DIN2
       (_____________22088), .Q (_____9__22720));
  and2s1 __9____512708(.DIN1 (____0___22364), .DIN2
       (_____________________21672), .Q (________22719));
  nor2s1 __9____512709(.DIN1 (____0___23697), .DIN2 (________22717), .Q
       (________22718));
  nor2s1 __9____512710(.DIN1 (___0____22325), .DIN2 (____0___23412), .Q
       (________22716));
  nor2s1 __9__9_512711(.DIN1 (____0___23697), .DIN2 (____09__22848), .Q
       (________23443));
  nnd2s1 __9_9_512712(.DIN1 (________22715), .DIN2 (____0___22846), .Q
       (___0____23254));
  and2s1 __9_9__512713(.DIN1 (________22715), .DIN2
       (_____________________21694), .Q (________23421));
  nnd2s1 __9_9__512714(.DIN1 (________24544), .DIN2 (________22678), .Q
       (___0_0__23263));
  nor2s1 __9_9_512715(.DIN1 (___0____22320), .DIN2 (________22871), .Q
       (____99__23406));
  or2s1 __9_90_512716(.DIN1 (______________________21700), .DIN2
       (____9___22542), .Q (___0____23257));
  nnd2s1 __9____512717(.DIN1 (________25569), .DIN2 (________22535), .Q
       (___9____23177));
  nor2s1 __9___512718(.DIN1 (___9____26912), .DIN2 (________25438), .Q
       (________23023));
  nnd2s1 __9_90_512719(.DIN1 (________22698), .DIN2 (________22532), .Q
       (________23439));
  nnd2s1 __9_0__512720(.DIN1 (____9___26583), .DIN2 (________22714), .Q
       (________23020));
  nnd2s1 __9___512721(.DIN1 (___9____24123), .DIN2 (____9___26583), .Q
       (____0___23044));
  nnd2s1 __9____512722(.DIN1 (____9___22933), .DIN2 (________23089), .Q
       (___0____23239));
  and2s1 __9__9_512723(.DIN1 (________24884), .DIN2
       (_________________9___21696), .Q (_____0__23702));
  nnd2s1 __9_9__512724(.DIN1 (________22713), .DIN2 (________22712), .Q
       (______9__34068));
  nor2s1 __9_9__512725(.DIN1 (____90__24060), .DIN2 (_____0__22711), .Q
       (________23442));
  nor2s1 __9_9__512726(.DIN1 (________22530), .DIN2 (_____9__22710), .Q
       (____909__33345));
  nor2s1 __9_0__512727(.DIN1 (_____________________21735), .DIN2
       (________22606), .Q (________23012));
  nnd2s1 __9_9__512728(.DIN1 (________22709), .DIN2 (___0____22292), .Q
       (______0__32793));
  nor2s1 __9___512729(.DIN1 (____0___23697), .DIN2 (________22708), .Q
       (___9____25079));
  nor2s1 __9_0__512730(.DIN1 (___9____23150), .DIN2 (____9___22543), .Q
       (___9____23159));
  nnd2s1 __9____512731(.DIN1 (________22862), .DIN2 (_____9__22613), .Q
       (_____0__23009));
  nnd2s1 __9__0_512732(.DIN1 (___0____23292), .DIN2 (________22707), .Q
       (____00__23039));
  nor2s1 __9_9__512733(.DIN1 (____0___22846), .DIN2 (________22706), .Q
       (________23431));
  nnd2s1 __9_9__512734(.DIN1 (_____0__23095), .DIN2 (________22705), .Q
       (________23424));
  nnd2s1 __9_0__512735(.DIN1 (________25931), .DIN2
       (____0________________21721), .Q (___9_9));
  nnd2s1 __9_0__512736(.DIN1 (________22473), .DIN2
       (_____________________21735), .Q (___0____23267));
  and2s1 __9__512737(.DIN1 (________23006), .DIN2 (_____9__25368), .Q
       (_____0__24487));
  nor2s1 __9_9_512738(.DIN1 (____99__22838), .DIN2 (________22704), .Q
       (________23523));
  or2s1 __9_9__512739(.DIN1 (______22153), .DIN2 (________22717), .Q
       (________23724));
  and2s1 __9____512740(.DIN1 (________22762), .DIN2
       (_____________________21691), .Q (________23566));
  and2s1 __9___512741(.DIN1 (____9___26583), .DIN2 (________22855), .Q
       (___9_0__25095));
  nor2s1 __9__512742(.DIN1 (________24300), .DIN2 (____0___22845), .Q
       (____9___23588));
  nnd2s1 __9_0__512743(.DIN1 (________22703), .DIN2 (____0____37167),
       .Q (________23452));
  nor2s1 __9___512744(.DIN1 (________26419), .DIN2 (_____0__26149), .Q
       (________23953));
  nnd2s1 __9_0__512745(.DIN1 (____0___22366), .DIN2
       (____0_____________0_), .Q (________23418));
  nnd2s1 __9____512746(.DIN1 (________22862), .DIN2 (___9____23167), .Q
       (________25356));
  nor2s1 __9___512747(.DIN1 (___0____23252), .DIN2 (______22153), .Q
       (____0___23509));
  nnd2s1 __9___512748(.DIN1 (_____9__22383), .DIN2 (________22885), .Q
       (_____9__25280));
  nnd2s1 __9_9__512749(.DIN1 (________23006), .DIN2 (________22727), .Q
       (________23347));
  nor2s1 __9_9_512750(.DIN1 (____9___23032), .DIN2 (____99__22838), .Q
       (________23440));
  nnd2s1 __9_9_512751(.DIN1 (________22534), .DIN2 (________22714), .Q
       (________23759));
  nor2s1 __9_9__512752(.DIN1 (_________________9___21711), .DIN2
       (________22695), .Q (________23427));
  nnd2s1 __9_9_512753(.DIN1 (____9___23786), .DIN2 (________22389), .Q
       (________25726));
  nor2s1 __9____512754(.DIN1 (_____________________21678), .DIN2
       (________22381), .Q (___90___24076));
  nnd2s1 __9__9_512755(.DIN1 (________22702), .DIN2 (________22818), .Q
       (________23805));
  and2s1 __9__0_512756(.DIN1 (___9____23152), .DIN2
       (_____________________21669), .Q (________23434));
  nnd2s1 __9__9_512757(.DIN1 (____0___22847), .DIN2 (____9___23970), .Q
       (________24341));
  and2s1 __9_9__512758(.DIN1 (____9___23786), .DIN2
       (_____________________21680), .Q (_____0__24411));
  nnd2s1 __9_9__512759(.DIN1 (________22973), .DIN2 (________23024), .Q
       (________23583));
  nnd2s1 __9_9__512760(.DIN1 (________26618), .DIN2 (________26431), .Q
       (___0____23268));
  nor2s1 __9__512761(.DIN1 (_____9__23842), .DIN2 (_________35677), .Q
       (________23450));
  and2s1 __9_9__512762(.DIN1 (___90____39055), .DIN2 (________22872),
       .Q (____0___24269));
  or2s1 __9_9__512763(.DIN1 (____0___22555), .DIN2 (________23080), .Q
       (____09__25871));
  or2s1 __9_9__512764(.DIN1 (____0_____________0___21723), .DIN2
       (_____0__22701), .Q (________23932));
  nor2s1 __9_0_512765(.DIN1 (_____9__23900), .DIN2 (____9___22837), .Q
       (____9___23500));
  nor2s1 __9__9_512766(.DIN1 (_____9__23842), .DIN2 (____9___22547), .Q
       (_____0__23910));
  nor2s1 __9_9__512767(.DIN1 (_____________________21694), .DIN2
       (_____9__22478), .Q (____9___23400));
  or2s1 __9_9__512768(.DIN1 (____________________), .DIN2
       (________26419), .Q (________23485));
  nor2s1 __9__9_512769(.DIN1 (_____9__24635), .DIN2 (___990), .Q
       (___0____23299));
  nor2s1 __9____512770(.DIN1 (________22852), .DIN2 (____0___22942), .Q
       (________24699));
  nor2s1 __9____512771(.DIN1 (________22852), .DIN2 (________24300), .Q
       (____0___23603));
  or2s1 __9_0_512772(.DIN1 (____0___22843), .DIN2 (_____9__22623), .Q
       (________25510));
  nor2s1 __9_0__512773(.DIN1 (_____________________21694), .DIN2
       (________22795), .Q (________24351));
  nnd2s1 __9_99_512774(.DIN1 (_____9__22700), .DIN2
       (_____________________21729), .Q (______0__35181));
  or2s1 __9_990(.DIN1 (____0________________21719), .DIN2
       (___9____23147), .Q (_____9__23425));
  and2s1 __9_9__512775(.DIN1 (________22699), .DIN2 (________22698), .Q
       (________23752));
  nnd2s1 __9____512776(.DIN1 (________22629), .DIN2 (___99___26049), .Q
       (________24632));
  nnd2s1 __9____512777(.DIN1 (________22862), .DIN2 (____0___22847), .Q
       (___9_9__25047));
  nor2s1 __9____512778(.DIN1 (________22697), .DIN2 (________25744), .Q
       (____0___25229));
  nnd2s1 __9_00_512779(.DIN1 (___90____39055), .DIN2 (________22696),
       .Q (____00__24267));
  nnd2s1 __9___512780(.DIN1 (________22862), .DIN2 (____9___23782), .Q
       (___9____26019));
  nor2s1 __9___512781(.DIN1 (____0_________________21725), .DIN2
       (___0___22276), .Q (___0____26064));
  nor2s1 __9_0__512782(.DIN1 (________22695), .DIN2 (_______22251), .Q
       (________23667));
  nnd2s1 __9_9__512783(.DIN1 (________22818), .DIN2 (________22699), .Q
       (________24711));
  nnd2s1 __9_00_512784(.DIN1 (____0___23311), .DIN2 (____9___22833), .Q
       (________23860));
  nnd2s1 __9_0__512785(.DIN1 (________24884), .DIN2 (________22380), .Q
       (________24280));
  nnd2s1 __9_0_512786(.DIN1 (________22762), .DIN2
       (_____________________21689), .Q (_____9__23482));
  nnd2s1 __9_0__512787(.DIN1 (________22864), .DIN2 (___00__22272), .Q
       (________23538));
  nnd2s1 __9_512788(.DIN1 (________22715), .DIN2
       (_____________________21695), .Q (____9___24455));
  and2s1 __9_0__512789(.DIN1 (____09__22458), .DIN2
       (_____________________21679), .Q (___9____24134));
  and2s1 __9___512790(.DIN1 (________22694), .DIN2 (________26618), .Q
       (________25343));
  nnd2s1 __9_00_512791(.DIN1 (________22702), .DIN2 (________22698), .Q
       (________23946));
  or2s1 __9____512792(.DIN1 (________26431), .DIN2 (________23391), .Q
       (________24791));
  nnd2s1 __9____512793(.DIN1 (_____9__22700), .DIN2 (_____9__25368), .Q
       (________24659));
  nnd2s1 __9_0__512794(.DIN1 (____9___24062), .DIN2 (_____0__22691), .Q
       (________23451));
  or2s1 __9_0__512795(.DIN1 (____0________________21719), .DIN2
       (____9___23037), .Q (_____0__25319));
  nor2s1 __9_0__512796(.DIN1 (________22704), .DIN2 (_____9__23900), .Q
       (________24398));
  and2s1 __9_0__512797(.DIN1 (_____0__23095), .DIN2
       (____0________________21719), .Q (________24415));
  nor2s1 __9____512798(.DIN1 (_____________________21684), .DIN2
       (________22693), .Q (____0___23413));
  nnd2s1 __9_0__512799(.DIN1 (____90__23962), .DIN2 (________22387), .Q
       (________25327));
  nnd2s1 __9____512800(.DIN1 (___9_9__25977), .DIN2 (________22694), .Q
       (_____9__25632));
  nnd2s1 __9_0_512801(.DIN1 (_____0__22624), .DIN2 (____0___23412), .Q
       (____0___24564));
  nor2s1 __9_0_512802(.DIN1 (____0________________21714), .DIN2
       (________22856), .Q (________23423));
  or2s1 __9_0__512803(.DIN1 (________24475), .DIN2 (________23618), .Q
       (________23715));
  nnd2s1 __9_0__512804(.DIN1 (________22702), .DIN2 (________22399), .Q
       (________24338));
  and2s1 __9_0__512805(.DIN1 (________22630), .DIN2 (________23618), .Q
       (____9_9__37984));
  nor2s1 __9____512806(.DIN1 (_____9__22518), .DIN2 (________24544), .Q
       (_____9___35917));
  nor2s1 __9____512807(.DIN1 (_____________________21683), .DIN2
       (______22153), .Q (________23580));
  nnd2s1 __9_0__512808(.DIN1 (____9___22832), .DIN2 (________22692), .Q
       (_________36527));
  nnd2s1 __9_0__512809(.DIN1 (_____9__23028), .DIN2 (_____0__22810), .Q
       (________24883));
  nnd2s1 __9_0__512810(.DIN1 (____0___22845), .DIN2 (____9___22832), .Q
       (____0____36215));
  nnd2s1 __9_0__512811(.DIN1 (________22626), .DIN2 (________23021), .Q
       (_________38533));
  nnd2s1 __9___512812(.DIN1 (________22955), .DIN2
       (____0________________21662), .Q (________24727));
  nor2s1 __9____512813(.DIN1 (____0____37167), .DIN2 (________22434),
       .Q (_________38583));
  nor2s1 __9____512814(.DIN1 (________22618), .DIN2 (_____9__22918), .Q
       (____0___24466));
  nor2s1 __9_0__512815(.DIN1 (______________________21752), .DIN2
       (_____0__22691), .Q (_________34145));
  or2s1 __9_0_512816(.DIN1 (____0________________21721), .DIN2
       (________23092), .Q (_____9__25927));
  nor2s1 __9____512817(.DIN1 (_____9__24635), .DIN2 (____0___22942), .Q
       (________23518));
  nnd2s1 __9_0__512818(.DIN1 (_____9__22690), .DIN2 (________22689), .Q
       (____0____33482));
  and2s1 __9__9_512819(.DIN1 (___9____23156), .DIN2 (_____0__22810), .Q
       (________25332));
  nnd2s1 __9____512820(.DIN1 (____0___22845), .DIN2 (____0___23599), .Q
       (_________36349));
  nnd2s1 __9__0_512821(.DIN1 (_____9__23028), .DIN2 (___9____23152), .Q
       (________26576));
  nor2s1 __9___512822(.DIN1 (____0________________21662), .DIN2
       (________22866), .Q (________25373));
  nnd2s1 __9_0__512823(.DIN1 (________24625), .DIN2 (___9____26912), .Q
       (___0____26067));
  nnd2s1 __9_09_512824(.DIN1 (________22533), .DIN2
       (______________________21701), .Q (______0__38256));
  nnd2s1 __9_0_512825(.DIN1 (____0___23414), .DIN2 (________22495), .Q
       (_________35663));
  hi1s1 __9_9__512826(.DIN (___9_____39627), .Q (______0__34897));
  hi1s1 __9____512827(.DIN (________25740), .Q (________27288));
  nnd2s1 __9_0__512828(.DIN1 (________22864), .DIN2
       (____0________________21714), .Q (___9_____39746));
  nnd2s1 __9_0__512829(.DIN1 (_____9__22442), .DIN2 (________22496), .Q
       (___9__9__39659));
  nor2s1 __9__0_512830(.DIN1 (________22851), .DIN2 (________22965), .Q
       (___90___25034));
  nor2s1 __9_0__512831(.DIN1 (________22594), .DIN2 (________23469), .Q
       (_________35680));
  nnd2s1 __9_09_512832(.DIN1 (____90__23962), .DIN2 (______22147), .Q
       (______0__37673));
  hi1s1 __9____512833(.DIN (___900__24070), .Q (________25944));
  nor2s1 __9_0__512834(.DIN1 (_____0__22691), .DIN2 (_____9__22828), .Q
       (___9_9___39339));
  nor2s1 __9___512835(.DIN1 (_________________9_), .DIN2
       (________24703), .Q (________22688));
  xor2s1 __9__9_512836(.DIN1
       (_________________________________________0___21840), .DIN2
       (_________37245), .Q (________22687));
  nnd2s1 __9____512837(.DIN1 (___0____23248), .DIN2 (________24602), .Q
       (________22686));
  and2s1 __9____512838(.DIN1 (____0___23311), .DIN2
       (____0________________21719), .Q (________22685));
  hi1s1 __9___512839(.DIN (________22683), .Q (________22684));
  nnd2s1 __9____512840(.DIN1 (_____0__22681), .DIN2 (_____22117), .Q
       (________22682));
  nnd2s1 __9____512841(.DIN1 (________22679), .DIN2 (________22678), .Q
       (_____9__22680));
  nor2s1 __9____512842(.DIN1 (____00__23597), .DIN2 (____0___23311), .Q
       (________22677));
  nor2s1 __9___512843(.DIN1 (____0__22235), .DIN2 (________22675), .Q
       (________22676));
  and2s1 __9____512844(.DIN1 (____9___22734), .DIN2
       (_____________________21704), .Q (________22674));
  nor2s1 __9____512845(.DIN1 (___0____23252), .DIN2 (________22672), .Q
       (________22673));
  nor2s1 __9____512846(.DIN1 (_____0__22384), .DIN2 (____9___24062), .Q
       (_____0__22671));
  or2s1 __9___512847(.DIN1 (________22669), .DIN2 (____9___25949), .Q
       (________22670));
  hi1s1 __9____512848(.DIN (________22667), .Q (________22668));
  xor2s1 __9__9_512849(.DIN1
       (_____________________________________________21810), .DIN2
       (___0_____30948), .Q (________22665));
  nor2s1 __9____512850(.DIN1 (___0_____40515), .DIN2 (_______22210), .Q
       (________22664));
  nor2s1 __9_9__512851(.DIN1 (_____9__22662), .DIN2 (________22661), .Q
       (_____0__22663));
  xor2s1 __9___512852(.DIN1
       (_________________________________________9___21855), .DIN2
       (_________36762), .Q (________22660));
  xor2s1 __9____512853(.DIN1 (_________22042), .DIN2 (_____00__35736),
       .Q (________22659));
  xor2s1 __9____512854(.DIN1 (___0_____30948), .DIN2 (_________36761),
       .Q (________22658));
  nnd2s1 __9____512855(.DIN1 (__9___22166), .DIN2
       (_________________________________________________________________22001),
       .Q (________22657));
  and2s1 __9___512856(.DIN1 (_________38649), .DIN2 (___9___22194), .Q
       (________22656));
  or2s1 __9_900(.DIN1 (________22513), .DIN2 (____9___22734), .Q
       (________22655));
  xor2s1 __9____512857(.DIN1 (_________22042), .DIN2 (_________37245),
       .Q (____09__22653));
  nor2s1 __9____512858(.DIN1 (_____________________21682), .DIN2
       (____90__22539), .Q (____0___22652));
  and2s1 __9____512859(.DIN1 (___0____23248), .DIN2
       (_____________________21709), .Q (____0___22651));
  hi1s1 __9____512860(.DIN (_____9__22858), .Q (____0___22650));
  nor2s1 __9____512861(.DIN1 (____09__23048), .DIN2 (____0___22648), .Q
       (____0___22649));
  nor2s1 __9__9_512862(.DIN1 (_________35727), .DIN2 (___0___22197), .Q
       (____0___22647));
  and2s1 __9___512863(.DIN1 (___9____23150), .DIN2
       (____0________________21720), .Q (____0___22646));
  xor2s1 __9___512864(.DIN1
       (____________________________________________21866), .DIN2
       (______9__32959), .Q (____0___22645));
  nnd2s1 __9___512865(.DIN1 (____0__22225), .DIN2 (clk), .Q
       (____00__22644));
  hi1s1 __9____512866(.DIN (________22818), .Q (____99__22643));
  or2s1 __9____512867(.DIN1 (_________35727), .DIN2 (____9___22641), .Q
       (____9___22642));
  and2s1 __9____512868(.DIN1 (________25942), .DIN2 (___0____25161), .Q
       (____9___22640));
  nor2s1 __9___512869(.DIN1 (_______22245), .DIN2 (___9___22190), .Q
       (____9___22639));
  hi1s1 __9___512870(.DIN (___9____23147), .Q (____9___22638));
  xor2s1 __9___512871(.DIN1 (____9___22636), .DIN2 (___0_____40575), .Q
       (____9___22637));
  hi1s1 __9____512872(.DIN (________22693), .Q (____9___22635));
  xor2s1 __9____512873(.DIN1 (___0_____40448), .DIN2 (_____9__22633),
       .Q (____90__22634));
  hi1s1 __9___512874(.DIN (________22632), .Q (________23015));
  hi1s1 __9____512875(.DIN (________22631), .Q (________23087));
  nor2s1 __9_9__512876(.DIN1 (________22388), .DIN2 (____0___23042), .Q
       (_____9__23104));
  hi1s1 __9___512877(.DIN (________22630), .Q (___9____23162));
  hi1s1 __9____512878(.DIN (________22629), .Q (____9___23031));
  and2s1 __9_90_512879(.DIN1 (____0___25498), .DIN2
       (_________________0___21687), .Q (________23111));
  and2s1 __9____512880(.DIN1 (____0___23412), .DIN2
       (_________________9___21737), .Q (___9____23161));
  or2s1 __9_9__512881(.DIN1 (____0________________21721), .DIN2
       (________25756), .Q (___9____23146));
  nor2s1 __9_9_512882(.DIN1 (________22628), .DIN2 (____9___24062), .Q
       (________23335));
  nor2s1 __9__9_512883(.DIN1 (________22627), .DIN2 (_____9__23376), .Q
       (________23010));
  hi1s1 __9____512884(.DIN (________22626), .Q (________23013));
  hi1s1 __9_9__512885(.DIN (___9_____39461), .Q (________23025));
  nnd2s1 __9_9__512886(.DIN1 (____0___25498), .DIN2 (________22884), .Q
       (____0___23045));
  and2s1 __9_9__512887(.DIN1 (________22625), .DIN2 (________22679), .Q
       (___9____24083));
  nor2s1 __9_9__512888(.DIN1 (________24602), .DIN2 (_____9__23900), .Q
       (___0____23247));
  nnd2s1 __9_9__512889(.DIN1 (________25942), .DIN2 (________26431), .Q
       (________23894));
  hi1s1 __9___512890(.DIN (_____0__22624), .Q (____9___23033));
  or2s1 __9__0_512891(.DIN1 (________22860), .DIN2 (________24703), .Q
       (____0___23600));
  hi1s1 __9_9__512892(.DIN (________23092), .Q (________23072));
  hi1s1 __9____512893(.DIN (_____0__22849), .Q (____99__23133));
  hi1s1 __9____512894(.DIN (___0____26080), .Q (___9_9__26020));
  nor2s1 __9_9_512895(.DIN1 (_____9___37752), .DIN2 (________22689), .Q
       (___9____23160));
  hi1s1 __9____512896(.DIN (____0___22845), .Q (________23083));
  hi1s1 __9____512897(.DIN (_____9__22623), .Q (___9____23148));
  hi1s1 __9____512898(.DIN (________22708), .Q (____0___24464));
  and2s1 __9_99_512899(.DIN1 (___0____23248), .DIN2 (____9___23032), .Q
       (___9____23207));
  hi1s1 __9_90_512900(.DIN (________22622), .Q (________23081));
  or2s1 __9_9_512901(.DIN1 (_____________________21735), .DIN2
       (________22472), .Q (___9____23144));
  hi1s1 __9_90_512902(.DIN (________22621), .Q (___0____23228));
  hi1s1 __9____512903(.DIN (____0___23504), .Q (___9____23169));
  hi1s1 __9____512904(.DIN (____9___23036), .Q (___999));
  or2s1 __9____512905(.DIN1 (___9____23149), .DIN2 (________22672), .Q
       (___9____23197));
  hi1s1 __9___512906(.DIN (____9___24360), .Q (________24013));
  hi1s1 __9____512907(.DIN (________22620), .Q (___9____23170));
  nnd2s1 __9____512908(.DIN1 (____0_______________), .DIN2
       (____90__24060), .Q (________23330));
  hi1s1 __9_512909(.DIN (________22619), .Q (________24768));
  hi1s1 __9____512910(.DIN (________25744), .Q (____0___26415));
  hi1s1 __9_90_512911(.DIN (________22618), .Q (___9____23158));
  hi1s1 __9_9__512912(.DIN (____0___22841), .Q (________25508));
  hi1s1 __9____512913(.DIN (________22617), .Q (________25352));
  hi1s1 __9_9__512914(.DIN (______9__36337), .Q (________24760));
  hi1s1 __9_9__512915(.DIN (________22955), .Q (___99_));
  hi1s1 __9____512916(.DIN (________22865), .Q (________23075));
  hi1s1 __9_9_512917(.DIN (________22697), .Q (________25605));
  nor2s1 __9_0__512918(.DIN1 (_____________________21684), .DIN2
       (________22672), .Q (________23327));
  hi1s1 __9_9__512919(.DIN (________22616), .Q (________23662));
  nor2s1 __9____512920(.DIN1 (_________________9___21737), .DIN2
       (________22689), .Q (________23552));
  hi1s1 __9____512921(.DIN (________22977), .Q (_____0__23852));
  hi1s1 __9____512922(.DIN (________22615), .Q (________23517));
  hi1s1 __9__9_512923(.DIN (________22973), .Q (________23726));
  hi1s1 __9__512924(.DIN (___990), .Q (________23535));
  hi1s1 __9____512925(.DIN (____0___23602), .Q (___99___26045));
  hi1s1 __9___512926(.DIN (_____0__22614), .Q (___99___23210));
  hi1s1 __9____512927(.DIN (_____9__22613), .Q (____0___26410));
  nor2s1 __9_0__512928(.DIN1 (_____________________21704), .DIN2
       (_______22227), .Q (___00___25129));
  xor2s1 __9____512929(.DIN1 (________22611), .DIN2
       (______________________________________0_______21890), .Q
       (________22612));
  hi1s1 __9____512930(.DIN (________22609), .Q (________22610));
  hi1s1 __9____512931(.DIN (________22606), .Q (________22607));
  xor2s1 __9____512932(.DIN1 (___0____23297), .DIN2 (______9__32959),
       .Q (_____0__22605));
  nnd2s1 __9__9_512933(.DIN1 (________22672), .DIN2 (___9____23149), .Q
       (_____9__22604));
  xor2s1 __9____512934(.DIN1 (_____9__23492), .DIN2 (_________22038),
       .Q (________22603));
  nnd2s1 __9____512935(.DIN1 (________22599), .DIN2 (_______22241), .Q
       (________22600));
  xor2s1 __9____512936(.DIN1 (___0_____40479), .DIN2
       (______________22066), .Q (________22598));
  and2s1 __9___512937(.DIN1 (____0___25498), .DIN2
       (_____________________21690), .Q (_____0__22597));
  xor2s1 __9____512938(.DIN1
       (_____________________________________________21796), .DIN2
       (_________33591), .Q (_____9__22596));
  nnd2s1 __9____512939(.DIN1 (________22594), .DIN2 (________26426), .Q
       (________22595));
  hi1s1 __9____512940(.DIN (________22592), .Q (________22593));
  nor2s1 __9_9_512941(.DIN1 (________22590), .DIN2 (________22589), .Q
       (________22591));
  xor2s1 __9___512942(.DIN1
       (__________________________________________0___21935), .DIN2
       (___0_____40045), .Q (________22588));
  and2s1 __9____512943(.DIN1 (_____0__22899), .DIN2 (____09__23048), .Q
       (_____9__22587));
  or2s1 __9___512944(.DIN1 (_________________0___21728), .DIN2
       (____0___22743), .Q (________22586));
  nnd2s1 __9___512945(.DIN1 (____9___22546), .DIN2
       (______________________21699), .Q (________22585));
  hi1s1 __9____512946(.DIN (________22583), .Q (________22584));
  hi1s1 __9___512947(.DIN (________22581), .Q (________22582));
  nnd2s1 __9____512948(.DIN1 (_____9___38319), .DIN2
       (_____________________21747), .Q (________22580));
  nor2s1 __9____512949(.DIN1 (________26530), .DIN2 (______22160), .Q
       (________22579));
  xor2s1 __9___512950(.DIN1 (_____9__22577), .DIN2 (___0__0__40421), .Q
       (_____0__22578));
  xor2s1 __9____512951(.DIN1 (______________22064), .DIN2
       (_________32918), .Q (________22576));
  xor2s1 __9____512952(.DIN1 (___0_____40523), .DIN2 (________27043),
       .Q (________22575));
  hi1s1 __9____512953(.DIN (___9____23152), .Q (________22574));
  nor2s1 __9____512954(.DIN1 (___0__9__40430), .DIN2 (_________38838),
       .Q (________22573));
  nor2s1 __9___512955(.DIN1 (_____9__22868), .DIN2 (________24300), .Q
       (________22572));
  nnd2s1 __9__9_512956(.DIN1 (________22860), .DIN2 (____0___23042), .Q
       (________22571));
  hi1s1 __9___512957(.DIN (________22876), .Q (________22570));
  or2s1 __9___512958(.DIN1 (_______22218), .DIN2 (________22984), .Q
       (________22569));
  xor2s1 __9__512959(.DIN1 (_____9__22567), .DIN2
       (__________9___22107), .Q (_____0__22568));
  or2s1 __9____512960(.DIN1 (_____________________21744), .DIN2
       (____0___22648), .Q (________22566));
  hi1s1 __9____512961(.DIN (________22564), .Q (________22565));
  nor2s1 __9____512962(.DIN1 (______9__22030), .DIN2 (________28146),
       .Q (________22563));
  xor2s1 __9___512963(.DIN1 (___0__9__40510), .DIN2 (________22561), .Q
       (________22562));
  nor2s1 __9__9_512964(.DIN1 (_____0__22559), .DIN2 (____09__22558), .Q
       (________22560));
  and2s1 __9____512965(.DIN1 (_____9__23028), .DIN2
       (_____________________21672), .Q (____0___22557));
  nor2s1 __9____512966(.DIN1 (____90__24060), .DIN2 (____0___22555), .Q
       (____0___22556));
  hi1s1 __9____512967(.DIN (________23080), .Q (____0___22554));
  xor2s1 __9____512968(.DIN1 (_______________22074), .DIN2
       (_________37789), .Q (____0___22553));
  nnd2s1 __9____512969(.DIN1 (___0___22200), .DIN2
       (______________________________________________21912), .Q
       (____0___22552));
  xor2s1 __9____512970(.DIN1 (______________22064), .DIN2
       (_________32611), .Q (____0___22551));
  nnd2s1 __9__9_512971(.DIN1 (________22689), .DIN2
       (_________________9___21737), .Q (____0___22550));
  xor2s1 __9____512972(.DIN1
       (____________________________________________21791), .DIN2
       (_____0___33534), .Q (____00__22549));
  nnd2s1 __9_0_512973(.DIN1 (____99__22548), .DIN2 (_____9__22402), .Q
       (____9___22836));
  nor2s1 __9_9__512974(.DIN1 (________23449), .DIN2 (____9___22546), .Q
       (________23011));
  or2s1 __9_9__512975(.DIN1 (____0________________21721), .DIN2
       (___9____23150), .Q (_____9__23008));
  hi1s1 __9_9__512976(.DIN (________25931), .Q (________23093));
  nnd2s1 __9_9__512977(.DIN1 (________22696), .DIN2 (____9___22545), .Q
       (___9____23166));
  hi1s1 __9__9_512978(.DIN (________23066), .Q (____0___23601));
  nor2s1 __9_9__512979(.DIN1 (_____________________21743), .DIN2
       (____0___22648), .Q (_____9__22760));
  nnd2s1 __9_9__512980(.DIN1 (____0___23412), .DIN2 (_____9___37752),
       .Q (_____0__22879));
  hi1s1 __9_9__512981(.DIN (____9___22547), .Q (___090__23301));
  nor2s1 __9__512982(.DIN1 (_____________________21730), .DIN2
       (________23384), .Q (________22877));
  hi1s1 __9_9__512983(.DIN (____9___22547), .Q (________23513));
  and2s1 __9__9_512984(.DIN1 (________22679), .DIN2
       (____0_____________0_), .Q (____9___23035));
  nnd2s1 __9____512985(.DIN1 (____9___22544), .DIN2 (______22155), .Q
       (________23069));
  nnd2s1 __9_9_512986(.DIN1 (___9____24088), .DIN2 (________23734), .Q
       (___0____23269));
  hi1s1 __9__9_512987(.DIN (____9___22543), .Q (____9___23030));
  nor2s1 __9_9__512988(.DIN1 (________23734), .DIN2 (________23384), .Q
       (________23903));
  nor2s1 __9_99_512989(.DIN1 (______________________21699), .DIN2
       (____9___22546), .Q (________23022));
  hi1s1 __9____512990(.DIN (____9___23592), .Q (________23065));
  nnd2s1 __9_0_512991(.DIN1 (____9___22933), .DIN2
       (____0________________21662), .Q (___900__24070));
  or2s1 __9____512992(.DIN1 (________26431), .DIN2 (____0___22648), .Q
       (________23515));
  nnd2s1 __9__0_512993(.DIN1 (____9___23782), .DIN2 (___9____23151), .Q
       (___9_0));
  nor2s1 __9_9__512994(.DIN1 (_____________________21682), .DIN2
       (_____9__23376), .Q (________24824));
  hi1s1 __9____512995(.DIN (____9___22542), .Q (___9_9__23172));
  or2s1 __9_9__512996(.DIN1 (_____________________21690), .DIN2
       (____0___22843), .Q (________23481));
  hi1s1 __9____512997(.DIN (____9___22541), .Q (___9____23190));
  hi1s1 __9___512998(.DIN (____9___22540), .Q (___9____23165));
  hi1s1 __9_9__512999(.DIN (____9___22547), .Q (___00____41368));
  nor2s1 __9_0_513000(.DIN1 (___9____23149), .DIN2 (____90__22539), .Q
       (___0____23236));
  hi1s1 __9____513001(.DIN (_____9__22538), .Q (_____0__23077));
  and2s1 __9_00_513002(.DIN1 (___0____23248), .DIN2
       (_____________________21707), .Q (___9_9__23154));
  nor2s1 __9_9__513003(.DIN1 (_____9__24325), .DIN2 (________23384), .Q
       (___9____23143));
  nnd2s1 __9_99_513004(.DIN1 (_________38301), .DIN2 (_____9__23842),
       .Q (________23916));
  hi1s1 __9____513005(.DIN (________22537), .Q (_________32663));
  nnd2s1 __9_0__513006(.DIN1 (____99__22548), .DIN2
       (_____________________21704), .Q (___0_0__25155));
  and2s1 __9_0__513007(.DIN1 (_____0__22899), .DIN2
       (_____________________21743), .Q (________25337));
  nor2s1 __9_0__513008(.DIN1 (___0____23252), .DIN2 (____90__22539), .Q
       (___9____23175));
  hi1s1 __9____513009(.DIN (_____0__22859), .Q (___99___23213));
  nnd2s1 __9_0_513010(.DIN1 (_______22187), .DIN2
       (____0________________21668), .Q (_________38591));
  nor2s1 __9____513011(.DIN1 (________22536), .DIN2 (____0___22555), .Q
       (________25740));
  hi1s1 __9_9__513012(.DIN (________22535), .Q (___0____25163));
  hi1s1 __9____513013(.DIN (___9____23167), .Q (____9___26581));
  or2s1 __9_0__513014(.DIN1 (____9___23032), .DIN2 (_____9__23900), .Q
       (___99___24165));
  hi1s1 __9___513015(.DIN (________22798), .Q (________23101));
  hi1s1 __9____513016(.DIN (________22534), .Q (___00___26054));
  hi1s1 __9__9_513017(.DIN (________22533), .Q (_____99__36913));
  hi1s1 __9_9__513018(.DIN (________25925), .Q (________26433));
  hi1s1 __9____513019(.DIN (________22853), .Q (________26272));
  nnd2s1 __9_0__513020(.DIN1 (________22390), .DIN2 (________22532), .Q
       (_____9___38412));
  nor2s1 __9____513021(.DIN1 (___9_____39397), .DIN2
       (___________________), .Q (___9_____39627));
  hi1s1 __9____513022(.DIN (________22530), .Q (________22531));
  nor2s1 __9____513023(.DIN1 (____0_0__38093), .DIN2 (_________36883),
       .Q (_____0__22529));
  xor2s1 __9____513024(.DIN1
       (_____________________________________________21787), .DIN2
       (_________________________________________9_), .Q
       (_____9__22528));
  nor2s1 __9____513025(.DIN1 (___0____22300), .DIN2
       (______________22105), .Q (________22527));
  nor2s1 __9____513026(.DIN1 (_____9__23444), .DIN2
       (_________________0___21687), .Q (________22526));
  nor2s1 __9____513027(.DIN1 (________22524), .DIN2 (___0_____40495),
       .Q (________22525));
  xor2s1 __9____513028(.DIN1 (_______________22076), .DIN2
       (_____________________________________________21859), .Q
       (________22523));
  nnd2s1 __9_9__513029(.DIN1 (_________37412), .DIN2 (________27043),
       .Q (________22522));
  nnd2s1 __9_9__513030(.DIN1 (_____9___37752), .DIN2 (inData[27]), .Q
       (________22521));
  xor2s1 __9____513031(.DIN1 (___0_____40417), .DIN2 (___0_____40418),
       .Q (________22520));
  nor2s1 __9_99_513032(.DIN1 (___0____22346), .DIN2
       (______________22111), .Q (_____0__22519));
  nor2s1 __9____513033(.DIN1 (________22678), .DIN2
       (____0____________9_), .Q (_____9__22518));
  and2s1 __9__0_513034(.DIN1 (_________________0___21728), .DIN2
       (_____9__24325), .Q (________22517));
  xnr2s1 __9____513035(.DIN1
       (_____________________________________________21974), .DIN2
       (___0_____40417), .Q (________22516));
  nnd2s1 __9_0__513036(.DIN1 (_____0___32287), .DIN2 (_____9___33157),
       .Q (________22515));
  nnd2s1 __9__9_513037(.DIN1 (_____________________21704), .DIN2
       (________22513), .Q (________22514));
  nor2s1 __9_0__513038(.DIN1 (_________34538), .DIN2
       (_______________22069), .Q (________22512));
  nnd2s1 __9_0__513039(.DIN1 (_____9__23492), .DIN2 (_________22038),
       .Q (________22511));
  nnd2s1 __9____513040(.DIN1 (_____________________21670), .DIN2
       (____9__22261), .Q (________22510));
  xor2s1 __9__513041(.DIN1
       (_______________________________________________________________0),
       .DIN2 (___0_____40449), .Q (_____0__22509));
  nor2s1 __9___513042(.DIN1
       (____________________________________________21866), .DIN2
       (______9__32959), .Q (_____9__22508));
  nor2s1 __9___513043(.DIN1
       (__________________________________________________________________21985),
       .DIN2 (_________35587), .Q (________22507));
  xnr2s1 __9____513044(.DIN1
       (_________________________________________0___21939), .DIN2
       (___0__0__40431), .Q (________22506));
  nor2s1 __9__513045(.DIN1 (___0_9___40455), .DIN2 (________22504), .Q
       (________22505));
  nnd2s1 __9____513046(.DIN1 (___0_____40447), .DIN2 (________22502),
       .Q (________22503));
  nnd2s1 __9_0__513047(.DIN1 (_____22115), .DIN2 (___0_0___40568), .Q
       (________22501));
  nor2s1 __9____513048(.DIN1 (_____0__22499), .DIN2 (___0_____40611),
       .Q (________22500));
  nnd2s1 __9_9__513049(.DIN1 (_______________22072), .DIN2
       (_________37321), .Q (_____9__22498));
  nnd2s1 __9_0__513050(.DIN1 (_____________________21742), .DIN2
       (________22754), .Q (________22497));
  nnd2s1 __9___513051(.DIN1 (________22857), .DIN2
       (____0____________0___21713), .Q (________22496));
  or2s1 __9___513052(.DIN1 (_________________0___21740), .DIN2
       (________26426), .Q (________22495));
  xnr2s1 __9__0_513053(.DIN1
       (__________________________________________________________________21999),
       .DIN2 (__________________________________________9___21934), .Q
       (________22494));
  nor2s1 __9_0_513054(.DIN1 (___0_____40620), .DIN2 (______22124), .Q
       (________22493));
  xnr2s1 __9__9_513055(.DIN1
       (______________________________________________21922), .DIN2
       (______________________________________________21916), .Q
       (________22492));
  nnd2s1 __9_0__513056(.DIN1
       (_________________________________________________________________________________________22091),
       .DIN2 (_________36556), .Q (________22491));
  nnd2s1 __9_00_513057(.DIN1 (____9___25676), .DIN2 (inData[18]), .Q
       (________22490));
  nor2s1 __9_0__513058(.DIN1 (_________37867), .DIN2 (_________35844),
       .Q (_____0__22489));
  nor2s1 __9____513059(.DIN1 (___0_____40589), .DIN2 (___9), .Q
       (_____9__22488));
  xor2s1 __9__9_513060(.DIN1 (___0_____40519), .DIN2 (___0_____40506),
       .Q (________22487));
  nor2s1 __9_9__513061(.DIN1 (________22485), .DIN2 (_____0___32287),
       .Q (________22486));
  xor2s1 __9____513062(.DIN1 (_____9___22050), .DIN2
       (_____________________________________0______21756), .Q
       (________22484));
  xor2s1 __9____513063(.DIN1 (___0__0__40521), .DIN2
       (_______________22075), .Q (________22483));
  xor2s1 __9___513064(.DIN1 (outData[17]), .DIN2 (outData[19]), .Q
       (________22482));
  and2s1 __9____513065(.DIN1 (___0_____40582), .DIN2 (________22480),
       .Q (________22481));
  nor2s1 __9_9__513066(.DIN1 (_________36761), .DIN2
       (_________________________________________________________________________________________22091),
       .Q (_____0__22479));
  nnd2s1 __9_9__513067(.DIN1 (________23362), .DIN2 (________23026), .Q
       (_____9__22478));
  nor2s1 __9_9__513068(.DIN1 (_________34538), .DIN2
       (_________________________________________________________________________________________22091),
       .Q (________22477));
  xnr2s1 __9____513069(.DIN1 (___0_____40503), .DIN2
       (____________________________________________21830), .Q
       (________22476));
  nnd2s1 __9_0__513070(.DIN1 (______22135), .DIN2
       (__________________________________________0___21919), .Q
       (________22475));
  nor2s1 __9_9_513071(.DIN1 (_________37789), .DIN2
       (_______________22074), .Q (________22474));
  hi1s1 __9____513072(.DIN (________22472), .Q (________22473));
  nor2s1 __9____513073(.DIN1 (________22470), .DIN2
       (_________________________________________________________________21991),
       .Q (________22471));
  xor2s1 __9____513074(.DIN1 (___0_____40512), .DIN2 (_________22038),
       .Q (_____0__22469));
  xnr2s1 __9____513075(.DIN1 (______________22110), .DIN2
       (______________22108), .Q (_____9__22468));
  nnd2s1 __9_9__513076(.DIN1 (_______________22075), .DIN2
       (______9__34981), .Q (________22467));
  nnd2s1 __9_9__513077(.DIN1
       (_________________________________________________________________________________________22095),
       .DIN2 (_________34538), .Q (________22466));
  xnr2s1 __9____513078(.DIN1
       (_____________________________________________21785), .DIN2
       (_________________________________________9___21803), .Q
       (________22465));
  xor2s1 __9__0_513079(.DIN1 (___0_____40579), .DIN2 (___0__0__40491),
       .Q (________22464));
  nnd2s1 __9_9__513080(.DIN1 (_____9___33157), .DIN2
       (____________________________________________21867), .Q
       (________22463));
  nnd2s1 __9_0_513081(.DIN1 (____0___22846), .DIN2 (________22461), .Q
       (________22462));
  nor2s1 __9_0__513082(.DIN1 (___0_9__22343), .DIN2 (_____9__22567), .Q
       (________22460));
  or2s1 __9_0__513083(.DIN1 (_______22280), .DIN2
       (______________22109), .Q (_____0__22459));
  nor2s1 __9_9__513084(.DIN1 (________22924), .DIN2 (____0___22457), .Q
       (____09__22458));
  nor2s1 __9_99_513085(.DIN1 (_____9__23492), .DIN2 (______9__31640),
       .Q (____0___22456));
  xor2s1 __9__0_513086(.DIN1
       (____________________________________________21792), .DIN2
       (___0__0__40511), .Q (____0___22455));
  nnd2s1 __9_9__513087(.DIN1 (_____9__24635), .DIN2 (_______22254), .Q
       (____0___22454));
  xor2s1 __9____513088(.DIN1 (___0_____40478), .DIN2
       (_______________22070), .Q (____0___22453));
  nnd2s1 __9____513089(.DIN1 (___0____22317), .DIN2
       (______________________________________________21938), .Q
       (____0___22452));
  nnd2s1 __9____513090(.DIN1 (_______________0), .DIN2 (____99), .Q
       (____0___22451));
  nor2s1 __9___513091(.DIN1 (____99), .DIN2 (_______________0), .Q
       (____00__22450));
  xor2s1 __9____513092(.DIN1 (_________22014), .DIN2 (___0_____40594),
       .Q (____9___22449));
  nor2s1 __9_0__513093(.DIN1 (____9___22447), .DIN2 (_________34167),
       .Q (____9___22448));
  xnr2s1 __9____513094(.DIN1 (___0__9__40420), .DIN2
       (_____________________________________________21969), .Q
       (____9___22446));
  nor2s1 __9_9__513095(.DIN1 (________22727), .DIN2 (________23734), .Q
       (____9___22445));
  xnr2s1 __9__513096(.DIN1
       (_____________________________________0______21755), .DIN2
       (_____________________________________________21852), .Q
       (____9___22444));
  xor2s1 __9____513097(.DIN1
       (______________________________________0_______21891), .DIN2
       (______________________________________0_______21889), .Q
       (____9___22443));
  xor2s1 __9____513098(.DIN1
       (_____________________________________________21770), .DIN2
       (___0_____40535), .Q (____9_));
  nor2s1 __9_9__513099(.DIN1 (______9__32959), .DIN2 (___0____23297),
       .Q (____90));
  or2s1 __9____513100(.DIN1 (____0________________21715), .DIN2
       (________22857), .Q (_____9__22442));
  and2s1 __9____513101(.DIN1 (___0_____40502), .DIN2 (_____0___33161),
       .Q (________22441));
  nor2s1 __9_0__513102(.DIN1
       (______________________________________________21930), .DIN2
       (________22439), .Q (________22440));
  xor2s1 __9____513103(.DIN1
       (__________________________________________________________________21996),
       .DIN2 (_____________22101), .Q (________22438));
  xor2s1 __9__0_513104(.DIN1 (___0_____40483), .DIN2 (___0_0___40464),
       .Q (________22437));
  xor2s1 __9___513105(.DIN1
       (______________________________________________________________________________________0__22093),
       .DIN2 (_______________22077), .Q (________22436));
  xnr2s1 __9___513106(.DIN1 (___0_____40512), .DIN2 (___0__9__40530),
       .Q (________22435));
  nor2s1 __9__9_513107(.DIN1 (____90__26673), .DIN2
       (_____________________21748), .Q (________22434));
  nor2s1 __9____513108(.DIN1 (_________33206), .DIN2 (___0_____40546),
       .Q (_____0__22433));
  nor2s1 __9_9__513109(.DIN1
       (______________________________________0__0_), .DIN2
       (______22126), .Q (_____9__22432));
  xor2s1 __9__9_513110(.DIN1 (_________0_), .DIN2 (_____________22083),
       .Q (________22431));
  xor2s1 __9____513111(.DIN1 (___0__0__40491), .DIN2
       (__________________________________________), .Q
       (________22430));
  nnd2s1 __9___513112(.DIN1 (___0_____40503), .DIN2 (________24514), .Q
       (________22429));
  xnr2s1 __9____513113(.DIN1
       (_____________________________________________21787), .DIN2
       (____________________________________________21772), .Q
       (________22428));
  nor2s1 __9____513114(.DIN1 (___0__0__40531), .DIN2 (___0), .Q
       (________22427));
  nnd2s1 __9_9_513115(.DIN1 (___________9___22071), .DIN2
       (____9___22447), .Q (________22426));
  nor2s1 __9__0_513116(.DIN1 (___0_____40573), .DIN2 (________22424),
       .Q (________22425));
  nor2s1 __9_9__513117(.DIN1 (_________36402), .DIN2
       (______________________________________________________________________________________0),
       .Q (_____0__22423));
  nor2s1 __9____513118(.DIN1 (___0_____40428), .DIN2 (____9___23878),
       .Q (_____9__22422));
  nor2s1 __9____513119(.DIN1 (________22420), .DIN2
       (_________________________________________0___21798), .Q
       (________22421));
  nor2s1 __9____513120(.DIN1 (________22678), .DIN2
       (____0________________21668), .Q (________22419));
  xor2s1 __9____513121(.DIN1 (___0_____40524), .DIN2
       (_____________________________________________21838), .Q
       (________22418));
  nor2s1 __9____513122(.DIN1 (______________22103), .DIN2 (_____22116),
       .Q (________22417));
  nor2s1 __9____513123(.DIN1 (________23026), .DIN2 (____0___22846), .Q
       (________22416));
  and2s1 __9__9_513124(.DIN1 (______9__32959), .DIN2
       (____________________________________________21866), .Q
       (________22415));
  nor2s1 __9____513125(.DIN1
       (__________________________________________0___21981), .DIN2
       (______22138), .Q (________22414));
  xnr2s1 __9__9_513126(.DIN1 (_____________22080), .DIN2
       (___0_____40588), .Q (_____0__22413));
  nor2s1 __9____513127(.DIN1 (_________33293), .DIN2 (_________32918),
       .Q (_____9__22412));
  and2s1 __9_0__513128(.DIN1 (___0_____40509), .DIN2 (________22396),
       .Q (________22411));
  nnd2s1 __9_0_513129(.DIN1 (_________32918), .DIN2
       (______________22066), .Q (________22410));
  xor2s1 __9__9_513130(.DIN1 (___0_____40597), .DIN2 (___0_____40596),
       .Q (________22409));
  nor2s1 __9__9_513131(.DIN1 (________22884), .DIN2
       (_____________________21688), .Q (________22408));
  and2s1 __9_00_513132(.DIN1 (_________36583), .DIN2 (___0__9__40500),
       .Q (________22407));
  xor2s1 __9____513133(.DIN1
       (_____________________________________________21796), .DIN2
       (___0_9___40552), .Q (________22406));
  xnr2s1 __9____513134(.DIN1
       (_____________________________________0______21755), .DIN2
       (_____90__22048), .Q (________22405));
  or2s1 __9_0__513135(.DIN1 (________22485), .DIN2
       (_____________________________________________21823), .Q
       (________22404));
  nor2s1 __9_09_513136(.DIN1 (_________33117), .DIN2 (_________33973),
       .Q (_____9__22710));
  nnd2s1 __9___513137(.DIN1 (________22401), .DIN2
       (_____________________21733), .Q (________22606));
  nnd2s1 __9____513138(.DIN1 (___9__22133), .DIN2
       (______________________________________________21955), .Q
       (________22766));
  hi1s1 __9____513139(.DIN (________25756), .Q (_____0__22999));
  nnd2s1 __9___513140(.DIN1 (__________________0___21712), .DIN2
       (________22532), .Q (________22626));
  nor2s1 __9_0__513141(.DIN1 (____9___22447), .DIN2 (___0__9__40412),
       .Q (________22874));
  nnd2s1 __9___513142(.DIN1 (_____________________21742), .DIN2
       (________26431), .Q (________22619));
  nnd2s1 __9____513143(.DIN1 (_________________9___21737), .DIN2
       (___9_9__23163), .Q (_____9__22690));
  or2s1 __9__9_513144(.DIN1 (_____0__22403), .DIN2
       (_____________________________________________21845), .Q
       (_____9__23123));
  nor2s1 __9____513145(.DIN1 (___0_____40445), .DIN2 (______22144), .Q
       (________22963));
  nor2s1 __9____513146(.DIN1 (____00__23597), .DIN2
       (____0________________21719), .Q (_____0__22614));
  or2s1 __9____513147(.DIN1 (____0________________21665), .DIN2
       (____0___23599), .Q (________22692));
  xnr2s1 __9__0_513148(.DIN1 (_____________22083), .DIN2
       (___0_____40449), .Q (________22601));
  nnd2s1 __9____513149(.DIN1 (_________________0___21728), .DIN2
       (________22727), .Q (________22617));
  nor2s1 __9____513150(.DIN1 (________22513), .DIN2 (_____9__22402), .Q
       (________22616));
  nnd2s1 __9_0__513151(.DIN1 (___9___22263), .DIN2 (________22401), .Q
       (________22583));
  nor2s1 __9____513152(.DIN1 (____0____37167), .DIN2
       (_____________________21743), .Q (________22629));
  hi1s1 __9_90_513153(.DIN (_____9__23635), .Q (____0___22844));
  nnd2s1 __9_09_513154(.DIN1 (___9____23151), .DIN2 (________22400), .Q
       (_____0__22711));
  nnd2s1 __9__9_513155(.DIN1 (___0_____40528), .DIN2 (___0__22134), .Q
       (________23052));
  nnd2s1 __9_0__513156(.DIN1 (____9___22447), .DIN2 (_____0___32287),
       .Q (_____0__28128));
  hi1s1 __9____513157(.DIN (________22399), .Q (________22695));
  nnd2s1 __9___513158(.DIN1 (___0_____30727), .DIN2 (___0_____40515),
       .Q (________22970));
  xor2s1 __9____513159(.DIN1 (___0_____40597), .DIN2
       (_____________22098), .Q (___0____24250));
  nor2s1 __9____513160(.DIN1 (________22398), .DIN2 (___0_____40589),
       .Q (___9____23203));
  xor2s1 __9__9_513161(.DIN1 (___0_____40588), .DIN2 (_________22016),
       .Q (________22602));
  nnd2s1 __9_0__513162(.DIN1 (_______________22072), .DIN2
       (_________36493), .Q (________24984));
  nor2s1 __9____513163(.DIN1 (________22397), .DIN2
       (_____________________21747), .Q (________22703));
  nor2s1 __9____513164(.DIN1 (________22396), .DIN2 (___0_____40509),
       .Q (____9___22935));
  and2s1 __9____513165(.DIN1 (_________________0___21740), .DIN2
       (_____________________21742), .Q (________22753));
  nnd2s1 __9____513166(.DIN1 (____0______________), .DIN2
       (_____9__22868), .Q (________22615));
  nnd2s1 __9____513167(.DIN1 (_____________________21703), .DIN2
       (________22513), .Q (________22631));
  nnd2s1 __9_0__513168(.DIN1 (_______________22072), .DIN2
       (_________36556), .Q (___9____23171));
  and2s1 __9_0_513169(.DIN1 (___0_____40595), .DIN2 (________22395), .Q
       (________22725));
  nor2s1 __9____513170(.DIN1 (________23449), .DIN2
       (______________________21700), .Q (________22533));
  xnr2s1 __9___513171(.DIN1 (_________0_), .DIN2 (___0__9__40450), .Q
       (_________38239));
  nnd2s1 __9__0_513172(.DIN1 (________22395), .DIN2
       (_________________________________________0___21952), .Q
       (________22608));
  nnd2s1 __9___513173(.DIN1 (____9___23970), .DIN2
       (____0________________21721), .Q (____9___22543));
  nnd2s1 __9_09_513174(.DIN1
       (______________________________________________________________________________________0),
       .DIN2 (______9__34981), .Q (____0___23043));
  nor2s1 __9____513175(.DIN1 (________22394), .DIN2 (________24494), .Q
       (___9_0__23192));
  nor2s1 __9_0__513176(.DIN1 (________23021), .DIN2 (________22532), .Q
       (____09__23416));
  nor2s1 __9__0_513177(.DIN1 (______9__32360), .DIN2
       (______________22064), .Q (_____90__33241));
  nor2s1 __9_09_513178(.DIN1 (______9__34981), .DIN2
       (______________________________________________________________________________________0),
       .Q (________22564));
  nnd2s1 __9_0__513179(.DIN1 (_______________22069), .DIN2
       (_________34538), .Q (___9____26879));
  nor2s1 __9_0_513180(.DIN1 (_________36493), .DIN2
       (_________________________________________________________________________________________22094),
       .Q (________22873));
  nor2s1 __9_0__513181(.DIN1 (________22395), .DIN2 (___0_____40595),
       .Q (________22724));
  nnd2s1 __9____513182(.DIN1 (_________37321), .DIN2 (_________36556),
       .Q (________22712));
  nor2s1 __9_0__513183(.DIN1 (_________37320), .DIN2
       (_______________22076), .Q (________22609));
  nor2s1 __9____513184(.DIN1 (_____0__22393), .DIN2
       (_____________________21706), .Q (_____9__22538));
  nor2s1 __9____513185(.DIN1 (________22400), .DIN2
       (____0_________________21727), .Q (_____9__22613));
  nor2s1 __9_0_513186(.DIN1 (_____________22086), .DIN2
       (_____9__22633), .Q (________23004));
  nor2s1 __9_0_513187(.DIN1 (______9__31640), .DIN2 (______9__32360),
       .Q (_____0__22869));
  nor2s1 __9__0_513188(.DIN1 (_________32611), .DIN2 (____________), .Q
       (____99__23038));
  hi1s1 __9__9_513189(.DIN (________22381), .Q (________22666));
  xnr2s1 __9__513190(.DIN1 (___0_____40587), .DIN2
       (______________22105), .Q (_____0__22654));
  nor2s1 __9____513191(.DIN1 (_____9__22392), .DIN2
       (_____________________________________________21768), .Q
       (________22913));
  nor2s1 __9_0__513192(.DIN1 (_________36761), .DIN2 (_________34538),
       .Q (_____0__28424));
  nor2s1 __9____513193(.DIN1 (___0____22340), .DIN2 (___0_____40572),
       .Q (________22927));
  nnd2s1 __9____513194(.DIN1 (_____________________21748), .DIN2
       (________23555), .Q (________22853));
  nnd2s1 __9___513195(.DIN1 (__________________0___21738), .DIN2
       (___9_9__23163), .Q (____9___23034));
  hi1s1 __9__9_513196(.DIN (________22391), .Q (____9___22833));
  hi1s1 __9_90_513197(.DIN (________22625), .Q (________23709));
  nor2s1 __9____513198(.DIN1 (________23611), .DIN2
       (____0_________________21725), .Q (___9____23168));
  hi1s1 __9____513199(.DIN (________22390), .Q (________22698));
  hi1s1 __9____513200(.DIN (___0____25161), .Q (___9____25060));
  nnd2s1 __9____513201(.DIN1 (______22154), .DIN2
       (_____________________21732), .Q (________23066));
  hi1s1 __9____513202(.DIN (________22389), .Q (________22717));
  nor2s1 __9____513203(.DIN1 (________22388), .DIN2
       (_____________________21674), .Q (________22865));
  nnd2s1 __9____513204(.DIN1 (_____________________21680), .DIN2
       (____0___22457), .Q (_____0__22849));
  nor2s1 __9____513205(.DIN1 (_____0__23445), .DIN2
       (_________________9___21696), .Q (________22921));
  nor2s1 __9____513206(.DIN1 (________22754), .DIN2
       (_________________0___21740), .Q (________22981));
  and2s1 __9____513207(.DIN1 (__________________0___21686), .DIN2
       (___9____23149), .Q (___0____23276));
  hi1s1 __9__9_513208(.DIN (________22387), .Q (________22854));
  and2s1 __9____513209(.DIN1 (_____0__23445), .DIN2
       (______________________21700), .Q (________22872));
  nnd2s1 __9___513210(.DIN1 (_____________________21681), .DIN2
       (_____9__23842), .Q (________22708));
  nor2s1 __9____513211(.DIN1 (________23555), .DIN2
       (_____________________21745), .Q (________22861));
  nor2s1 __9__9_513212(.DIN1 (________23474), .DIN2 (_____9__22868), .Q
       (________22955));
  nnd2s1 __9____513213(.DIN1 (________26426), .DIN2 (________22754), .Q
       (____0___23414));
  nor2s1 __9____513214(.DIN1 (___9____26912), .DIN2
       (__________________0___21750), .Q (________23669));
  nnd2s1 __9__9_513215(.DIN1 (______________________21752), .DIN2
       (________22754), .Q (________23391));
  nor2s1 __9___513216(.DIN1 (________22727), .DIN2
       (_________________0___21728), .Q (_____9__25368));
  hi1s1 __9__9_513217(.DIN (________22386), .Q (________22762));
  nnd2s1 __9__0_513218(.DIN1 (_____________________21680), .DIN2
       (____0___23697), .Q (___9_0__23201));
  nor2s1 __9____513219(.DIN1 (___0____23256), .DIN2
       (_____________________21691), .Q (________23800));
  nnd2s1 __9__9_513220(.DIN1 (____________________), .DIN2
       (_____0__23445), .Q (________22950));
  hi1s1 __9__9_513221(.DIN (_________38301), .Q (_________35677));
  hi1s1 __9_90_513222(.DIN (________22536), .Q (________24302));
  or2s1 __9__0_513223(.DIN1 (____0________________21666), .DIN2
       (____0___23599), .Q (____9___22832));
  hi1s1 __9__513224(.DIN (________22385), .Q (_____0__22810));
  hi1s1 __9_9__513225(.DIN (____0___22555), .Q (____0___22847));
  hi1s1 __9____513226(.DIN (___9____24088), .Q (________22851));
  nnd2s1 __9___513227(.DIN1 (_____________________21744), .DIN2
       (____09__23048), .Q (________22850));
  nnd2s1 __9___513228(.DIN1 (____90__26673), .DIN2 (________22397), .Q
       (________23372));
  nor2s1 __9____513229(.DIN1 (_____9__22868), .DIN2
       (____0______________), .Q (________23364));
  nnd2s1 __9____513230(.DIN1 (___0____26120), .DIN2
       (____0_____________0___21723), .Q (________23092));
  nnd2s1 __9____513231(.DIN1 (____0________________21715), .DIN2
       (_______22258), .Q (________22876));
  nor2s1 __9____513232(.DIN1 (________22382), .DIN2
       (____0________________21666), .Q (____9___23036));
  nor2s1 __9____513233(.DIN1 (________22628), .DIN2 (_____0__22384), .Q
       (____0___22842));
  hi1s1 __9____513234(.DIN (_____9__22383), .Q (________24418));
  hi1s1 __9_9__513235(.DIN (____0___23311), .Q (____9___23037));
  hi1s1 __9___513236(.DIN (________26440), .Q (________26601));
  nor2s1 __9___513237(.DIN1 (______22127), .DIN2
       (____0________________21668), .Q (________24544));
  nnd2s1 __9____513238(.DIN1 (_____0__22384), .DIN2 (________22628), .Q
       (___0____23292));
  nnd2s1 __9____513239(.DIN1 (_____________________21673), .DIN2
       (_______22260), .Q (_____9__22858));
  hi1s1 __9_9_513240(.DIN (____0___22840), .Q (________26419));
  nor2s1 __9____513241(.DIN1 (________22754), .DIN2
       (______________________21752), .Q (____0___25502));
  nor2s1 __9____513242(.DIN1 (________23021), .DIN2
       (__________________0___21712), .Q (________22818));
  nnd2s1 __9__9_513243(.DIN1 (________24602), .DIN2 (____9___23032), .Q
       (____9___23591));
  nor2s1 __9___513244(.DIN1 (______22123), .DIN2
       (__________________0_), .Q (____90__23962));
  nnd2s1 __9__9_513245(.DIN1 (_____________________21743), .DIN2
       (________26431), .Q (________22953));
  nor2s1 __9____513246(.DIN1 (_____________________21742), .DIN2
       (_________________0___21740), .Q (________23469));
  nnd2s1 __9____513247(.DIN1 (___9_9___39790), .DIN2
       (_________________0___21676), .Q (___9_____39461));
  nnd2s1 __9____513248(.DIN1 (____0________________21666), .DIN2
       (________22382), .Q (____0___22845));
  nor2s1 __9____513249(.DIN1 (___9____23151), .DIN2
       (____0_________________21724), .Q (________22862));
  nor2s1 __9____513250(.DIN1 (________22380), .DIN2
       (_________________9___21696), .Q (____9___26583));
  nnd2s1 __9___513251(.DIN1 (_________________0___21740), .DIN2
       (_____0__22384), .Q (___0____26080));
  nor2s1 __9__0_513252(.DIN1 (____0_____________0___21723), .DIN2
       (___0____26120), .Q (________25931));
  hi1s1 __9_9__513253(.DIN (________22379), .Q (____9___24358));
  nnd2s1 __9_9__513254(.DIN1
       (_________________________________________________________________________________________22094),
       .DIN2 (_________36556), .Q (________22378));
  nor2s1 __9_9__513255(.DIN1 (_________34538), .DIN2
       (_________________________________________________________________________________________22095),
       .Q (________22377));
  nnd2s1 __9_9_513256(.DIN1 (____________), .DIN2 (_____9__23492), .Q
       (________22376));
  nor2s1 __9__0_513257(.DIN1 (____90__26673), .DIN2 (____0____37167),
       .Q (_____0__22375));
  xnr2s1 __9___513258(.DIN1
       (__________________________________________________________________21983),
       .DIN2
       (_______________________________________________________________9),
       .Q (_____9));
  xor2s1 __9____513259(.DIN1 (___0_9___40459), .DIN2 (___0_____40589),
       .Q (________22374));
  xor2s1 __9____513260(.DIN1 (___0_____40478), .DIN2 (___0__0__40413),
       .Q (________22373));
  nnd2s1 __9___513261(.DIN1 (___0__0__40521), .DIN2 (______22142), .Q
       (________22372));
  nnd2s1 __9__0_513262(.DIN1 (__________9_), .DIN2 (______9__32360), .Q
       (________22371));
  or2s1 __9____513263(.DIN1
       (______________________________________________21938), .DIN2
       (________22369), .Q (________22370));
  nor2s1 __9_9_513264(.DIN1 (_________36402), .DIN2
       (_________________________________________________________________________________________22090),
       .Q (________22368));
  nnd2s1 __9_0_513265(.DIN1 (___09___22357), .DIN2
       (______________22104), .Q (_____0));
  xnr2s1 __9__9_513266(.DIN1
       (_____________________________________________21941), .DIN2
       (_________________________________________9___21943), .Q
       (____09));
  nor2s1 __9__9_513267(.DIN1 (___09___22355), .DIN2
       (_____________22083), .Q (____0___22367));
  hi1s1 __9____513268(.DIN (____0___22365), .Q (____0___22366));
  or2s1 __9____513269(.DIN1 (_____________________21673), .DIN2
       (________24475), .Q (____0___22364));
  and2s1 __9__0_513270(.DIN1 (_____________________21703), .DIN2
       (________23754), .Q (____0___22363));
  nnd2s1 __9_9__513271(.DIN1 (___9____23151), .DIN2 (________23611), .Q
       (____0___22362));
  nnd2s1 __9_0_513272(.DIN1 (_________32918), .DIN2 (_________33293),
       .Q (____0___22361));
  or2s1 __9____513273(.DIN1 (____00), .DIN2 (___0__0__40531), .Q
       (____0_));
  nor2s1 __9___513274(.DIN1 (___09___22360), .DIN2 (____9___22447), .Q
       (___099));
  or2s1 __9____513275(.DIN1 (___9_0__29602), .DIN2
       (__________________________________________9___21934), .Q
       (___09___22359));
  nor2s1 __9_00_513276(.DIN1 (______________22104), .DIN2
       (___09___22357), .Q (___09___22358));
  nnd2s1 __9__0_513277(.DIN1 (_____________22083), .DIN2
       (___09___22355), .Q (___09___22356));
  nnd2s1 __9__9_513278(.DIN1 (_____________________21729), .DIN2
       (_____9__24325), .Q (___09___22354));
  nor2s1 __9___513279(.DIN1 (____9___22447), .DIN2 (_____0___32287), .Q
       (___09_));
  xnr2s1 __9__0_513280(.DIN1
       (_____________________________________________21842), .DIN2
       (___0__0__40521), .Q (___090));
  nor2s1 __9_00_513281(.DIN1 (_____9__23444), .DIN2 (___0____23256), .Q
       (___0_9__22353));
  nor2s1 __9_9__513282(.DIN1 (__0), .DIN2 (___0_____40446), .Q
       (___0____22352));
  xor2s1 __9____513283(.DIN1
       (_______________________________________________________________0__21998),
       .DIN2 (_____________________________________________21924), .Q
       (___0____22351));
  nnd2s1 __9____513284(.DIN1
       (_________________________________________9___21779), .DIN2
       (____0___28017), .Q (___0____22350));
  nnd2s1 __9____513285(.DIN1 (_________34167), .DIN2 (_____9___33157),
       .Q (___0____22349));
  xnr2s1 __9__9_513286(.DIN1
       (____________________________________________21793), .DIN2
       (___0_____40528), .Q (___0____22348));
  nnd2s1 __9__0_513287(.DIN1 (___0_____40584), .DIN2 (___0____22346),
       .Q (___0____22347));
  xor2s1 __9___513288(.DIN1
       (____________________________________________21792), .DIN2
       (___0_9___40554), .Q (___0____22345));
  nor2s1 __9___513289(.DIN1 (___0_9__22343), .DIN2 (_________0_), .Q
       (___0_0__22344));
  nnd2s1 __9_09_513290(.DIN1 (___009), .DIN2
       (_____________________________________9_______21881), .Q
       (___0____22342));
  nnd2s1 __9____513291(.DIN1 (___0_____40572), .DIN2 (___0____22340),
       .Q (___0____22341));
  nnd2s1 __9____513292(.DIN1 (___0__9__40420), .DIN2 (_____22113), .Q
       (___0____22339));
  xnr2s1 __9____513293(.DIN1 (_____________22101), .DIN2
       (_____________22100), .Q (___0____22338));
  nor2s1 __9_9_513294(.DIN1 (_________37321), .DIN2
       (_______________22072), .Q (___0____22337));
  nor2s1 __9_9__513295(.DIN1 (____________), .DIN2 (___0____23297), .Q
       (___0____22336));
  nnd2s1 __9_0__513296(.DIN1 (_________36761), .DIN2 (_________34538),
       .Q (___0____22335));
  xnr2s1 __9___513297(.DIN1
       (_____________________________________________21899), .DIN2
       (__________________________________________________________________21988),
       .Q (___0_0__22334));
  nor2s1 __9_9_513298(.DIN1 (_________35844), .DIN2
       (_______________22075), .Q (___0_9__22333));
  nor2s1 __9____513299(.DIN1 (______9__32360), .DIN2 (__________9_), .Q
       (___0____22332));
  xnr2s1 __9____513300(.DIN1
       (_____________________________________________21970), .DIN2
       (___0__9__40420), .Q (___0____22331));
  nor2s1 __9____513301(.DIN1 (_____0__22384), .DIN2
       (______________________21751), .Q (___0____22330));
  nnd2s1 __9___513302(.DIN1 (______22121), .DIN2
       (____________________________________________21764), .Q
       (___0____22329));
  xnr2s1 __9____513303(.DIN1 (___0_9___40558), .DIN2 (___0_____40539),
       .Q (___0____22328));
  xnr2s1 __9__9_513304(.DIN1
       (______________________________________0______21887), .DIN2
       (______________________________________0____), .Q
       (___0____22327));
  xor2s1 __9____513305(.DIN1
       (______________________________________________21979), .DIN2
       (___0_____40414), .Q (___0____22326));
  nor2s1 __9_00_513306(.DIN1 (___9_9__23163), .DIN2 (_____9___37752),
       .Q (___0____22325));
  nor2s1 __9_0__513307(.DIN1 (_________36493), .DIN2
       (_______________22070), .Q (___0_0__22324));
  nor2s1 __9____513308(.DIN1 (_____0__22499), .DIN2 (________22398), .Q
       (___0_9__22323));
  nnd2s1 __9_0__513309(.DIN1 (______22132), .DIN2
       (_____________________________________________21839), .Q
       (___0____22322));
  nnd2s1 __9_9__513310(.DIN1 (_____________________21743), .DIN2
       (___9____26912), .Q (___0____22321));
  nor2s1 __9_0__513311(.DIN1 (________22380), .DIN2 (_____0__23445), .Q
       (___0____22320));
  xor2s1 __9____513312(.DIN1 (___0_____40446), .DIN2
       (_________________________________________0___21895), .Q
       (___0____22319));
  nor2s1 __9___513313(.DIN1
       (______________________________________________21938), .DIN2
       (___0____22317), .Q (___0____22318));
  nnd2s1 __9____513314(.DIN1 (___9_9___39696), .DIN2
       (_____________________________________________21907), .Q
       (___0_9__22316));
  nor2s1 __9____513315(.DIN1 (___0__0__40599), .DIN2 (___0__22149), .Q
       (___0____22315));
  nor2s1 __9__9_513316(.DIN1 (___0____22313), .DIN2
       (_______________22070), .Q (___0____22314));
  xnr2s1 __9___513317(.DIN1 (___0__0__40531), .DIN2 (___0_____40547),
       .Q (___0____22312));
  nor2s1 __9____513318(.DIN1 (________22502), .DIN2 (___0_____40447),
       .Q (___0____22311));
  nnd2s1 __9_513319(.DIN1 (________23362), .DIN2 (________22461), .Q
       (___0____22310));
  xor2s1 __9__0_513320(.DIN1
       (____________________________________________21848), .DIN2
       (____________________________________________21831), .Q
       (___0____22309));
  nnd2s1 __9___513321(.DIN1 (______22136), .DIN2
       (______________________________________0_______21892), .Q
       (___0____22308));
  xor2s1 __9____513322(.DIN1 (___0__9__40580), .DIN2 (___0_____40493),
       .Q (___0_0__22307));
  nor2s1 __9__513323(.DIN1 (________22504), .DIN2 (_____________22088),
       .Q (___0_9__22306));
  nnd2s1 __9_0__513324(.DIN1 (________22480), .DIN2 (inData[2]), .Q
       (___0____22305));
  nor2s1 __9__513325(.DIN1 (_________34167), .DIN2 (___0_____40478), .Q
       (___0____22304));
  nor2s1 __9_0__513326(.DIN1 (_________36556), .DIN2 (_________36493),
       .Q (___0____22303));
  or2s1 __9__0_513327(.DIN1 (___99____39814), .DIN2
       (_____________________________________________21969), .Q
       (___0____22302));
  nnd2s1 __9____513328(.DIN1 (______________22105), .DIN2
       (___0____22300), .Q (___0____22301));
  xor2s1 __9____513329(.DIN1
       (_____________________________________________21811), .DIN2
       (_________________________________________________________________________________________22089),
       .Q (___0____22299));
  xor2s1 __9___513330(.DIN1
       (_____________________________________________21853), .DIN2
       (_____________________________________0______21756), .Q
       (___0____22298));
  nor2s1 __9___513331(.DIN1 (___0_____40423), .DIN2 (_________35587),
       .Q (___0_0__22297));
  nnd2s1 __9_9__513332(.DIN1 (______________22067), .DIN2
       (_____9___33157), .Q (___0_9));
  xor2s1 __9____513333(.DIN1
       (______________________________________________21913), .DIN2
       (______________________________________________21916), .Q
       (___0____22296));
  xnr2s1 __9____513334(.DIN1 (______________22110), .DIN2
       (______________22109), .Q (___0____22295));
  xor2s1 __9__513335(.DIN1 (___0_____40546), .DIN2 (___0_0___40564), .Q
       (___0____22294));
  nnd2s1 __9_0__513336(.DIN1 (___0__9__40412), .DIN2 (_________36762),
       .Q (___0____22293));
  hi1s1 __9____513337(.DIN (___0____22291), .Q (___0____22292));
  nor2s1 __9_9_513338(.DIN1 (_________37320), .DIN2
       (_________________________________________________________________________________________22089),
       .Q (___0____22290));
  nor2s1 __9___513339(.DIN1 (________22627), .DIN2 (___9____23149), .Q
       (___0__));
  nor2s1 __9___513340(.DIN1 (___009), .DIN2 (___0__9__40450), .Q
       (___0_0));
  or2s1 __9__0_513341(.DIN1 (_____9__22402), .DIN2
       (_____________________21703), .Q (___00___22289));
  xnr2s1 __9____513342(.DIN1
       (____________________________________________21846), .DIN2
       (____________________________________________21847), .Q
       (___00___22288));
  nnd2s1 __9_0__513343(.DIN1 (______22140), .DIN2
       (____________________________________________21762), .Q
       (___00_));
  xor2s1 __9____513344(.DIN1 (___0_____40547), .DIN2
       (____________________________________________21818), .Q
       (__9____22287));
  nor2s1 __9____513345(.DIN1 (________26530), .DIN2 (___0_____40425),
       .Q (__9__));
  nor2s1 __9_0__513346(.DIN1 (_____________22097), .DIN2 (____99), .Q
       (_______22286));
  xor2s1 __9__513347(.DIN1
       (_____________________________________________21845), .DIN2
       (___0__9__40480), .Q (_______22285));
  nnd2s1 __9_9__513348(.DIN1 (___0_____40598), .DIN2 (_________32918),
       .Q (_______22284));
  and2s1 __9_9__513349(.DIN1 (____99), .DIN2 (_____________22097), .Q
       (_______22283));
  or2s1 __9__9_513350(.DIN1 (________22513), .DIN2
       (_____________________21703), .Q (_______22282));
  nor2s1 __9____513351(.DIN1 (_____________22085), .DIN2
       (_______22280), .Q (____0__22281));
  nor2s1 __9_513352(.DIN1 (________22628), .DIN2 (________26217), .Q
       (_______22279));
  nor2s1 __9_513353(.DIN1 (_________35727), .DIN2
       (______________22066), .Q (_______22278));
  nnd2s1 __9_0__513354(.DIN1 (_________36762), .DIN2 (inData[18]), .Q
       (_______22277));
  nnd2s1 __9__513355(.DIN1 (____0_________________21724), .DIN2
       (________23611), .Q (___0___22276));
  nor2s1 __9_9__513356(.DIN1 (___9____25102), .DIN2 (_____9__23492), .Q
       (___0___22275));
  xor2s1 __9___513357(.DIN1 (__________9_), .DIN2
       (______________22067), .Q (___0___22274));
  xor2s1 __9____513358(.DIN1 (___0_____40446), .DIN2 (___0_____40582),
       .Q (___0___22273));
  or2s1 __9____513359(.DIN1 (____0____________0___21713), .DIN2
       (________22857), .Q (___00__22272));
  nor2s1 __9__0_513360(.DIN1 (___0_____40443), .DIN2 (______22141), .Q
       (___99__22271));
  nnd2s1 __9_9__513361(.DIN1 (__________9_), .DIN2 (_________32918), .Q
       (___9___22270));
  nor2s1 __9_9__513362(.DIN1 (_________37412), .DIN2
       (_______________22077), .Q (___9___22269));
  nnd2s1 __9____513363(.DIN1 (_________34601), .DIN2 (inData[24]), .Q
       (___9___22268));
  nnd2s1 __9__0_513364(.DIN1 (_____9__22577), .DIN2
       (______________________________________________21967), .Q
       (___9___22267));
  nnd2s1 __9_9__513365(.DIN1 (___0_____40411), .DIN2 (_________37412),
       .Q (___9___22266));
  nnd2s1 __9____513366(.DIN1
       (_________________________________________0___21798), .DIN2
       (________22420), .Q (___9___22265));
  or2s1 __9_0__513367(.DIN1 (___9__22137), .DIN2 (___0__9__40440), .Q
       (___9___22264));
  nnd2s1 __9___513368(.DIN1 (____9___23970), .DIN2 (____90__24060), .Q
       (________22621));
  or2s1 __9__9_513369(.DIN1 (_________37424), .DIN2
       (_____________________________________________21924), .Q
       (___90___23137));
  nnd2s1 __9____513370(.DIN1 (___9___22263), .DIN2
       (_____________________21734), .Q (________22667));
  nnd2s1 __9__0_513371(.DIN1 (____________), .DIN2 (_________32611), .Q
       (________22592));
  nnd2s1 __9__9_513372(.DIN1 (______________________21701), .DIN2
       (________23449), .Q (____9___22542));
  nnd2s1 __9____513373(.DIN1 (____0________________21664), .DIN2
       (_____9__22868), .Q (________22875));
  nnd2s1 __9___513374(.DIN1 (___________________), .DIN2
       (_________________0_), .Q (________22630));
  nnd2s1 __9__513375(.DIN1
       (_________________________________________________________________________________________22089),
       .DIN2 (___90__22262), .Q (___90___23134));
  nnd2s1 __9____513376(.DIN1 (_____________________21689), .DIN2
       (___9_9__23181), .Q (____9___22540));
  xor2s1 __9__9_513377(.DIN1 (_____________22088), .DIN2
       (___0_____40447), .Q (___9__9__39098));
  nor2s1 __9___513378(.DIN1 (________23362), .DIN2
       (_____________________21694), .Q (________22620));
  nor2s1 __9_0__513379(.DIN1 (_____9__23492), .DIN2 (______9__32360),
       .Q (____0___22747));
  nnd2s1 __9____513380(.DIN1 (____9__22261), .DIN2 (_______22260), .Q
       (________22618));
  nor2s1 __9_0__513381(.DIN1 (_________34167), .DIN2 (___0__9__40412),
       .Q (________23115));
  nor2s1 __9____513382(.DIN1 (____9___26770), .DIN2
       (__________________________________________0___21935), .Q
       (________22996));
  nor2s1 __9____513383(.DIN1 (___0__9__40500), .DIN2 (_________36583),
       .Q (________22960));
  nor2s1 __9__513384(.DIN1 (_______22259), .DIN2 (____0____________9_),
       .Q (________22863));
  xnr2s1 __9____513385(.DIN1 (___0_9___40454), .DIN2
       (_______________0), .Q (________22537));
  nor2s1 __9____513386(.DIN1 (________22627), .DIN2
       (__________________0___21686), .Q (____9___22834));
  nnd2s1 __9____513387(.DIN1 (______________________21751), .DIN2
       (_____0__22384), .Q (________22707));
  nnd2s1 __9_0__513388(.DIN1 (________22678), .DIN2 (_______22259), .Q
       (________22683));
  nor2s1 __9____513389(.DIN1 (_________________9___21737), .DIN2
       (______22154), .Q (_____0__22624));
  nor2s1 __9____513390(.DIN1 (___0_9___40454), .DIN2 (____), .Q
       (________22788));
  nor2s1 __9_0__513391(.DIN1 (_______22258), .DIN2 (_______22250), .Q
       (____9___22831));
  and2s1 __9_09_513392(.DIN1 (_____9__22633), .DIN2
       (_____________22086), .Q (________23003));
  nnd2s1 __9____513393(.DIN1 (____0________________21719), .DIN2
       (________23959), .Q (________22632));
  nor2s1 __9____513394(.DIN1 (___9_____39773), .DIN2
       (______________________________________________21937), .Q
       (___000___39893));
  nor2s1 __9____513395(.DIN1 (________22994), .DIN2
       (__________________0___21697), .Q (________22534));
  nnd2s1 __9__513396(.DIN1 (_____________________21690), .DIN2
       (________22884), .Q (_____9__22623));
  nnd2s1 __9____513397(.DIN1 (_____________________21692), .DIN2
       (________23026), .Q (________22706));
  nor2s1 __9___513398(.DIN1 (_________37789), .DIN2 (____99___36174),
       .Q (________22890));
  hi1s1 __9____513399(.DIN (_______22257), .Q (________26516));
  and2s1 __9____513400(.DIN1 (___0_____40546), .DIN2 (_________33206),
       .Q (________22782));
  nor2s1 __9__0_513401(.DIN1 (____0___22846), .DIN2
       (_____________________21692), .Q (____9___22541));
  hi1s1 __9_513402(.DIN (________22855), .Q (___9____23145));
  nor2s1 __9__9_513403(.DIN1 (____09__23048), .DIN2 (____0____37167),
       .Q (________22535));
  nnd2s1 __9_0_513404(.DIN1 (_______________22076), .DIN2
       (_________37320), .Q (___9____23174));
  nor2s1 __9____513405(.DIN1 (________22400), .DIN2 (___9____23151), .Q
       (________22622));
  nor2s1 __9_0__513406(.DIN1 (_________36556), .DIN2
       (_______________22072), .Q (________22581));
  hi1s1 __9__513407(.DIN (_______22256), .Q (________22714));
  nnd2s1 __9___513408(.DIN1 (________23754), .DIN2 (____9___23032), .Q
       (________22704));
  nnd2s1 __9___513409(.DIN1 (________23026), .DIN2 (________22461), .Q
       (________22795));
  nor2s1 __9____513410(.DIN1 (_________37320), .DIN2 (_________36762),
       .Q (________25597));
  hi1s1 __9__9_513411(.DIN (_______22255), .Q (___0____23289));
  nor2s1 __9____513412(.DIN1 (_______22254), .DIN2 (_____9__24635), .Q
       (____9___22932));
  nor2s1 __9___513413(.DIN1 (____0___26590), .DIN2 (________26426), .Q
       (________23911));
  nor2s1 __9____513414(.DIN1 (___0_____40607), .DIN2 (______22122), .Q
       (________23117));
  nnd2s1 __9___513415(.DIN1 (________26217), .DIN2 (____90__26673), .Q
       (____0___22841));
  hi1s1 __9__9_513416(.DIN (_______22253), .Q (________22887));
  and2s1 __9____513417(.DIN1 (_________________0___21740), .DIN2
       (________22754), .Q (___0____23251));
  nnd2s1 __9____513418(.DIN1 (______________________21753), .DIN2
       (________22628), .Q (_____9__22828));
  xor2s1 __9____513419(.DIN1 (___0_____40624), .DIN2 (___0_9___40455),
       .Q (___9____26034));
  nnd2s1 __9____513420(.DIN1 (__________________0___21686), .DIN2
       (________22627), .Q (________22693));
  nnd2s1 __9___513421(.DIN1 (_____________________21674), .DIN2
       (________22388), .Q (_____0__22859));
  hi1s1 __9_9__513422(.DIN (_________38203), .Q (____0____36245));
  nnd2s1 __9____513423(.DIN1 (____0___26590), .DIN2 (________26217), .Q
       (_____0__22691));
  nor2s1 __9____513424(.DIN1 (_______22252), .DIN2 (________23959), .Q
       (________23071));
  hi1s1 __9_9__513425(.DIN (____9___22933), .Q (________22866));
  hi1s1 __9__9_513426(.DIN (_______22251), .Q (________22699));
  nnd2s1 __9___513427(.DIN1 (____0________________21720), .DIN2
       (_______22252), .Q (_____0__22701));
  nnd2s1 __9__0_513428(.DIN1 (_____________________21743), .DIN2
       (____0____37167), .Q (________22697));
  nor2s1 __9____513429(.DIN1 (________22884), .DIN2
       (_____________________21690), .Q (____9___22835));
  hi1s1 __9_9_513430(.DIN (____0___22743), .Q (_____9__22700));
  nnd2s1 __9____513431(.DIN1 (_____________________21681), .DIN2
       (________22924), .Q (____09__22848));
  nnd2s1 __9____513432(.DIN1 (_____________________21705), .DIN2
       (____9___23032), .Q (____9___22837));
  nnd2s1 __9___513433(.DIN1 (_______22250), .DIN2 (_______22258), .Q
       (________22856));
  nnd2s1 __9__513434(.DIN1 (____0______________), .DIN2
       (_____9__24635), .Q (____0___22943));
  hi1s1 __9_9__513435(.DIN (___99___26049), .Q (________25438));
  nor2s1 __9____513436(.DIN1 (______22130), .DIN2
       (_________________9_), .Q (________22798));
  nor2s1 __9____513437(.DIN1 (________23026), .DIN2
       (_____________________21692), .Q (________22792));
  nor2s1 __9__0_513438(.DIN1 (___9_9__23181), .DIN2
       (_____________________21689), .Q (________22885));
  nor2s1 __9____513439(.DIN1 (_______22252), .DIN2 (____9___23970), .Q
       (____9___24360));
  nor2s1 __9__0_513440(.DIN1 (________22532), .DIN2
       (_____________________21709), .Q (________22702));
  nnd2s1 __9___513441(.DIN1 (_____00__35736), .DIN2 (___9_____39397),
       .Q (________23618));
  hi1s1 __9_9__513442(.DIN (___9____23156), .Q (___09___23306));
  hi1s1 __9_90_513443(.DIN (_______22249), .Q (________22852));
  hi1s1 __9_9__513444(.DIN (____9___23782), .Q (________23438));
  nor2s1 __9____513445(.DIN1 (________22461), .DIN2 (________23026), .Q
       (________22715));
  and2s1 __9__0_513446(.DIN1 (____0________________21663), .DIN2
       (_____9__24635), .Q (________23089));
  hi1s1 __9_9__513447(.DIN (________23384), .Q (____00__22839));
  nor2s1 __9____513448(.DIN1 (_____0__22384), .DIN2
       (_________________0___21740), .Q (____0___23602));
  nor2s1 __9__513449(.DIN1 (________23024), .DIN2
       (____0________________21718), .Q (________23014));
  nnd2s1 __9__9_513450(.DIN1 (_____________________21706), .DIN2
       (_____0__22393), .Q (____99__22838));
  nor2s1 __9____513451(.DIN1 (____0___26590), .DIN2
       (_____________________21742), .Q (________24625));
  nor2s1 __9____513452(.DIN1 (_____________________21732), .DIN2
       (______22154), .Q (____9___23592));
  or2s1 __9___513453(.DIN1 (________23356), .DIN2
       (_____________________21670), .Q (_____9__22918));
  nor2s1 __9____513454(.DIN1 (________26217), .DIN2
       (_____________________21747), .Q (________25925));
  nnd2s1 __9____513455(.DIN1 (____9___23970), .DIN2
       (____0_________________21724), .Q (________23080));
  nnd2s1 __9____513456(.DIN1 (_____________________21670), .DIN2
       (________23356), .Q (____0___23504));
  nor2s1 __9____513457(.DIN1 (_____9___37752), .DIN2
       (__________________0___21738), .Q (________22977));
  nor2s1 __9____513458(.DIN1 (________23611), .DIN2
       (____0_________________21726), .Q (___9____23167));
  nor2s1 __9____513459(.DIN1 (____00__23407), .DIN2
       (_____________________21695), .Q (___9____24123));
  nor2s1 __9___513460(.DIN1 (____9___24066), .DIN2 (______22154), .Q
       (___0_9__24217));
  nnd2s1 __9___513461(.DIN1 (____0________________21663), .DIN2
       (______22151), .Q (___990));
  nnd2s1 __9____513462(.DIN1 (____0____________0___21713), .DIN2
       (_______22250), .Q (________22864));
  nor2s1 __9____513463(.DIN1 (________23734), .DIN2
       (_____________________21731), .Q (________23006));
  nor2s1 __9____513464(.DIN1 (________22628), .DIN2 (________22754), .Q
       (________26618));
  nor2s1 __9____513465(.DIN1 (____0____37167), .DIN2
       (_____________________21748), .Q (________24882));
  nor2s1 __9____513466(.DIN1 (____0___23697), .DIN2 (_____9__23842), .Q
       (____9___23786));
  nnd2s1 __9____513467(.DIN1 (____00__23597), .DIN2 (________22705), .Q
       (________22867));
  or2s1 __9___513468(.DIN1 (_________________0___21676), .DIN2
       (___9_9___39790), .Q (____9___22547));
  nor2s1 __9____513469(.DIN1 (________22705), .DIN2
       (____0________________21716), .Q (________22973));
  hi1s1 __9_9_513470(.DIN (________26421), .Q (___9_9__25977));
  nnd2s1 __9____513471(.DIN1 (_____________________21695), .DIN2
       (____00__23407), .Q (_____0__26149));
  nor2s1 __9____513472(.DIN1 (_____0__23445), .DIN2
       (____________________), .Q (________24884));
  nnd2s1 __9____513473(.DIN1 (_____________________21746), .DIN2
       (________22397), .Q (________25744));
  nor2s1 __9____513474(.DIN1 (_______22260), .DIN2
       (_____________________21673), .Q (___9____23152));
  nnd2s1 __9____513475(.DIN1 (____0___26590), .DIN2 (___9____26912), .Q
       (________25644));
  hi1s1 __9_9__513476(.DIN (________22786), .Q (________22871));
  nnd2s1 __9____513477(.DIN1 (____0________________21718), .DIN2
       (________23024), .Q (___9____23147));
  hi1s1 __9_9__513478(.DIN (________22694), .Q (________26174));
  nnd2s1 __9___513479(.DIN1 (___________________), .DIN2
       (___9_____39397), .Q (______9__36337));
  hi1s1 __9_9__513480(.DIN (_________38838), .Q (___90____38993));
  nor2s1 __9__9_513481(.DIN1 (____90__26673), .DIN2
       (______________________21751), .Q (________25569));
  hi1s1 __9_9__513482(.DIN (_______22248), .Q (____09__26331));
  hi1s1 __9_9__513483(.DIN (_____9___36725), .Q (___90____39055));
  nnd2s1 __9____513484(.DIN1 (_____9__24325), .DIN2 (________23734), .Q
       (________22965));
  nnd2s1 __9____513485(.DIN1 (____0________________21664), .DIN2
       (_______22254), .Q (____0___22942));
  hi1s1 __9_9_513486(.DIN (____0__22247), .Q (_____0__23095));
  and2s1 __9__0_513487(.DIN1 (___0_____40512), .DIN2 (inData[20]), .Q
       (____9__22246));
  and2s1 __9_0__513488(.DIN1 (_________________9___21749), .DIN2
       (_____________________________________________21768), .Q
       (_______22245));
  and2s1 __9____513489(.DIN1 (_________22014), .DIN2 (___0_____40594),
       .Q (_______22244));
  nor2s1 __9____513490(.DIN1 (___0__0__40619), .DIN2
       (______________________________________0_______21889), .Q
       (_______22243));
  or2s1 __9__0_513491(.DIN1 (___0_____40523), .DIN2
       (_____________________________________________21823), .Q
       (_______22242));
  or2s1 __9____513492(.DIN1
       (_____________________________________0_______21759), .DIN2
       (___0_____40539), .Q (_______22241));
  nor2s1 __9____513493(.DIN1 (______________22108), .DIN2
       (_____________22084), .Q (_______22240));
  and2s1 __9____513494(.DIN1 (___0__9__40450), .DIN2 (inData[0]), .Q
       (_______22239));
  and2s1 __9__0_513495(.DIN1 (___0__0__40431), .DIN2
       (_____________________________________________21940), .Q
       (_______22238));
  nnd2s1 __9__513496(.DIN1
       (______________________________________________21979), .DIN2
       (______________________________________________21980), .Q
       (_______22237));
  and2s1 __9____513497(.DIN1 (___0_____40584), .DIN2
       (______________22110), .Q (_______22236));
  nor2s1 __9____513498(.DIN1
       (_____________________________________________21770), .DIN2
       (___0_____40549), .Q (____0__22235));
  and2s1 __9_0_513499(.DIN1
       (_________________________________________0___21814), .DIN2
       (___0_0___40565), .Q (____9__22234));
  nnd2s1 __9____513500(.DIN1
       (__________________________________________9___21977), .DIN2
       (______________________________________________21976), .Q
       (_______22233));
  and2s1 __9____513501(.DIN1 (___0__0__40501), .DIN2 (inData[14]), .Q
       (_______22232));
  nor2s1 __9___513502(.DIN1 (_________9_), .DIN2 (___0__0__40591), .Q
       (_______22231));
  nnd2s1 __9_9__513503(.DIN1 (__________9_), .DIN2
       (_______________22070), .Q (_______22230));
  nor2s1 __9_09_513504(.DIN1 (___0_____40418), .DIN2 (___0_____40611),
       .Q (_______22229));
  nor2s1 __9_9__513505(.DIN1 (___0_____40598), .DIN2
       (______________22064), .Q (_______22228));
  nnd2s1 __9_0_513506(.DIN1 (_____________________21703), .DIN2
       (_________________0___21702), .Q (_______22227));
  and2s1 __9____513507(.DIN1 (___0_____40485), .DIN2 (inData[18]), .Q
       (_______22226));
  or2s1 __9_0__513508(.DIN1 (___0_____40504), .DIN2 (___0_____40516),
       .Q (____0__22225));
  and2s1 __9____513509(.DIN1 (___0_____40504), .DIN2 (inData[10]), .Q
       (____9__22224));
  nor2s1 __9__0_513510(.DIN1 (_____________22098), .DIN2
       (___0_____40597), .Q (_______22223));
  nor2s1 __9____513511(.DIN1 (___0_0___40466), .DIN2
       (_________________________________________0___21840), .Q
       (_______22222));
  nor2s1 __9_0_513512(.DIN1
       (______________________________________________________________________________________0__22093),
       .DIN2 (_______________22077), .Q (_______22221));
  nor2s1 __9____513513(.DIN1 (___0_99__40560), .DIN2 (___0_____40542),
       .Q (_______22220));
  and2s1 __9_0__513514(.DIN1 (___0_____40446), .DIN2 (___0_____40582),
       .Q (_______22219));
  and2s1 __9_99_513515(.DIN1 (___0_____40437), .DIN2 (___0_____40438),
       .Q (_______22218));
  nor2s1 __9__0_513516(.DIN1
       (_____________________________________________21784), .DIN2
       (___0_____40536), .Q (_______22217));
  nnd2s1 __9____513517(.DIN1
       (__________________________________________________________________21996),
       .DIN2 (_____________22102), .Q (_______22216));
  and2s1 __9__0_513518(.DIN1 (___0_____40597), .DIN2
       (_____________22098), .Q (____0__22215));
  nor2s1 __9_0__513519(.DIN1 (___0_____40582), .DIN2 (___0_____40446),
       .Q (____9__22214));
  and2s1 __9____513520(.DIN1 (____0________________21667), .DIN2
       (____0________________21666), .Q (_______22213));
  or2s1 __9_0__513521(.DIN1
       (____________________________________________21790), .DIN2
       (_____________________________________________21783), .Q
       (_______22212));
  or2s1 __9____513522(.DIN1
       (__________________________________________________________________21986),
       .DIN2 (___0_____40617), .Q (_______22211));
  nor2s1 __9_0__513523(.DIN1
       (____________________________________________21804), .DIN2
       (____________________________________________21832), .Q
       (_______22210));
  nnd2s1 __9_0__513524(.DIN1
       (_____________________________________________21899), .DIN2
       (_____________________________________________21900), .Q
       (_______22209));
  and2s1 __9_0__513525(.DIN1 (___0_____40594), .DIN2 (___0_____40595),
       .Q (_______22208));
  and2s1 __9__9_513526(.DIN1
       (_________________________________________0___21824), .DIN2
       (_____________________________________________21841), .Q
       (_______22207));
  nnd2s1 __9___513527(.DIN1
       (______________________________________________21967), .DIN2
       (inData[18]), .Q (_______22206));
  nnd2s1 __9____513528(.DIN1 (_____________22084), .DIN2
       (______________22108), .Q (____0__22205));
  nnd2s1 __9_9_513529(.DIN1
       (__________________________________________9_), .DIN2
       (inData[12]), .Q (___09));
  or2s1 __9____513530(.DIN1
       (_____________________________________________21795), .DIN2
       (___________________________________________), .Q
       (___0___22204));
  nnd2s1 __9__0_513531(.DIN1 (___0__0__40431), .DIN2 (___0_____40612),
       .Q (___0___22203));
  nor2s1 __9_0__513532(.DIN1 (____0________________21664), .DIN2
       (____0________________21662), .Q (___0___22202));
  or2s1 __9____513533(.DIN1
       (_________________________________________9___21803), .DIN2
       (___0_0___40565), .Q (___0___22201));
  or2s1 __9__9_513534(.DIN1 (___0_____40436), .DIN2
       (__________________________________________0_), .Q
       (___0___22200));
  nor2s1 __9____513535(.DIN1
       (__________________________________________________________________21985),
       .DIN2
       (__________________________________________________________________21983),
       .Q (___0___22199));
  and2s1 __9____513536(.DIN1 (___0__9__40530), .DIN2 (___0__0__40501),
       .Q (___0___22198));
  and2s1 __9____513537(.DIN1 (___0_____40598), .DIN2 (_________22038),
       .Q (___0___22197));
  nor2s1 __9____513538(.DIN1 (___0_____40534), .DIN2
       (_____________________________________________21787), .Q
       (___00__22196));
  and2s1 __9__513539(.DIN1 (____0________________21720), .DIN2
       (____0_____________0___21723), .Q (___99));
  and2s1 __9_9__513540(.DIN1 (_____________________21684), .DIN2
       (__________________0___21686), .Q (___9___22195));
  nnd2s1 __9_0_513541(.DIN1 (_____________________21734), .DIN2
       (_____________________21733), .Q (________22472));
  nnd2s1 __9____513542(.DIN1 (_________________0___21687), .DIN2
       (_____________________21688), .Q (________22386));
  nor2s1 __9__0_513543(.DIN1 (_____________________21743), .DIN2
       (_________________9___21749), .Q (_______22248));
  nor2s1 __9____513544(.DIN1 (___0_____40598), .DIN2
       (_________________________________________________________________________________________22092),
       .Q (________22986));
  nnd2s1 __9____513545(.DIN1 (_____________________21677), .DIN2
       (_________________0___21676), .Q (________22381));
  nnd2s1 __9____513546(.DIN1 (_____________________21672), .DIN2
       (_____________________21673), .Q (________22385));
  nor2s1 __9____513547(.DIN1
       (____________________________________________21867), .DIN2
       (______________________________________________________________________________________0__22096),
       .Q (_____0__22559));
  nnd2s1 __9___513548(.DIN1 (___0__0__40413), .DIN2
       (_________________________________________________________________________________________22095),
       .Q (________22709));
  nnd2s1 __9____513549(.DIN1 (____0________________21717), .DIN2
       (____0________________21718), .Q (____0__22247));
  nnd2s1 __9____513550(.DIN1 (___0_____40621), .DIN2
       (_____________________________________9_______21882), .Q
       (____9___22544));
  and2s1 __9____513551(.DIN1 (__________9_), .DIN2 (___0_____40479), .Q
       (________22589));
  nnd2s1 __9____513552(.DIN1 (____0________________21720), .DIN2
       (____0________________21719), .Q (________22391));
  nor2s1 __9____513553(.DIN1 (_____________________21680), .DIN2
       (_____________________21681), .Q (________22389));
  nor2s1 __9____513554(.DIN1
       (______________________________________________21912), .DIN2
       (___0_____40436), .Q (_____0__22681));
  and2s1 __9____513555(.DIN1 (_______________22077), .DIN2
       (___0_0___40466), .Q (_____9__22662));
  nor2s1 __9____513556(.DIN1
       (__________________________________________________________________21999),
       .DIN2 (__________________________________________9___21934), .Q
       (_____0__22771));
  and2s1 __9____513557(.DIN1 (___0_____40549), .DIN2
       (_____________________________________________21770), .Q
       (________22675));
  and2s1 __9___513558(.DIN1
       (______________________________________________________________________________________0__22096),
       .DIN2 (____________________________________________21867), .Q
       (____09__22558));
  nnd2s1 __9____513559(.DIN1 (_____________________21709), .DIN2
       (_____________________21707), .Q (_______22253));
  nor2s1 __9____513560(.DIN1 (_____________________21675), .DIN2
       (_____________________21674), .Q (________22387));
  nor2s1 __9_513561(.DIN1
       (_________________________________________________________________________________________22095),
       .DIN2 (___0__0__40413), .Q (___0____22291));
  nor2s1 __9____513562(.DIN1 (_________22038), .DIN2
       (______________22065), .Q (____0___22746));
  nor2s1 __9____513563(.DIN1 (___0_____40438), .DIN2 (___0_____40437),
       .Q (________22984));
  or2s1 __9____513564(.DIN1 (______________________21700), .DIN2
       (______________________21701), .Q (____9___22546));
  nor2s1 __9____513565(.DIN1 (_________________0___21702), .DIN2
       (_____________________21703), .Q (____99__22548));
  nor2s1 __9____513566(.DIN1 (___0_____40602), .DIN2 (___0_____40415),
       .Q (________28146));
  nnd2s1 __9____513567(.DIN1 (____0_________________21724), .DIN2
       (____0_________________21725), .Q (________22536));
  nor2s1 __9__513568(.DIN1 (_________________0___21740), .DIN2
       (______________________21753), .Q (________22694));
  nnd2s1 __9__9_513569(.DIN1 (____0_________________21727), .DIN2
       (____0_________________21726), .Q (____0___22555));
  or2s1 __9____513570(.DIN1 (__________________0___21686), .DIN2
       (_____________________21684), .Q (_____9__23376));
  nor2s1 __9__9_513571(.DIN1 (_____________________21670), .DIN2
       (_____________________21671), .Q (___9____23156));
  nor2s1 __9____513572(.DIN1 (_____________________21746), .DIN2
       (_____________________21745), .Q (_____0__22899));
  nor2s1 __9__0_513573(.DIN1 (____0____________9_), .DIN2
       (____0________________21668), .Q (________22679));
  nnd2s1 __9____513574(.DIN1 (____0________________21665), .DIN2
       (____0________________21666), .Q (_____9__23635));
  nnd2s1 __9____513575(.DIN1 (_____________________21730), .DIN2
       (_____________________21731), .Q (____0___22743));
  or2s1 __9____513576(.DIN1 (__________________0___21738), .DIN2
       (______________________21739), .Q (________22689));
  nor2s1 __9__0_513577(.DIN1 (____0_________________21726), .DIN2
       (____0_________________21727), .Q (____9___23782));
  and2s1 __9____513578(.DIN1 (_____________________21671), .DIN2
       (_____________________21670), .Q (_____9__23028));
  nnd2s1 __9____513579(.DIN1 (__________________0_), .DIN2
       (_________________9_), .Q (________22860));
  or2s1 __9____513580(.DIN1 (_________________9_), .DIN2
       (__________________0_), .Q (____0___23042));
  and2s1 __9____513581(.DIN1 (______________________21739), .DIN2
       (__________________0___21738), .Q (____0___23412));
  nnd2s1 __9____513582(.DIN1 (_____________________21747), .DIN2
       (______________________21751), .Q (________26421));
  and2s1 __9___513583(.DIN1 (_____________________21708), .DIN2
       (_____________________21706), .Q (___0____23248));
  nor2s1 __9____513584(.DIN1 (_________________0___21728), .DIN2
       (_____________________21729), .Q (___9____24088));
  nnd2s1 __9___513585(.DIN1 (____0____________9___21722), .DIN2
       (____0_____________0___21723), .Q (________25756));
  nnd2s1 __9__513586(.DIN1 (__________________0___21750), .DIN2
       (______________________21751), .Q (____9___24062));
  nor2s1 __9____513587(.DIN1 (_____________________21688), .DIN2
       (_____________________21689), .Q (____0___25498));
  nor2s1 __9____513588(.DIN1 (_________________0___21676), .DIN2
       (_____________________21677), .Q (_________38301));
  nor2s1 __9____513589(.DIN1 (____0________________21718), .DIN2
       (____0________________21717), .Q (____0___23311));
  or2s1 __9_9_513590(.DIN1 (_____________22086), .DIN2
       (_____________________________________9_______21883), .Q
       (___9___22194));
  and2s1 __9__0_513591(.DIN1 (___0__0__40491), .DIN2 (___0_____40579),
       .Q (___9___22193));
  nnd2s1 __9_9__513592(.DIN1
       (_______________________________________________________________0__22010),
       .DIN2 (_____________________________________________21953), .Q
       (___9___22192));
  or2s1 __9__0_513593(.DIN1
       (____________________________________________21866), .DIN2
       (____________________________________________21831), .Q
       (___9___22191));
  nor2s1 __9_00_513594(.DIN1 (_________________9___21749), .DIN2
       (_________________________________________________________________________________________22089),
       .Q (___9___22190));
  or2s1 __9_0__513595(.DIN1
       (____________________________________________21820), .DIN2
       (____________________________________________21791), .Q (___9_));
  and2s1 __9____513596(.DIN1 (___0_____40417), .DIN2 (inData[26]), .Q
       (___90));
  nnd2s1 __9____513597(.DIN1 (___0_____40592), .DIN2
       (_____________22101), .Q (____9__22189));
  nor2s1 __9_99_513598(.DIN1
       (______________________________________________________________________________________0__22096),
       .DIN2 (_______________22070), .Q (_______22188));
  nnd2s1 __9_99_513599(.DIN1 (____0_____________0_), .DIN2
       (____0____________9_), .Q (_______22187));
  nor2s1 __9____513600(.DIN1 (_____________22101), .DIN2
       (___0_____40592), .Q (_______22186));
  nor2s1 __9____513601(.DIN1 (___0_____40576), .DIN2
       (_____________________________________________21796), .Q
       (_______22185));
  and2s1 __9____513602(.DIN1 (___0_____40586), .DIN2 (inData[6]), .Q
       (_______22184));
  nnd2s1 __9____513603(.DIN1
       (______________________________________________21931), .DIN2
       (inData[10]), .Q (_______22183));
  and2s1 __9_9__513604(.DIN1 (___0_____40588), .DIN2 (_________22016),
       .Q (_______22182));
  nnd2s1 __9_0__513605(.DIN1
       (______________________________________________________________________________________0__22096),
       .DIN2 (_______________22070), .Q (_______22181));
  nor2s1 __9____513606(.DIN1 (______________22110), .DIN2
       (___0_____40584), .Q (____0));
  and2s1 __9_00_513607(.DIN1
       (_________________________________________9___21861), .DIN2
       (inData[30]), .Q (____9));
  and2s1 __9____513608(.DIN1 (___0_____40596), .DIN2
       (_____________22099), .Q (_______22180));
  and2s1 __9____513609(.DIN1 (___0__0__40591), .DIN2 (_________9_), .Q
       (_______22179));
  or2s1 __9_9__513610(.DIN1 (_________22016), .DIN2 (___0_____40588),
       .Q (_______22178));
  nor2s1 __9_0__513611(.DIN1 (___0__9__40412), .DIN2
       (___________9___22071), .Q (_______22177));
  nnd2s1 __9_9__513612(.DIN1
       (_____________________________________________21940), .DIN2
       (inData[4]), .Q (_______22176));
  nnd2s1 __9_0__513613(.DIN1
       (______________________________________________21975), .DIN2
       (inData[30]), .Q (_______22175));
  or2s1 __9_0_513614(.DIN1 (_________________0___21740), .DIN2
       (_____________________21741), .Q (_______22174));
  nnd2s1 __9___513615(.DIN1 (___0_____40586), .DIN2
       (__________9___22107), .Q (_______22173));
  or2s1 __9____513616(.DIN1 (_________22014), .DIN2 (___0_____40594),
       .Q (_______22172));
  nor2s1 __9_0__513617(.DIN1 (______________22064), .DIN2
       (______________22067), .Q (_____));
  nnd2s1 __9_99_513618(.DIN1
       (_____________________________________0_______21759), .DIN2
       (inData[6]), .Q (___0___22171));
  nnd2s1 __9____513619(.DIN1
       (_____________________________________________21839), .DIN2
       (clk), .Q (___0___22170));
  nor2s1 __9___513620(.DIN1 (_____________22099), .DIN2
       (___0_____40596), .Q (___0_));
  or2s1 __9_0__513621(.DIN1
       (____________________________________________21807), .DIN2
       (____________________________________________21792), .Q (___00));
  nor2s1 __9_0__513622(.DIN1 (_______________22070), .DIN2
       (_________________________________________________________________________________________22094),
       .Q (__9___22169));
  nnd2s1 __9_0__513623(.DIN1 (____0________________21716), .DIN2
       (____0________________21719), .Q (__9___22168));
  nnd2s1 __9_0__513624(.DIN1 (__________9_), .DIN2
       (______________________________________________________________________________________0__22096),
       .Q (__9___22167));
  nnd2s1 __9_0__513625(.DIN1
       (______________________________________________21955), .DIN2
       (_________________________________________________________________22000),
       .Q (__9___22166));
  nor2s1 __9___513626(.DIN1 (__________9___22107), .DIN2
       (___0_____40586), .Q (__9_));
  nnd2s1 __9_0__513627(.DIN1 (_______________22075), .DIN2
       (_______________________________________________________________________________________),
       .Q (__90));
  nnd2s1 __9_99_513628(.DIN1
       (_____________________________________________21907), .DIN2
       (inData[6]), .Q (___9__22165));
  nnd2s1 __9_00_513629(.DIN1
       (_____________________________________9_____), .DIN2
       (inData[4]), .Q (______22164));
  and2s1 __9____513630(.DIN1 (___0_____40507), .DIN2 (inData[16]), .Q
       (______22163));
  nor2s1 __9____513631(.DIN1 (___0_____40622), .DIN2
       (_____________22080), .Q (______22162));
  nnd2s1 __9___513632(.DIN1 (___0_9___40556), .DIN2
       (_____________________________________________21782), .Q
       (______22161));
  nor2s1 __9__513633(.DIN1
       (______________________________________0_______21893), .DIN2
       (___0_____40617), .Q (______22160));
  or2s1 __9_9__513634(.DIN1 (___0__9__40520), .DIN2
       (_________________________________________0___21798), .Q
       (______22159));
  nnd2s1 __9_513635(.DIN1
       (______________________________________0_____), .DIN2
       (inData[16]), .Q (______22158));
  nnd2s1 __9__0_513636(.DIN1 (__________), .DIN2 (___0_99__40460), .Q
       (___0__22157));
  and2s1 __9_0__513637(.DIN1 (___0_0___40565), .DIN2
       (_________________________________________9___21803), .Q
       (___9__22156));
  or2s1 __9__513638(.DIN1
       (_____________________________________9_______21882), .DIN2
       (___0_____40621), .Q (______22155));
  nor2s1 __9____513639(.DIN1
       (_________________________________________________________________________________________22089),
       .DIN2 (_______________22076), .Q (________22891));
  nor2s1 __9____513640(.DIN1 (_______________22069), .DIN2
       (_________________________________________________________________________________________22095),
       .Q (________22530));
  nor2s1 __9_513641(.DIN1 (______________22064), .DIN2
       (_________________________________________________________________________________________22092),
       .Q (________22870));
  nor2s1 __9____513642(.DIN1 (___0_____40479), .DIN2 (__________9_), .Q
       (________22590));
  nnd2s1 __9_09_513643(.DIN1 (___________9___22071), .DIN2
       (_______________22073), .Q (________22713));
  nnd2s1 __9_0_513644(.DIN1 (______________22067), .DIN2
       (______________22064), .Q (____9___22641));
  nor2s1 __9___513645(.DIN1 (__________________0___21712), .DIN2
       (_____________________21710), .Q (________22399));
  nor2s1 __9____513646(.DIN1 (_______________22072), .DIN2
       (_______________22074), .Q (_______22257));
  nor2s1 __9____513647(.DIN1 (_________________9___21685), .DIN2
       (_____________________21684), .Q (_______22255));
  nnd2s1 __9___513648(.DIN1 (____0________________21664), .DIN2
       (____0________________21663), .Q (________22379));
  and2s1 __9_0__513649(.DIN1 (_____________________21741), .DIN2
       (_________________0___21740), .Q (________22594));
  nnd2s1 __9____513650(.DIN1 (___0_____40539), .DIN2
       (_____________________________________0_______21759), .Q
       (________22599));
  nor2s1 __9____513651(.DIN1 (___0_0___40466), .DIN2
       (_______________22077), .Q (________22661));
  nor2s1 __9____513652(.DIN1 (_________________0___21687), .DIN2
       (_____________________21690), .Q (_____9__22383));
  nor2s1 __9____513653(.DIN1 (____0________________21666), .DIN2
       (____0________________21665), .Q (_______22249));
  nnd2s1 __9____513654(.DIN1 (_____________________21710), .DIN2
       (__________________0___21712), .Q (________22390));
  nnd2s1 __9___513655(.DIN1 (_____________________21695), .DIN2
       (____________________), .Q (_______22256));
  nnd2s1 __9____513656(.DIN1 (_____________________21709), .DIN2
       (_________________9___21711), .Q (_______22251));
  nnd2s1 __9_0__513657(.DIN1 (____0________________21668), .DIN2
       (____0____________9_), .Q (____0___22365));
  and2s1 __9____513658(.DIN1 (___0_0___40464), .DIN2 (___0_____40483),
       .Q (_____0__22909));
  or2s1 __9____513659(.DIN1 (_________________9___21685), .DIN2
       (__________________0___21686), .Q (____90__22539));
  nnd2s1 __9__0_513660(.DIN1 (_________________9___21696), .DIN2
       (__________________0___21697), .Q (________22786));
  and2s1 __9____513661(.DIN1 (___0_____40504), .DIN2 (___0_____40516),
       .Q (____9___25949));
  nor2s1 __9__513662(.DIN1 (__________________0___21697), .DIN2
       (_________________9___21696), .Q (____0___22840));
  nor2s1 __9____513663(.DIN1 (____0_____________0_), .DIN2
       (____0________________21667), .Q (________22625));
  nnd2s1 __9____513664(.DIN1 (___0_____40536), .DIN2
       (_____________________________________________21784), .Q
       (________25354));
  and2s1 __9____513665(.DIN1 (______________________21698), .DIN2
       (______________________21700), .Q (________22696));
  nor2s1 __9____513666(.DIN1 (_____________________21695), .DIN2
       (____________________), .Q (________22855));
  nnd2s1 __9____513667(.DIN1
       (_____________________________________9_______21883), .DIN2
       (_____________22086), .Q (_________38649));
  nnd2s1 __9____513668(.DIN1 (_____________________21705), .DIN2
       (_____________________21703), .Q (____9___22734));
  nnd2s1 __9__9_513669(.DIN1 (_____________________21689), .DIN2
       (_____________________21688), .Q (____0___22843));
  hi1s1 __9____513670(.DIN (______22154), .Q (________24282));
  nnd2s1 __9____513671(.DIN1 (_____________________21745), .DIN2
       (_____________________21746), .Q (____0___22648));
  nor2s1 __9____513672(.DIN1 (____0______________), .DIN2
       (____0____________0_), .Q (____9___22933));
  nnd2s1 __9____513673(.DIN1 (_________________9___21685), .DIN2
       (__________________0___21686), .Q (________22672));
  or2s1 __9___513674(.DIN1 (____0_____________0___21723), .DIN2
       (____0____________9___21722), .Q (___9____23150));
  nor2s1 __9___513675(.DIN1 (______________________21752), .DIN2
       (_____________________21741), .Q (___0____25161));
  nnd2s1 __9____513676(.DIN1 (______________________21699), .DIN2
       (______________________21701), .Q (_____9___36725));
  nnd2s1 __9____513677(.DIN1 (____0________________21667), .DIN2
       (____0________________21665), .Q (_________38203));
  nnd2s1 __9__0_513678(.DIN1 (_____________________21729), .DIN2
       (_________________0___21728), .Q (________23384));
  nnd2s1 __9____513679(.DIN1 (____0____________9___21722), .DIN2
       (____0________________21721), .Q (_________38838));
  nor2s1 __9__0_513680(.DIN1 (_____________________21748), .DIN2
       (_____________________21746), .Q (___99___26049));
  nnd2s1 __9__0_513681(.DIN1 (_________________9___21749), .DIN2
       (_____________________21748), .Q (_____9___38319));
  or2s1 __9____513682(.DIN1 (____0________________21663), .DIN2
       (____0________________21664), .Q (________24300));
  nnd2s1 __9__9_513683(.DIN1 (_____________________21674), .DIN2
       (_____________________21675), .Q (________24703));
  nnd2s1 __9___513684(.DIN1 (_____________________21746), .DIN2
       (_____________________21748), .Q (________26440));
  or2s1 __9__513685(.DIN1 (_____________________21708), .DIN2
       (_____________________21706), .Q (_____9__23900));
  and2s1 __9___513686(.DIN1 (______________________21753), .DIN2
       (_________________0___21740), .Q (________25942));
  hi1s1 __9__513687(.DIN (__________________________________________),
       .Q (______22152));
  hi1s1 __9____513688(.DIN (____0________________21664), .Q
       (______22151));
  hi1s1 __9____513689(.DIN (______0__22040), .Q (______22150));
  hi1s1 __9__513690(.DIN
       (_____________________________________________21941), .Q
       (___0__22149));
  hi1s1 __9____513691(.DIN (___0_____40506), .Q (______22148));
  hi1s1 __9____513692(.DIN (_____________________21674), .Q
       (______22147));
  hi1s1 __9___513693(.DIN (___0_____40516), .Q (______22146));
  hi1s1 __9__9_513694(.DIN
       (_________________________________________0___21824), .Q
       (______22145));
  hi1s1 __9___513695(.DIN (___0_____40446), .Q (______22144));
  hi1s1 __9____513696(.DIN (___0_____40527), .Q (___9__22143));
  hi1s1 __9__9_513697(.DIN
       (_____________________________________________21825), .Q
       (______22142));
  hi1s1 __9____513698(.DIN
       (______________________________________0______21887), .Q
       (______22141));
  hi1s1 __9____513699(.DIN
       (_____________________________________________21852), .Q
       (______22140));
  hi1s1 __9___513700(.DIN
       (_____________________________________________21799), .Q
       (______22139));
  hi1s1 __9____513701(.DIN (___0_____40607), .Q (______22138));
  hi1s1 __9____513702(.DIN (___0_____40617), .Q (___9__22137));
  hi1s1 __9____513703(.DIN
       (______________________________________0_______21890), .Q
       (______22136));
  hi1s1 __9____513704(.DIN
       (______________________________________________21916), .Q
       (______22135));
  hi1s1 __9__0_513705(.DIN
       (____________________________________________21793), .Q
       (___0__22134));
  hi1s1 __9__9_513706(.DIN
       (_________________________________________________________________22001),
       .Q (___9__22133));
  hi1s1 __9____513707(.DIN
       (_____________________________________________21810), .Q
       (______22132));
  hi1s1 __9____513708(.DIN
       (_____________________________________0______21754), .Q
       (______22131));
  hi1s1 __9____513709(.DIN (__________________0_), .Q (______22130));
  hi1s1 __9____513710(.DIN
       (_____________________________________________21928), .Q
       (________22439));
  hi1s1 __9__0_513711(.DIN (____0________________21665), .Q
       (________22382));
  hi1s1 __9____513712(.DIN (_____________________21734), .Q
       (________22401));
  hi1s1 __9____513713(.DIN (_____________________21673), .Q
       (____9__22261));
  hi1s1 __9____513714(.DIN
       (_____________________________________________21897), .Q
       (____0___27923));
  hi1s1 __9___513715(.DIN (_________0_), .Q (___009));
  hi1s1 __9____513716(.DIN (___0_____40478), .Q (___0____22313));
  hi1s1 __9____513717(.DIN
       (__________________________________________0___21935), .Q
       (________22470));
  hi1s1 __9____513718(.DIN (_____________________21682), .Q
       (______22153));
  hi1s1 __9____513719(.DIN
       (_____________________________________________21769), .Q
       (________24055));
  hi1s1 __9____513720(.DIN (___0__9__40450), .Q (___0_9__22343));
  hi1s1 __9___513721(.DIN
       (_____________________________________________21837), .Q
       (________22561));
  hi1s1 __9__9_513722(.DIN (_____________22080), .Q (___09___22357));
  hi1s1 __9__9_513723(.DIN (___0_____40524), .Q (________22396));
  hi1s1 __9__0_513724(.DIN
       (______________________________________________21937), .Q
       (________23476));
  hi1s1 __9____513725(.DIN (___0_____40517), .Q (________22524));
  hi1s1 __9____513726(.DIN (_____________22085), .Q (___0____22346));
  hi1s1 __9__0_513727(.DIN (___0__9__40540), .Q (________22424));
  hi1s1 __9____513728(.DIN (___0_9___40453), .Q (________22395));
  hi1s1 __9____513729(.DIN
       (_________________________________________________________________21991),
       .Q (____9___26770));
  hi1s1 __9___513730(.DIN (___0_9___40459), .Q (________22398));
  hi1s1 __9____513731(.DIN (inData[0]), .Q (________22485));
  hi1s1 __9____513732(.DIN
       (______________________________________0_______21894), .Q
       (________24431));
  hi1s1 __9____513733(.DIN (___0_____40624), .Q (________22504));
  hi1s1 __9____513734(.DIN (inData[16]), .Q (_____0__22499));
  hi1s1 __9____513735(.DIN (_____________________21672), .Q
       (_______22260));
  hi1s1 __9__513736(.DIN (_____________22088), .Q (________22502));
  hi1s1 __9____513737(.DIN
       (_____________________________________9_______21884), .Q
       (________22480));
  hi1s1 __9___513738(.DIN (___0__9__40580), .Q (________24494));
  hi1s1 __9____513739(.DIN (____0____________0___21713), .Q
       (_______22258));
  hi1s1 __9__513740(.DIN (_____________________21681), .Q
       (____0___22457));
  hi1s1 __9____513741(.DIN
       (____________________________________________21850), .Q
       (________24514));
  hi1s1 __9____513742(.DIN
       (____________________________________________21832), .Q
       (___0_____30727));
  hi1s1 __9__0_513743(.DIN (___0_____40486), .Q (_________36583));
  hi1s1 __9____513744(.DIN
       (_____________________________________________21767), .Q
       (____0____36194));
  hi1s1 __9____513745(.DIN
       (_____________________________________________21766), .Q
       (____0____35320));
  hi1s1 __9___513746(.DIN (____0________________21721), .Q
       (_______22252));
  hi1s1 __9____513747(.DIN
       (_________________________________________9___21901), .Q
       (_________38767));
  hi1s1 __9____513748(.DIN (___0_____40508), .Q (___0_____30948));
  hi1s1 __9____513749(.DIN
       (____________________________________________21864), .Q
       (_________33293));
  hi1s1 __9___513750(.DIN (__________), .Q (____99));
  hi1s1 __9____513751(.DIN (_________________9___21696), .Q
       (________22994));
  hi1s1 __9____513752(.DIN (___0_00__40561), .Q (_________33591));
  hi1s1 __9____513753(.DIN
       (_____________________________________0_____), .Q
       (_________34601));
  hi1s1 __9____513754(.DIN (____0________________21719), .Q
       (________22705));
  hi1s1 __9__513755(.DIN (____0_________________21726), .Q
       (________22400));
  hi1s1 __9____513756(.DIN (_____________________21688), .Q
       (___9_9__23181));
  hi1s1 __9___513757(.DIN (_____________________21748), .Q
       (________22397));
  hi1s1 __9__0_513758(.DIN (___0_____40529), .Q (_____0___33534));
  hi1s1 __9____513759(.DIN (___0__9__40520), .Q (____0___28017));
  hi1s1 __9____513760(.DIN (______________22066), .Q (___0____23297));
  hi1s1 __9__0_513761(.DIN (____0_____________0_), .Q (________22678));
  hi1s1 __9____513762(.DIN (______________22064), .Q (______9__31640));
  hi1s1 __9____513763(.DIN (___0_____40505), .Q (_________37748));
  hi1s1 __9__9_513764(.DIN (_____________________21692), .Q
       (________22461));
  hi1s1 __9__513765(.DIN (___0_____40487), .Q (_________36852));
  hi1s1 __9____513766(.DIN (_________________9___21711), .Q
       (________22532));
  hi1s1 __9____513767(.DIN
       (_________________________________________________________________________________________22095),
       .Q (_________33117));
  hi1s1 __9__9_513768(.DIN (_________________0___21702), .Q
       (________22513));
  hi1s1 __9____513769(.DIN (___0_____40432), .Q (___9_____39773));
  hi1s1 __9____513770(.DIN
       (_______________________________________________________________________________________),
       .Q (________27043));
  hi1s1 __9____513771(.DIN (_____________________21695), .Q
       (________23362));
  hi1s1 __9___513772(.DIN (_________________0___21687), .Q
       (________22884));
  hi1s1 __9____513773(.DIN (____0____________0_), .Q (_____9__22868));
  hi1s1 __9____513774(.DIN (______________________21753), .Q
       (_____0__22384));
  hi1s1 __9___513775(.DIN (inData[10]), .Q (_____00__34847));
  hi1s1 __9____513776(.DIN (___0_0___40566), .Q (_________36883));
  hi1s1 __9____513777(.DIN (_____________________21684), .Q
       (___9____23149));
  hi1s1 __9____513778(.DIN (_____________________21693), .Q
       (________23026));
  hi1s1 __9____513779(.DIN (_________________0_), .Q (___9_____39397));
  hi1s1 __9____513780(.DIN (____0________________21714), .Q
       (________22857));
  hi1s1 __9____513781(.DIN (______________________21751), .Q
       (________26217));
  hi1s1 __9__0_513782(.DIN (_____________________21707), .Q
       (____9___23032));
  hi1s1 __9____513783(.DIN (____0____________9___21722), .Q
       (___0____26120));
  hi1s1 __9___513784(.DIN (inData[28]), .Q (_________35587));
  hi1s1 __9____513785(.DIN (___0_____40411), .Q (______9__34981));
  hi1s1 __9____513786(.DIN (inData[6]), .Q (___9_0__29602));
  hi1s1 __9____513787(.DIN (_____________________21741), .Q
       (________22754));
  hi1s1 __9____513788(.DIN (_____________________21709), .Q
       (________24602));
  hi1s1 __9____513789(.DIN (inData[12]), .Q (________26530));
  hi1s1 __9__9_513790(.DIN (_______________22070), .Q (_________34167));
  hi1s1 __9____513791(.DIN (______________________21698), .Q
       (_____0__23445));
  hi1s1 __9____513792(.DIN (______________22065), .Q (_________32611));
  hi1s1 __9___513793(.DIN (_____________________21705), .Q
       (________23754));
  hi1s1 __9____513794(.DIN (_____________________21731), .Q
       (_____9__24325));
  hi1s1 __9____513795(.DIN
       (______________________________________________________________________________________0__22093),
       .Q (_________37867));
  hi1s1 __9____513796(.DIN (inData[31]), .Q (_________32159));
  hi1s1 __9__513797(.DIN (_______________22069), .Q (_________33973));
  hi1s1 __9____513798(.DIN (____0________________21662), .Q
       (_____9__24635));
  hi1s1 __9___513799(.DIN (_______________22077), .Q (_________35844));
  hi1s1 __9____513800(.DIN (_________________9___21737), .Q
       (_____9___37752));
  hi1s1 __9____513801(.DIN
       (_________________________________________________________________________________________22089),
       .Q (_________37789));
  hi1s1 __9____513802(.DIN (_______________22072), .Q (_________36762));
  hi1s1 __9____513803(.DIN (_____________________21691), .Q
       (________23989));
  hi1s1 __9____513804(.DIN
       (_________________________________________________________________________________________22091),
       .Q (_________36402));
  hi1s1 __9____513805(.DIN (_______________22074), .Q (_________37320));
  hi1s1 __9__9_513806(.DIN (_______________22076), .Q (____99___36174));
  hi1s1 __9____513807(.DIN (_________________9___21749), .Q
       (____0____37167));
  hi1s1 __9____513808(.DIN (_____________________21742), .Q
       (________26426));
  hi1s1 __9__9_513809(.DIN (____0________________21720), .Q
       (________23959));
  hi1s1 __9___513810(.DIN (_____________________21736), .Q
       (______22154));
  hi1s1 __9____513811(.DIN (_____________________21745), .Q
       (___9____26912));
  hi1s1 __9____513812(.DIN (_______________22073), .Q (_________37321));
  hi1s1 __9____513813(.DIN
       (______________________________________________________________________________________0),
       .Q (_________36761));
  hi1s1 __9___513814(.DIN
       (_____________________________________0______21757), .Q
       (______22129));
  hi1s1 __9____513815(.DIN
       (____________________________________________21820), .Q
       (______22128));
  hi1s1 __9___513816(.DIN (____0____________9_), .Q (______22127));
  hi1s1 __9____513817(.DIN
       (______________________________________0______21886), .Q
       (______22126));
  hi1s1 __9____513818(.DIN
       (__________________________________________9___21918), .Q
       (______22125));
  hi1s1 __9__9_513819(.DIN (______________22103), .Q (___9));
  hi1s1 __9__0_513820(.DIN (___0_____40597), .Q (______22124));
  hi1s1 __9___513821(.DIN (_________________9_), .Q (______22123));
  hi1s1 __9____513822(.DIN
       (__________________________________________0___21981), .Q
       (______22122));
  hi1s1 __9____513823(.DIN
       (_____________________________________________21853), .Q
       (______22121));
  hi1s1 __9___513824(.DIN (___0_____40537), .Q (______22120));
  hi1s1 __9__9_513825(.DIN
       (____________________________________________21848), .Q
       (______22119));
  hi1s1 __9____513826(.DIN (_______________0), .Q (____));
  hi1s1 __9__9_513827(.DIN (___0_____40547), .Q (___0));
  hi1s1 __9___513828(.DIN (___0_____40492), .Q (_____22118));
  hi1s1 __9____513829(.DIN
       (__________________________________________0_), .Q (_____22117));
  hi1s1 __9____513830(.DIN (___0_____40589), .Q (_____22116));
  hi1s1 __9____513831(.DIN
       (_____________________________________________21768), .Q
       (_____22115));
  hi1s1 __9____513832(.DIN
       (____________________________________________21833), .Q
       (_____22114));
  hi1s1 __9____513833(.DIN
       (_____________________________________________21969), .Q
       (_____22113));
  hi1s1 __9____513834(.DIN
       (_________________________________________________________________22000),
       .Q (___));
  hi1s1 __9___513835(.DIN (___0_____40445), .Q (__0));
  hi1s1 __9____513836(.DIN (___0_____40493), .Q (________22394));
  hi1s1 __9____513837(.DIN (___0_____40587), .Q (___0____22300));
  hi1s1 __9___513838(.DIN (___0_____40579), .Q (_________33187));
  hi1s1 __9__513839(.DIN (_____________22084), .Q (____9___22930));
  hi1s1 __9____513840(.DIN
       (_____________________________________________21811), .Q
       (___90__22262));
  hi1s1 __9____513841(.DIN (______0___22054), .Q (____9___22636));
  hi1s1 __9____513842(.DIN (______________22111), .Q (_______22280));
  hi1s1 __9____513843(.DIN (inData[4]), .Q (____00));
  hi1s1 __9____513844(.DIN (___0_____40525), .Q (____9___24637));
  hi1s1 __9____513845(.DIN (____0________________21668), .Q
       (_______22259));
  hi1s1 __9____513846(.DIN (___0_____40532), .Q (________25248));
  hi1s1 __9____513847(.DIN (___0_____40536), .Q (________25838));
  hi1s1 __9__9_513848(.DIN (______________________21701), .Q
       (____9___22545));
  hi1s1 __9__9_513849(.DIN (___0_____40484), .Q (___0____22340));
  hi1s1 __9____513850(.DIN
       (_________________________________________0___21814), .Q
       (_____9__23871));
  hi1s1 __9____513851(.DIN (___0_____40449), .Q (___09___22355));
  hi1s1 __9____513852(.DIN
       (_____________________________________________21953), .Q
       (___0____22317));
  hi1s1 __9____513853(.DIN (___0__9__40510), .Q (___9____23140));
  hi1s1 __9____513854(.DIN
       (____________________________________________21774), .Q
       (____9____32454));
  hi1s1 __9____513855(.DIN
       (______________________________________0___0_), .Q
       (________22611));
  hi1s1 __9____513856(.DIN (___0_00__40461), .Q (_____9__22392));
  hi1s1 __9____513857(.DIN
       (____________________________________________), .Q
       (____9____37062));
  hi1s1 __9____513858(.DIN (_____________________21733), .Q
       (___9___22263));
  hi1s1 __9___513859(.DIN (___0__9__40480), .Q (_____0__22403));
  hi1s1 __9___513860(.DIN (___0_09__40570), .Q (______9__35974));
  hi1s1 __9___513861(.DIN
       (______________________________________________21933), .Q
       (________22772));
  hi1s1 __9____513862(.DIN
       (_______________________________________________________________0__22010),
       .Q (________22369));
  hi1s1 __9___513863(.DIN
       (____________________________________________21851), .Q
       (____9___23131));
  hi1s1 __9____513864(.DIN (inData[24]), .Q (___09___22360));
  hi1s1 __9____513865(.DIN (__________22059), .Q (________22669));
  hi1s1 __9____513866(.DIN (_____9___22051), .Q (_____00__33066));
  hi1s1 __9____513867(.DIN (__________________0___21697), .Q
       (________22380));
  hi1s1 __9___513868(.DIN (___0_____40548), .Q (_________32032));
  hi1s1 __9____513869(.DIN (_____________________21675), .Q
       (________22388));
  hi1s1 __9__9_513870(.DIN
       (____________________________________________21806), .Q
       (_____0___33161));
  hi1s1 __9____513871(.DIN
       (______________________________________________21960), .Q
       (_____9__22577));
  hi1s1 __9__9_513872(.DIN
       (_______________________________________________________________0),
       .Q (_____9__22567));
  hi1s1 __9__0_513873(.DIN (____0________________21663), .Q
       (_______22254));
  hi1s1 __9____513874(.DIN (_____________________21704), .Q
       (_____9__22402));
  hi1s1 __9___513875(.DIN (___0_9___40559), .Q (________26819));
  hi1s1 __9____513876(.DIN (___0_____40427), .Q (________26698));
  hi1s1 __9____513877(.DIN
       (_________________________________________9___21779), .Q
       (________22420));
  hi1s1 __9____513878(.DIN (_____________________21708), .Q
       (_____0__22393));
  hi1s1 __9____513879(.DIN
       (_____________________________________________21910), .Q
       (____9___25676));
  hi1s1 __9___513880(.DIN (____0________________21715), .Q
       (_______22250));
  hi1s1 __9__0_513881(.DIN (____0______________), .Q (________23474));
  hi1s1 __9____513882(.DIN (inData[2]), .Q (________25850));
  hi1s1 __9____513883(.DIN (_____________________21680), .Q
       (________22924));
  hi1s1 __9____513884(.DIN (inData[18]), .Q (____9____38963));
  hi1s1 __9__0_513885(.DIN
       (_____________________________________________21858), .Q
       (____0____36220));
  hi1s1 __9____513886(.DIN (___0__0__40541), .Q (____9____35264));
  hi1s1 __9__9_513887(.DIN (___0__9__40590), .Q (________27071));
  hi1s1 __9___513888(.DIN (____________________), .Q (____00__23407));
  hi1s1 __9____513889(.DIN
       (_______________________________________________________________0__21998),
       .Q (_________37424));
  hi1s1 __9____513890(.DIN (______________22112), .Q (_____9__22633));
  hi1s1 __9____513891(.DIN (_____________________21710), .Q
       (________23021));
  hi1s1 __9____513892(.DIN
       (_____________________________________________21857), .Q
       (_________37245));
  hi1s1 __9____513893(.DIN (inData[8]), .Q (__99____30501));
  hi1s1 __9____513894(.DIN
       (_____________________________________0____), .Q
       (_________33206));
  hi1s1 __9____513895(.DIN (_________________9___21685), .Q
       (________22627));
  hi1s1 __9___513896(.DIN
       (__________________________________________________________________21993),
       .Q (___0_____40045));
  hi1s1 __9____513897(.DIN (______________________21739), .Q
       (___9_9__23163));
  hi1s1 __9____513898(.DIN (inData[26]), .Q (____9___23878));
  hi1s1 __9__9_513899(.DIN
       (_____________________________________________21801), .Q
       (____0_0__36258));
  hi1s1 __9____513900(.DIN (____0________________21717), .Q
       (________23024));
  hi1s1 __9____513901(.DIN (inData[20]), .Q (___9____25102));
  hi1s1 __9___513902(.DIN (____________), .Q (_________35727));
  hi1s1 __9____513903(.DIN (_____________________21743), .Q
       (____09__23048));
  hi1s1 __9__0_513904(.DIN (_____________________21729), .Q
       (________22727));
  hi1s1 __9____513905(.DIN (_____________________21690), .Q
       (___0____23256));
  hi1s1 __9____513906(.DIN (_____________________21671), .Q
       (________23356));
  hi1s1 __9__0_513907(.DIN (______________________21699), .Q
       (________23449));
  hi1s1 __9__0_513908(.DIN (____0_________________21727), .Q
       (________23611));
  hi1s1 __9____513909(.DIN
       (_________________________________________________________________________________________22094),
       .Q (____9___22447));
  hi1s1 __9____513910(.DIN (_____________________21689), .Q
       (_____9__23444));
  hi1s1 __9____513911(.DIN (______________________21752), .Q
       (________22628));
  hi1s1 __9__513912(.DIN (_____________________21694), .Q
       (____0___22846));
  hi1s1 __9____513913(.DIN (___________________), .Q (_____00__35736));
  hi1s1 __9___513914(.DIN (_____________________21746), .Q
       (________23555));
  hi1s1 __9____513915(.DIN (inData[22]), .Q (____0_0__38093));
  hi1s1 __9____513916(.DIN (___0_____40598), .Q (_____9__23492));
  hi1s1 __9____513917(.DIN (_____________________21730), .Q
       (________23734));
  hi1s1 __9____513918(.DIN (____0________________21716), .Q
       (____00__23597));
  hi1s1 __9___513919(.DIN (clk), .Q (___99____39814));
  hi1s1 __9___513920(.DIN (_____________________21747), .Q
       (____90__26673));
  hi1s1 __9___513921(.DIN
       (______________________________________________21906), .Q
       (___9_9___39696));
  hi1s1 __9____513922(.DIN (inData[14]), .Q (__99_9__30508));
  hi1s1 __9____513923(.DIN (____0_________________21725), .Q
       (___9____23151));
  hi1s1 __9____513924(.DIN (_____________________21683), .Q
       (___0____23252));
  hi1s1 __9____513925(.DIN
       (_________________________________________________________________________________________22090),
       .Q (_________34538));
  hi1s1 __9___513926(.DIN (_____________________21679), .Q
       (____0___23697));
  hi1s1 __9____513927(.DIN (____0_________________21724), .Q
       (____90__24060));
  hi1s1 __9____513928(.DIN (_____________________21678), .Q
       (_____9__23842));
  hi1s1 __9____513929(.DIN
       (_________________________________________________________________________________________22092),
       .Q (______9__32360));
  hi1s1 __9____513930(.DIN (_____________________21732), .Q
       (____9___24066));
  hi1s1 __9____513931(.DIN (____0________________21667), .Q
       (____0___23599));
  hi1s1 __9____513932(.DIN (___0__0__40413), .Q (______9__32959));
  hi1s1 __9____513933(.DIN (______________22067), .Q (_________32918));
  hi1s1 __9__9_513934(.DIN
       (______________________________________________________________________________________0__22096),
       .Q (_____0___32287));
  hi1s1 __9____513935(.DIN (___0__9__40412), .Q (_________36493));
  hi1s1 __9___513936(.DIN (_____________________21744), .Q
       (________26431));
  hi1s1 __9___513937(.DIN (__________9_), .Q (_____9___33157));
  hi1s1 __9____513938(.DIN (_______________22075), .Q (_________37412));
  ib1s1 __9__9_513939(.DIN (____0_______________), .Q (____9___23970));
  hi1s1 __9___513940(.DIN (___________9___22071), .Q (_________36556));
  hi1s1 __9__9_513941(.DIN (_____________________21677), .Q
       (___9_9___39790));
  hi1s1 __9___513942(.DIN (_____________________21669), .Q
       (________24475));
  hi1s1 __9__9_513943(.DIN (__________________0___21750), .Q
       (____0___26590));
  or2s1 __(.DIN1 (___0__0__40629), .DIN2 (_________35635), .Q
       (___0_____40630));
  xnr2s1 __513944(.DIN1 (___9_____39301), .DIN2 (_________35661), .Q
       (___0__0__40629));
  nor2s1 __9____513945(.DIN1 (___0_____40631), .DIN2 (_________34733),
       .Q (___0_____40632));
  xnr2s1 __9___513946(.DIN1 (___909___39065), .DIN2 (______9__34705),
       .Q (___0_____40631));
  and2s1 __9___513947(.DIN1 (___0_____40633), .DIN2 (____9____33380),
       .Q (___0_____40634));
  xor2s1 __9____513948(.DIN1 (_________33318), .DIN2 (___00____39910),
       .Q (___0_____40633));
  nor2s1 __9____513949(.DIN1 (___0_____40635), .DIN2 (_________33260),
       .Q (___0_____40636));
  xnr2s1 __9____513950(.DIN1 (___9_____39372), .DIN2 (_________33214),
       .Q (___0_____40635));
  and2s1 __9____513951(.DIN1 (___0_____40637), .DIN2 (___0_____31038),
       .Q (___0__9__40638));
  xnr2s1 __9____513952(.DIN1 (____0____36215), .DIN2 (___0_0___31220),
       .Q (___0_____40637));
  or2s1 __9____513953(.DIN1 (___0__0__40639), .DIN2 (________28939), .Q
       (___0_____40640));
  xor2s1 __9____513954(.DIN1 (_________33973), .DIN2 (________28165),
       .Q (___0__0__40639));
  or2s1 __9____513955(.DIN1 (___0_____40641), .DIN2 (___99___26043), .Q
       (___0_____40642));
  xnr2s1 __9___513956(.DIN1 (_____0___32287), .DIN2 (____9___26222), .Q
       (___0_____40641));
  or2s1 __9___513957(.DIN1 (___0_____40643), .DIN2 (________25898), .Q
       (___0_____40644));
  xnr2s1 __9____513958(.DIN1 (_________36761), .DIN2 (________25897),
       .Q (___0_____40643));
  ib1s1 _________9____(.DIN (____9____38953), .Q (____9____38965));
  ib1s1 _________9__9_(.DIN (___9_00__39527), .Q (___0_9___40645));
  ib1s1 _________9__09(.DIN (___0_____40647), .Q (___0_____40646));
  ib1s1 _________9___0(.DIN (_________36079), .Q (___0_____40647));
  ib1s1 _________9____513959(.DIN (______________22068), .Q
       (_________33321));
  ib1s1 _________9____513960(.DIN (___0_____40649), .Q
       (___0__0__40648));
  ib1s1 _________9____513961(.DIN (___00____39970), .Q
       (___0_____40649));
  ib1s1 _________9____513962(.DIN (___0_____40651), .Q
       (___0_____40650));
  ib1s1 _________9____513963(.DIN (___9_____39332), .Q
       (___0_____40651));
  ib1s1 _________9____513964(.DIN (_________35799), .Q
       (___0_____40652));
  ib1s1 _________9____513965(.DIN (_________35847), .Q
       (_________35799));
  ib1s1 _________9____513966(.DIN (___0_9___40654), .Q
       (___0_9___40653));
  ib1s1 _________9____513967(.DIN (___9__0__39136), .Q
       (___0_9___40654));
  nb1s1 _________9__0_(.DIN (___0_____31037), .Q (___0909__40655));
  xnr2s1 __9____513968(.DIN1 (___9_9___39696), .DIN2 (___9_____39752),
       .Q (___09____40657));
  and2s1 __9____513969(.DIN1
       (__________________________________________0___21959), .DIN2
       (___0__0__40283), .Q (___09____40658));
  or2s1 __9____513970(.DIN1 (___00____39962), .DIN2 (___99____39866),
       .Q (___09____40659));
  and2s1 __9____513971(.DIN1 (___09____40657), .DIN2 (___9_____39758),
       .Q (___09_9__40660));
  xnr2s1 __9____513972(.DIN1 (___9_____39685), .DIN2 (___9_9___39701),
       .Q (___09_0__40661));
  xnr2s1 __9____513973(.DIN1 (___9_____39444), .DIN2 (___9_____39464),
       .Q (___09____40662));
  xnr2s1 __9____513974(.DIN1 (___0__0__40609), .DIN2 (___0_____40428),
       .Q (___09____40663));
  xnr2s1 __9____513975(.DIN1
       (_____________________________________________21828), .DIN2
       (_____9__23123), .Q (___09____40664));
  xnr2s1 __9___513976(.DIN1 (_________38716), .DIN2 (_________38735),
       .Q (___09____40665));
  xnr2s1 __9___513977(.DIN1 (_____0___38333), .DIN2 (______0__38527),
       .Q (___09____40666));
  xnr2s1 __9____513978(.DIN1 (____9____37989), .DIN2 (____999__38037),
       .Q (___09____40667));
  xnr2s1 __9____513979(.DIN1 (_________37922), .DIN2 (____0____40764),
       .Q (___09____40668));
  or2s1 __9____513980(.DIN1 (_____99__37759), .DIN2 (________28979), .Q
       (___09____40669));
  xnr2s1 __9____513981(.DIN1 (_________37695), .DIN2 (___9_____39312),
       .Q (___09_9__40670));
  and2s1 __9____513982(.DIN1 (_________37510), .DIN2 (_________37502),
       .Q (___09_0__40671));
  xnr2s1 __9____513983(.DIN1 (___0_0___40468), .DIN2 (_________37412),
       .Q (___09____40672));
  and2s1 __9____513984(.DIN1 (_________36771), .DIN2 (_________36899),
       .Q (___09____40673));
  or2s1 __9____513985(.DIN1 (______0__36784), .DIN2 (____9____35235),
       .Q (___09____40674));
  xnr2s1 __9___513986(.DIN1 (___0_____40473), .DIN2 (___0_____40474),
       .Q (___09____40675));
  xnr2s1 __9___513987(.DIN1 (______9__36295), .DIN2 (_____9___37367),
       .Q (___09____40676));
  xnr2s1 __9____513988(.DIN1 (____9_9__36130), .DIN2 (______9__35906),
       .Q (___09____40677));
  xnr2s1 __9____513989(.DIN1 (___0_____40543), .DIN2 (______9__35627),
       .Q (___09____40678));
  xnr2s1 __9____513990(.DIN1
       (_____________________________________________21822), .DIN2
       (______9__34997), .Q (___09____40679));
  xnr2s1 __9____513991(.DIN1 (_____99__22053), .DIN2
       (_____________________________________0___0_), .Q
       (___09_9__40680));
  xnr2s1 __9____513992(.DIN1 (___0_____40529), .DIN2 (_________22047),
       .Q (___09_0__40681));
  xor2s1 __9____513993(.DIN1 (______0__34622), .DIN2 (_____9___33150),
       .Q (___09____40682));
  xnr2s1 __9____513994(.DIN1 (__90____29684), .DIN2 (_________38587),
       .Q (_________38729));
  or2s1 __9____513995(.DIN1 (_____9__28488), .DIN2 (___9_9__25996), .Q
       (___09____40683));
  and2s1 __9___513996(.DIN1 (________26357), .DIN2 (________27584), .Q
       (___09____40684));
  and2s1 __9___513997(.DIN1 (_____9__26563), .DIN2 (________26366), .Q
       (___09____40685));
  xnr2s1 __9____513998(.DIN1 (_____0__22654), .DIN2 (____9____37088),
       .Q (___09____40686));
  xnr2s1 __9____513999(.DIN1 (_________22014), .DIN2 (________22608),
       .Q (___09____40687));
  xnr2s1 __9____514000(.DIN1 (________22602), .DIN2 (_____9___36907),
       .Q (___09____40688));
  xor2s1 __9____514001(.DIN1 (_________38364), .DIN2 (________22601),
       .Q (___09_9__40689));
  xnr2s1 __9____514002(.DIN1
       (__________________________________________________________________21996),
       .DIN2 (___00____39959), .Q (___09_0__40690));
  and2s1 __9____514003(.DIN1 (___09____40691), .DIN2 (___9_____39515),
       .Q (___09____40692));
  xor2s1 __9____514004(.DIN1 (___0_____40323), .DIN2 (___0_____40324),
       .Q (___09____40691));
  nor2s1 __9____514005(.DIN1 (___09____40693), .DIN2 (___9_____39445),
       .Q (___09____40694));
  xnr2s1 __9___514006(.DIN1 (___0_____40308), .DIN2 (___0_____40307),
       .Q (___09____40693));
  and2s1 __9___514007(.DIN1 (___09____40695), .DIN2 (___0_____40219),
       .Q (___09____40696));
  nor2s1 __9____514008(.DIN1 (___0__9__40098), .DIN2 (___9__0__39561),
       .Q (___09____40695));
  or2s1 __9____514009(.DIN1 (___09____40697), .DIN2 (___9__0__39643),
       .Q (___09____40698));
  nor2s1 __9____514010(.DIN1 (___9_____39665), .DIN2 (___0_____40205),
       .Q (___09____40697));
  and2s1 __9____514011(.DIN1 (___09_9__40699), .DIN2 (_____0___38427),
       .Q (___09_0__40700));
  nnd2s1 __9____514012(.DIN1 (___0_____40163), .DIN2 (_________38450),
       .Q (___09_9__40699));
  or2s1 __9____514013(.DIN1 (___09____40701), .DIN2 (___0_____40026),
       .Q (___09____40702));
  nnd2s1 __9____514014(.DIN1 (___0_9___40070), .DIN2 (______0__22027),
       .Q (___09____40701));
  or2s1 __9____514015(.DIN1 (___09____40703), .DIN2 (___99____39843),
       .Q (___09____40704));
  xnr2s1 __9___514016(.DIN1 (___00____39929), .DIN2 (___00____39928),
       .Q (___09____40703));
  or2s1 __9___514017(.DIN1 (___09____40705), .DIN2 (___9_____39769), .Q
       (___09____40706));
  xnr2s1 __9____514018(.DIN1 (___99_9__39836), .DIN2 (___99_0__39837),
       .Q (___09____40705));
  or2s1 __9____514019(.DIN1 (___09____40707), .DIN2 (___9_____39545),
       .Q (___09____40708));
  nor2s1 __9____514020(.DIN1 (___9_____39564), .DIN2 (___9_____39762),
       .Q (___09____40707));
  and2s1 __9____514021(.DIN1 (___09_9__40709), .DIN2 (___9_____39138),
       .Q (___0990__40710));
  xor2s1 __9____514022(.DIN1 (___9_____39688), .DIN2 (___9__0__39687),
       .Q (___09_9__40709));
  and2s1 __9____514023(.DIN1 (___099___40711), .DIN2 (___9__0__39536),
       .Q (___099___40712));
  xor2s1 __9____514024(.DIN1 (___9_0___39624), .DIN2 (___9_09__39625),
       .Q (___099___40711));
  and2s1 __9____514025(.DIN1 (___099___40713), .DIN2 (___9_____39090),
       .Q (___099___40714));
  xor2s1 __9___514026(.DIN1 (___9_0___39619), .DIN2 (___9_0___39620),
       .Q (___099___40713));
  or2s1 __9__514027(.DIN1 (___099___40715), .DIN2 (___9_____39486), .Q
       (___099___40716));
  xnr2s1 __9__9_514028(.DIN1 (___9_____39554), .DIN2 (___9__0__39553),
       .Q (___099___40715));
  or2s1 __9__9_514029(.DIN1 (___099___40717), .DIN2
       (__________________________________________________________________22004),
       .Q (___099___40718));
  xnr2s1 __9__9_514030(.DIN1 (_________38733), .DIN2 (___9_0___39619),
       .Q (___099___40717));
  and2s1 __9__9_514031(.DIN1 (___0999__40719), .DIN2 (___9_0___39350),
       .Q (____000__40720));
  xor2s1 __9__9_514032(.DIN1 (___9_____39384), .DIN2 (___9_____39385),
       .Q (___0999__40719));
  or2s1 __9__9_514033(.DIN1 (____00___40721), .DIN2 (___9_____39137),
       .Q (____00___40722));
  xnr2s1 __9__9_514034(.DIN1 (___9_____39301), .DIN2 (___9_____39302),
       .Q (____00___40721));
  or2s1 __9__9_514035(.DIN1 (____00___40723), .DIN2 (___9_9___39156),
       .Q (____00___40724));
  xnr2s1 __9__514036(.DIN1 (_____9___41303), .DIN2 (___9_9___39249), .Q
       (____00___40723));
  and2s1 __9__514037(.DIN1 (____00___40725), .DIN2 (___9_____39150), .Q
       (____00___40726));
  xor2s1 __9__0_514038(.DIN1 (___9_____39231), .DIN2 (___9_____39229),
       .Q (____00___40725));
  or2s1 __9__0_514039(.DIN1 (____00___40727), .DIN2 (_________38442),
       .Q (____00___40728));
  xnr2s1 __9__0_514040(.DIN1 (___9_____39206), .DIN2 (___9_____39205),
       .Q (____00___40727));
  and2s1 __9__0_514041(.DIN1 (____009__40729), .DIN2 (___9_____39095),
       .Q (____0_0__40730));
  xor2s1 __9__0_514042(.DIN1 (___9_____39123), .DIN2 (___9_____39122),
       .Q (____009__40729));
  and2s1 __9__0_514043(.DIN1 (____0____40731), .DIN2 (____9____38958),
       .Q (____0____40732));
  xor2s1 __9__0_514044(.DIN1 (___90____39055), .DIN2 (___90____39056),
       .Q (____0____40731));
  or2s1 __9__0_514045(.DIN1 (____0____40733), .DIN2 (____99___38970),
       .Q (____0____40734));
  xnr2s1 __9__514046(.DIN1 (___90____39001), .DIN2 (___90____39002), .Q
       (____0____40733));
  and2s1 __9___514047(.DIN1 (____0____40735), .DIN2 (____9____38907),
       .Q (____0____40736));
  xor2s1 __9____514048(.DIN1 (____9_9__38931), .DIN2 (____9____38930),
       .Q (____0____40735));
  and2s1 __9____514049(.DIN1 (____0____40737), .DIN2 (_________38829),
       .Q (____0____40738));
  xor2s1 __9____514050(.DIN1 (_________38876), .DIN2 (_________38877),
       .Q (____0____40737));
  or2s1 __9____514051(.DIN1 (____0_9__40739), .DIN2 (_________38763),
       .Q (____0_0__40740));
  xnr2s1 __9____514052(.DIN1 (_________38871), .DIN2 (_________38872),
       .Q (____0_9__40739));
  or2s1 __9____514053(.DIN1 (____0____40741), .DIN2 (______9__38720),
       .Q (____0____40742));
  xnr2s1 __9____514054(.DIN1 (_________38842), .DIN2 (_________38841),
       .Q (____0____40741));
  or2s1 __9____514055(.DIN1 (____0____40743), .DIN2 (_____9___38696),
       .Q (____0____40744));
  xnr2s1 __9___514056(.DIN1 (_________38842), .DIN2 (_________38822),
       .Q (____0____40743));
  or2s1 __9___514057(.DIN1 (____0____40745), .DIN2 (____9___25949), .Q
       (____0____40746));
  nnd2s1 __9____514058(.DIN1 (_________38435), .DIN2 (__________22060),
       .Q (____0____40745));
  and2s1 __9____514059(.DIN1 (____0____40747), .DIN2 (___0____26098),
       .Q (____0____40748));
  nor2s1 __9____514060(.DIN1 (______0__22035), .DIN2 (_________38649),
       .Q (____0____40747));
  or2s1 __9____514061(.DIN1 (____0_9__40749), .DIN2 (_________38300),
       .Q (____0_0__40750));
  xnr2s1 __9____514062(.DIN1 (_____0___38422), .DIN2 (_________38337),
       .Q (____0_9__40749));
  and2s1 __9____514063(.DIN1 (____0____40751), .DIN2 (____0____38068),
       .Q (____0____40752));
  xor2s1 __9____514064(.DIN1 (_________38214), .DIN2 (_________38168),
       .Q (____0____40751));
  and2s1 __9____514065(.DIN1 (____0____40753), .DIN2 (_________37925),
       .Q (____0____40754));
  xor2s1 __9___514066(.DIN1 (____9____38007), .DIN2 (____9____37999),
       .Q (____0____40753));
  or2s1 __9___514067(.DIN1 (____0____40755), .DIN2 (____9____37997), .Q
       (____0____40756));
  nor2s1 __9____514068(.DIN1 (____9_0__38019), .DIN2 (____0____38053),
       .Q (____0____40755));
  or2s1 __9____514069(.DIN1 (____0____40757), .DIN2 (____009__38047),
       .Q (____0____40758));
  nnd2s1 __9____514070(.DIN1
       (____________________________________________21846), .DIN2
       (___0_0___40465), .Q (____0____40757));
  or2s1 __9____514071(.DIN1 (____0_9__40759), .DIN2 (_________37338),
       .Q (____0_0__40760));
  nnd2s1 __9____514072(.DIN1 (____90___37952), .DIN2 (_____0___34938),
       .Q (____0_9__40759));
  and2s1 __9____514073(.DIN1 (____0____40761), .DIN2 (______0__37863),
       .Q (____0____40762));
  nnd2s1 __9____514074(.DIN1
       (_____________________________________________21802), .DIN2
       (_________37748), .Q (____0____40761));
  and2s1 __9____514075(.DIN1 (____0____40763), .DIN2 (_________37639),
       .Q (____0____40764));
  xor2s1 __9___514076(.DIN1 (___9_0___39705), .DIN2 (_____0___37762),
       .Q (____0____40763));
  and2s1 __9___514077(.DIN1 (____0____40765), .DIN2 (_____0___36915),
       .Q (____0____40766));
  nor2s1 __9____514078(.DIN1 (___0__9__40098), .DIN2 (_________37356),
       .Q (____0____40765));
  and2s1 __9____514079(.DIN1 (____0____40767), .DIN2 (____9____37075),
       .Q (____0____40768));
  xor2s1 __9____514080(.DIN1 (____9____38948), .DIN2 (____0____37157),
       .Q (____0____40767));
  or2s1 __9____514081(.DIN1 (____0_9__40769), .DIN2 (____0____40776),
       .Q (____0_0__40770));
  nnd2s1 __9____514082(.DIN1 (______9__37353), .DIN2 (_________35430),
       .Q (____0_9__40769));
  and2s1 __9____514083(.DIN1 (____0____40771), .DIN2 (____0____36253),
       .Q (____0____40772));
  xor2s1 __9____514084(.DIN1 (_________41252), .DIN2 (____0____37149),
       .Q (____0____40771));
  and2s1 __9____514085(.DIN1 (____0____40773), .DIN2 (_________36954),
       .Q (____0____40774));
  xor2s1 __9___514086(.DIN1 (____0____37113), .DIN2 (____0____37114),
       .Q (____0____40773));
  and2s1 __9___514087(.DIN1 (____0____40775), .DIN2 (____0_0__35350),
       .Q (____0____40776));
  xor2s1 __9____514088(.DIN1 (___90____39008), .DIN2 (____9____37059),
       .Q (____0____40775));
  or2s1 __9____514089(.DIN1 (____0____40777), .DIN2 (_________36863),
       .Q (____0____40778));
  nor2s1 __9____514090(.DIN1 (_________36884), .DIN2 (____9____37016),
       .Q (____0____40777));
  and2s1 __9____514091(.DIN1 (____0_9__40779), .DIN2 (_________36880),
       .Q (____0_0__40780));
  xor2s1 __9____514092(.DIN1 (_________36973), .DIN2 (_________36972),
       .Q (____0_9__40779));
  and2s1 __9____514093(.DIN1 (____0____40781), .DIN2 (______9__36783),
       .Q (____0____40782));
  xor2s1 __9____514094(.DIN1 (_________36928), .DIN2 (_________36929),
       .Q (____0____40781));
  and2s1 __9____514095(.DIN1 (____0____40783), .DIN2 (______0__36707),
       .Q (____0____40784));
  xor2s1 __9___514096(.DIN1 (_________38876), .DIN2 (_________36895),
       .Q (____0____40783));
  and2s1 __9___514097(.DIN1 (____0____40785), .DIN2 (______0__36842),
       .Q (____0____40786));
  nnd2s1 __9____514098(.DIN1 (___09____40674), .DIN2 (___0_____40485),
       .Q (____0____40785));
  and2s1 __9____514099(.DIN1 (____0____40787), .DIN2 (_________34547),
       .Q (____0____40788));
  xor2s1 __9____514100(.DIN1 (_________38680), .DIN2 (_________36674),
       .Q (____0____40787));
  and2s1 __9____514101(.DIN1 (____0_9__40789), .DIN2 (_________35074),
       .Q (____0_0__40790));
  xor2s1 __9____514102(.DIN1 (______0__36598), .DIN2 (______9__36597),
       .Q (____0_9__40789));
  or2s1 __9____514103(.DIN1 (____0____40791), .DIN2 (____09___34473),
       .Q (____0____40792));
  xnr2s1 __9____514104(.DIN1 (______0__37673), .DIN2 (_________36599),
       .Q (____0____40791));
  or2s1 __9____514105(.DIN1 (____0____40793), .DIN2
       (_____________________________________________21781), .Q
       (____0____40794));
  and2s1 __9___514106(.DIN1 (____0_0__36258), .DIN2 (____0____36194),
       .Q (____0____40793));
  and2s1 __9___514107(.DIN1 (____0____40795), .DIN2 (_____0___36369),
       .Q (____0____40796));
  xor2s1 __9____514108(.DIN1 (_________36512), .DIN2 (_________36511),
       .Q (____0____40795));
  or2s1 __9____514109(.DIN1 (____0____40797), .DIN2 (_________36468),
       .Q (____0____40798));
  xnr2s1 __9____514110(.DIN1 (_________41341), .DIN2 (_________36496),
       .Q (____0____40797));
  or2s1 __9____514111(.DIN1 (____0_9__40799), .DIN2 (____0_9__34413),
       .Q (____0_0__40800));
  xnr2s1 __9____514112(.DIN1 (_________36480), .DIN2 (_________36479),
       .Q (____0_9__40799));
  or2s1 __9____514113(.DIN1 (____0____40801), .DIN2 (______9__35992),
       .Q (____0____40802));
  xnr2s1 __9____514114(.DIN1 (_____99__37662), .DIN2 (_________36408),
       .Q (____0____40801));
  or2s1 __9____514115(.DIN1 (____0____40803), .DIN2 (_____9___34924),
       .Q (____0____40804));
  xnr2s1 __9___514116(.DIN1 (______0__36697), .DIN2 (_________36409),
       .Q (____0____40803));
  or2s1 __9___514117(.DIN1 (____0____40805), .DIN2 (______0__35509), .Q
       (____0____40806));
  xnr2s1 __9____514118(.DIN1 (____9___23594), .DIN2 (_________36307),
       .Q (____0____40805));
  or2s1 __9____514119(.DIN1 (____0____40807), .DIN2 (____09___36269),
       .Q (____0____40808));
  xnr2s1 __9____514120(.DIN1 (_________36301), .DIN2 (_________36300),
       .Q (____0____40807));
  and2s1 __9____514121(.DIN1 (____0_9__40809), .DIN2 (____0____36205),
       .Q (____090__40810));
  xor2s1 __9____514122(.DIN1 (_________36291), .DIN2 (_____0___36282),
       .Q (____0_9__40809));
  and2s1 __9____514123(.DIN1 (____09___40811), .DIN2 (______9__35852),
       .Q (____09___40812));
  xor2s1 __9____514124(.DIN1 (___________________), .DIN2
       (____9____36158), .Q (____09___40811));
  or2s1 __9____514125(.DIN1 (____09___40813), .DIN2 (______9__34133),
       .Q (____09___40814));
  xnr2s1 __9___514126(.DIN1 (____9___23594), .DIN2 (____9____36120), .Q
       (____09___40813));
  and2s1 __9__514127(.DIN1 (____09___40815), .DIN2 (_____0___36014), .Q
       (____09___40816));
  xor2s1 __9__9_514128(.DIN1 (_________38680), .DIN2 (_________36074),
       .Q (____09___40815));
  or2s1 __9__9_514129(.DIN1 (____09___40817), .DIN2 (_________36030),
       .Q (____09___40818));
  xnr2s1 __9__9_514130(.DIN1 (_________36087), .DIN2 (_________36086),
       .Q (____09___40817));
  and2s1 __9__9_514131(.DIN1 (____099__40819), .DIN2 (_____9___35650),
       .Q (_____00__40820));
  nor2s1 __9__9_514132(.DIN1 (_____9___36094), .DIN2 (_____9___36095),
       .Q (____099__40819));
  and2s1 __9__9_514133(.DIN1 (_____0___40821), .DIN2 (_________36046),
       .Q (_____0___40822));
  xor2s1 __9__9_514134(.DIN1 (_________37547), .DIN2 (_________36063),
       .Q (_____0___40821));
  or2s1 __9__9_514135(.DIN1 (_____0___40823), .DIN2 (_________35672),
       .Q (_____0___40824));
  xnr2s1 __9__514136(.DIN1 (___0__9__40158), .DIN2 (_____00__36010), .Q
       (_____0___40823));
  or2s1 __9__514137(.DIN1 (_____0___40825), .DIN2 (_________35705), .Q
       (_____0___40826));
  or2s1 __9__0_514138(.DIN1 (_____9___36006), .DIN2 (______9__35764),
       .Q (_____0___40825));
  or2s1 __9__0_514139(.DIN1 (_____0___40827), .DIN2 (_________35911),
       .Q (_____0___40828));
  xnr2s1 __9__0_514140(.DIN1 (_________36871), .DIN2 (______0__35942),
       .Q (_____0___40827));
  and2s1 __9__0_514141(.DIN1 (_____09__40829), .DIN2 (_____9___34566),
       .Q (______0__40830));
  xor2s1 __9__0_514142(.DIN1 (_____9___35917), .DIN2 (_____9___35918),
       .Q (_____09__40829));
  and2s1 __9__0_514143(.DIN1 (_________40831), .DIN2 (_________33670),
       .Q (_________40832));
  xor2s1 __9__0_514144(.DIN1 (_________38876), .DIN2 (_________35894),
       .Q (_________40831));
  and2s1 __9__0_514145(.DIN1 (_________40833), .DIN2 (_________35797),
       .Q (_________40834));
  xor2s1 __9__514146(.DIN1 (_________38680), .DIN2 (_________35878), .Q
       (_________40833));
  or2s1 __9___514147(.DIN1 (_________40835), .DIN2 (_____9___33809), .Q
       (_________40836));
  xnr2s1 __9____514148(.DIN1 (_________35867), .DIN2 (_________35868),
       .Q (_________40835));
  and2s1 __9____514149(.DIN1 (_________40837), .DIN2 (____00__28471),
       .Q (_________40838));
  nor2s1 __9____514150(.DIN1 (_________35943), .DIN2 (___0_____40626),
       .Q (_________40837));
  or2s1 __9____514151(.DIN1 (______9__40839), .DIN2 (_____9___34564),
       .Q (______0__40840));
  xnr2s1 __9____514152(.DIN1 (_____0___35660), .DIN2 (_____0___35659),
       .Q (______9__40839));
  and2s1 __9____514153(.DIN1 (_________40841), .DIN2 (_________35487),
       .Q (_________40842));
  xor2s1 __9____514154(.DIN1 (_________37452), .DIN2 (_________35639),
       .Q (_________40841));
  and2s1 __9____514155(.DIN1 (_________40843), .DIN2 (_____0___34195),
       .Q (_________40844));
  xor2s1 __9___514156(.DIN1 (_________35622), .DIN2 (_________35623),
       .Q (_________40843));
  and2s1 __9___514157(.DIN1 (_________40845), .DIN2 (______0__35545),
       .Q (_________40846));
  xor2s1 __9____514158(.DIN1 (_________38301), .DIN2 (_________35616),
       .Q (_________40845));
  or2s1 __9____514159(.DIN1 (_________40847), .DIN2 (_________35635),
       .Q (_________40848));
  and2s1 __9____514160(.DIN1 (_________35661), .DIN2 (_________37789),
       .Q (_________40847));
  or2s1 __9____514161(.DIN1 (______9__40849), .DIN2 (_____0___35385),
       .Q (______0__40850));
  xnr2s1 __9____514162(.DIN1 (_________35526), .DIN2 (_________35525),
       .Q (______9__40849));
  or2s1 __9____514163(.DIN1 (_________40851), .DIN2 (____0____35327),
       .Q (_________40852));
  nnd2s1 __9____514164(.DIN1 (_________35392), .DIN2 (inData[28]), .Q
       (_________40851));
  and2s1 __9____514165(.DIN1 (_________40853), .DIN2 (____0_0__35298),
       .Q (_________40854));
  xor2s1 __9___514166(.DIN1 (___9_0___39705), .DIN2 (_____0___35384),
       .Q (_________40853));
  or2s1 __9___514167(.DIN1 (_________40855), .DIN2 (___0____22313), .Q
       (_________40856));
  nnd2s1 __9____514168(.DIN1 (___0_____40477), .DIN2 (______0__35537),
       .Q (_________40855));
  and2s1 __9____514169(.DIN1 (_________40857), .DIN2 (_________34770),
       .Q (_________40858));
  xor2s1 __9____514170(.DIN1 (_________41252), .DIN2 (____0____35301),
       .Q (_________40857));
  or2s1 __9____514171(.DIN1 (______9__40859), .DIN2 (____9____34312),
       .Q (______0__40860));
  xnr2s1 __9____514172(.DIN1 (_________35806), .DIN2 (____9____35229),
       .Q (______9__40859));
  nor2s1 __9____514173(.DIN1 (_________40861), .DIN2 (_________35120),
       .Q (_________40862));
  xnr2s1 __9____514174(.DIN1 (_________35968), .DIN2 (____9____35231),
       .Q (_________40861));
  or2s1 __9____514175(.DIN1 (_________40863), .DIN2 (_____9___34183),
       .Q (_________40864));
  xnr2s1 __9___514176(.DIN1 (_________36349), .DIN2 (____9____35212),
       .Q (_________40863));
  or2s1 __9___514177(.DIN1 (_________40865), .DIN2 (______0__35024), .Q
       (_________40866));
  xnr2s1 __9____514178(.DIN1 (____9____38909), .DIN2 (_____9___35097),
       .Q (_________40865));
  or2s1 __9____514179(.DIN1 (_________40867), .DIN2 (______0__35059),
       .Q (_________40868));
  nor2s1 __9____514180(.DIN1
       (_______________________________________________________________________________________),
       .DIN2 (_________35031), .Q (_________40867));
  or2s1 __9____514181(.DIN1 (_________40869), .DIN2 (_________33788),
       .Q (_________40870));
  xnr2s1 __9____514182(.DIN1 (_____00__35736), .DIN2 (_________34979),
       .Q (_________40869));
  or2s1 __9___514183(.DIN1 (_________40871), .DIN2 (____9____32453), .Q
       (_________40872));
  xnr2s1 __9____514184(.DIN1 (___00____39929), .DIN2 (_________34918),
       .Q (_________40871));
  or2s1 __9____514185(.DIN1 (_________40873), .DIN2 (_________34590),
       .Q (_________40874));
  xnr2s1 __9____514186(.DIN1 (_________37614), .DIN2 (_________34899),
       .Q (_________40873));
  or2s1 __9____514187(.DIN1 (_________40875), .DIN2 (_________34767),
       .Q (_________40876));
  xnr2s1 __9____514188(.DIN1 (___9_____39542), .DIN2 (_____0___34849),
       .Q (_________40875));
  or2s1 __9____514189(.DIN1 (_________40877), .DIN2 (_________34066),
       .Q (_________40878));
  xnr2s1 __9___514190(.DIN1 (___90____39001), .DIN2 (______0__34819),
       .Q (_________40877));
  or2s1 __9___514191(.DIN1 (_________40879), .DIN2 (_____0___33067), .Q
       (_________40880));
  xnr2s1 __9____514192(.DIN1 (_________34775), .DIN2 (_________34776),
       .Q (_________40879));
  and2s1 __9____514193(.DIN1 (_________40881), .DIN2 (________26346),
       .Q (_________40882));
  nor2s1 __9____514194(.DIN1 (_____9___34650), .DIN2 (________25903),
       .Q (_________40881));
  and2s1 __9____514195(.DIN1 (______9__40883), .DIN2 (_________33762),
       .Q (______0__40884));
  xor2s1 __9____514196(.DIN1 (_________35084), .DIN2 (_____0___34573),
       .Q (______9__40883));
  and2s1 __9____514197(.DIN1 (_________40885), .DIN2 (____0____33507),
       .Q (_________40886));
  xor2s1 __9____514198(.DIN1 (______9__34553), .DIN2 (_________34647),
       .Q (_________40885));
  and2s1 __9____514199(.DIN1 (_________40887), .DIN2 (____0____31538),
       .Q (_________40888));
  xor2s1 __9___514200(.DIN1 (______0__34517), .DIN2 (______9__34516),
       .Q (_________40887));
  and2s1 __9___514201(.DIN1 (_________40889), .DIN2 (____9____32455),
       .Q (_________40890));
  xor2s1 __9____514202(.DIN1 (_________35523), .DIN2 (_________34512),
       .Q (_________40889));
  and2s1 __9____514203(.DIN1 (_________40891), .DIN2 (______9__34276),
       .Q (_________40892));
  xor2s1 __9____514204(.DIN1 (_________38395), .DIN2 (____0____34422),
       .Q (_________40891));
  or2s1 __9____514205(.DIN1 (______9__40893), .DIN2 (____90___34288),
       .Q (______0__40894));
  xnr2s1 __9____514206(.DIN1 (_____09__35744), .DIN2 (____0____34404),
       .Q (______9__40893));
  and2s1 __9____514207(.DIN1 (_________40895), .DIN2 (___0__9__31167),
       .Q (_________40896));
  nor2s1 __9____514208(.DIN1 (___0_____30937), .DIN2 (_________34156),
       .Q (_________40895));
  and2s1 __9____514209(.DIN1 (_________40897), .DIN2 (_____0___34007),
       .Q (_________40898));
  xor2s1 __9___514210(.DIN1 (_________35523), .DIN2 (______0__34117),
       .Q (_________40897));
  and2s1 __9___514211(.DIN1 (_________40899), .DIN2 (_________34126),
       .Q (_________40900));
  nnd2s1 __9____514212(.DIN1 (______9__34143), .DIN2
       (____________________________________________21791), .Q
       (_________40899));
  or2s1 __9____514213(.DIN1 (_________40901), .DIN2 (____0____32511),
       .Q (_________40902));
  xnr2s1 __9____514214(.DIN1 (____90___36104), .DIN2 (_____0___34005),
       .Q (_________40901));
  or2s1 __9____514215(.DIN1 (______9__40903), .DIN2 (______0__33649),
       .Q (_____90__40904));
  xnr2s1 __9____514216(.DIN1 (_________38200), .DIN2 (_____0___33916),
       .Q (______9__40903));
  and2s1 __9____514217(.DIN1 (_____9___40905), .DIN2 (_________33853),
       .Q (_____9___40906));
  nor2s1 __9____514218(.DIN1 (___09____31451), .DIN2 (___999__29637),
       .Q (_____9___40905));
  or2s1 __9____514219(.DIN1 (_____9___40907), .DIN2 (________26810), .Q
       (_____9___40908));
  nnd2s1 __9___514220(.DIN1 (_________33853), .DIN2 (________27168), .Q
       (_____9___40907));
  or2s1 __9__514221(.DIN1 (_____9___40909), .DIN2 (____0____33505), .Q
       (_____9___40910));
  xnr2s1 __9__9_514222(.DIN1 (_________33702), .DIN2 (_________35968),
       .Q (_____9___40909));
  or2s1 __9__9_514223(.DIN1 (_____9___40911), .DIN2 (____09___32570),
       .Q (_____9___40912));
  nor2s1 __9__9_514224(.DIN1 (_________32617), .DIN2 (_____0___33624),
       .Q (_____9___40911));
  or2s1 __9__9_514225(.DIN1 (_____99__40913), .DIN2 (____0_0__33500),
       .Q (_____00__40914));
  nnd2s1 __9__9_514226(.DIN1 (___09___27916), .DIN2 (___0____26106), .Q
       (_____99__40913));
  or2s1 __9__9_514227(.DIN1 (_____0___40915), .DIN2 (____0____33503),
       .Q (_____0___40916));
  nnd2s1 __9__9_514228(.DIN1 (__99_0__30469), .DIN2 (_____0__26276), .Q
       (_____0___40915));
  or2s1 __9__9_514229(.DIN1 (_____0___40917), .DIN2 (___00_9__30583),
       .Q (_____0___40918));
  nnd2s1 __9__514230(.DIN1 (____0____33501), .DIN2 (________24907), .Q
       (_____0___40917));
  and2s1 __9__514231(.DIN1 (_____0___40919), .DIN2 (_____0___40922), .Q
       (_____0___40920));
  nor2s1 __9__0_514232(.DIN1 (_____9__27204), .DIN2 (__9__9__30073), .Q
       (_____0___40919));
  and2s1 __9__0_514233(.DIN1 (_____0___40921), .DIN2 (___0__9__30898),
       .Q (_____0___40922));
  nor2s1 __9__0_514234(.DIN1 (____00___33440), .DIN2 (___099___31499),
       .Q (_____0___40921));
  and2s1 __9__0_514235(.DIN1 (_____09__40923), .DIN2 (_________33215),
       .Q (______0__40924));
  xor2s1 __9__0_514236(.DIN1 (___________________), .DIN2
       (_________33279), .Q (_____09__40923));
  or2s1 __9__0_514237(.DIN1 (_________40925), .DIN2 (_____0___33251),
       .Q (_________40926));
  nnd2s1 __9__0_514238(.DIN1 (__9__0__29832), .DIN2 (____9___29365), .Q
       (_________40925));
  and2s1 __9__0_514239(.DIN1 (_________40927), .DIN2 (________26260),
       .Q (_________40928));
  xor2s1 __9__514240(.DIN1 (_____90__33241), .DIN2 (______9__33240), .Q
       (_________40927));
  or2s1 __9___514241(.DIN1 (_________40929), .DIN2 (_________31856), .Q
       (_________40930));
  nnd2s1 __9____514242(.DIN1 (_________33136), .DIN2 (_____9__28626),
       .Q (_________40929));
  and2s1 __9____514243(.DIN1 (_________40931), .DIN2 (________27708),
       .Q (_________40932));
  xor2s1 __9____514244(.DIN1 (_________36527), .DIN2 (_____99__33065),
       .Q (_________40931));
  and2s1 __9____514245(.DIN1 (______9__40933), .DIN2 (_________32985),
       .Q (______0__40934));
  xor2s1 __9____514246(.DIN1 (______9__34088), .DIN2 (_________33044),
       .Q (______9__40933));
  and2s1 __9____514247(.DIN1 (_________40935), .DIN2 (_____9___32279),
       .Q (_________40936));
  xor2s1 __9____514248(.DIN1 (___90____39055), .DIN2 (______9__32921),
       .Q (_________40935));
  and2s1 __9____514249(.DIN1 (_________40937), .DIN2 (_________32604),
       .Q (_________40938));
  nor2s1 __9___514250(.DIN1 (________29293), .DIN2 (_____9___32771), .Q
       (_________40937));
  or2s1 __9___514251(.DIN1 (_________40939), .DIN2 (_________32025), .Q
       (_________40940));
  xnr2s1 __9____514252(.DIN1 (_________33924), .DIN2 (_________32314),
       .Q (_________40939));
  nor2s1 __9____514253(.DIN1 (_________40941), .DIN2 (_____0___31707),
       .Q (_________40942));
  nnd2s1 __9____514254(.DIN1 (________29341), .DIN2 (________26809), .Q
       (_________40941));
  or2s1 __9____514255(.DIN1 (______9__40943), .DIN2 (________28526), .Q
       (______0__40944));
  nnd2s1 __9____514256(.DIN1 (_________31687), .DIN2 (________28889),
       .Q (______9__40943));
  and2s1 __9____514257(.DIN1 (_________40945), .DIN2 (___0_____31385),
       .Q (_________40946));
  and2s1 __9____514258(.DIN1 (_________32140), .DIN2 (____0____31534),
       .Q (_________40945));
  nor2s1 __9___514259(.DIN1 (___9____28675), .DIN2 (______0__40953), .Q
       (_________40947));
  and2s1 __9___514260(.DIN1 (_________40948), .DIN2 (___0_____31038),
       .Q (_________40949));
  or2s1 __9____514261(.DIN1 (_____9___33157), .DIN2 (___0_0___31220),
       .Q (_________40948));
  nnd2s1 __9____514262(.DIN1 (_________40950), .DIN2 (___0_____30781),
       .Q (_________40951));
  nor2s1 __9____514263(.DIN1 (__9__0__30394), .DIN2 (___0_____31282),
       .Q (_________40950));
  or2s1 __9____514264(.DIN1 (______9__40952), .DIN2 (_________31870),
       .Q (______0__40953));
  or2s1 __9____514265(.DIN1 (___099___31496), .DIN2 (___0_____30767),
       .Q (______9__40952));
  and2s1 __9____514266(.DIN1 (_________40954), .DIN2 (_________40979),
       .Q (_________40955));
  nor2s1 __9____514267(.DIN1 (________28077), .DIN2 (__9__0__29824), .Q
       (_________40954));
  nnd2s1 __9____514268(.DIN1 (_________40956), .DIN2 (__99____30486),
       .Q (_________40957));
  nor2s1 __9___514269(.DIN1 (________26333), .DIN2 (___0_____31345), .Q
       (_________40956));
  and2s1 __9___514270(.DIN1 (_________40958), .DIN2 (___0__0__30796),
       .Q (_________40959));
  nor2s1 __9____514271(.DIN1 (________29025), .DIN2 (__9_____30428), .Q
       (_________40958));
  and2s1 __9____514272(.DIN1 (_________40960), .DIN2 (__90____29675),
       .Q (_________40961));
  nor2s1 __9____514273(.DIN1 (__9_____29855), .DIN2 (__9_____30232), .Q
       (_________40960));
  and2s1 __9____514274(.DIN1 (______9__40962), .DIN2 (__9_____30068),
       .Q (______0__40963));
  nor2s1 __9____514275(.DIN1 (__990___30461), .DIN2 (__9__0__30438), .Q
       (______9__40962));
  nor2s1 __9____514276(.DIN1 (_________40964), .DIN2 (___9____28667),
       .Q (_________40965));
  nnd2s1 __9____514277(.DIN1 (___0_____30803), .DIN2 (____0___27302),
       .Q (_________40964));
  and2s1 __9____514278(.DIN1 (_________40966), .DIN2 (__9_____30117),
       .Q (_________40967));
  nor2s1 __9___514279(.DIN1 (__9_____29745), .DIN2 (__9_____30441), .Q
       (_________40966));
  nor2s1 __9___514280(.DIN1 (_________40968), .DIN2 (__9_____30036), .Q
       (_________40969));
  nnd2s1 __9____514281(.DIN1 (___0_____31173), .DIN2 (____9___29367),
       .Q (_________40968));
  or2s1 __9____514282(.DIN1 (_________40970), .DIN2 (__9_____29884), .Q
       (_________40971));
  nnd2s1 __9____514283(.DIN1 (________27712), .DIN2 (________28169), .Q
       (_________40970));
  or2s1 __9____514284(.DIN1 (______9__40972), .DIN2 (__9_____29844), .Q
       (______0__40973));
  nnd2s1 __9____514285(.DIN1 (________29395), .DIN2 (________29389), .Q
       (______9__40972));
  or2s1 __9____514286(.DIN1 (_________40974), .DIN2 (_________36618),
       .Q (_________40975));
  nnd2s1 __9____514287(.DIN1 (inData[30]), .DIN2
       (_____________________________________________21808), .Q
       (_________40974));
  and2s1 __9____514288(.DIN1 (_________40976), .DIN2 (________28139),
       .Q (_________40977));
  xor2s1 __9___514289(.DIN1 (__9_____29971), .DIN2 (__9_____29970), .Q
       (_________40976));
  and2s1 __9___514290(.DIN1 (_________40978), .DIN2 (________29391), .Q
       (_________40979));
  nor2s1 __9____514291(.DIN1 (______0__41082), .DIN2 (___9____29578),
       .Q (_________40978));
  and2s1 __9____514292(.DIN1 (_________40980), .DIN2 (___0____27007),
       .Q (_________40981));
  nor2s1 __9____514293(.DIN1 (__9_____30400), .DIN2 (__90____29648), .Q
       (_________40980));
  and2s1 __9____514294(.DIN1 (______9__40982), .DIN2 (________29339),
       .Q (______0__40983));
  nor2s1 __9____514295(.DIN1 (____9___29364), .DIN2 (________28412), .Q
       (______9__40982));
  or2s1 __9____514296(.DIN1 (_________40984), .DIN2 (________29499), .Q
       (_________40985));
  nnd2s1 __9____514297(.DIN1 (____9___28289), .DIN2 (__9__9__30300), .Q
       (_________40984));
  nor2s1 __9___514298(.DIN1 (____9___29092), .DIN2 (____0___29467), .Q
       (_________40986));
  and2s1 __9___514299(.DIN1 (_________40987), .DIN2 (________29494), .Q
       (_________40988));
  nor2s1 __9____514300(.DIN1 (________28160), .DIN2 (__9_9___29892), .Q
       (_________40987));
  or2s1 __9____514301(.DIN1 (_________40989), .DIN2 (__9_____29835), .Q
       (_________40990));
  nnd2s1 __9____514302(.DIN1 (____9___29367), .DIN2 (__9_99__29895), .Q
       (_________40989));
  and2s1 __9____514303(.DIN1 (______9__40991), .DIN2 (__9_____29748),
       .Q (______0__40992));
  nor2s1 __9____514304(.DIN1 (__9_____30109), .DIN2 (________29216), .Q
       (______9__40991));
  or2s1 __9____514305(.DIN1 (_________40993), .DIN2 (___0_____31262),
       .Q (_________40994));
  or2s1 __9____514306(.DIN1 (__9_____29742), .DIN2 (_________41078), .Q
       (_________40993));
  or2s1 __9____514307(.DIN1 (_________40995), .DIN2 (___9____26913), .Q
       (_________40996));
  nnd2s1 __9___514308(.DIN1 (____9___29277), .DIN2 (________25732), .Q
       (_________40995));
  or2s1 __9___514309(.DIN1 (_________40997), .DIN2 (_________41345), .Q
       (_________40998));
  and2s1 __9____514310(.DIN1 (________29162), .DIN2 (inData[22]), .Q
       (_________40997));
  nnd2s1 __9____514311(.DIN1 (_________40999), .DIN2 (_____9__29027),
       .Q (_________41000));
  nor2s1 __9____514312(.DIN1 (________27049), .DIN2 (____0___27482), .Q
       (_________40999));
  nor2s1 __9____514313(.DIN1 (______9__41001), .DIN2 (____0___28292),
       .Q (_____90__41002));
  nnd2s1 __9____514314(.DIN1 (________28877), .DIN2 (__9__9__30056), .Q
       (______9__41001));
  or2s1 __9____514315(.DIN1 (_____9___41003), .DIN2 (___09___26134), .Q
       (_____9___41004));
  nnd2s1 __9____514316(.DIN1 (________28980), .DIN2 (_____0__27978), .Q
       (_____9___41003));
  nnd2s1 __9____514317(.DIN1 (_____9___41005), .DIN2 (_____0__28890),
       .Q (_____9___41006));
  nor2s1 __9___514318(.DIN1 (__9_9___29991), .DIN2 (___9____29573), .Q
       (_____9___41005));
  or2s1 __9__514319(.DIN1 (_____9___41007), .DIN2 (_____0___41112), .Q
       (_____9___41008));
  nnd2s1 __9__9_514320(.DIN1 (___9____29592), .DIN2 (________29523), .Q
       (_____9___41007));
  and2s1 __9__9_514321(.DIN1 (_____9___41009), .DIN2 (________29420),
       .Q (_____9___41010));
  nor2s1 __9__9_514322(.DIN1 (________26353), .DIN2 (________29409), .Q
       (_____9___41009));
  and2s1 __9__9_514323(.DIN1 (_____99__41011), .DIN2 (_____9__27471),
       .Q (_____00__41012));
  or2s1 __9__9_514324(.DIN1 (__9_9___29892), .DIN2 (_____9___41108), .Q
       (_____99__41011));
  or2s1 __9__9_514325(.DIN1 (_____0___41013), .DIN2 (________28588), .Q
       (_____0___41014));
  nnd2s1 __9__9_514326(.DIN1 (__9__9__29859), .DIN2 (____99__27208), .Q
       (_____0___41013));
  or2s1 __9__9_514327(.DIN1 (_____0___41015), .DIN2 (____9___28915), .Q
       (_____0___41016));
  nnd2s1 __9__514328(.DIN1 (________28487), .DIN2 (________29031), .Q
       (_____0___41015));
  nnd2s1 __9__514329(.DIN1 (_____0___41017), .DIN2 (_____0__29227), .Q
       (_____0___41018));
  nor2s1 __9__0_514330(.DIN1 (__9_____29754), .DIN2 (_____9__28492), .Q
       (_____0___41017));
  and2s1 __9__0_514331(.DIN1 (_____0___41019), .DIN2 (________27500),
       .Q (_____0___41020));
  nor2s1 __9__0_514332(.DIN1 (__9_0___29897), .DIN2 (__9__0__29824), .Q
       (_____0___41019));
  and2s1 __9__0_514333(.DIN1 (_____09__41021), .DIN2 (________28491),
       .Q (______0__41022));
  nor2s1 __9__0_514334(.DIN1 (__9_____29750), .DIN2 (________29217), .Q
       (_____09__41021));
  or2s1 __9__0_514335(.DIN1 (_________41023), .DIN2 (___99___27824), .Q
       (_________41024));
  nnd2s1 __9__0_514336(.DIN1 (________28489), .DIN2 (____9___27478), .Q
       (_________41023));
  or2s1 __9__0_514337(.DIN1 (_________41025), .DIN2 (__9_____30071), .Q
       (_________41026));
  nnd2s1 __9__514338(.DIN1 (_________41138), .DIN2 (________29405), .Q
       (_________41025));
  and2s1 __9___514339(.DIN1 (_________41027), .DIN2 (_____0__27610), .Q
       (_________41028));
  nor2s1 __9____514340(.DIN1 (__9_0___29995), .DIN2 (________28490), .Q
       (_________41027));
  or2s1 __9____514341(.DIN1 (_________41029), .DIN2 (________27378), .Q
       (_________41030));
  nnd2s1 __9____514342(.DIN1 (_____9__28546), .DIN2 (_____9__27996), .Q
       (_________41029));
  nor2s1 __9____514343(.DIN1 (______9__41031), .DIN2 (________29229),
       .Q (______0__41032));
  nnd2s1 __9____514344(.DIN1 (____9___28547), .DIN2 (__9_0___29899), .Q
       (______9__41031));
  nor2s1 __9____514345(.DIN1 (_________41033), .DIN2 (______0__41260),
       .Q (_________41034));
  nnd2s1 __9____514346(.DIN1 (_________34136), .DIN2 (___0_____40594),
       .Q (_________41033));
  and2s1 __9____514347(.DIN1 (_________41035), .DIN2 (____9___28375),
       .Q (_________41036));
  nor2s1 __9___514348(.DIN1 (____0___28202), .DIN2 (_____0__27723), .Q
       (_________41035));
  nor2s1 __9___514349(.DIN1 (_________41037), .DIN2 (________28541), .Q
       (_________41038));
  nnd2s1 __9____514350(.DIN1 (____9___28288), .DIN2 (___9____29590), .Q
       (_________41037));
  and2s1 __9____514351(.DIN1 (_________41039), .DIN2 (____9___28372),
       .Q (_________41040));
  nor2s1 __9____514352(.DIN1 (________28187), .DIN2 (____9___29093), .Q
       (_________41039));
  nor2s1 __9____514353(.DIN1 (______9__41041), .DIN2 (___00___28741),
       .Q (______0__41042));
  nnd2s1 __9____514354(.DIN1 (___9____28716), .DIN2 (___900__29553), .Q
       (______9__41041));
  and2s1 __9____514355(.DIN1 (_________41043), .DIN2 (________29056),
       .Q (_________41044));
  nor2s1 __9____514356(.DIN1 (________29268), .DIN2 (___99___27824), .Q
       (_________41043));
  nor2s1 __9____514357(.DIN1 (_________41045), .DIN2 (____00__28291),
       .Q (_________41046));
  nnd2s1 __9___514358(.DIN1 (________29246), .DIN2 (________29533), .Q
       (_________41045));
  nnd2s1 __9___514359(.DIN1 (_________41047), .DIN2 (______0__32108),
       .Q (_________41048));
  nor2s1 __9____514360(.DIN1 (________29531), .DIN2 (_____0__29037), .Q
       (_________41047));
  or2s1 __9____514361(.DIN1 (_________41049), .DIN2 (___0____28757), .Q
       (_________41050));
  nnd2s1 __9____514362(.DIN1 (____9___28290), .DIN2 (________28252), .Q
       (_________41049));
  nor2s1 __9____514363(.DIN1 (______9__41051), .DIN2 (________27165),
       .Q (______0__41052));
  nnd2s1 __9____514364(.DIN1 (____00__28376), .DIN2 (__9_____29843), .Q
       (______9__41051));
  nnd2s1 __9____514365(.DIN1 (_________41053), .DIN2 (_____0__29213),
       .Q (_________41054));
  nor2s1 __9____514366(.DIN1 (_________41273), .DIN2 (____0___28292),
       .Q (_________41053));
  nor2s1 __9____514367(.DIN1 (_________41055), .DIN2 (_____0__28168),
       .Q (_________41056));
  nnd2s1 __9___514368(.DIN1 (________28895), .DIN2 (________29498), .Q
       (_________41055));
  or2s1 __9___514369(.DIN1 (_________41057), .DIN2 (________28991), .Q
       (_________41058));
  nnd2s1 __9____514370(.DIN1 (________28176), .DIN2 (________25834), .Q
       (_________41057));
  nnd2s1 __9____514371(.DIN1 (_________41059), .DIN2 (________28889),
       .Q (_________41060));
  nor2s1 __9____514372(.DIN1 (________29500), .DIN2 (________28179), .Q
       (_________41059));
  and2s1 __9____514373(.DIN1 (______9__41061), .DIN2 (________28982),
       .Q (______0__41062));
  nor2s1 __9____514374(.DIN1 (___0____27868), .DIN2 (________28175), .Q
       (______9__41061));
  nor2s1 __9____514375(.DIN1 (_________41063), .DIN2 (________28936),
       .Q (_________41064));
  nnd2s1 __9____514376(.DIN1 (____0___28297), .DIN2 (____09___31598),
       .Q (_________41063));
  or2s1 __9____514377(.DIN1 (_________41065), .DIN2 (____99__27391), .Q
       (_________41066));
  nnd2s1 __9___514378(.DIN1 (________28300), .DIN2 (________29066), .Q
       (_________41065));
  or2s1 __9___514379(.DIN1 (_________41067), .DIN2 (________28857), .Q
       (_________41068));
  nnd2s1 __9____514380(.DIN1 (_____0__29495), .DIN2 (____0___28020), .Q
       (_________41067));
  or2s1 __9____514381(.DIN1 (_________41069), .DIN2 (________28625), .Q
       (_________41070));
  nnd2s1 __9____514382(.DIN1 (____0___27302), .DIN2 (___00___26956), .Q
       (_________41069));
  or2s1 __9____514383(.DIN1 (______9__41071), .DIN2 (___99___27823), .Q
       (______0__41072));
  nnd2s1 __9____514384(.DIN1 (________28507), .DIN2 (____90__29272), .Q
       (______9__41071));
  and2s1 __9____514385(.DIN1 (_________41073), .DIN2 (________28537),
       .Q (_________41074));
  nor2s1 __9____514386(.DIN1 (__9__0__30394), .DIN2 (____9___28915), .Q
       (_________41073));
  or2s1 __9____514387(.DIN1 (_________41075), .DIN2 (___0____27880), .Q
       (_________41076));
  nnd2s1 __9___514388(.DIN1 (________29223), .DIN2 (___99___27826), .Q
       (_________41075));
  nnd2s1 __9___514389(.DIN1 (_________41077), .DIN2 (___9____27779), .Q
       (_________41078));
  nor2s1 __9____514390(.DIN1 (_____0__28168), .DIN2 (________27615), .Q
       (_________41077));
  and2s1 __9____514391(.DIN1 (_________41079), .DIN2 (________28408),
       .Q (_________41080));
  nor2s1 __9____514392(.DIN1 (_________41176), .DIN2 (___0____28806),
       .Q (_________41079));
  or2s1 __9____514393(.DIN1 (______9__41081), .DIN2 (___9____29573), .Q
       (______0__41082));
  nnd2s1 __9____514394(.DIN1 (_____9___31694), .DIN2 (___0__9__31260),
       .Q (______9__41081));
  nnd2s1 __9____514395(.DIN1 (_________41083), .DIN2 (________27236),
       .Q (_________41084));
  nor2s1 __9____514396(.DIN1 (________29088), .DIN2 (____0___27655), .Q
       (_________41083));
  and2s1 __9____514397(.DIN1 (_________41085), .DIN2 (________27591),
       .Q (_________41086));
  nor2s1 __9___514398(.DIN1 (________29508), .DIN2 (________27592), .Q
       (_________41085));
  and2s1 __9___514399(.DIN1 (_________41087), .DIN2 (________27710), .Q
       (_________41088));
  nor2s1 __9____514400(.DIN1 (________26639), .DIN2 (___0____26096), .Q
       (_________41087));
  or2s1 __9____514401(.DIN1 (_________41089), .DIN2 (_____9__27176), .Q
       (_________41090));
  nnd2s1 __9____514402(.DIN1 (___909__27751), .DIN2 (________28454), .Q
       (_________41089));
  or2s1 __9____514403(.DIN1 (______9__41091), .DIN2 (________28343), .Q
       (______0__41092));
  nnd2s1 __9____514404(.DIN1 (_____0__28966), .DIN2 (________27591), .Q
       (______9__41091));
  or2s1 __9____514405(.DIN1 (_________41093), .DIN2 (____0___28377), .Q
       (_________41094));
  nnd2s1 __9____514406(.DIN1 (________28364), .DIN2 (________28537), .Q
       (_________41093));
  nor2s1 __9____514407(.DIN1 (_________41095), .DIN2 (____0___27122),
       .Q (_________41096));
  nnd2s1 __9___514408(.DIN1 (____0___28926), .DIN2 (___00___26957), .Q
       (_________41095));
  or2s1 __9____514409(.DIN1 (_________41097), .DIN2 (________29217), .Q
       (_________41098));
  nnd2s1 __9____514410(.DIN1 (____00__27654), .DIN2 (________29523), .Q
       (_________41097));
  or2s1 __9____514411(.DIN1 (______9__41099), .DIN2 (____00__27480), .Q
       (_____90__41100));
  nnd2s1 __9____514412(.DIN1 (__90____29657), .DIN2 (________28628), .Q
       (______9__41099));
  nor2s1 __9____514413(.DIN1 (_____9___41101), .DIN2 (________27681),
       .Q (_____9___41102));
  nnd2s1 __9____514414(.DIN1 (________29311), .DIN2 (___9____28722), .Q
       (_____9___41101));
  or2s1 __9____514415(.DIN1 (_____9___41103), .DIN2 (________27951), .Q
       (_____9___41104));
  nnd2s1 __9___514416(.DIN1 (___99___28730), .DIN2 (________26358), .Q
       (_____9___41103));
  or2s1 __9__514417(.DIN1 (_____9___41105), .DIN2 (_____9__27222), .Q
       (_____9___41106));
  nnd2s1 __9__9_514418(.DIN1 (_____9__27996), .DIN2 (____9___29007), .Q
       (_____9___41105));
  or2s1 __9__9_514419(.DIN1 (_____9___41107), .DIN2 (________27341), .Q
       (_____9___41108));
  nnd2s1 __9__9_514420(.DIN1 (_____0__28395), .DIN2 (________27954), .Q
       (_____9___41107));
  and2s1 __9__9_514421(.DIN1 (_____99__41109), .DIN2 (_____9__27075),
       .Q (_____00__41110));
  nor2s1 __9__9_514422(.DIN1 (________27935), .DIN2 (___9_0__28655), .Q
       (_____99__41109));
  or2s1 __9__9_514423(.DIN1 (_____0___41111), .DIN2 (____9_0__33415),
       .Q (_____0___41112));
  nnd2s1 __9__9_514424(.DIN1 (___09___27920), .DIN2 (____0___28109), .Q
       (_____0___41111));
  or2s1 __9__9_514425(.DIN1 (_____0___41113), .DIN2 (___9_9__27813), .Q
       (_____0___41114));
  nnd2s1 __9__514426(.DIN1 (____9___28550), .DIN2 (________29079), .Q
       (_____0___41113));
  or2s1 __9_514427(.DIN1 (_____0___41115), .DIN2 (___0____27880), .Q
       (_____0___41116));
  nnd2s1 __9_90_514428(.DIN1 (____9___28642), .DIN2 (________27440), .Q
       (_____0___41115));
  or2s1 __9_90_514429(.DIN1 (_____0___41117), .DIN2 (_____0__27941), .Q
       (_____0___41118));
  nnd2s1 __9_90_514430(.DIN1 (________28596), .DIN2 (____9___27295), .Q
       (_____0___41117));
  and2s1 __9_90_514431(.DIN1 (_____09__41119), .DIN2 (________28364),
       .Q (______0__41120));
  nor2s1 __9_90_514432(.DIN1 (___0_____30764), .DIN2 (________27547),
       .Q (_____09__41119));
  or2s1 __9_90_514433(.DIN1 (_________41121), .DIN2 (___9____27809), .Q
       (_________41122));
  nnd2s1 __9_90_514434(.DIN1 (________27203), .DIN2 (________28533), .Q
       (_________41121));
  or2s1 __9_90_514435(.DIN1 (_________41123), .DIN2 (________27197), .Q
       (_________41124));
  nnd2s1 __9_514436(.DIN1 (________28519), .DIN2 (_____0__26390), .Q
       (_________41123));
  or2s1 __9_9_514437(.DIN1 (_________41125), .DIN2 (________27504), .Q
       (_________41126));
  nnd2s1 __9_9__514438(.DIN1 (________27156), .DIN2 (___0_99__30832),
       .Q (_________41125));
  or2s1 __9_9__514439(.DIN1 (_________41127), .DIN2 (___0_____30801),
       .Q (_________41128));
  nnd2s1 __9_9__514440(.DIN1 (________27439), .DIN2 (__9_____30058), .Q
       (_________41127));
  and2s1 __9_9__514441(.DIN1 (______9__41129), .DIN2 (________27707),
       .Q (______0__41130));
  nor2s1 __9_9__514442(.DIN1 (________29359), .DIN2 (_____9__27986), .Q
       (______9__41129));
  nnd2s1 __9_9__514443(.DIN1 (_________41131), .DIN2 (___0_99__30926),
       .Q (_________41132));
  nor2s1 __9_9__514444(.DIN1 (________27284), .DIN2 (________28310), .Q
       (_________41131));
  nor2s1 __9_9__514445(.DIN1 (_________41133), .DIN2 (____9___27651),
       .Q (_________41134));
  nnd2s1 __9_9_514446(.DIN1 (________29379), .DIN2 (________28242), .Q
       (_________41133));
  or2s1 __9_9_514447(.DIN1 (_________41135), .DIN2 (______0__41250), .Q
       (_________41136));
  nnd2s1 __9_9__514448(.DIN1 (________28034), .DIN2 (________27526), .Q
       (_________41135));
  and2s1 __9_9__514449(.DIN1 (_________41137), .DIN2 (________27605),
       .Q (_________41138));
  nor2s1 __9_9__514450(.DIN1 (________28153), .DIN2 (___0_____30656),
       .Q (_________41137));
  and2s1 __9_9__514451(.DIN1 (______9__41139), .DIN2 (________24768),
       .Q (______0__41140));
  nor2s1 __9_9__514452(.DIN1 (________26421), .DIN2 (___0____26993), .Q
       (______9__41139));
  or2s1 __9_9__514453(.DIN1 (_________41141), .DIN2 (_____9__26447), .Q
       (_________41142));
  nnd2s1 __9_9__514454(.DIN1 (__9_9___30267), .DIN2 (________27353), .Q
       (_________41141));
  and2s1 __9_9__514455(.DIN1 (_________41143), .DIN2 (____0___27393),
       .Q (_________41144));
  nor2s1 __9_9_514456(.DIN1 (_____0__25778), .DIN2 (________26423), .Q
       (_________41143));
  and2s1 __9_9_514457(.DIN1 (_________41145), .DIN2 (____0____31517),
       .Q (_________41146));
  nor2s1 __9_9__514458(.DIN1 (_________32755), .DIN2 (________26807),
       .Q (_________41145));
  and2s1 __9_9__514459(.DIN1 (_________41147), .DIN2 (_____0__27419),
       .Q (_________41148));
  nor2s1 __9_9__514460(.DIN1 (________26656), .DIN2 (___0____27873), .Q
       (_________41147));
  or2s1 __9_9__514461(.DIN1 (______9__41149), .DIN2 (________27221), .Q
       (______0__41150));
  nnd2s1 __9_9__514462(.DIN1 (____0____33459), .DIN2 (________25733),
       .Q (______9__41149));
  or2s1 __9_9__514463(.DIN1 (_________41151), .DIN2 (________27582), .Q
       (_________41152));
  nnd2s1 __9_9__514464(.DIN1 (_________32140), .DIN2 (________26369),
       .Q (_________41151));
  nor2s1 __9_9__514465(.DIN1 (_________41153), .DIN2 (____0___27214),
       .Q (_________41154));
  nnd2s1 __9_9_514466(.DIN1 (___0__9__30880), .DIN2 (____0____31517),
       .Q (_________41153));
  nnd2s1 __9_9_514467(.DIN1 (_________41155), .DIN2 (___0_____30894),
       .Q (_________41156));
  nor2s1 __9_9__514468(.DIN1 (________26481), .DIN2 (_________32071),
       .Q (_________41155));
  nnd2s1 __9_9__514469(.DIN1 (_________41157), .DIN2 (________27256),
       .Q (_________41158));
  nor2s1 __9_9__514470(.DIN1 (_____9___41301), .DIN2 (________27220),
       .Q (_________41157));
  or2s1 __9_9__514471(.DIN1 (______9__41159), .DIN2 (______0__41270),
       .Q (______0__41160));
  nnd2s1 __9_9__514472(.DIN1 (____9___26404), .DIN2 (________27173), .Q
       (______9__41159));
  or2s1 __9_9__514473(.DIN1 (_________41161), .DIN2 (________28131), .Q
       (_________41162));
  nnd2s1 __9_9__514474(.DIN1 (_____9__27967), .DIN2 (____09___31598),
       .Q (_________41161));
  and2s1 __9_9__514475(.DIN1 (_________41163), .DIN2 (_____0__26547),
       .Q (_________41164));
  nor2s1 __9_9_514476(.DIN1 (________27627), .DIN2 (___9____26942), .Q
       (_________41163));
  and2s1 __9_9_514477(.DIN1 (_________41165), .DIN2 (________27726), .Q
       (_________41166));
  nor2s1 __9_9__514478(.DIN1 (________29359), .DIN2 (________27608), .Q
       (_________41165));
  nnd2s1 __9_9__514479(.DIN1 (_________41167), .DIN2 (____0___27035),
       .Q (_________41168));
  nor2s1 __9_9__514480(.DIN1 (____0____32521), .DIN2 (________26730),
       .Q (_________41167));
  nnd2s1 __9_9__514481(.DIN1 (______9__41169), .DIN2 (___0_0__26960),
       .Q (______0__41170));
  nor2s1 __9_9__514482(.DIN1 (_____9__26635), .DIN2 (________27964), .Q
       (______9__41169));
  and2s1 __9_9__514483(.DIN1 (_________41171), .DIN2 (________28497),
       .Q (_________41172));
  nor2s1 __9_9__514484(.DIN1 (____0___27925), .DIN2 (________27554), .Q
       (_________41171));
  and2s1 __9_9__514485(.DIN1 (_________41173), .DIN2 (_____9__27084),
       .Q (_________41174));
  nor2s1 __9_9_514486(.DIN1 (___0_0__26122), .DIN2 (___9____27774), .Q
       (_________41173));
  or2s1 __9_9_514487(.DIN1 (_________41175), .DIN2 (________27242), .Q
       (_________41176));
  or2s1 __9_9__514488(.DIN1 (____99__26682), .DIN2 (________26662), .Q
       (_________41175));
  and2s1 __9_9__514489(.DIN1 (_________41177), .DIN2 (______0__31825),
       .Q (_________41178));
  nor2s1 __9_9__514490(.DIN1 (____0____31545), .DIN2 (___0_0___30649),
       .Q (_________41177));
  nor2s1 __9_9__514491(.DIN1 (______9__41179), .DIN2 (___09___27028),
       .Q (______0__41180));
  nnd2s1 __9_9__514492(.DIN1 (____9____33353), .DIN2 (____9___25854),
       .Q (______9__41179));
  or2s1 __9_9__514493(.DIN1 (_________41181), .DIN2 (_________41351),
       .Q (_________41182));
  nnd2s1 __9_9__514494(.DIN1 (___0____26070), .DIN2 (________27468), .Q
       (_________41181));
  and2s1 __9_9__514495(.DIN1 (_________41183), .DIN2
       (______________________________________________21930), .Q
       (_________41184));
  nor2s1 __9_9_514496(.DIN1 (________26787), .DIN2 (____0_0__38093), .Q
       (_________41183));
  nor2s1 __9_9_514497(.DIN1 (_________41185), .DIN2 (___0_____40574),
       .Q (_________41186));
  nnd2s1 __9_9__514498(.DIN1 (________26514), .DIN2 (___0_9___40559),
       .Q (_________41185));
  nor2s1 __9_9__514499(.DIN1 (_________41187), .DIN2 (________24489),
       .Q (_________41188));
  nnd2s1 __9_9__514500(.DIN1 (___0____26073), .DIN2 (_____0__27411), .Q
       (_________41187));
  or2s1 __9_9__514501(.DIN1 (______9__41189), .DIN2 (___0____26118), .Q
       (______0__41190));
  nnd2s1 __9_9__514502(.DIN1 (________27365), .DIN2 (________26242), .Q
       (______9__41189));
  nor2s1 __9_9__514503(.DIN1 (_________41191), .DIN2 (___9____27798),
       .Q (_________41192));
  nnd2s1 __9_9__514504(.DIN1 (________27309), .DIN2 (________25694), .Q
       (_________41191));
  or2s1 __9_9__514505(.DIN1 (_________41193), .DIN2 (___0_____31198),
       .Q (_________41194));
  or2s1 __9_9_514506(.DIN1 (___9____27771), .DIN2 (___99___26042), .Q
       (_________41193));
  and2s1 __9_9_514507(.DIN1 (_________41195), .DIN2 (________25706), .Q
       (_________41196));
  nor2s1 __9_9__514508(.DIN1 (___9____26885), .DIN2 (___9____26942), .Q
       (_________41195));
  nor2s1 __9_9__514509(.DIN1 (_________41197), .DIN2 (_____9__26812),
       .Q (_________41198));
  nnd2s1 __9_9__514510(.DIN1 (___0_____31164), .DIN2 (____9____33362),
       .Q (_________41197));
  or2s1 __9_9__514511(.DIN1 (______9__41199), .DIN2 (________26764), .Q
       (_____90__41200));
  nnd2s1 __9_9__514512(.DIN1 (___90___25966), .DIN2 (________26190), .Q
       (______9__41199));
  or2s1 __9_9__514513(.DIN1 (_____9___41201), .DIN2 (___0__0__40571),
       .Q (_____9___41202));
  nnd2s1 __9_9__514514(.DIN1 (___0_0__26069), .DIN2 (____0_0__37159),
       .Q (_____9___41201));
  nor2s1 __9_9__514515(.DIN1 (_____9___41203), .DIN2 (____0___27488),
       .Q (_____9___41204));
  nnd2s1 __9_9_514516(.DIN1 (_________31831), .DIN2 (________25709), .Q
       (_____9___41203));
  and2s1 __9_514517(.DIN1 (_____9___41205), .DIN2 (___9____26900), .Q
       (_____9___41206));
  nor2s1 __9_99_514518(.DIN1 (________24814), .DIN2 (________27161), .Q
       (_____9___41205));
  or2s1 __9_99_514519(.DIN1 (_____9___41207), .DIN2 (___0____23270), .Q
       (_____9___41208));
  nnd2s1 __9_99_514520(.DIN1 (________24596), .DIN2 (________26299), .Q
       (_____9___41207));
  and2s1 __9_99_514521(.DIN1 (_____99__41209), .DIN2 (______0___22056),
       .Q (_____00__41210));
  nor2s1 __9_99_514522(.DIN1 (________27052), .DIN2 (________22927), .Q
       (_____99__41209));
  or2s1 __9_99_514523(.DIN1 (_____0___41211), .DIN2 (___90___25961), .Q
       (_____0___41212));
  nnd2s1 __9_99_514524(.DIN1 (___________), .DIN2 (________27071), .Q
       (_____0___41211));
  and2s1 __9_99_514525(.DIN1 (_____0___41213), .DIN2 (________24823),
       .Q (_____0___41214));
  nor2s1 __9_514526(.DIN1 (________26561), .DIN2 (________27042), .Q
       (_____0___41213));
  or2s1 __9_514527(.DIN1 (_____0___41215), .DIN2 (________26472), .Q
       (_____0___41216));
  nnd2s1 __9_00_514528(.DIN1 (_____0__27039), .DIN2 (________25246), .Q
       (_____0___41215));
  nnd2s1 __9_00_514529(.DIN1 (_____0___41217), .DIN2 (___9____25969),
       .Q (_____0___41218));
  nor2s1 __9_00_514530(.DIN1 (________26760), .DIN2 (________26289), .Q
       (_____0___41217));
  or2s1 __9_00_514531(.DIN1 (_____09__41219), .DIN2 (_____9__27176), .Q
       (______0__41220));
  nnd2s1 __9_00_514532(.DIN1 (________25345), .DIN2 (________25552), .Q
       (_____09__41219));
  and2s1 __9_00_514533(.DIN1 (_________41221), .DIN2 (__9__0__30234),
       .Q (_________41222));
  nor2s1 __9_00_514534(.DIN1 (__9_____30115), .DIN2 (________26613), .Q
       (_________41221));
  and2s1 __9_00_514535(.DIN1 (_________41223), .DIN2 (________27602),
       .Q (_________41224));
  nor2s1 __9_514536(.DIN1 (____0___27484), .DIN2 (________28860), .Q
       (_________41223));
  or2s1 __9_0_514537(.DIN1 (_________41225), .DIN2 (________26337), .Q
       (_________41226));
  nnd2s1 __9_0__514538(.DIN1 (________29181), .DIN2 (____9___29190), .Q
       (_________41225));
  or2s1 __9_0__514539(.DIN1 (_________41227), .DIN2 (__90_9__29708), .Q
       (_________41228));
  nnd2s1 __9_0__514540(.DIN1 (inData[24]), .DIN2 (______________22106),
       .Q (_________41227));
  or2s1 __9_0__514541(.DIN1 (______9__41229), .DIN2 (____0___25413), .Q
       (______0__41230));
  nnd2s1 __9_0__514542(.DIN1 (_____9__25757), .DIN2 (_____0__26832), .Q
       (______9__41229));
  nor2s1 __9_0__514543(.DIN1 (_________41231), .DIN2 (_____9__25738),
       .Q (_________41232));
  nnd2s1 __9_0__514544(.DIN1 (___0_____40549), .DIN2 (_____9__26765),
       .Q (_________41231));
  nnd2s1 __9_0__514545(.DIN1 (_________41233), .DIN2 (________26181),
       .Q (_________41234));
  nor2s1 __9_0_514546(.DIN1 (________29354), .DIN2 (____9___25580), .Q
       (_________41233));
  or2s1 __9_0_514547(.DIN1 (_________41235), .DIN2 (___0_0__26102), .Q
       (_________41236));
  nnd2s1 __9_0__514548(.DIN1 (____0___27398), .DIN2 (________24888), .Q
       (_________41235));
  nor2s1 __9_0__514549(.DIN1 (_________41237), .DIN2 (________26198),
       .Q (_________41238));
  nnd2s1 __9_0__514550(.DIN1 (__9_____30239), .DIN2 (________28870), .Q
       (_________41237));
  or2s1 __9_0__514551(.DIN1 (______9__41239), .DIN2 (___0____22294), .Q
       (______0__41240));
  nnd2s1 __9_0__514552(.DIN1 (________25525), .DIN2 (_________33596),
       .Q (______9__41239));
  and2s1 __9_0__514553(.DIN1 (_________41241), .DIN2 (____9___25494),
       .Q (_________41242));
  nor2s1 __9_0__514554(.DIN1 (___9____26942), .DIN2 (________27378), .Q
       (_________41241));
  and2s1 __9_0__514555(.DIN1 (_________41243), .DIN2 (____9___25764),
       .Q (_________41244));
  nor2s1 __9_0_514556(.DIN1 (___9____27774), .DIN2 (____0___28479), .Q
       (_________41243));
  and2s1 __9_0_514557(.DIN1 (_________41245), .DIN2 (___9____26915), .Q
       (_________41246));
  nor2s1 __9_0__514558(.DIN1 (_________31942), .DIN2 (________28310),
       .Q (_________41245));
  and2s1 __9_0__514559(.DIN1 (_________41247), .DIN2 (________23658),
       .Q (_________41248));
  and2s1 __9_0__514560(.DIN1 (___0____23239), .DIN2 (_____9__25397), .Q
       (_________41247));
  and2s1 __9_0__514561(.DIN1 (______9__41249), .DIN2 (________25515),
       .Q (______0__41250));
  nor2s1 __9_0__514562(.DIN1 (_____0__25417), .DIN2 (___9____26019), .Q
       (______9__41249));
  and2s1 __9_0__514563(.DIN1 (_________41251), .DIN2 (____9___25024),
       .Q (_________41252));
  nor2s1 __9_0__514564(.DIN1 (________25549), .DIN2 (________25448), .Q
       (_________41251));
  and2s1 __9_0__514565(.DIN1 (_________41253), .DIN2 (_____9__24924),
       .Q (_________41254));
  nor2s1 __9_0_514566(.DIN1 (________23840), .DIN2 (____0___26501), .Q
       (_________41253));
  or2s1 __9_0_514567(.DIN1 (_________41255), .DIN2 (_________34644), .Q
       (_________41256));
  nor2s1 __9_0__514568(.DIN1
       (____________________________________________21832), .DIN2
       (________25831), .Q (_________41255));
  or2s1 __9_0__514569(.DIN1 (_________41257), .DIN2 (___9____25091), .Q
       (_________41258));
  nnd2s1 __9_0__514570(.DIN1 (___9____25975), .DIN2 (_____9__26727), .Q
       (_________41257));
  and2s1 __9_0__514571(.DIN1 (______9__41259), .DIN2 (_____0__25010),
       .Q (______0__41260));
  nor2s1 __9_0__514572(.DIN1 (___0____23278), .DIN2 (________26450), .Q
       (______9__41259));
  nor2s1 __9_0__514573(.DIN1 (_________41261), .DIN2 (________23920),
       .Q (_________41262));
  nnd2s1 __9_0__514574(.DIN1 (________25749), .DIN2 (________25690), .Q
       (_________41261));
  or2s1 __9_0__514575(.DIN1 (_________41263), .DIN2 (________24609), .Q
       (_________41264));
  or2s1 __9_0_514576(.DIN1 (________24950), .DIN2 (____9___24454), .Q
       (_________41263));
  or2s1 __9_0_514577(.DIN1 (_________41265), .DIN2 (_____0__26149), .Q
       (_________41266));
  nnd2s1 __9_0__514578(.DIN1 (________24816), .DIN2 (____9___26316), .Q
       (_________41265));
  and2s1 __9_0__514579(.DIN1 (_________41267), .DIN2 (________26429),
       .Q (_________41268));
  nor2s1 __9_0__514580(.DIN1 (___9_0__25978), .DIN2 (_____9__24857), .Q
       (_________41267));
  and2s1 __9_0__514581(.DIN1 (______9__41269), .DIN2 (________25547),
       .Q (______0__41270));
  nor2s1 __9_0__514582(.DIN1 (________25391), .DIN2
       (_____________________21682), .Q (______9__41269));
  and2s1 __9_0__514583(.DIN1 (______0__41366), .DIN2 (________23953),
       .Q (_________41271));
  and2s1 __9_0__514584(.DIN1 (_________41272), .DIN2 (________25690),
       .Q (_________41273));
  nor2s1 __9_0_514585(.DIN1 (_____9__24954), .DIN2 (_____0__24316), .Q
       (_________41272));
  and2s1 __9_0_514586(.DIN1 (_________41274), .DIN2 (____0___25229), .Q
       (_________41275));
  nor2s1 __9_0__514587(.DIN1 (________23451), .DIN2 (________24852), .Q
       (_________41274));
  and2s1 __9_0__514588(.DIN1 (_________41276), .DIN2
       (_____________________________________________21900), .Q
       (_________41277));
  nor2s1 __9_0__514589(.DIN1 (___9_90__39245), .DIN2 (________24880),
       .Q (_________41276));
  or2s1 __9_0__514590(.DIN1 (______9__41278), .DIN2 (________24873), .Q
       (______0__41279));
  nnd2s1 __9_0__514591(.DIN1 (________25640), .DIN2 (____0___26146), .Q
       (______9__41278));
  or2s1 __9_0__514592(.DIN1 (_________41280), .DIN2 (________25466), .Q
       (_________41281));
  nnd2s1 __9_0__514593(.DIN1 (________27150), .DIN2 (____0___26146), .Q
       (_________41280));
  and2s1 __9_0__514594(.DIN1 (_________41282), .DIN2 (________25508),
       .Q (_________41283));
  nor2s1 __9_0_514595(.DIN1 (___0____26067), .DIN2 (________24417), .Q
       (_________41282));
  and2s1 __9_0_514596(.DIN1 (_________41284), .DIN2 (________24875), .Q
       (_________41285));
  nor2s1 __9_0__514597(.DIN1 (___9_9__25057), .DIN2 (________25018), .Q
       (_________41284));
  and2s1 __9_0__514598(.DIN1 (_________41286), .DIN2 (________25270),
       .Q (_________41287));
  nor2s1 __9_0__514599(.DIN1 (_____________________21683), .DIN2
       (_____9__24735), .Q (_________41286));
  or2s1 __9_0__514600(.DIN1 (______9__41288), .DIN2 (___9____23175), .Q
       (______0__41289));
  or2s1 __9_0__514601(.DIN1 (____9___25023), .DIN2 (________23947), .Q
       (______9__41288));
  and2s1 __9_0__514602(.DIN1 (_________41290), .DIN2 (_____9__23944),
       .Q (_________41291));
  nor2s1 __9_0__514603(.DIN1 (________26280), .DIN2 (___9_9__25057), .Q
       (_________41290));
  and2s1 __9_0__514604(.DIN1 (_________41292), .DIN2 (___0_0__24248),
       .Q (_________41293));
  nor2s1 __9_0_514605(.DIN1 (____09__26331), .DIN2 (________23948), .Q
       (_________41292));
  and2s1 __9_0_514606(.DIN1 (_________41294), .DIN2 (________24875), .Q
       (_________41295));
  nor2s1 __9_0__514607(.DIN1 (________24910), .DIN2 (___900__25958), .Q
       (_________41294));
  and2s1 __9_0__514608(.DIN1 (_________41296), .DIN2 (____09__24467),
       .Q (_________41297));
  nor2s1 __9_0__514609(.DIN1 (________25371), .DIN2 (________24901), .Q
       (_________41296));
  and2s1 __9_0__514610(.DIN1 (______9__41298), .DIN2 (___90___25034),
       .Q (_____90__41299));
  nor2s1 __9_0__514611(.DIN1 (____9___25578), .DIN2 (________24658), .Q
       (______9__41298));
  and2s1 __9_0__514612(.DIN1 (_____9___41300), .DIN2 (___9____24136),
       .Q (_____9___41301));
  nor2s1 __9_0__514613(.DIN1 (_____9__24964), .DIN2 (________25278), .Q
       (_____9___41300));
  or2s1 __9_0__514614(.DIN1 (_____9___41302), .DIN2 (________23828), .Q
       (_____9___41303));
  or2s1 __9_0_514615(.DIN1 (________22956), .DIN2 (___0____24229), .Q
       (_____9___41302));
  and2s1 __9_514616(.DIN1 (_____9___41304), .DIN2 (________25354), .Q
       (_____9___41305));
  nor2s1 __9_09_514617(.DIN1 (__________22061), .DIN2 (______0__37872),
       .Q (_____9___41304));
  or2s1 __9_09_514618(.DIN1 (_____9___41306), .DIN2 (______9__37314),
       .Q (_____9___41307));
  nor2s1 __9_09_514619(.DIN1
       (_____________________________________________21825), .DIN2
       (________23533), .Q (_____9___41306));
  or2s1 __9_09_514620(.DIN1 (_____99__41308), .DIN2 (____9___24640), .Q
       (_____00__41309));
  nnd2s1 __9_09_514621(.DIN1 (inData[0]), .DIN2 (___0_____40526), .Q
       (_____99__41308));
  nor2s1 __9_09_514622(.DIN1 (_____0___41310), .DIN2
       (_________________________________________0___21862), .Q
       (_____0___41311));
  nnd2s1 __9_09_514623(.DIN1 (________24044), .DIN2 (___0_0___40566),
       .Q (_____0___41310));
  nnd2s1 __9_09_514624(.DIN1 (_____0___41312), .DIN2 (____9___23687),
       .Q (_____0___41313));
  nor2s1 __9_514625(.DIN1 (_____9__25632), .DIN2 (________24632), .Q
       (_____0___41312));
  and2s1 __9__514626(.DIN1 (_____0___41314), .DIN2 (____00__23788), .Q
       (_____0___41315));
  nor2s1 __9__0_514627(.DIN1 (________26174), .DIN2 (___00___25132), .Q
       (_____0___41314));
  nor2s1 __9__0_514628(.DIN1 (_____0___41316), .DIN2 (_____9__24525),
       .Q (_____0___41317));
  nnd2s1 __9__0_514629(.DIN1 (________24395), .DIN2 (________25569), .Q
       (_____0___41316));
  or2s1 __9__0_514630(.DIN1 (_____09__41318), .DIN2 (_____0__24326), .Q
       (______0__41319));
  nnd2s1 __9__0_514631(.DIN1 (___0____25176), .DIN2 (____9___23588), .Q
       (_____09__41318));
  or2s1 __9__0_514632(.DIN1 (_________41320), .DIN2 (____9___24830), .Q
       (_________41321));
  nnd2s1 __9__0_514633(.DIN1 (_____9__23928), .DIN2 (___9_0___39344),
       .Q (_________41320));
  nnd2s1 __9__0_514634(.DIN1 (_________41322), .DIN2 (___0____24201),
       .Q (_________41323));
  nor2s1 __9__514635(.DIN1
       (____________________________________________21807), .DIN2
       (____0_0__38093), .Q (_________41322));
  or2s1 __9___514636(.DIN1 (_________41324), .DIN2 (_____0__24393), .Q
       (_________41325));
  nnd2s1 __9____514637(.DIN1 (___9____25984), .DIN2 (_____0__24478), .Q
       (_________41324));
  and2s1 __9____514638(.DIN1 (_________41326), .DIN2 (___0_0__24248),
       .Q (_________41327));
  nor2s1 __9____514639(.DIN1 (___00___25132), .DIN2 (________23672), .Q
       (_________41326));
  and2s1 __9____514640(.DIN1 (______9__41328), .DIN2 (________23933),
       .Q (______0__41329));
  nor2s1 __9____514641(.DIN1 (________25371), .DIN2 (________23946), .Q
       (______9__41328));
  nnd2s1 __9____514642(.DIN1 (_________41330), .DIN2 (________23669),
       .Q (_________41331));
  nor2s1 __9____514643(.DIN1 (___0____25204), .DIN2 (___9____23177), .Q
       (_________41330));
  and2s1 __9____514644(.DIN1 (_________41332), .DIN2 (___9____23144),
       .Q (_________41333));
  nor2s1 __9___514645(.DIN1 (____9___24066), .DIN2 (________23430), .Q
       (_________41332));
  or2s1 __9___514646(.DIN1 (_________41334), .DIN2 (________23903), .Q
       (_________41335));
  nnd2s1 __9____514647(.DIN1 (________23984), .DIN2 (_____0__25556), .Q
       (_________41334));
  or2s1 __9____514648(.DIN1 (_________41336), .DIN2 (___0_0__23235), .Q
       (_________41337));
  nnd2s1 __9____514649(.DIN1 (___9____23150), .DIN2 (___909), .Q
       (_________41336));
  and2s1 __9____514650(.DIN1 (______9__41338), .DIN2 (___0____22310),
       .Q (______0__41339));
  nor2s1 __9____514651(.DIN1 (________24351), .DIN2 (____9___23400), .Q
       (______9__41338));
  or2s1 __9____514652(.DIN1 (_________41340), .DIN2 (_____0__23702), .Q
       (_________41341));
  nnd2s1 __9____514653(.DIN1 (________24280), .DIN2 (___9____23142), .Q
       (_________41340));
  or2s1 __9____514654(.DIN1 (_________41342), .DIN2 (________22904), .Q
       (_________41343));
  or2s1 __9___514655(.DIN1 (___099__23309), .DIN2 (_____9__22888), .Q
       (_________41342));
  and2s1 __9___514656(.DIN1 (_________41344), .DIN2 (_____0__23086), .Q
       (_________41345));
  or2s1 __9____514657(.DIN1 (________23383), .DIN2 (________22976), .Q
       (_________41344));
  or2s1 __9____514658(.DIN1 (_________41346), .DIN2 (____9____34370),
       .Q (_________41347));
  nnd2s1 __9____514659(.DIN1 (inData[26]), .DIN2
       (____________________________________________21789), .Q
       (_________41346));
  and2s1 __9____514660(.DIN1 (______9__41348), .DIN2 (_____9___37656),
       .Q (______0__41349));
  nnd2s1 __9____514661(.DIN1 (___0_0___40464), .DIN2 (inData[8]), .Q
       (______9__41348));
  and2s1 __9____514662(.DIN1 (_________41350), .DIN2 (________23523),
       .Q (_________41351));
  and2s1 __9____514663(.DIN1 (___00___25129), .DIN2 (________23667), .Q
       (_________41350));
  and2s1 __9____514664(.DIN1 (_________41352), .DIN2 (_____0__22701),
       .Q (_________41353));
  or2s1 __9___514665(.DIN1 (___0____26120), .DIN2 (________23959), .Q
       (_________41352));
  or2s1 __9___514666(.DIN1 (_________41354), .DIN2 (_________34232), .Q
       (_________41355));
  xor2s1 __9____514667(.DIN1 (_____9___38512), .DIN2 (_________34989),
       .Q (_________41354));
  or2s1 __9____514668(.DIN1 (_________41356), .DIN2 (_________33672),
       .Q (_________41357));
  xor2s1 __9____514669(.DIN1 (___9__9__39125), .DIN2 (_________34956),
       .Q (_________41356));
  or2s1 __9____514670(.DIN1 (______9__41358), .DIN2 (_________32907),
       .Q (______0__41359));
  xor2s1 __9____514671(.DIN1 (_____9___36721), .DIN2 (_________34864),
       .Q (______9__41358));
  or2s1 __9____514672(.DIN1 (_________41360), .DIN2 (________28457), .Q
       (_________41361));
  nnd2s1 __9____514673(.DIN1 (____90__28285), .DIN2 (_________40947),
       .Q (_________41360));
  nor2s1 __9____514674(.DIN1 (_________41362), .DIN2 (_________41194),
       .Q (_________41363));
  nnd2s1 __9___514675(.DIN1 (___9____28674), .DIN2 (_________40986), .Q
       (_________41362));
  and2s1 __9___514676(.DIN1 (_________41364), .DIN2 (___99___23212), .Q
       (_________41365));
  xnr2s1 __9____514677(.DIN1 (____0___27657), .DIN2 (____90___36104),
       .Q (_________41364));
  nor2s1 __9____514678(.DIN1 (___0____26087), .DIN2 (________24804), .Q
       (______0__41366));
  xnr2s1 __9____514679(.DIN1 (____9____38919), .DIN2 (___9_0___39705),
       .Q (_________41372));
endmodule

