
module fir_core_obf(inData, clk, reset, outData);
  input [31:0] inData;
  input clk, reset;
  output [31:0] outData;
  wire [31:0] inData;
  wire clk, reset;
  wire [31:0] outData;
  wire __0, __9, __9_0, __9_00, __9_00__26419, __9_00__26514,
       __9_00__26702, __9_00__26798;
  wire __9_00__26892, __9_00__26989, __9_0_, __9_0___26334,
       __9_0___26335, __9_0___26336, __9_0___26337, __9_0___26338;
  wire __9_0___26339, __9_0___26340, __9_0___26420, __9_0___26421,
       __9_0___26422, __9_0___26423, __9_0___26424, __9_0___26425;
  wire __9_0___26426, __9_0___26427, __9_0___26515, __9_0___26516,
       __9_0___26517, __9_0___26518, __9_0___26519, __9_0___26520;
  wire __9_0___26521, __9_0___26609, __9_0___26610, __9_0___26611,
       __9_0___26612, __9_0___26613, __9_0___26614, __9_0___26615;
  wire __9_0___26616, __9_0___26703, __9_0___26704, __9_0___26705,
       __9_0___26706, __9_0___26707, __9_0___26708, __9_0___26709;
  wire __9_0___26710, __9_0___26799, __9_0___26800, __9_0___26801,
       __9_0___26802, __9_0___26803, __9_0___26804, __9_0___26805;
  wire __9_0___26806, __9_0___26893, __9_0___26894, __9_0___26895,
       __9_0___26896, __9_0___26897, __9_0___26898, __9_0___26899;
  wire __9_0___26900, __9_0___26990, __9_0___26991, __9_0___26992,
       __9_0___26993, __9_0___26994, __9_09, __9_09__26428;
  wire __9_09__26522, __9_09__26617, __9_09__26711, __9_09__26807,
       __9_09__26901, __9_09__26995, __9_9_, __9_9___26413;
  wire __9_9___26414, __9_9___26415, __9_9___26416, __9_9___26417,
       __9_9___26418, __9_9___26505, __9_9___26506, __9_9___26507;
  wire __9_9___26508, __9_9___26509, __9_9___26510, __9_9___26511,
       __9_9___26512, __9_9___26600, __9_9___26601, __9_9___26602;
  wire __9_9___26603, __9_9___26604, __9_9___26605, __9_9___26606,
       __9_9___26607, __9_9___26693, __9_9___26694, __9_9___26695;
  wire __9_9___26696, __9_9___26697, __9_9___26698, __9_9___26699,
       __9_9___26700, __9_9___26789, __9_9___26790, __9_9___26791;
  wire __9_9___26792, __9_9___26793, __9_9___26794, __9_9___26795,
       __9_9___26796, __9_9___26884, __9_9___26885, __9_9___26886;
  wire __9_9___26887, __9_9___26888, __9_9___26889, __9_9___26890,
       __9_9___26980, __9_9___26981, __9_9___26982, __9_9___26983;
  wire __9_9___26984, __9_9___26985, __9_9___26986, __9_9___26987,
       __9_9___27075, __9_9___27076, __9_9___27077, __9_9___27078;
  wire __9_9___27079, __9_9___27080, __9_9___27081, __9_90,
       __9_90__26504, __9_90__26599, __9_90__26692, __9_90__26788;
  wire __9_90__26883, __9_90__26979, __9_90__27074, __9_99,
       __9_99__26513, __9_99__26608, __9_99__26701, __9_99__26797;
  wire __9_99__26891, __9_99__26988, __9_99__27082, __9__0,
       __9__0__26346, __9__0__26356, __9__0__26366, __9__0__26376;
  wire __9__0__26394, __9__0__26403, __9__0__26429, __9__0__26439,
       __9__0__26449, __9__0__26459, __9__0__26467, __9__0__26477;
  wire __9__0__26485, __9__0__26494, __9__0__26523, __9__0__26532,
       __9__0__26541, __9__0__26551, __9__0__26560, __9__0__26570;
  wire __9__0__26589, __9__0__26618, __9__0__26628, __9__0__26637,
       __9__0__26645, __9__0__26654, __9__0__26664, __9__0__26674;
  wire __9__0__26683, __9__0__26712, __9__0__26720, __9__0__26729,
       __9__0__26739, __9__0__26749, __9__0__26758, __9__0__26768;
  wire __9__0__26778, __9__0__26816, __9__0__26825, __9__0__26834,
       __9__0__26844, __9__0__26854, __9__0__26864, __9__0__26873;
  wire __9__0__26902, __9__0__26912, __9__0__26922, __9__0__26931,
       __9__0__26941, __9__0__26951, __9__0__26961, __9__0__26969;
  wire __9__0__26996, __9__0__27005, __9__0__27015, __9__0__27025,
       __9__0__27035, __9__0__27044, __9__0__27054, __9__0__27064;
  wire __9__9, __9__9__26355, __9__9__26365, __9__9__26375,
       __9__9__26384, __9__9__26393, __9__9__26412, __9__9__26438;
  wire __9__9__26448, __9__9__26458, __9__9__26476, __9__9__26484,
       __9__9__26493, __9__9__26503, __9__9__26531, __9__9__26540;
  wire __9__9__26550, __9__9__26559, __9__9__26569, __9__9__26579,
       __9__9__26588, __9__9__26598, __9__9__26627, __9__9__26636;
  wire __9__9__26644, __9__9__26653, __9__9__26663, __9__9__26673,
       __9__9__26682, __9__9__26691, __9__9__26719, __9__9__26738;
  wire __9__9__26748, __9__9__26757, __9__9__26767, __9__9__26777,
       __9__9__26787, __9__9__26815, __9__9__26824, __9__9__26833;
  wire __9__9__26843, __9__9__26853, __9__9__26863, __9__9__26872,
       __9__9__26882, __9__9__26911, __9__9__26921, __9__9__26930;
  wire __9__9__26940, __9__9__26950, __9__9__26960, __9__9__26968,
       __9__9__26978, __9__9__27014, __9__9__27024, __9__9__27034;
  wire __9__9__27043, __9__9__27053, __9__9__27063, __9__9__27073,
       __9___, __9_____26341, __9_____26342, __9_____26343;
  wire __9_____26344, __9_____26345, __9_____26347, __9_____26348,
       __9_____26349, __9_____26350, __9_____26351, __9_____26352;
  wire __9_____26353, __9_____26354, __9_____26357, __9_____26358,
       __9_____26359, __9_____26360, __9_____26361, __9_____26362;
  wire __9_____26363, __9_____26364, __9_____26367, __9_____26368,
       __9_____26369, __9_____26370, __9_____26371, __9_____26372;
  wire __9_____26373, __9_____26374, __9_____26377, __9_____26378,
       __9_____26379, __9_____26380, __9_____26381, __9_____26382;
  wire __9_____26383, __9_____26385, __9_____26386, __9_____26387,
       __9_____26388, __9_____26389, __9_____26390, __9_____26391;
  wire __9_____26392, __9_____26395, __9_____26396, __9_____26397,
       __9_____26398, __9_____26399, __9_____26400, __9_____26401;
  wire __9_____26402, __9_____26404, __9_____26405, __9_____26406,
       __9_____26407, __9_____26408, __9_____26409, __9_____26410;
  wire __9_____26411, __9_____26430, __9_____26431, __9_____26432,
       __9_____26433, __9_____26434, __9_____26435, __9_____26436;
  wire __9_____26437, __9_____26440, __9_____26441, __9_____26442,
       __9_____26443, __9_____26444, __9_____26445, __9_____26446;
  wire __9_____26447, __9_____26450, __9_____26451, __9_____26452,
       __9_____26453, __9_____26454, __9_____26455, __9_____26456;
  wire __9_____26457, __9_____26460, __9_____26461, __9_____26462,
       __9_____26463, __9_____26464, __9_____26465, __9_____26466;
  wire __9_____26468, __9_____26469, __9_____26470, __9_____26471,
       __9_____26472, __9_____26473, __9_____26474, __9_____26475;
  wire __9_____26478, __9_____26479, __9_____26480, __9_____26481,
       __9_____26482, __9_____26483, __9_____26486, __9_____26487;
  wire __9_____26488, __9_____26489, __9_____26490, __9_____26491,
       __9_____26492, __9_____26495, __9_____26496, __9_____26497;
  wire __9_____26498, __9_____26499, __9_____26500, __9_____26501,
       __9_____26502, __9_____26524, __9_____26525, __9_____26526;
  wire __9_____26527, __9_____26528, __9_____26529, __9_____26530,
       __9_____26533, __9_____26534, __9_____26535, __9_____26536;
  wire __9_____26537, __9_____26538, __9_____26539, __9_____26542,
       __9_____26543, __9_____26544, __9_____26545, __9_____26546;
  wire __9_____26547, __9_____26548, __9_____26549, __9_____26552,
       __9_____26553, __9_____26554, __9_____26555, __9_____26556;
  wire __9_____26557, __9_____26558, __9_____26561, __9_____26562,
       __9_____26563, __9_____26564, __9_____26565, __9_____26566;
  wire __9_____26567, __9_____26568, __9_____26571, __9_____26572,
       __9_____26573, __9_____26574, __9_____26575, __9_____26576;
  wire __9_____26577, __9_____26578, __9_____26580, __9_____26581,
       __9_____26582, __9_____26583, __9_____26584, __9_____26585;
  wire __9_____26586, __9_____26587, __9_____26590, __9_____26591,
       __9_____26592, __9_____26593, __9_____26594, __9_____26595;
  wire __9_____26596, __9_____26597, __9_____26619, __9_____26620,
       __9_____26621, __9_____26622, __9_____26623, __9_____26624;
  wire __9_____26625, __9_____26626, __9_____26629, __9_____26630,
       __9_____26631, __9_____26632, __9_____26633, __9_____26634;
  wire __9_____26635, __9_____26638, __9_____26639, __9_____26640,
       __9_____26641, __9_____26642, __9_____26643, __9_____26646;
  wire __9_____26647, __9_____26648, __9_____26649, __9_____26650,
       __9_____26651, __9_____26652, __9_____26655, __9_____26656;
  wire __9_____26657, __9_____26658, __9_____26659, __9_____26660,
       __9_____26661, __9_____26662, __9_____26665, __9_____26666;
  wire __9_____26667, __9_____26668, __9_____26669, __9_____26670,
       __9_____26671, __9_____26672, __9_____26675, __9_____26676;
  wire __9_____26677, __9_____26678, __9_____26679, __9_____26680,
       __9_____26681, __9_____26684, __9_____26685, __9_____26686;
  wire __9_____26687, __9_____26688, __9_____26689, __9_____26690,
       __9_____26713, __9_____26714, __9_____26715, __9_____26716;
  wire __9_____26717, __9_____26718, __9_____26721, __9_____26722,
       __9_____26723, __9_____26724, __9_____26725, __9_____26726;
  wire __9_____26727, __9_____26728, __9_____26730, __9_____26731,
       __9_____26732, __9_____26733, __9_____26734, __9_____26735;
  wire __9_____26736, __9_____26737, __9_____26740, __9_____26741,
       __9_____26742, __9_____26743, __9_____26744, __9_____26745;
  wire __9_____26746, __9_____26747, __9_____26750, __9_____26751,
       __9_____26752, __9_____26753, __9_____26754, __9_____26755;
  wire __9_____26756, __9_____26759, __9_____26760, __9_____26761,
       __9_____26762, __9_____26763, __9_____26764, __9_____26765;
  wire __9_____26766, __9_____26769, __9_____26770, __9_____26771,
       __9_____26772, __9_____26773, __9_____26774, __9_____26775;
  wire __9_____26776, __9_____26779, __9_____26780, __9_____26781,
       __9_____26782, __9_____26783, __9_____26784, __9_____26785;
  wire __9_____26786, __9_____26808, __9_____26809, __9_____26810,
       __9_____26811, __9_____26812, __9_____26813, __9_____26814;
  wire __9_____26817, __9_____26818, __9_____26819, __9_____26820,
       __9_____26821, __9_____26822, __9_____26823, __9_____26826;
  wire __9_____26827, __9_____26828, __9_____26829, __9_____26830,
       __9_____26831, __9_____26832, __9_____26835, __9_____26836;
  wire __9_____26837, __9_____26838, __9_____26839, __9_____26840,
       __9_____26841, __9_____26842, __9_____26845, __9_____26846;
  wire __9_____26847, __9_____26848, __9_____26849, __9_____26850,
       __9_____26851, __9_____26852, __9_____26855, __9_____26856;
  wire __9_____26857, __9_____26858, __9_____26859, __9_____26860,
       __9_____26861, __9_____26862, __9_____26865, __9_____26866;
  wire __9_____26867, __9_____26868, __9_____26869, __9_____26870,
       __9_____26871, __9_____26874, __9_____26875, __9_____26876;
  wire __9_____26877, __9_____26878, __9_____26879, __9_____26880,
       __9_____26881, __9_____26903, __9_____26904, __9_____26905;
  wire __9_____26906, __9_____26907, __9_____26908, __9_____26909,
       __9_____26910, __9_____26913, __9_____26914, __9_____26915;
  wire __9_____26916, __9_____26917, __9_____26918, __9_____26919,
       __9_____26920, __9_____26923, __9_____26924, __9_____26925;
  wire __9_____26926, __9_____26927, __9_____26928, __9_____26929,
       __9_____26932, __9_____26933, __9_____26934, __9_____26935;
  wire __9_____26936, __9_____26937, __9_____26938, __9_____26939,
       __9_____26942, __9_____26943, __9_____26944, __9_____26945;
  wire __9_____26946, __9_____26947, __9_____26948, __9_____26949,
       __9_____26952, __9_____26953, __9_____26954, __9_____26955;
  wire __9_____26956, __9_____26957, __9_____26958, __9_____26959,
       __9_____26962, __9_____26963, __9_____26964, __9_____26965;
  wire __9_____26966, __9_____26967, __9_____26970, __9_____26971,
       __9_____26972, __9_____26973, __9_____26974, __9_____26975;
  wire __9_____26976, __9_____26977, __9_____26997, __9_____26998,
       __9_____26999, __9_____27000, __9_____27001, __9_____27002;
  wire __9_____27003, __9_____27004, __9_____27006, __9_____27007,
       __9_____27008, __9_____27009, __9_____27010, __9_____27011;
  wire __9_____27012, __9_____27013, __9_____27016, __9_____27017,
       __9_____27018, __9_____27019, __9_____27020, __9_____27021;
  wire __9_____27022, __9_____27023, __9_____27026, __9_____27027,
       __9_____27028, __9_____27029, __9_____27030, __9_____27031;
  wire __9_____27032, __9_____27033, __9_____27036, __9_____27037,
       __9_____27038, __9_____27039, __9_____27040, __9_____27041;
  wire __9_____27042, __9_____27045, __9_____27046, __9_____27047,
       __9_____27048, __9_____27049, __9_____27050, __9_____27051;
  wire __9_____27052, __9_____27055, __9_____27056, __9_____27057,
       __9_____27058, __9_____27059, __9_____27060, __9_____27061;
  wire __9_____27062, __9_____27065, __9_____27066, __9_____27067,
       __9_____27068, __9_____27069, __9_____27070, __9_____27071;
  wire __9_____27072, __90_0, __90_0__26261, __90_0__26271,
       __90_0__26281, __90_0__26291, __90_0__26300, __90_0__26309;
  wire __90_0__26318, __90_9, __90_9__26270, __90_9__26280,
       __90_9__26290, __90_9__26299, __90_9__26308, __90_9__26317;
  wire __90_9__26327, __90__, __90____26254, __90____26255,
       __90____26256, __90____26257, __90____26258, __90____26259;
  wire __90____26260, __90____26262, __90____26263, __90____26264,
       __90____26265, __90____26266, __90____26267, __90____26268;
  wire __90____26269, __90____26272, __90____26273, __90____26274,
       __90____26275, __90____26276, __90____26277, __90____26278;
  wire __90____26279, __90____26282, __90____26283, __90____26284,
       __90____26285, __90____26286, __90____26287, __90____26288;
  wire __90____26289, __90____26292, __90____26293, __90____26294,
       __90____26295, __90____26296, __90____26297, __90____26298;
  wire __90____26301, __90____26302, __90____26303, __90____26304,
       __90____26305, __90____26306, __90____26307, __90____26310;
  wire __90____26311, __90____26312, __90____26313, __90____26314,
       __90____26315, __90____26316, __90____26319, __90____26320;
  wire __90____26321, __90____26322, __90____26323, __90____26324,
       __90____26325, __90____26326, __99_0, __99_0__27097;
  wire __99_0__27107, __99_0__27117, __99_0__27126, __99_0__27134,
       __99_0__27144, __99_0__27154, __99_9, __99_9__27106;
  wire __99_9__27116, __99_9__27125, __99_9__27133, __99_9__27143,
       __99_9__27153, __99_9__27162, __99__, __99____27090;
  wire __99____27091, __99____27092, __99____27093, __99____27094,
       __99____27095, __99____27096, __99____27098, __99____27099;
  wire __99____27100, __99____27101, __99____27102, __99____27103,
       __99____27104, __99____27105, __99____27108, __99____27109;
  wire __99____27110, __99____27111, __99____27112, __99____27113,
       __99____27114, __99____27115, __99____27118, __99____27119;
  wire __99____27120, __99____27121, __99____27122, __99____27123,
       __99____27124, __99____27127, __99____27128, __99____27129;
  wire __99____27130, __99____27131, __99____27132, __99____27135,
       __99____27136, __99____27137, __99____27138, __99____27139;
  wire __99____27140, __99____27141, __99____27142, __99____27145,
       __99____27146, __99____27147, __99____27148, __99____27149;
  wire __99____27150, __99____27151, __99____27152, __99____27155,
       __99____27156, __99____27157, __99____27158, __99____27159;
  wire __99____27160, __99____27161, __900_, __900___26247,
       __900___26248, __900___26249, __900___26250, __900___26251;
  wire __900___26252, __900___26253, __909, __909_, __909___26328,
       __909___26329, __909___26330, __909___26331;
  wire __909___26332, __909___26333, __990_, __990___27083,
       __990___27084, __990___27085, __990___27086, __990___27087;
  wire __990___27088, __990___27089, __999_, __999___27163,
       __999___27164, __999___27165, __999___27166, __999___27167;
  wire __999___27168, __999___27169, __9000, __9009, __9090, __9099,
       __9900, __9909;
  wire __9990, ___, ___0, ___00, ___000, ___0000__27170, ___000__20699,
       ___000__21633;
  wire ___000__22536, ___000__23437, ___000__24333, ___000__25271,
       ___000___27171, ___000___27172, ___000___27173, ___000___27174;
  wire ___000___27175, ___000___27176, ___000___27177, ___00_,
       ___00_0__27179, ___00_0__27189, ___00_0__27199, ___00_0__27208;
  wire ___00_0__27218, ___00_0__27228, ___00_0__27238, ___00_0__27247,
       ___00_9__27188, ___00_9__27198, ___00_9__27217, ___00_9__27227;
  wire ___00_9__27237, ___00_9__27246, ___00_9__27256, ___00__19033,
       ___00___19771, ___00___19772, ___00___19773, ___00___19774;
  wire ___00___19775, ___00___19776, ___00___19777, ___00___20700,
       ___00___20701, ___00___20702, ___00___20703, ___00___20704;
  wire ___00___20705, ___00___20706, ___00___21634, ___00___21635,
       ___00___21636, ___00___21637, ___00___21638, ___00___21639;
  wire ___00___21640, ___00___22537, ___00___22538, ___00___22539,
       ___00___22540, ___00___22541, ___00___22542, ___00___22543;
  wire ___00___23438, ___00___23439, ___00___23440, ___00___23441,
       ___00___23442, ___00___23443, ___00___23444, ___00___24334;
  wire ___00___24335, ___00___24336, ___00___24337, ___00___24338,
       ___00___24339, ___00___24340, ___00___24341, ___00___25272;
  wire ___00___25273, ___00___25274, ___00___25275, ___00___25276,
       ___00___25277, ___00___25278, ___00___25279, ___00____27180;
  wire ___00____27181, ___00____27182, ___00____27183, ___00____27184,
       ___00____27185, ___00____27186, ___00____27187, ___00____27190;
  wire ___00____27191, ___00____27192, ___00____27193, ___00____27194,
       ___00____27195, ___00____27196, ___00____27197, ___00____27200;
  wire ___00____27201, ___00____27202, ___00____27203, ___00____27204,
       ___00____27205, ___00____27206, ___00____27207, ___00____27209;
  wire ___00____27210, ___00____27211, ___00____27212, ___00____27213,
       ___00____27214, ___00____27215, ___00____27216, ___00____27219;
  wire ___00____27220, ___00____27221, ___00____27222, ___00____27223,
       ___00____27224, ___00____27225, ___00____27226, ___00____27229;
  wire ___00____27230, ___00____27231, ___00____27232, ___00____27233,
       ___00____27234, ___00____27235, ___00____27236, ___00____27239;
  wire ___00____27240, ___00____27241, ___00____27242, ___00____27243,
       ___00____27244, ___00____27245, ___00____27248, ___00____27249;
  wire ___00____27250, ___00____27251, ___00____27252, ___00____27253,
       ___00____27254, ___00____27255, ___0_, ___0_0;
  wire ___0_00__27267, ___0_00__27364, ___0_00__27461, ___0_00__27656,
       ___0_00__27753, ___0_00__27850, ___0_0__19785, ___0_0__19793;
  wire ___0_0__19810, ___0_0__19826, ___0_0__19835, ___0_0__20708,
       ___0_0__20724, ___0_0__20733, ___0_0__20743, ___0_0__20752;
  wire ___0_0__20762, ___0_0__20771, ___0_0__21641, ___0_0__21649,
       ___0_0__21658, ___0_0__21667, ___0_0__21676, ___0_0__21686;
  wire ___0_0__21696, ___0_0__21705, ___0_0__22554, ___0_0__22564,
       ___0_0__22573, ___0_0__22582, ___0_0__22600, ___0_0__22608;
  wire ___0_0__23455, ___0_0__23464, ___0_0__23473, ___0_0__23481,
       ___0_0__23490, ___0_0__23500, ___0_0__23509, ___0_0__24343;
  wire ___0_0__24352, ___0_0__24362, ___0_0__24372, ___0_0__24382,
       ___0_0__24391, ___0_0__24410, ___0_0__25281, ___0_0__25290;
  wire ___0_0__25300, ___0_0__25310, ___0_0__25319, ___0_0__25328,
       ___0_0__25338, ___0_0__25347, ___0_0___27268, ___0_0___27269;
  wire ___0_0___27270, ___0_0___27271, ___0_0___27272, ___0_0___27273,
       ___0_0___27274, ___0_0___27275, ___0_0___27365, ___0_0___27366;
  wire ___0_0___27367, ___0_0___27368, ___0_0___27369, ___0_0___27370,
       ___0_0___27371, ___0_0___27372, ___0_0___27462, ___0_0___27463;
  wire ___0_0___27464, ___0_0___27465, ___0_0___27466, ___0_0___27467,
       ___0_0___27468, ___0_0___27469, ___0_0___27560, ___0_0___27561;
  wire ___0_0___27562, ___0_0___27563, ___0_0___27564, ___0_0___27565,
       ___0_0___27566, ___0_0___27567, ___0_0___27657, ___0_0___27658;
  wire ___0_0___27659, ___0_0___27660, ___0_0___27661, ___0_0___27662,
       ___0_0___27663, ___0_0___27664, ___0_0___27754, ___0_0___27755;
  wire ___0_0___27756, ___0_0___27757, ___0_0___27758, ___0_0___27759,
       ___0_0___27760, ___0_0___27851, ___0_0___27852, ___0_0___27853;
  wire ___0_0___27854, ___0_0___27855, ___0_0___27856, ___0_0___27857,
       ___0_0___27858, ___0_0___27948, ___0_0___27949, ___0_0___27950;
  wire ___0_0___27951, ___0_0___27952, ___0_0___27953, ___0_09__27276,
       ___0_09__27373, ___0_09__27470, ___0_09__27568, ___0_09__27665;
  wire ___0_09__27761, ___0_09__27859, ___0_09__27954, ___0_9,
       ___0_9__19802, ___0_9__19809, ___0_9__19817, ___0_9__19825;
  wire ___0_9__19834, ___0_9__19844, ___0_9__20715, ___0_9__20723,
       ___0_9__20732, ___0_9__20742, ___0_9__20751, ___0_9__20761;
  wire ___0_9__20770, ___0_9__20779, ___0_9__21648, ___0_9__21657,
       ___0_9__21666, ___0_9__21675, ___0_9__21685, ___0_9__21695;
  wire ___0_9__22553, ___0_9__22563, ___0_9__22572, ___0_9__22581,
       ___0_9__22599, ___0_9__23454, ___0_9__23463, ___0_9__23472;
  wire ___0_9__23489, ___0_9__23499, ___0_9__23517, ___0_9__24351,
       ___0_9__24361, ___0_9__24371, ___0_9__24381, ___0_9__24390;
  wire ___0_9__24400, ___0_9__24409, ___0_9__24418, ___0_9__25289,
       ___0_9__25299, ___0_9__25309, ___0_9__25318, ___0_9__25327;
  wire ___0_9__25337, ___0_9__25346, ___0_9__25356, ___0_9___27355,
       ___0_9___27356, ___0_9___27357, ___0_9___27358, ___0_9___27359;
  wire ___0_9___27360, ___0_9___27361, ___0_9___27362, ___0_9___27454,
       ___0_9___27455, ___0_9___27456, ___0_9___27457, ___0_9___27458;
  wire ___0_9___27459, ___0_9___27552, ___0_9___27553, ___0_9___27554,
       ___0_9___27555, ___0_9___27556, ___0_9___27557, ___0_9___27558;
  wire ___0_9___27559, ___0_9___27647, ___0_9___27648, ___0_9___27649,
       ___0_9___27650, ___0_9___27651, ___0_9___27652, ___0_9___27653;
  wire ___0_9___27654, ___0_9___27744, ___0_9___27745, ___0_9___27746,
       ___0_9___27747, ___0_9___27748, ___0_9___27749, ___0_9___27750;
  wire ___0_9___27751, ___0_9___27841, ___0_9___27842, ___0_9___27843,
       ___0_9___27844, ___0_9___27845, ___0_9___27846, ___0_9___27847;
  wire ___0_9___27848, ___0_9___27939, ___0_9___27940, ___0_9___27941,
       ___0_9___27942, ___0_9___27943, ___0_9___27944, ___0_9___27945;
  wire ___0_9___27946, ___0_9___28033, ___0_9___28034, ___0_9___28035,
       ___0_9___28036, ___0_9___28037, ___0_9___28038, ___0_9___28039;
  wire ___0_9___28040, ___0_90__27354, ___0_90__27453, ___0_90__27551,
       ___0_90__27646, ___0_90__27743, ___0_90__27840, ___0_90__27938;
  wire ___0_90__28032, ___0_99__27363, ___0_99__27460, ___0_99__27655,
       ___0_99__27752, ___0_99__27849, ___0_99__27947, ___0_99__28041;
  wire ___0__, ___0__0__27277, ___0__0__27287, ___0__0__27297,
       ___0__0__27307, ___0__0__27316, ___0__0__27325, ___0__0__27335;
  wire ___0__0__27345, ___0__0__27374, ___0__0__27384, ___0__0__27393,
       ___0__0__27403, ___0__0__27413, ___0__0__27423, ___0__0__27433;
  wire ___0__0__27443, ___0__0__27471, ___0__0__27481, ___0__0__27491,
       ___0__0__27501, ___0__0__27511, ___0__0__27521, ___0__0__27531;
  wire ___0__0__27541, ___0__0__27569, ___0__0__27579, ___0__0__27589,
       ___0__0__27599, ___0__0__27609, ___0__0__27618, ___0__0__27628;
  wire ___0__0__27637, ___0__0__27666, ___0__0__27676, ___0__0__27685,
       ___0__0__27694, ___0__0__27704, ___0__0__27714, ___0__0__27724;
  wire ___0__0__27733, ___0__0__27762, ___0__0__27772, ___0__0__27782,
       ___0__0__27792, ___0__0__27802, ___0__0__27810, ___0__0__27820;
  wire ___0__0__27830, ___0__0__27860, ___0__0__27870, ___0__0__27880,
       ___0__0__27890, ___0__0__27899, ___0__0__27909, ___0__0__27919;
  wire ___0__0__27929, ___0__0__27955, ___0__0__27965, ___0__0__27984,
       ___0__0__27994, ___0__0__28004, ___0__0__28014, ___0__0__28022;
  wire ___0__9__27286, ___0__9__27296, ___0__9__27306, ___0__9__27315,
       ___0__9__27324, ___0__9__27334, ___0__9__27344, ___0__9__27353;
  wire ___0__9__27383, ___0__9__27392, ___0__9__27402, ___0__9__27412,
       ___0__9__27422, ___0__9__27432, ___0__9__27442, ___0__9__27452;
  wire ___0__9__27480, ___0__9__27490, ___0__9__27500, ___0__9__27510,
       ___0__9__27520, ___0__9__27530, ___0__9__27540, ___0__9__27550;
  wire ___0__9__27578, ___0__9__27588, ___0__9__27598, ___0__9__27608,
       ___0__9__27617, ___0__9__27627, ___0__9__27636, ___0__9__27645;
  wire ___0__9__27675, ___0__9__27684, ___0__9__27693, ___0__9__27703,
       ___0__9__27713, ___0__9__27723, ___0__9__27732, ___0__9__27742;
  wire ___0__9__27771, ___0__9__27781, ___0__9__27791, ___0__9__27801,
       ___0__9__27819, ___0__9__27829, ___0__9__27839, ___0__9__27869;
  wire ___0__9__27879, ___0__9__27889, ___0__9__27898, ___0__9__27908,
       ___0__9__27918, ___0__9__27928, ___0__9__27937, ___0__9__27964;
  wire ___0__9__27974, ___0__9__27983, ___0__9__27993, ___0__9__28003,
       ___0__9__28013, ___0__9__28021, ___0__9__28031, ___0__18915;
  wire ___0__18921, ___0__18931, ___0__18935, ___0__18943,
       ___0___18982, ___0___18983, ___0___18984, ___0___18985;
  wire ___0___18986, ___0___18987, ___0___18988, ___0___19034,
       ___0___19042, ___0____19778, ___0____19779, ___0____19780;
  wire ___0____19781, ___0____19782, ___0____19783, ___0____19784,
       ___0____19786, ___0____19787, ___0____19788, ___0____19789;
  wire ___0____19790, ___0____19791, ___0____19792, ___0____19794,
       ___0____19795, ___0____19796, ___0____19797, ___0____19798;
  wire ___0____19799, ___0____19800, ___0____19801, ___0____19803,
       ___0____19804, ___0____19805, ___0____19806, ___0____19807;
  wire ___0____19808, ___0____19811, ___0____19812, ___0____19813,
       ___0____19814, ___0____19815, ___0____19816, ___0____19818;
  wire ___0____19819, ___0____19820, ___0____19821, ___0____19822,
       ___0____19823, ___0____19824, ___0____19827, ___0____19828;
  wire ___0____19829, ___0____19830, ___0____19831, ___0____19832,
       ___0____19833, ___0____19836, ___0____19837, ___0____19838;
  wire ___0____19839, ___0____19840, ___0____19841, ___0____19842,
       ___0____19843, ___0____20709, ___0____20710, ___0____20711;
  wire ___0____20712, ___0____20713, ___0____20714, ___0____20716,
       ___0____20717, ___0____20718, ___0____20719, ___0____20720;
  wire ___0____20721, ___0____20722, ___0____20725, ___0____20726,
       ___0____20727, ___0____20728, ___0____20729, ___0____20730;
  wire ___0____20731, ___0____20734, ___0____20735, ___0____20736,
       ___0____20737, ___0____20738, ___0____20739, ___0____20740;
  wire ___0____20741, ___0____20744, ___0____20745, ___0____20746,
       ___0____20747, ___0____20748, ___0____20749, ___0____20750;
  wire ___0____20753, ___0____20754, ___0____20755, ___0____20756,
       ___0____20757, ___0____20758, ___0____20759, ___0____20760;
  wire ___0____20763, ___0____20764, ___0____20765, ___0____20766,
       ___0____20767, ___0____20768, ___0____20769, ___0____20772;
  wire ___0____20773, ___0____20774, ___0____20775, ___0____20776,
       ___0____20777, ___0____20778, ___0____21642, ___0____21643;
  wire ___0____21644, ___0____21645, ___0____21646, ___0____21647,
       ___0____21650, ___0____21651, ___0____21652, ___0____21653;
  wire ___0____21654, ___0____21655, ___0____21656, ___0____21659,
       ___0____21660, ___0____21661, ___0____21662, ___0____21663;
  wire ___0____21664, ___0____21665, ___0____21668, ___0____21669,
       ___0____21670, ___0____21671, ___0____21672, ___0____21673;
  wire ___0____21674, ___0____21677, ___0____21678, ___0____21679,
       ___0____21680, ___0____21681, ___0____21682, ___0____21683;
  wire ___0____21684, ___0____21687, ___0____21688, ___0____21689,
       ___0____21690, ___0____21691, ___0____21692, ___0____21693;
  wire ___0____21694, ___0____21697, ___0____21698, ___0____21699,
       ___0____21700, ___0____21701, ___0____21702, ___0____21703;
  wire ___0____21704, ___0____21706, ___0____21707, ___0____21708,
       ___0____21709, ___0____21710, ___0____22545, ___0____22546;
  wire ___0____22547, ___0____22548, ___0____22549, ___0____22550,
       ___0____22551, ___0____22552, ___0____22555, ___0____22556;
  wire ___0____22557, ___0____22558, ___0____22559, ___0____22560,
       ___0____22561, ___0____22562, ___0____22565, ___0____22566;
  wire ___0____22567, ___0____22568, ___0____22569, ___0____22570,
       ___0____22571, ___0____22574, ___0____22575, ___0____22576;
  wire ___0____22577, ___0____22578, ___0____22579, ___0____22580,
       ___0____22583, ___0____22584, ___0____22585, ___0____22586;
  wire ___0____22587, ___0____22588, ___0____22589, ___0____22590,
       ___0____22591, ___0____22592, ___0____22593, ___0____22594;
  wire ___0____22595, ___0____22596, ___0____22597, ___0____22598,
       ___0____22601, ___0____22602, ___0____22603, ___0____22604;
  wire ___0____22605, ___0____22606, ___0____22607, ___0____22609,
       ___0____22610, ___0____22611, ___0____22612, ___0____22613;
  wire ___0____22614, ___0____22615, ___0____22616, ___0____23446,
       ___0____23447, ___0____23448, ___0____23449, ___0____23450;
  wire ___0____23451, ___0____23452, ___0____23453, ___0____23456,
       ___0____23457, ___0____23458, ___0____23459, ___0____23460;
  wire ___0____23461, ___0____23462, ___0____23465, ___0____23466,
       ___0____23467, ___0____23468, ___0____23469, ___0____23470;
  wire ___0____23471, ___0____23474, ___0____23475, ___0____23476,
       ___0____23477, ___0____23478, ___0____23479, ___0____23480;
  wire ___0____23482, ___0____23483, ___0____23484, ___0____23485,
       ___0____23486, ___0____23487, ___0____23488, ___0____23491;
  wire ___0____23492, ___0____23493, ___0____23494, ___0____23495,
       ___0____23496, ___0____23497, ___0____23498, ___0____23501;
  wire ___0____23502, ___0____23503, ___0____23504, ___0____23505,
       ___0____23506, ___0____23507, ___0____23508, ___0____23510;
  wire ___0____23511, ___0____23512, ___0____23513, ___0____23514,
       ___0____23515, ___0____23516, ___0____24344, ___0____24345;
  wire ___0____24346, ___0____24347, ___0____24348, ___0____24349,
       ___0____24350, ___0____24353, ___0____24354, ___0____24355;
  wire ___0____24356, ___0____24357, ___0____24358, ___0____24359,
       ___0____24360, ___0____24363, ___0____24364, ___0____24365;
  wire ___0____24366, ___0____24367, ___0____24368, ___0____24369,
       ___0____24370, ___0____24373, ___0____24374, ___0____24375;
  wire ___0____24376, ___0____24377, ___0____24378, ___0____24379,
       ___0____24380, ___0____24383, ___0____24384, ___0____24385;
  wire ___0____24386, ___0____24387, ___0____24388, ___0____24389,
       ___0____24392, ___0____24393, ___0____24394, ___0____24395;
  wire ___0____24396, ___0____24397, ___0____24398, ___0____24399,
       ___0____24401, ___0____24402, ___0____24403, ___0____24404;
  wire ___0____24405, ___0____24406, ___0____24407, ___0____24408,
       ___0____24411, ___0____24412, ___0____24413, ___0____24414;
  wire ___0____24415, ___0____24416, ___0____24417, ___0____25282,
       ___0____25283, ___0____25284, ___0____25285, ___0____25286;
  wire ___0____25287, ___0____25288, ___0____25291, ___0____25292,
       ___0____25293, ___0____25294, ___0____25295, ___0____25296;
  wire ___0____25297, ___0____25298, ___0____25301, ___0____25302,
       ___0____25303, ___0____25304, ___0____25305, ___0____25306;
  wire ___0____25307, ___0____25308, ___0____25311, ___0____25312,
       ___0____25313, ___0____25314, ___0____25315, ___0____25316;
  wire ___0____25317, ___0____25320, ___0____25321, ___0____25322,
       ___0____25323, ___0____25324, ___0____25325, ___0____25326;
  wire ___0____25329, ___0____25330, ___0____25331, ___0____25332,
       ___0____25333, ___0____25334, ___0____25335, ___0____25336;
  wire ___0____25339, ___0____25340, ___0____25341, ___0____25342,
       ___0____25343, ___0____25344, ___0____25345, ___0____25348;
  wire ___0____25349, ___0____25350, ___0____25351, ___0____25352,
       ___0____25353, ___0____25354, ___0____25355, ___0_____27278;
  wire ___0_____27279, ___0_____27280, ___0_____27281, ___0_____27282,
       ___0_____27283, ___0_____27284, ___0_____27285, ___0_____27288;
  wire ___0_____27289, ___0_____27290, ___0_____27291, ___0_____27292,
       ___0_____27293, ___0_____27294, ___0_____27295, ___0_____27298;
  wire ___0_____27299, ___0_____27300, ___0_____27301, ___0_____27302,
       ___0_____27303, ___0_____27304, ___0_____27305, ___0_____27308;
  wire ___0_____27309, ___0_____27310, ___0_____27311, ___0_____27312,
       ___0_____27313, ___0_____27314, ___0_____27317, ___0_____27318;
  wire ___0_____27319, ___0_____27320, ___0_____27321, ___0_____27322,
       ___0_____27323, ___0_____27326, ___0_____27327, ___0_____27328;
  wire ___0_____27329, ___0_____27330, ___0_____27331, ___0_____27332,
       ___0_____27333, ___0_____27336, ___0_____27337, ___0_____27338;
  wire ___0_____27339, ___0_____27340, ___0_____27341, ___0_____27342,
       ___0_____27343, ___0_____27346, ___0_____27347, ___0_____27348;
  wire ___0_____27349, ___0_____27350, ___0_____27351, ___0_____27352,
       ___0_____27375, ___0_____27376, ___0_____27377, ___0_____27378;
  wire ___0_____27379, ___0_____27380, ___0_____27381, ___0_____27382,
       ___0_____27385, ___0_____27386, ___0_____27387, ___0_____27388;
  wire ___0_____27389, ___0_____27390, ___0_____27391, ___0_____27394,
       ___0_____27395, ___0_____27396, ___0_____27397, ___0_____27398;
  wire ___0_____27399, ___0_____27400, ___0_____27401, ___0_____27404,
       ___0_____27405, ___0_____27406, ___0_____27407, ___0_____27408;
  wire ___0_____27409, ___0_____27410, ___0_____27411, ___0_____27414,
       ___0_____27415, ___0_____27416, ___0_____27417, ___0_____27418;
  wire ___0_____27419, ___0_____27420, ___0_____27421, ___0_____27424,
       ___0_____27425, ___0_____27426, ___0_____27427, ___0_____27428;
  wire ___0_____27429, ___0_____27430, ___0_____27431, ___0_____27434,
       ___0_____27435, ___0_____27436, ___0_____27437, ___0_____27438;
  wire ___0_____27439, ___0_____27440, ___0_____27441, ___0_____27444,
       ___0_____27445, ___0_____27446, ___0_____27447, ___0_____27448;
  wire ___0_____27449, ___0_____27450, ___0_____27451, ___0_____27472,
       ___0_____27473, ___0_____27474, ___0_____27475, ___0_____27476;
  wire ___0_____27477, ___0_____27478, ___0_____27479, ___0_____27482,
       ___0_____27483, ___0_____27484, ___0_____27485, ___0_____27486;
  wire ___0_____27487, ___0_____27488, ___0_____27489, ___0_____27492,
       ___0_____27493, ___0_____27494, ___0_____27495, ___0_____27496;
  wire ___0_____27497, ___0_____27498, ___0_____27499, ___0_____27502,
       ___0_____27503, ___0_____27504, ___0_____27505, ___0_____27506;
  wire ___0_____27507, ___0_____27508, ___0_____27509, ___0_____27512,
       ___0_____27513, ___0_____27514, ___0_____27515, ___0_____27516;
  wire ___0_____27517, ___0_____27518, ___0_____27519, ___0_____27522,
       ___0_____27523, ___0_____27524, ___0_____27525, ___0_____27526;
  wire ___0_____27527, ___0_____27528, ___0_____27529, ___0_____27532,
       ___0_____27533, ___0_____27534, ___0_____27535, ___0_____27536;
  wire ___0_____27537, ___0_____27538, ___0_____27539, ___0_____27542,
       ___0_____27543, ___0_____27544, ___0_____27545, ___0_____27546;
  wire ___0_____27547, ___0_____27548, ___0_____27549, ___0_____27570,
       ___0_____27571, ___0_____27572, ___0_____27573, ___0_____27574;
  wire ___0_____27575, ___0_____27576, ___0_____27577, ___0_____27580,
       ___0_____27581, ___0_____27582, ___0_____27583, ___0_____27584;
  wire ___0_____27585, ___0_____27586, ___0_____27587, ___0_____27590,
       ___0_____27591, ___0_____27592, ___0_____27593, ___0_____27594;
  wire ___0_____27595, ___0_____27596, ___0_____27597, ___0_____27600,
       ___0_____27601, ___0_____27602, ___0_____27603, ___0_____27604;
  wire ___0_____27605, ___0_____27606, ___0_____27607, ___0_____27610,
       ___0_____27611, ___0_____27612, ___0_____27613, ___0_____27614;
  wire ___0_____27615, ___0_____27616, ___0_____27619, ___0_____27620,
       ___0_____27621, ___0_____27622, ___0_____27623, ___0_____27624;
  wire ___0_____27625, ___0_____27626, ___0_____27629, ___0_____27630,
       ___0_____27631, ___0_____27632, ___0_____27633, ___0_____27634;
  wire ___0_____27635, ___0_____27638, ___0_____27639, ___0_____27640,
       ___0_____27641, ___0_____27642, ___0_____27643, ___0_____27644;
  wire ___0_____27667, ___0_____27668, ___0_____27669, ___0_____27670,
       ___0_____27671, ___0_____27672, ___0_____27673, ___0_____27674;
  wire ___0_____27677, ___0_____27678, ___0_____27679, ___0_____27680,
       ___0_____27681, ___0_____27682, ___0_____27683, ___0_____27686;
  wire ___0_____27687, ___0_____27688, ___0_____27689, ___0_____27690,
       ___0_____27691, ___0_____27692, ___0_____27695, ___0_____27696;
  wire ___0_____27697, ___0_____27698, ___0_____27699, ___0_____27700,
       ___0_____27701, ___0_____27702, ___0_____27705, ___0_____27706;
  wire ___0_____27707, ___0_____27708, ___0_____27709, ___0_____27710,
       ___0_____27711, ___0_____27712, ___0_____27715, ___0_____27716;
  wire ___0_____27717, ___0_____27718, ___0_____27719, ___0_____27720,
       ___0_____27721, ___0_____27722, ___0_____27725, ___0_____27726;
  wire ___0_____27727, ___0_____27728, ___0_____27729, ___0_____27730,
       ___0_____27731, ___0_____27734, ___0_____27735, ___0_____27736;
  wire ___0_____27737, ___0_____27738, ___0_____27739, ___0_____27740,
       ___0_____27741, ___0_____27763, ___0_____27764, ___0_____27765;
  wire ___0_____27766, ___0_____27767, ___0_____27768, ___0_____27769,
       ___0_____27770, ___0_____27773, ___0_____27774, ___0_____27775;
  wire ___0_____27776, ___0_____27777, ___0_____27778, ___0_____27779,
       ___0_____27780, ___0_____27783, ___0_____27784, ___0_____27785;
  wire ___0_____27786, ___0_____27787, ___0_____27788, ___0_____27789,
       ___0_____27790, ___0_____27793, ___0_____27794, ___0_____27795;
  wire ___0_____27796, ___0_____27797, ___0_____27798, ___0_____27799,
       ___0_____27800, ___0_____27803, ___0_____27804, ___0_____27805;
  wire ___0_____27806, ___0_____27807, ___0_____27808, ___0_____27809,
       ___0_____27811, ___0_____27812, ___0_____27813, ___0_____27814;
  wire ___0_____27815, ___0_____27816, ___0_____27817, ___0_____27818,
       ___0_____27821, ___0_____27822, ___0_____27823, ___0_____27824;
  wire ___0_____27825, ___0_____27826, ___0_____27827, ___0_____27828,
       ___0_____27831, ___0_____27832, ___0_____27833, ___0_____27834;
  wire ___0_____27835, ___0_____27836, ___0_____27837, ___0_____27838,
       ___0_____27861, ___0_____27862, ___0_____27863, ___0_____27864;
  wire ___0_____27865, ___0_____27866, ___0_____27867, ___0_____27868,
       ___0_____27871, ___0_____27872, ___0_____27873, ___0_____27874;
  wire ___0_____27875, ___0_____27876, ___0_____27877, ___0_____27878,
       ___0_____27881, ___0_____27882, ___0_____27883, ___0_____27884;
  wire ___0_____27885, ___0_____27886, ___0_____27887, ___0_____27888,
       ___0_____27891, ___0_____27892, ___0_____27893, ___0_____27894;
  wire ___0_____27895, ___0_____27896, ___0_____27897, ___0_____27900,
       ___0_____27901, ___0_____27902, ___0_____27903, ___0_____27904;
  wire ___0_____27905, ___0_____27906, ___0_____27907, ___0_____27910,
       ___0_____27911, ___0_____27912, ___0_____27913, ___0_____27914;
  wire ___0_____27915, ___0_____27916, ___0_____27917, ___0_____27920,
       ___0_____27921, ___0_____27922, ___0_____27923, ___0_____27924;
  wire ___0_____27925, ___0_____27926, ___0_____27927, ___0_____27930,
       ___0_____27931, ___0_____27932, ___0_____27933, ___0_____27934;
  wire ___0_____27935, ___0_____27936, ___0_____27956, ___0_____27957,
       ___0_____27958, ___0_____27959, ___0_____27960, ___0_____27961;
  wire ___0_____27962, ___0_____27963, ___0_____27966, ___0_____27967,
       ___0_____27968, ___0_____27969, ___0_____27970, ___0_____27971;
  wire ___0_____27972, ___0_____27973, ___0_____27975, ___0_____27976,
       ___0_____27977, ___0_____27978, ___0_____27979, ___0_____27980;
  wire ___0_____27981, ___0_____27982, ___0_____27985, ___0_____27986,
       ___0_____27987, ___0_____27988, ___0_____27989, ___0_____27990;
  wire ___0_____27991, ___0_____27992, ___0_____27995, ___0_____27996,
       ___0_____27997, ___0_____27998, ___0_____27999, ___0_____28000;
  wire ___0_____28001, ___0_____28002, ___0_____28005, ___0_____28006,
       ___0_____28007, ___0_____28008, ___0_____28009, ___0_____28010;
  wire ___0_____28011, ___0_____28012, ___0_____28015, ___0_____28016,
       ___0_____28017, ___0_____28018, ___0_____28019, ___0_____28020;
  wire ___0_____28023, ___0_____28024, ___0_____28025, ___0_____28026,
       ___0_____28027, ___0_____28028, ___0_____28029, ___0_____28030;
  wire ___0009__27178, ___009, ___009__20707, ___009__22544,
       ___009__23445, ___009__24342, ___009__25280, ___009___27258;
  wire ___009___27259, ___009___27260, ___009___27261, ___009___27262,
       ___009___27263, ___009___27264, ___009___27265, ___09;
  wire ___09_, ___09_0__28051, ___09_0__28061, ___09_0__28071,
       ___09_0__28081, ___09_0__28091, ___09_0__28101, ___09_0__28111;
  wire ___09_0__28120, ___09_9__28060, ___09_9__28070, ___09_9__28080,
       ___09_9__28090, ___09_9__28100, ___09_9__28110, ___09_9__28119;
  wire ___09___19845, ___09___19846, ___09___19847, ___09___19848,
       ___09___19849, ___09___19850, ___09___19851, ___09___20781;
  wire ___09___20782, ___09___20783, ___09___20784, ___09___20785,
       ___09___20786, ___09___20787, ___09___20788, ___09___21712;
  wire ___09___21713, ___09___21714, ___09___21715, ___09___21716,
       ___09___21717, ___09___22618, ___09___22619, ___09___22620;
  wire ___09___22621, ___09___22622, ___09___22623, ___09___22624,
       ___09___23519, ___09___23520, ___09___23521, ___09___23522;
  wire ___09___23523, ___09___23524, ___09___23525, ___09___23526,
       ___09___24420, ___09___24421, ___09___24422, ___09___24423;
  wire ___09___24424, ___09___24425, ___09___24426, ___09___24427,
       ___09___25358, ___09___25359, ___09___25360, ___09___25361;
  wire ___09___25362, ___09___25363, ___09___25364, ___09___25365,
       ___09____28052, ___09____28053, ___09____28054, ___09____28055;
  wire ___09____28056, ___09____28057, ___09____28058, ___09____28059,
       ___09____28062, ___09____28063, ___09____28064, ___09____28065;
  wire ___09____28066, ___09____28067, ___09____28068, ___09____28069,
       ___09____28072, ___09____28073, ___09____28074, ___09____28075;
  wire ___09____28076, ___09____28077, ___09____28078, ___09____28079,
       ___09____28082, ___09____28083, ___09____28084, ___09____28085;
  wire ___09____28086, ___09____28087, ___09____28088, ___09____28089,
       ___09____28092, ___09____28093, ___09____28094, ___09____28095;
  wire ___09____28096, ___09____28097, ___09____28098, ___09____28099,
       ___09____28102, ___09____28103, ___09____28104, ___09____28105;
  wire ___09____28106, ___09____28107, ___09____28108, ___09____28109,
       ___09____28112, ___09____28113, ___09____28114, ___09____28115;
  wire ___09____28116, ___09____28117, ___09____28118, ___09____28121,
       ___09____28122, ___09____28123, ___09____28124, ___09____28125;
  wire ___09____28126, ___09____28127, ___9, ___9_, ___9_0,
       ___9_0__19698, ___9_0__19707, ___9_0__19717;
  wire ___9_0__19727, ___9_0__19737, ___9_0__19745, ___9_0__19755,
       ___9_0__20614, ___9_0__20624, ___9_0__20634, ___9_0__20644;
  wire ___9_0__20654, ___9_0__20663, ___9_0__20672, ___9_0__20682,
       ___9_0__21553, ___9_0__21561, ___9_0__21571, ___9_0__21580;
  wire ___9_0__21590, ___9_0__21599, ___9_0__21608, ___9_0__21617,
       ___9_0__22455, ___9_0__22465, ___9_0__22472, ___9_0__22481;
  wire ___9_0__22491, ___9_0__22500, ___9_0__22508, ___9_0__22517,
       ___9_0__23356, ___9_0__23366, ___9_0__23376, ___9_0__23386;
  wire ___9_0__23405, ___9_0__23413, ___9_0__24249, ___9_0__24257,
       ___9_0__24267, ___9_0__24276, ___9_0__24286, ___9_0__24296;
  wire ___9_0__24306, ___9_0__24316, ___9_0__25184, ___9_0__25194,
       ___9_0__25203, ___9_0__25211, ___9_0__25221, ___9_0__25231;
  wire ___9_0__25241, ___9_0__25251, ___9_0__26157, ___9_0__26167,
       ___9_0__26177, ___9_0__26187, ___9_0__26197, ___9_0__26207;
  wire ___9_0__26217, ___9_0__26227, ___9_9, ___9_9__19706,
       ___9_9__19716, ___9_9__19726, ___9_9__19736, ___9_9__19744;
  wire ___9_9__19754, ___9_9__20623, ___9_9__20633, ___9_9__20643,
       ___9_9__20653, ___9_9__20662, ___9_9__20671, ___9_9__20681;
  wire ___9_9__21560, ___9_9__21570, ___9_9__21579, ___9_9__21589,
       ___9_9__21598, ___9_9__21607, ___9_9__21616, ___9_9__21625;
  wire ___9_9__22464, ___9_9__22480, ___9_9__22490, ___9_9__22499,
       ___9_9__22507, ___9_9__22516, ___9_9__23365, ___9_9__23375;
  wire ___9_9__23385, ___9_9__23395, ___9_9__23404, ___9_9__23412,
       ___9_9__23422, ___9_9__24256, ___9_9__24266, ___9_9__24285;
  wire ___9_9__24295, ___9_9__24305, ___9_9__24315, ___9_9__24325,
       ___9_9__25193, ___9_9__25202, ___9_9__25210, ___9_9__25220;
  wire ___9_9__25230, ___9_9__25240, ___9_9__25250, ___9_9__25260,
       ___9_9__26166, ___9_9__26176, ___9_9__26186, ___9_9__26196;
  wire ___9_9__26206, ___9_9__26216, ___9_9__26226, ___9_9__26236,
       ___9__, ___9__18926, ___9__18930, ___9__18934;
  wire ___9__18942, ___9___18952, ___9___18953, ___9___18975,
       ___9___18976, ___9___18977, ___9___18978, ___9___18979;
  wire ___9___18980, ___9___18981, ___9___19030, ___9___19031,
       ___9___19032, ___9____19691, ___9____19692, ___9____19693;
  wire ___9____19694, ___9____19695, ___9____19696, ___9____19697,
       ___9____19699, ___9____19700, ___9____19701, ___9____19702;
  wire ___9____19703, ___9____19704, ___9____19705, ___9____19708,
       ___9____19709, ___9____19710, ___9____19711, ___9____19712;
  wire ___9____19713, ___9____19714, ___9____19715, ___9____19718,
       ___9____19719, ___9____19720, ___9____19721, ___9____19722;
  wire ___9____19723, ___9____19724, ___9____19725, ___9____19728,
       ___9____19729, ___9____19730, ___9____19731, ___9____19732;
  wire ___9____19733, ___9____19734, ___9____19735, ___9____19738,
       ___9____19739, ___9____19740, ___9____19741, ___9____19742;
  wire ___9____19743, ___9____19746, ___9____19747, ___9____19748,
       ___9____19749, ___9____19750, ___9____19751, ___9____19752;
  wire ___9____19753, ___9____19756, ___9____19757, ___9____19758,
       ___9____19759, ___9____19760, ___9____19761, ___9____19762;
  wire ___9____19763, ___9____20615, ___9____20616, ___9____20617,
       ___9____20618, ___9____20619, ___9____20620, ___9____20621;
  wire ___9____20622, ___9____20625, ___9____20626, ___9____20627,
       ___9____20628, ___9____20629, ___9____20630, ___9____20631;
  wire ___9____20632, ___9____20635, ___9____20636, ___9____20637,
       ___9____20638, ___9____20639, ___9____20640, ___9____20641;
  wire ___9____20642, ___9____20645, ___9____20646, ___9____20647,
       ___9____20648, ___9____20649, ___9____20650, ___9____20651;
  wire ___9____20652, ___9____20655, ___9____20656, ___9____20657,
       ___9____20658, ___9____20659, ___9____20660, ___9____20661;
  wire ___9____20664, ___9____20665, ___9____20666, ___9____20667,
       ___9____20668, ___9____20669, ___9____20670, ___9____20673;
  wire ___9____20674, ___9____20675, ___9____20676, ___9____20677,
       ___9____20678, ___9____20679, ___9____20680, ___9____20683;
  wire ___9____20684, ___9____20685, ___9____20686, ___9____20687,
       ___9____20688, ___9____20689, ___9____20690, ___9____21554;
  wire ___9____21555, ___9____21556, ___9____21557, ___9____21558,
       ___9____21559, ___9____21562, ___9____21563, ___9____21564;
  wire ___9____21565, ___9____21566, ___9____21567, ___9____21568,
       ___9____21569, ___9____21572, ___9____21573, ___9____21574;
  wire ___9____21575, ___9____21576, ___9____21577, ___9____21578,
       ___9____21581, ___9____21582, ___9____21583, ___9____21584;
  wire ___9____21585, ___9____21586, ___9____21587, ___9____21588,
       ___9____21591, ___9____21592, ___9____21593, ___9____21594;
  wire ___9____21595, ___9____21596, ___9____21597, ___9____21600,
       ___9____21601, ___9____21602, ___9____21603, ___9____21604;
  wire ___9____21605, ___9____21606, ___9____21609, ___9____21610,
       ___9____21611, ___9____21612, ___9____21613, ___9____21614;
  wire ___9____21615, ___9____21618, ___9____21619, ___9____21620,
       ___9____21621, ___9____21622, ___9____21623, ___9____21624;
  wire ___9____22456, ___9____22457, ___9____22458, ___9____22459,
       ___9____22460, ___9____22461, ___9____22462, ___9____22463;
  wire ___9____22466, ___9____22467, ___9____22468, ___9____22469,
       ___9____22470, ___9____22471, ___9____22473, ___9____22474;
  wire ___9____22475, ___9____22476, ___9____22477, ___9____22478,
       ___9____22479, ___9____22482, ___9____22483, ___9____22484;
  wire ___9____22485, ___9____22486, ___9____22487, ___9____22488,
       ___9____22489, ___9____22492, ___9____22493, ___9____22494;
  wire ___9____22495, ___9____22496, ___9____22497, ___9____22498,
       ___9____22501, ___9____22502, ___9____22503, ___9____22504;
  wire ___9____22505, ___9____22506, ___9____22509, ___9____22510,
       ___9____22511, ___9____22512, ___9____22513, ___9____22514;
  wire ___9____22515, ___9____22518, ___9____22519, ___9____22520,
       ___9____22521, ___9____22522, ___9____22523, ___9____22524;
  wire ___9____22525, ___9____23357, ___9____23358, ___9____23359,
       ___9____23360, ___9____23361, ___9____23362, ___9____23363;
  wire ___9____23364, ___9____23367, ___9____23368, ___9____23369,
       ___9____23370, ___9____23371, ___9____23372, ___9____23373;
  wire ___9____23374, ___9____23377, ___9____23378, ___9____23379,
       ___9____23380, ___9____23381, ___9____23382, ___9____23383;
  wire ___9____23384, ___9____23387, ___9____23388, ___9____23389,
       ___9____23390, ___9____23391, ___9____23392, ___9____23393;
  wire ___9____23394, ___9____23396, ___9____23397, ___9____23398,
       ___9____23399, ___9____23400, ___9____23401, ___9____23402;
  wire ___9____23403, ___9____23406, ___9____23407, ___9____23408,
       ___9____23409, ___9____23410, ___9____23411, ___9____23414;
  wire ___9____23415, ___9____23416, ___9____23417, ___9____23418,
       ___9____23419, ___9____23420, ___9____23421, ___9____23423;
  wire ___9____23424, ___9____23425, ___9____23426, ___9____24250,
       ___9____24251, ___9____24252, ___9____24253, ___9____24254;
  wire ___9____24255, ___9____24258, ___9____24259, ___9____24260,
       ___9____24261, ___9____24262, ___9____24263, ___9____24264;
  wire ___9____24265, ___9____24268, ___9____24269, ___9____24270,
       ___9____24271, ___9____24272, ___9____24273, ___9____24274;
  wire ___9____24275, ___9____24277, ___9____24278, ___9____24279,
       ___9____24280, ___9____24281, ___9____24282, ___9____24283;
  wire ___9____24284, ___9____24287, ___9____24288, ___9____24289,
       ___9____24290, ___9____24291, ___9____24292, ___9____24293;
  wire ___9____24294, ___9____24297, ___9____24298, ___9____24299,
       ___9____24300, ___9____24301, ___9____24302, ___9____24303;
  wire ___9____24304, ___9____24307, ___9____24308, ___9____24309,
       ___9____24310, ___9____24311, ___9____24312, ___9____24313;
  wire ___9____24314, ___9____24317, ___9____24318, ___9____24319,
       ___9____24320, ___9____24321, ___9____24322, ___9____24323;
  wire ___9____24324, ___9____25185, ___9____25186, ___9____25187,
       ___9____25188, ___9____25189, ___9____25190, ___9____25191;
  wire ___9____25192, ___9____25195, ___9____25196, ___9____25197,
       ___9____25198, ___9____25199, ___9____25200, ___9____25201;
  wire ___9____25204, ___9____25205, ___9____25206, ___9____25207,
       ___9____25208, ___9____25209, ___9____25212, ___9____25213;
  wire ___9____25214, ___9____25215, ___9____25216, ___9____25217,
       ___9____25218, ___9____25219, ___9____25222, ___9____25223;
  wire ___9____25224, ___9____25225, ___9____25226, ___9____25227,
       ___9____25228, ___9____25229, ___9____25232, ___9____25233;
  wire ___9____25234, ___9____25235, ___9____25236, ___9____25237,
       ___9____25238, ___9____25239, ___9____25242, ___9____25243;
  wire ___9____25244, ___9____25245, ___9____25246, ___9____25247,
       ___9____25248, ___9____25249, ___9____25252, ___9____25253;
  wire ___9____25254, ___9____25255, ___9____25256, ___9____25257,
       ___9____25258, ___9____25259, ___9____26158, ___9____26159;
  wire ___9____26160, ___9____26161, ___9____26162, ___9____26163,
       ___9____26164, ___9____26165, ___9____26168, ___9____26169;
  wire ___9____26170, ___9____26171, ___9____26172, ___9____26173,
       ___9____26174, ___9____26175, ___9____26178, ___9____26179;
  wire ___9____26180, ___9____26181, ___9____26182, ___9____26183,
       ___9____26184, ___9____26185, ___9____26188, ___9____26189;
  wire ___9____26190, ___9____26191, ___9____26192, ___9____26193,
       ___9____26194, ___9____26195, ___9____26198, ___9____26199;
  wire ___9____26200, ___9____26201, ___9____26202, ___9____26203,
       ___9____26204, ___9____26205, ___9____26208, ___9____26209;
  wire ___9____26210, ___9____26211, ___9____26212, ___9____26213,
       ___9____26214, ___9____26215, ___9____26218, ___9____26219;
  wire ___9____26220, ___9____26221, ___9____26222, ___9____26223,
       ___9____26224, ___9____26225, ___9____26228, ___9____26229;
  wire ___9____26230, ___9____26231, ___9____26232, ___9____26233,
       ___9____26234, ___9____26235, ___0090__27257, ___090;
  wire ___090__20780, ___090__21711, ___090__22617, ___090__23518,
       ___090__24419, ___090__25357, ___090___28043, ___090___28044;
  wire ___090___28045, ___090___28046, ___090___28047, ___090___28048,
       ___090___28049, ___90, ___90_, ___90___19686;
  wire ___90___19687, ___90___19688, ___90___19689, ___90___19690,
       ___90___20606, ___90___20607, ___90___20608, ___90___20609;
  wire ___90___20610, ___90___20611, ___90___20612, ___90___21544,
       ___90___21545, ___90___21546, ___90___21547, ___90___21548;
  wire ___90___21549, ___90___21550, ___90___21551, ___90___22447,
       ___90___22448, ___90___22449, ___90___22450, ___90___22451;
  wire ___90___22452, ___90___22453, ___90___23347, ___90___23348,
       ___90___23349, ___90___23350, ___90___23351, ___90___23352;
  wire ___90___23353, ___90___23354, ___90___24242, ___90___24243,
       ___90___24244, ___90___24245, ___90___24246, ___90___24247;
  wire ___90___25175, ___90___25176, ___90___25177, ___90___25178,
       ___90___25179, ___90___25180, ___90___25181, ___90___25182;
  wire ___90___26148, ___90___26149, ___90___26150, ___90___26151,
       ___90___26152, ___90___26153, ___90___26154, ___90___26155;
  wire ___0099__27266, ___099, ___099__20789, ___099__21718,
       ___099__22625, ___099__23527, ___099__24428, ___099__25366;
  wire ___099___28129, ___099___28130, ___099___28131, ___099___28132,
       ___099___28133, ___099___28134, ___099___28135, ___099___28136;
  wire ___99, ___99_, ___99___19764, ___99___19765, ___99___19766,
       ___99___19767, ___99___19768, ___99___19769;
  wire ___99___19770, ___99___20691, ___99___20692, ___99___20693,
       ___99___20694, ___99___20695, ___99___20696, ___99___20697;
  wire ___99___21626, ___99___21627, ___99___21628, ___99___21629,
       ___99___21630, ___99___21631, ___99___22527, ___99___22528;
  wire ___99___22529, ___99___22530, ___99___22531, ___99___22532,
       ___99___22533, ___99___22534, ___99___23428, ___99___23429;
  wire ___99___23430, ___99___23431, ___99___23432, ___99___23433,
       ___99___23434, ___99___23435, ___99___24327, ___99___24328;
  wire ___99___24329, ___99___24330, ___99___24331, ___99___25262,
       ___99___25263, ___99___25264, ___99___25265, ___99___25266;
  wire ___99___25267, ___99___25268, ___99___25269, ___99___26238,
       ___99___26239, ___99___26240, ___99___26241, ___99___26242;
  wire ___99___26243, ___99___26244, ___99___26245, ___0900__28042,
       ___900, ___900__20605, ___900__21543, ___900__22446;
  wire ___900__23346, ___900__24241, ___900__25174, ___900__26147,
       ___0909__28050, ___909, ___909__20613, ___909__21552;
  wire ___909__22454, ___909__23355, ___909__24248, ___909__25183,
       ___909__26156, ___0990__28128, ___990, ___990__22526;
  wire ___990__23427, ___990__24326, ___990__25261, ___990__26237,
       ___0999__28137, ___999, ___999__20698, ___999__21632;
  wire ___999__22535, ___999__23436, ___999__24332, ___999__25270,
       ___999__26246, ____, ____0, ____00;
  wire ____000__28138, ____000__29083, ____000__30000, ____000__30906,
       ____000__31808, ____000__32751, ____000__33674, ____000__34531;
  wire ____00__19114, ____00__19205, ____00__19302, ____00__19399,
       ____00__19496, ____00__19592, ____00__19852, ____00__19947;
  wire ____00__20040, ____00__20136, ____00__20226, ____00__20324,
       ____00__20420, ____00__20510, ____00__20790, ____00__20886;
  wire ____00__20982, ____00__21075, ____00__21166, ____00__21260,
       ____00__21355, ____00__21446, ____00__21719, ____00__21811;
  wire ____00__21904, ____00__21985, ____00__22081, ____00__22172,
       ____00__22261, ____00__22356, ____00__22626, ____00__22718;
  wire ____00__22807, ____00__22895, ____00__22989, ____00__23084,
       ____00__23171, ____00__23259, ____00__23528, ____00__23618;
  wire ____00__23802, ____00__23887, ____00__23974, ____00__24063,
       ____00__24429, ____00__24518, ____00__24608, ____00__24701;
  wire ____00__24792, ____00__24886, ____00__24984, ____00__25080,
       ____00__25367, ____00__25464, ____00__25558, ____00__25655;
  wire ____00__25751, ____00__25850, ____00__25948, ____00__26047,
       ____00___28139, ____00___28140, ____00___28141, ____00___28142;
  wire ____00___28143, ____00___28144, ____00___28145, ____00___28146,
       ____00___29084, ____00___29085, ____00___29086, ____00___29087;
  wire ____00___29088, ____00___29089, ____00___29090, ____00___30001,
       ____00___30002, ____00___30003, ____00___30004, ____00___30005;
  wire ____00___30006, ____00___30007, ____00___30907, ____00___30908,
       ____00___30909, ____00___30910, ____00___30911, ____00___30912;
  wire ____00___30913, ____00___30914, ____00___31809, ____00___31810,
       ____00___31811, ____00___31812, ____00___31813, ____00___31814;
  wire ____00___32752, ____00___32753, ____00___32754, ____00___32755,
       ____00___32756, ____00___32757, ____00___32758, ____00___32759;
  wire ____00___33675, ____00___33676, ____00___33677, ____00___33678,
       ____00___33679, ____00___33680, ____00___33681, ____00___33682;
  wire ____00___34532, ____00___34533, ____00___34534, ____00___34535,
       ____00___34536, ____00___34537, ____00___34538, ____00___34539;
  wire ____0_, ____0_0__28148, ____0_0__28158, ____0_0__28168,
       ____0_0__28177, ____0_0__28186, ____0_0__28196, ____0_0__28206;
  wire ____0_0__28215, ____0_0__29092, ____0_0__29101, ____0_0__29119,
       ____0_0__29128, ____0_0__29138, ____0_0__29146, ____0_0__29156;
  wire ____0_0__30009, ____0_0__30018, ____0_0__30028, ____0_0__30037,
       ____0_0__30047, ____0_0__30056, ____0_0__30064, ____0_0__30074;
  wire ____0_0__30916, ____0_0__30924, ____0_0__30932, ____0_0__30942,
       ____0_0__30952, ____0_0__30962, ____0_0__30972, ____0_0__30979;
  wire ____0_0__31824, ____0_0__31833, ____0_0__31842, ____0_0__31851,
       ____0_0__31861, ____0_0__31871, ____0_0__32761, ____0_0__32770;
  wire ____0_0__32780, ____0_0__32790, ____0_0__32800, ____0_0__32810,
       ____0_0__32820, ____0_0__32830, ____0_0__33684, ____0_0__33693;
  wire ____0_0__33702, ____0_0__33712, ____0_0__33722, ____0_0__33732,
       ____0_0__33741, ____0_0__34541, ____0_0__34550, ____0_0__34560;
  wire ____0_0__34570, ____0_0__34580, ____0_0__34588, ____0_0__34598,
       ____0_0__34608, ____0_9__28157, ____0_9__28167, ____0_9__28185;
  wire ____0_9__28195, ____0_9__28205, ____0_9__28214, ____0_9__28224,
       ____0_9__29100, ____0_9__29109, ____0_9__29118, ____0_9__29127;
  wire ____0_9__29137, ____0_9__29145, ____0_9__29155, ____0_9__29165,
       ____0_9__30017, ____0_9__30027, ____0_9__30036, ____0_9__30046;
  wire ____0_9__30055, ____0_9__30063, ____0_9__30073, ____0_9__30083,
       ____0_9__30923, ____0_9__30931, ____0_9__30941, ____0_9__30951;
  wire ____0_9__30961, ____0_9__30971, ____0_9__30987, ____0_9__31823,
       ____0_9__31832, ____0_9__31841, ____0_9__31850, ____0_9__31860;
  wire ____0_9__31870, ____0_9__31880, ____0_9__31889, ____0_9__32769,
       ____0_9__32779, ____0_9__32789, ____0_9__32799, ____0_9__32809;
  wire ____0_9__32819, ____0_9__32829, ____0_9__32839, ____0_9__33692,
       ____0_9__33701, ____0_9__33711, ____0_9__33721, ____0_9__33731;
  wire ____0_9__33740, ____0_9__33749, ____0_9__33758, ____0_9__34549,
       ____0_9__34559, ____0_9__34569, ____0_9__34579, ____0_9__34587;
  wire ____0_9__34597, ____0_9__34607, ____0_9__34617, ____0__18959,
       ____0__18967, ____0__18989, ____0__18997, ____0__19007;
  wire ____0__19016, ____0__19046, ____0___19054, ____0___19055,
       ____0___19056, ____0___19057, ____0___19058, ____0___19059;
  wire ____0___19115, ____0___19116, ____0___19117, ____0___19118,
       ____0___19119, ____0___19120, ____0___19121, ____0___19122;
  wire ____0___19206, ____0___19207, ____0___19208, ____0___19209,
       ____0___19210, ____0___19211, ____0___19212, ____0___19213;
  wire ____0___19303, ____0___19304, ____0___19305, ____0___19306,
       ____0___19307, ____0___19308, ____0___19309, ____0___19310;
  wire ____0___19400, ____0___19401, ____0___19402, ____0___19403,
       ____0___19404, ____0___19405, ____0___19406, ____0___19407;
  wire ____0___19497, ____0___19498, ____0___19499, ____0___19500,
       ____0___19501, ____0___19502, ____0___19503, ____0___19504;
  wire ____0___19593, ____0___19594, ____0___19595, ____0___19596,
       ____0___19597, ____0___19598, ____0___19599, ____0___19600;
  wire ____0___19853, ____0___19854, ____0___19855, ____0___19856,
       ____0___19857, ____0___19858, ____0___19859, ____0___19860;
  wire ____0___19948, ____0___19949, ____0___19950, ____0___19951,
       ____0___19952, ____0___19953, ____0___19954, ____0___20041;
  wire ____0___20042, ____0___20043, ____0___20044, ____0___20045,
       ____0___20046, ____0___20047, ____0___20137, ____0___20138;
  wire ____0___20139, ____0___20140, ____0___20141, ____0___20142,
       ____0___20143, ____0___20144, ____0___20227, ____0___20228;
  wire ____0___20229, ____0___20230, ____0___20231, ____0___20232,
       ____0___20233, ____0___20234, ____0___20325, ____0___20326;
  wire ____0___20327, ____0___20328, ____0___20329, ____0___20330,
       ____0___20421, ____0___20422, ____0___20423, ____0___20424;
  wire ____0___20425, ____0___20426, ____0___20427, ____0___20511,
       ____0___20512, ____0___20513, ____0___20514, ____0___20515;
  wire ____0___20516, ____0___20517, ____0___20518, ____0___20791,
       ____0___20792, ____0___20793, ____0___20794, ____0___20795;
  wire ____0___20796, ____0___20797, ____0___20887, ____0___20888,
       ____0___20889, ____0___20890, ____0___20891, ____0___20892;
  wire ____0___20893, ____0___20983, ____0___20984, ____0___20985,
       ____0___20986, ____0___20987, ____0___20988, ____0___20989;
  wire ____0___21076, ____0___21077, ____0___21078, ____0___21079,
       ____0___21080, ____0___21081, ____0___21082, ____0___21083;
  wire ____0___21167, ____0___21168, ____0___21169, ____0___21170,
       ____0___21171, ____0___21172, ____0___21261, ____0___21262;
  wire ____0___21263, ____0___21264, ____0___21265, ____0___21266,
       ____0___21267, ____0___21268, ____0___21356, ____0___21357;
  wire ____0___21358, ____0___21359, ____0___21360, ____0___21361,
       ____0___21362, ____0___21363, ____0___21447, ____0___21448;
  wire ____0___21449, ____0___21450, ____0___21451, ____0___21452,
       ____0___21453, ____0___21720, ____0___21721, ____0___21722;
  wire ____0___21723, ____0___21724, ____0___21725, ____0___21726,
       ____0___21727, ____0___21812, ____0___21813, ____0___21814;
  wire ____0___21815, ____0___21816, ____0___21817, ____0___21818,
       ____0___21819, ____0___21905, ____0___21906, ____0___21907;
  wire ____0___21908, ____0___21909, ____0___21910, ____0___21911,
       ____0___21912, ____0___21986, ____0___21987, ____0___21988;
  wire ____0___21989, ____0___21990, ____0___21991, ____0___21992,
       ____0___21993, ____0___22082, ____0___22083, ____0___22084;
  wire ____0___22085, ____0___22086, ____0___22087, ____0___22173,
       ____0___22174, ____0___22175, ____0___22176, ____0___22177;
  wire ____0___22178, ____0___22179, ____0___22180, ____0___22262,
       ____0___22263, ____0___22264, ____0___22265, ____0___22266;
  wire ____0___22267, ____0___22268, ____0___22269, ____0___22357,
       ____0___22358, ____0___22359, ____0___22360, ____0___22361;
  wire ____0___22362, ____0___22363, ____0___22364, ____0___22627,
       ____0___22628, ____0___22629, ____0___22630, ____0___22631;
  wire ____0___22632, ____0___22633, ____0___22719, ____0___22720,
       ____0___22721, ____0___22722, ____0___22723, ____0___22808;
  wire ____0___22809, ____0___22810, ____0___22811, ____0___22812,
       ____0___22813, ____0___22814, ____0___22896, ____0___22897;
  wire ____0___22898, ____0___22899, ____0___22900, ____0___22901,
       ____0___22902, ____0___22903, ____0___22990, ____0___22991;
  wire ____0___22992, ____0___22993, ____0___22994, ____0___22995,
       ____0___22996, ____0___22997, ____0___23085, ____0___23086;
  wire ____0___23087, ____0___23088, ____0___23089, ____0___23090,
       ____0___23172, ____0___23173, ____0___23174, ____0___23175;
  wire ____0___23176, ____0___23177, ____0___23178, ____0___23179,
       ____0___23260, ____0___23261, ____0___23262, ____0___23263;
  wire ____0___23264, ____0___23265, ____0___23266, ____0___23529,
       ____0___23530, ____0___23531, ____0___23532, ____0___23533;
  wire ____0___23534, ____0___23619, ____0___23620, ____0___23621,
       ____0___23622, ____0___23623, ____0___23624, ____0___23625;
  wire ____0___23626, ____0___23712, ____0___23713, ____0___23714,
       ____0___23715, ____0___23716, ____0___23717, ____0___23718;
  wire ____0___23719, ____0___23803, ____0___23804, ____0___23805,
       ____0___23806, ____0___23807, ____0___23808, ____0___23809;
  wire ____0___23810, ____0___23888, ____0___23889, ____0___23890,
       ____0___23891, ____0___23892, ____0___23893, ____0___23894;
  wire ____0___23895, ____0___23975, ____0___23976, ____0___23977,
       ____0___23978, ____0___23979, ____0___23980, ____0___23981;
  wire ____0___23982, ____0___24064, ____0___24065, ____0___24066,
       ____0___24067, ____0___24068, ____0___24069, ____0___24070;
  wire ____0___24155, ____0___24156, ____0___24157, ____0___24158,
       ____0___24159, ____0___24160, ____0___24161, ____0___24430;
  wire ____0___24431, ____0___24432, ____0___24433, ____0___24434,
       ____0___24435, ____0___24519, ____0___24520, ____0___24521;
  wire ____0___24522, ____0___24523, ____0___24609, ____0___24610,
       ____0___24611, ____0___24612, ____0___24613, ____0___24614;
  wire ____0___24702, ____0___24703, ____0___24704, ____0___24705,
       ____0___24706, ____0___24707, ____0___24708, ____0___24793;
  wire ____0___24794, ____0___24795, ____0___24796, ____0___24797,
       ____0___24798, ____0___24799, ____0___24800, ____0___24887;
  wire ____0___24888, ____0___24889, ____0___24890, ____0___24891,
       ____0___24892, ____0___24893, ____0___24894, ____0___24985;
  wire ____0___24986, ____0___24987, ____0___24988, ____0___24989,
       ____0___24990, ____0___24991, ____0___25081, ____0___25082;
  wire ____0___25083, ____0___25084, ____0___25085, ____0___25086,
       ____0___25087, ____0___25088, ____0___25368, ____0___25369;
  wire ____0___25370, ____0___25371, ____0___25372, ____0___25373,
       ____0___25374, ____0___25375, ____0___25465, ____0___25466;
  wire ____0___25467, ____0___25468, ____0___25469, ____0___25470,
       ____0___25471, ____0___25559, ____0___25560, ____0___25561;
  wire ____0___25562, ____0___25563, ____0___25564, ____0___25565,
       ____0___25566, ____0___25656, ____0___25657, ____0___25658;
  wire ____0___25659, ____0___25660, ____0___25661, ____0___25662,
       ____0___25663, ____0___25752, ____0___25753, ____0___25754;
  wire ____0___25755, ____0___25756, ____0___25757, ____0___25758,
       ____0___25759, ____0___25851, ____0___25852, ____0___25853;
  wire ____0___25854, ____0___25855, ____0___25856, ____0___25857,
       ____0___25858, ____0___25949, ____0___25950, ____0___25951;
  wire ____0___25952, ____0___25953, ____0___25954, ____0___25955,
       ____0___26048, ____0___26049, ____0___26050, ____0___26051;
  wire ____0___26052, ____0___26053, ____0___26054, ____0___26055,
       ____0____28149, ____0____28150, ____0____28151, ____0____28152;
  wire ____0____28153, ____0____28154, ____0____28155, ____0____28156,
       ____0____28159, ____0____28160, ____0____28161, ____0____28162;
  wire ____0____28163, ____0____28164, ____0____28165, ____0____28166,
       ____0____28169, ____0____28170, ____0____28171, ____0____28172;
  wire ____0____28173, ____0____28174, ____0____28175, ____0____28176,
       ____0____28178, ____0____28179, ____0____28180, ____0____28181;
  wire ____0____28182, ____0____28183, ____0____28184, ____0____28187,
       ____0____28188, ____0____28189, ____0____28190, ____0____28191;
  wire ____0____28192, ____0____28193, ____0____28194, ____0____28197,
       ____0____28198, ____0____28199, ____0____28200, ____0____28201;
  wire ____0____28202, ____0____28203, ____0____28204, ____0____28207,
       ____0____28208, ____0____28209, ____0____28210, ____0____28211;
  wire ____0____28212, ____0____28213, ____0____28216, ____0____28217,
       ____0____28218, ____0____28219, ____0____28220, ____0____28221;
  wire ____0____28222, ____0____28223, ____0____29093, ____0____29094,
       ____0____29095, ____0____29096, ____0____29097, ____0____29098;
  wire ____0____29099, ____0____29102, ____0____29103, ____0____29104,
       ____0____29105, ____0____29106, ____0____29107, ____0____29108;
  wire ____0____29110, ____0____29111, ____0____29112, ____0____29113,
       ____0____29114, ____0____29115, ____0____29116, ____0____29117;
  wire ____0____29120, ____0____29121, ____0____29122, ____0____29123,
       ____0____29124, ____0____29125, ____0____29126, ____0____29129;
  wire ____0____29130, ____0____29131, ____0____29132, ____0____29133,
       ____0____29134, ____0____29135, ____0____29136, ____0____29139;
  wire ____0____29140, ____0____29141, ____0____29142, ____0____29143,
       ____0____29144, ____0____29147, ____0____29148, ____0____29149;
  wire ____0____29150, ____0____29151, ____0____29152, ____0____29153,
       ____0____29154, ____0____29157, ____0____29158, ____0____29159;
  wire ____0____29160, ____0____29161, ____0____29162, ____0____29163,
       ____0____29164, ____0____30010, ____0____30011, ____0____30012;
  wire ____0____30013, ____0____30014, ____0____30015, ____0____30016,
       ____0____30019, ____0____30020, ____0____30021, ____0____30022;
  wire ____0____30023, ____0____30024, ____0____30025, ____0____30026,
       ____0____30029, ____0____30030, ____0____30031, ____0____30032;
  wire ____0____30033, ____0____30034, ____0____30035, ____0____30038,
       ____0____30039, ____0____30040, ____0____30041, ____0____30042;
  wire ____0____30043, ____0____30044, ____0____30045, ____0____30048,
       ____0____30049, ____0____30050, ____0____30051, ____0____30052;
  wire ____0____30053, ____0____30054, ____0____30057, ____0____30058,
       ____0____30059, ____0____30060, ____0____30061, ____0____30062;
  wire ____0____30065, ____0____30066, ____0____30067, ____0____30068,
       ____0____30069, ____0____30070, ____0____30071, ____0____30072;
  wire ____0____30075, ____0____30076, ____0____30077, ____0____30078,
       ____0____30079, ____0____30080, ____0____30081, ____0____30082;
  wire ____0____30917, ____0____30918, ____0____30919, ____0____30920,
       ____0____30921, ____0____30922, ____0____30925, ____0____30926;
  wire ____0____30927, ____0____30928, ____0____30929, ____0____30930,
       ____0____30933, ____0____30934, ____0____30935, ____0____30936;
  wire ____0____30937, ____0____30938, ____0____30939, ____0____30940,
       ____0____30943, ____0____30944, ____0____30945, ____0____30946;
  wire ____0____30947, ____0____30948, ____0____30949, ____0____30950,
       ____0____30953, ____0____30954, ____0____30955, ____0____30956;
  wire ____0____30957, ____0____30958, ____0____30959, ____0____30960,
       ____0____30963, ____0____30964, ____0____30965, ____0____30966;
  wire ____0____30967, ____0____30968, ____0____30969, ____0____30970,
       ____0____30973, ____0____30974, ____0____30975, ____0____30976;
  wire ____0____30977, ____0____30978, ____0____30980, ____0____30981,
       ____0____30982, ____0____30983, ____0____30984, ____0____30985;
  wire ____0____30986, ____0____31816, ____0____31817, ____0____31818,
       ____0____31819, ____0____31820, ____0____31821, ____0____31822;
  wire ____0____31825, ____0____31826, ____0____31827, ____0____31828,
       ____0____31829, ____0____31830, ____0____31831, ____0____31834;
  wire ____0____31835, ____0____31836, ____0____31837, ____0____31838,
       ____0____31839, ____0____31840, ____0____31843, ____0____31844;
  wire ____0____31845, ____0____31846, ____0____31847, ____0____31848,
       ____0____31849, ____0____31852, ____0____31853, ____0____31854;
  wire ____0____31855, ____0____31856, ____0____31857, ____0____31858,
       ____0____31859, ____0____31862, ____0____31863, ____0____31864;
  wire ____0____31865, ____0____31866, ____0____31867, ____0____31868,
       ____0____31869, ____0____31872, ____0____31873, ____0____31874;
  wire ____0____31875, ____0____31876, ____0____31877, ____0____31878,
       ____0____31879, ____0____31881, ____0____31882, ____0____31883;
  wire ____0____31884, ____0____31885, ____0____31886, ____0____31887,
       ____0____31888, ____0____32762, ____0____32763, ____0____32764;
  wire ____0____32765, ____0____32766, ____0____32767, ____0____32768,
       ____0____32771, ____0____32772, ____0____32773, ____0____32774;
  wire ____0____32775, ____0____32776, ____0____32777, ____0____32778,
       ____0____32781, ____0____32782, ____0____32783, ____0____32784;
  wire ____0____32785, ____0____32786, ____0____32787, ____0____32788,
       ____0____32791, ____0____32792, ____0____32793, ____0____32794;
  wire ____0____32795, ____0____32796, ____0____32797, ____0____32798,
       ____0____32801, ____0____32802, ____0____32803, ____0____32804;
  wire ____0____32805, ____0____32806, ____0____32807, ____0____32808,
       ____0____32811, ____0____32812, ____0____32813, ____0____32814;
  wire ____0____32815, ____0____32816, ____0____32817, ____0____32818,
       ____0____32821, ____0____32822, ____0____32823, ____0____32824;
  wire ____0____32825, ____0____32826, ____0____32827, ____0____32828,
       ____0____32831, ____0____32832, ____0____32833, ____0____32834;
  wire ____0____32835, ____0____32836, ____0____32837, ____0____32838,
       ____0____33685, ____0____33686, ____0____33687, ____0____33688;
  wire ____0____33689, ____0____33690, ____0____33691, ____0____33694,
       ____0____33695, ____0____33696, ____0____33697, ____0____33698;
  wire ____0____33699, ____0____33700, ____0____33703, ____0____33704,
       ____0____33705, ____0____33706, ____0____33707, ____0____33708;
  wire ____0____33709, ____0____33710, ____0____33713, ____0____33714,
       ____0____33715, ____0____33716, ____0____33717, ____0____33718;
  wire ____0____33719, ____0____33720, ____0____33723, ____0____33724,
       ____0____33725, ____0____33726, ____0____33727, ____0____33728;
  wire ____0____33729, ____0____33730, ____0____33733, ____0____33734,
       ____0____33735, ____0____33736, ____0____33737, ____0____33738;
  wire ____0____33739, ____0____33742, ____0____33743, ____0____33744,
       ____0____33745, ____0____33746, ____0____33747, ____0____33748;
  wire ____0____33750, ____0____33751, ____0____33752, ____0____33753,
       ____0____33754, ____0____33755, ____0____33756, ____0____33757;
  wire ____0____34542, ____0____34543, ____0____34544, ____0____34545,
       ____0____34546, ____0____34547, ____0____34548, ____0____34551;
  wire ____0____34552, ____0____34553, ____0____34554, ____0____34555,
       ____0____34556, ____0____34557, ____0____34558, ____0____34561;
  wire ____0____34562, ____0____34563, ____0____34564, ____0____34565,
       ____0____34566, ____0____34567, ____0____34568, ____0____34571;
  wire ____0____34572, ____0____34573, ____0____34574, ____0____34575,
       ____0____34576, ____0____34577, ____0____34578, ____0____34581;
  wire ____0____34582, ____0____34583, ____0____34584, ____0____34585,
       ____0____34586, ____0____34589, ____0____34590, ____0____34591;
  wire ____0____34592, ____0____34593, ____0____34594, ____0____34595,
       ____0____34596, ____0____34599, ____0____34600, ____0____34601;
  wire ____0____34602, ____0____34603, ____0____34604, ____0____34605,
       ____0____34606, ____0____34609, ____0____34610, ____0____34611;
  wire ____0____34612, ____0____34613, ____0____34614, ____0____34615,
       ____0____34616, ____0____________0_, ____0____________0___18645,
       ____0____________9_;
  wire ____0____________9___18654, ____0_____________0_,
       ____0_____________0___18655, ____0______________,
       ____0_______________, ____0________________18589,
       ____0________________18590, ____0________________18591;
  wire ____0________________18592, ____0________________18593,
       ____0________________18594, ____0________________18595,
       ____0________________18646, ____0________________18647,
       ____0________________18648, ____0________________18649;
  wire ____0________________18650, ____0________________18651,
       ____0________________18652, ____0________________18653,
       ____0_________________18596, ____0_________________18656,
       ____0_________________18657, ____0_________________18658;
  wire ____0_________________18659, ____009__28147, ____009__29091,
       ____009__30008, ____009__30915, ____009__31815, ____009__32760,
       ____009__33683;
  wire ____009__34540, ____09, ____09__19123, ____09__19214,
       ____09__19311, ____09__19408, ____09__19505, ____09__19601;
  wire ____09__19861, ____09__19955, ____09__20048, ____09__20145,
       ____09__20235, ____09__20331, ____09__20428, ____09__20519;
  wire ____09__20798, ____09__20894, ____09__20990, ____09__21084,
       ____09__21269, ____09__21364, ____09__21454, ____09__21728;
  wire ____09__21820, ____09__21913, ____09__21994, ____09__22088,
       ____09__22181, ____09__22270, ____09__22365, ____09__22634;
  wire ____09__22724, ____09__22815, ____09__22904, ____09__22998,
       ____09__23091, ____09__23180, ____09__23267, ____09__23535;
  wire ____09__23627, ____09__23896, ____09__23983, ____09__24071,
       ____09__24162, ____09__24436, ____09__24524, ____09__24615;
  wire ____09__24709, ____09__24801, ____09__24895, ____09__24992,
       ____09__25089, ____09__25376, ____09__25567, ____09__25664;
  wire ____09__25760, ____09__25859, ____09__25956, ____09__26056,
       ____09___28226, ____09___28227, ____09___28228, ____09___28229;
  wire ____09___28230, ____09___28231, ____09___28232, ____09___28233,
       ____09___29167, ____09___29168, ____09___29169, ____09___29170;
  wire ____09___29171, ____09___29172, ____09___29173, ____09___29174,
       ____09___30085, ____09___30086, ____09___30087, ____09___30088;
  wire ____09___30089, ____09___30090, ____09___30091, ____09___30092,
       ____09___30989, ____09___30990, ____09___30991, ____09___30992;
  wire ____09___30993, ____09___30994, ____09___30995, ____09___31891,
       ____09___31892, ____09___31893, ____09___31894, ____09___31895;
  wire ____09___31896, ____09___31897, ____09___31898, ____09___32841,
       ____09___32842, ____09___32843, ____09___32844, ____09___32845;
  wire ____09___32846, ____09___32847, ____09___33760, ____09___33761,
       ____09___33762, ____09___33763, ____09___33764, ____09___33765;
  wire ____09___33766, ____09___33767, ____09___34619, ____09___34620,
       ____09___34621, ____09___34622, ____09___34623, ____09___34624;
  wire ____09___34625, ____09___34626, ____9, ____9_, ____9_0__29002,
       ____9_0__29012, ____9_0__29019, ____9_0__29029;
  wire ____9_0__29038, ____9_0__29047, ____9_0__29055, ____9_0__29064,
       ____9_0__29920, ____9_0__29930, ____9_0__29940, ____9_0__29950;
  wire ____9_0__29960, ____9_0__29970, ____9_0__29980, ____9_0__30828,
       ____9_0__30838, ____9_0__30846, ____9_0__30854, ____9_0__30872;
  wire ____9_0__30881, ____9_0__30889, ____9_0__31733, ____9_0__31743,
       ____9_0__31750, ____9_0__31767, ____9_0__31782, ____9_0__31792;
  wire ____9_0__32665, ____9_0__32675, ____9_0__32685, ____9_0__32695,
       ____9_0__32705, ____9_0__32715, ____9_0__32725, ____9_0__33587;
  wire ____9_0__33597, ____9_0__33606, ____9_0__33616, ____9_0__33626,
       ____9_0__33635, ____9_0__33644, ____9_0__33654, ____9_9__29011;
  wire ____9_9__29018, ____9_9__29028, ____9_9__29037, ____9_9__29046,
       ____9_9__29054, ____9_9__29063, ____9_9__29072, ____9_9__29919;
  wire ____9_9__29929, ____9_9__29939, ____9_9__29949, ____9_9__29959,
       ____9_9__29969, ____9_9__29979, ____9_9__29989, ____9_9__30837;
  wire ____9_9__30845, ____9_9__30863, ____9_9__30871, ____9_9__30880,
       ____9_9__30888, ____9_9__30897, ____9_9__31742, ____9_9__31749;
  wire ____9_9__31757, ____9_9__31766, ____9_9__31774, ____9_9__31781,
       ____9_9__31791, ____9_9__31801, ____9_9__32674, ____9_9__32684;
  wire ____9_9__32694, ____9_9__32704, ____9_9__32714, ____9_9__32724,
       ____9_9__32734, ____9_9__32742, ____9_9__33596, ____9_9__33605;
  wire ____9_9__33615, ____9_9__33625, ____9_9__33634, ____9_9__33643,
       ____9_9__33653, ____9_9__33663, ____9_9__34520, ____9__18949;
  wire ____9__18955, ____9__18996, ____9__19006, ____9__19015,
       ____9__19035, ____9__19036, ____9__19041, ____9__19045;
  wire ____9___19053, ____9___19106, ____9___19107, ____9___19108,
       ____9___19109, ____9___19110, ____9___19111, ____9___19112;
  wire ____9___19197, ____9___19198, ____9___19199, ____9___19200,
       ____9___19201, ____9___19202, ____9___19203, ____9___19293;
  wire ____9___19294, ____9___19295, ____9___19296, ____9___19297,
       ____9___19298, ____9___19299, ____9___19300, ____9___19391;
  wire ____9___19392, ____9___19393, ____9___19394, ____9___19395,
       ____9___19396, ____9___19397, ____9___19488, ____9___19489;
  wire ____9___19490, ____9___19491, ____9___19492, ____9___19493,
       ____9___19494, ____9___19495, ____9___19583, ____9___19584;
  wire ____9___19585, ____9___19586, ____9___19587, ____9___19588,
       ____9___19589, ____9___19590, ____9___19678, ____9___19679;
  wire ____9___19680, ____9___19681, ____9___19682, ____9___19683,
       ____9___19684, ____9___19938, ____9___19939, ____9___19940;
  wire ____9___19941, ____9___19942, ____9___19943, ____9___19944,
       ____9___19945, ____9___20032, ____9___20033, ____9___20034;
  wire ____9___20035, ____9___20036, ____9___20037, ____9___20038,
       ____9___20127, ____9___20128, ____9___20129, ____9___20130;
  wire ____9___20131, ____9___20132, ____9___20133, ____9___20134,
       ____9___20218, ____9___20219, ____9___20220, ____9___20221;
  wire ____9___20222, ____9___20223, ____9___20224, ____9___20315,
       ____9___20316, ____9___20317, ____9___20318, ____9___20319;
  wire ____9___20320, ____9___20321, ____9___20322, ____9___20411,
       ____9___20412, ____9___20413, ____9___20414, ____9___20415;
  wire ____9___20416, ____9___20417, ____9___20418, ____9___20501,
       ____9___20502, ____9___20503, ____9___20504, ____9___20505;
  wire ____9___20506, ____9___20507, ____9___20508, ____9___20596,
       ____9___20597, ____9___20598, ____9___20599, ____9___20600;
  wire ____9___20601, ____9___20602, ____9___20603, ____9___20877,
       ____9___20878, ____9___20879, ____9___20880, ____9___20881;
  wire ____9___20882, ____9___20883, ____9___20884, ____9___20973,
       ____9___20974, ____9___20975, ____9___20976, ____9___20977;
  wire ____9___20978, ____9___20979, ____9___20980, ____9___21067,
       ____9___21068, ____9___21069, ____9___21070, ____9___21071;
  wire ____9___21072, ____9___21073, ____9___21157, ____9___21158,
       ____9___21159, ____9___21160, ____9___21161, ____9___21162;
  wire ____9___21163, ____9___21164, ____9___21251, ____9___21252,
       ____9___21253, ____9___21254, ____9___21255, ____9___21256;
  wire ____9___21257, ____9___21258, ____9___21346, ____9___21347,
       ____9___21348, ____9___21349, ____9___21350, ____9___21351;
  wire ____9___21352, ____9___21353, ____9___21439, ____9___21440,
       ____9___21441, ____9___21442, ____9___21443, ____9___21444;
  wire ____9___21534, ____9___21535, ____9___21536, ____9___21537,
       ____9___21538, ____9___21539, ____9___21540, ____9___21541;
  wire ____9___21802, ____9___21803, ____9___21804, ____9___21805,
       ____9___21806, ____9___21807, ____9___21808, ____9___21809;
  wire ____9___21896, ____9___21897, ____9___21898, ____9___21899,
       ____9___21900, ____9___21901, ____9___21902, ____9___21980;
  wire ____9___21981, ____9___21982, ____9___21983, ____9___21984,
       ____9___22072, ____9___22073, ____9___22074, ____9___22075;
  wire ____9___22076, ____9___22077, ____9___22078, ____9___22079,
       ____9___22163, ____9___22164, ____9___22165, ____9___22166;
  wire ____9___22167, ____9___22168, ____9___22169, ____9___22170,
       ____9___22252, ____9___22253, ____9___22254, ____9___22255;
  wire ____9___22256, ____9___22257, ____9___22258, ____9___22259,
       ____9___22347, ____9___22348, ____9___22349, ____9___22350;
  wire ____9___22351, ____9___22352, ____9___22353, ____9___22354,
       ____9___22437, ____9___22438, ____9___22439, ____9___22440;
  wire ____9___22441, ____9___22442, ____9___22443, ____9___22444,
       ____9___22710, ____9___22711, ____9___22712, ____9___22713;
  wire ____9___22714, ____9___22715, ____9___22716, ____9___22799,
       ____9___22800, ____9___22801, ____9___22802, ____9___22803;
  wire ____9___22804, ____9___22805, ____9___22886, ____9___22887,
       ____9___22888, ____9___22889, ____9___22890, ____9___22891;
  wire ____9___22892, ____9___22893, ____9___22982, ____9___22983,
       ____9___22984, ____9___22985, ____9___22986, ____9___22987;
  wire ____9___22988, ____9___23075, ____9___23076, ____9___23077,
       ____9___23078, ____9___23079, ____9___23080, ____9___23081;
  wire ____9___23082, ____9___23163, ____9___23164, ____9___23165,
       ____9___23166, ____9___23167, ____9___23168, ____9___23169;
  wire ____9___23251, ____9___23252, ____9___23253, ____9___23254,
       ____9___23255, ____9___23256, ____9___23257, ____9___23337;
  wire ____9___23338, ____9___23339, ____9___23340, ____9___23341,
       ____9___23342, ____9___23343, ____9___23344, ____9___23610;
  wire ____9___23611, ____9___23612, ____9___23613, ____9___23614,
       ____9___23615, ____9___23616, ____9___23705, ____9___23706;
  wire ____9___23707, ____9___23708, ____9___23709, ____9___23710,
       ____9___23793, ____9___23794, ____9___23795, ____9___23796;
  wire ____9___23797, ____9___23798, ____9___23799, ____9___23800,
       ____9___23878, ____9___23879, ____9___23880, ____9___23881;
  wire ____9___23882, ____9___23883, ____9___23884, ____9___23885,
       ____9___23966, ____9___23967, ____9___23968, ____9___23969;
  wire ____9___23970, ____9___23971, ____9___23972, ____9___23973,
       ____9___24054, ____9___24055, ____9___24056, ____9___24057;
  wire ____9___24058, ____9___24059, ____9___24060, ____9___24061,
       ____9___24148, ____9___24149, ____9___24150, ____9___24151;
  wire ____9___24152, ____9___24153, ____9___24154, ____9___24236,
       ____9___24237, ____9___24238, ____9___24239, ____9___24240;
  wire ____9___24509, ____9___24510, ____9___24511, ____9___24512,
       ____9___24513, ____9___24514, ____9___24515, ____9___24516;
  wire ____9___24599, ____9___24600, ____9___24601, ____9___24602,
       ____9___24603, ____9___24604, ____9___24605, ____9___24606;
  wire ____9___24694, ____9___24695, ____9___24696, ____9___24697,
       ____9___24698, ____9___24699, ____9___24783, ____9___24784;
  wire ____9___24785, ____9___24786, ____9___24787, ____9___24788,
       ____9___24789, ____9___24790, ____9___24878, ____9___24879;
  wire ____9___24880, ____9___24881, ____9___24882, ____9___24883,
       ____9___24884, ____9___24885, ____9___24975, ____9___24976;
  wire ____9___24977, ____9___24978, ____9___24979, ____9___24980,
       ____9___24981, ____9___24982, ____9___25072, ____9___25073;
  wire ____9___25074, ____9___25075, ____9___25076, ____9___25077,
       ____9___25078, ____9___25166, ____9___25167, ____9___25168;
  wire ____9___25169, ____9___25170, ____9___25171, ____9___25172,
       ____9___25456, ____9___25457, ____9___25458, ____9___25459;
  wire ____9___25460, ____9___25461, ____9___25462, ____9___25550,
       ____9___25551, ____9___25552, ____9___25553, ____9___25554;
  wire ____9___25555, ____9___25556, ____9___25646, ____9___25647,
       ____9___25648, ____9___25649, ____9___25650, ____9___25651;
  wire ____9___25652, ____9___25653, ____9___25742, ____9___25743,
       ____9___25744, ____9___25745, ____9___25746, ____9___25747;
  wire ____9___25748, ____9___25749, ____9___25841, ____9___25842,
       ____9___25843, ____9___25844, ____9___25845, ____9___25846;
  wire ____9___25847, ____9___25848, ____9___25940, ____9___25941,
       ____9___25942, ____9___25943, ____9___25944, ____9___25945;
  wire ____9___25946, ____9___26038, ____9___26039, ____9___26040,
       ____9___26041, ____9___26042, ____9___26043, ____9___26044;
  wire ____9___26045, ____9___26138, ____9___26139, ____9___26140,
       ____9___26141, ____9___26142, ____9___26143, ____9___26144;
  wire ____9___26145, ____9____29003, ____9____29004, ____9____29005,
       ____9____29006, ____9____29007, ____9____29008, ____9____29009;
  wire ____9____29010, ____9____29013, ____9____29014, ____9____29015,
       ____9____29016, ____9____29017, ____9____29020, ____9____29021;
  wire ____9____29022, ____9____29023, ____9____29024, ____9____29025,
       ____9____29026, ____9____29027, ____9____29030, ____9____29031;
  wire ____9____29032, ____9____29033, ____9____29034, ____9____29035,
       ____9____29036, ____9____29039, ____9____29040, ____9____29041;
  wire ____9____29042, ____9____29043, ____9____29044, ____9____29045,
       ____9____29048, ____9____29049, ____9____29050, ____9____29051;
  wire ____9____29052, ____9____29053, ____9____29056, ____9____29057,
       ____9____29058, ____9____29059, ____9____29060, ____9____29061;
  wire ____9____29062, ____9____29065, ____9____29066, ____9____29067,
       ____9____29068, ____9____29069, ____9____29070, ____9____29071;
  wire ____9____29911, ____9____29912, ____9____29913, ____9____29914,
       ____9____29915, ____9____29916, ____9____29917, ____9____29918;
  wire ____9____29921, ____9____29922, ____9____29923, ____9____29924,
       ____9____29925, ____9____29926, ____9____29927, ____9____29928;
  wire ____9____29931, ____9____29932, ____9____29933, ____9____29934,
       ____9____29935, ____9____29936, ____9____29937, ____9____29938;
  wire ____9____29941, ____9____29942, ____9____29943, ____9____29944,
       ____9____29945, ____9____29946, ____9____29947, ____9____29948;
  wire ____9____29951, ____9____29952, ____9____29953, ____9____29954,
       ____9____29955, ____9____29956, ____9____29957, ____9____29958;
  wire ____9____29961, ____9____29962, ____9____29963, ____9____29964,
       ____9____29965, ____9____29966, ____9____29967, ____9____29968;
  wire ____9____29971, ____9____29972, ____9____29973, ____9____29974,
       ____9____29975, ____9____29976, ____9____29977, ____9____29978;
  wire ____9____29981, ____9____29982, ____9____29983, ____9____29984,
       ____9____29985, ____9____29986, ____9____29987, ____9____29988;
  wire ____9____30829, ____9____30830, ____9____30831, ____9____30832,
       ____9____30833, ____9____30834, ____9____30835, ____9____30836;
  wire ____9____30839, ____9____30840, ____9____30841, ____9____30842,
       ____9____30843, ____9____30844, ____9____30847, ____9____30848;
  wire ____9____30849, ____9____30850, ____9____30851, ____9____30852,
       ____9____30853, ____9____30855, ____9____30856, ____9____30857;
  wire ____9____30858, ____9____30859, ____9____30860, ____9____30861,
       ____9____30862, ____9____30864, ____9____30865, ____9____30866;
  wire ____9____30867, ____9____30868, ____9____30869, ____9____30870,
       ____9____30873, ____9____30874, ____9____30875, ____9____30876;
  wire ____9____30877, ____9____30878, ____9____30879, ____9____30882,
       ____9____30883, ____9____30884, ____9____30885, ____9____30886;
  wire ____9____30887, ____9____30890, ____9____30891, ____9____30892,
       ____9____30893, ____9____30894, ____9____30895, ____9____30896;
  wire ____9____31734, ____9____31735, ____9____31736, ____9____31737,
       ____9____31738, ____9____31739, ____9____31740, ____9____31741;
  wire ____9____31744, ____9____31745, ____9____31746, ____9____31747,
       ____9____31748, ____9____31751, ____9____31752, ____9____31753;
  wire ____9____31754, ____9____31755, ____9____31756, ____9____31758,
       ____9____31759, ____9____31760, ____9____31761, ____9____31762;
  wire ____9____31763, ____9____31764, ____9____31765, ____9____31768,
       ____9____31769, ____9____31770, ____9____31771, ____9____31772;
  wire ____9____31773, ____9____31775, ____9____31776, ____9____31777,
       ____9____31778, ____9____31779, ____9____31780, ____9____31783;
  wire ____9____31784, ____9____31785, ____9____31786, ____9____31787,
       ____9____31788, ____9____31789, ____9____31790, ____9____31793;
  wire ____9____31794, ____9____31795, ____9____31796, ____9____31797,
       ____9____31798, ____9____31799, ____9____31800, ____9____32666;
  wire ____9____32667, ____9____32668, ____9____32669, ____9____32670,
       ____9____32671, ____9____32672, ____9____32673, ____9____32676;
  wire ____9____32677, ____9____32678, ____9____32679, ____9____32680,
       ____9____32681, ____9____32682, ____9____32683, ____9____32686;
  wire ____9____32687, ____9____32688, ____9____32689, ____9____32690,
       ____9____32691, ____9____32692, ____9____32693, ____9____32696;
  wire ____9____32697, ____9____32698, ____9____32699, ____9____32700,
       ____9____32701, ____9____32702, ____9____32703, ____9____32706;
  wire ____9____32707, ____9____32708, ____9____32709, ____9____32710,
       ____9____32711, ____9____32712, ____9____32713, ____9____32716;
  wire ____9____32717, ____9____32718, ____9____32719, ____9____32720,
       ____9____32721, ____9____32722, ____9____32723, ____9____32726;
  wire ____9____32727, ____9____32728, ____9____32729, ____9____32730,
       ____9____32731, ____9____32732, ____9____32733, ____9____32735;
  wire ____9____32736, ____9____32737, ____9____32738, ____9____32739,
       ____9____32740, ____9____32741, ____9____33588, ____9____33589;
  wire ____9____33590, ____9____33591, ____9____33592, ____9____33593,
       ____9____33594, ____9____33595, ____9____33598, ____9____33599;
  wire ____9____33600, ____9____33601, ____9____33602, ____9____33603,
       ____9____33604, ____9____33607, ____9____33608, ____9____33609;
  wire ____9____33610, ____9____33611, ____9____33612, ____9____33613,
       ____9____33614, ____9____33617, ____9____33618, ____9____33619;
  wire ____9____33620, ____9____33621, ____9____33622, ____9____33623,
       ____9____33624, ____9____33627, ____9____33628, ____9____33629;
  wire ____9____33630, ____9____33631, ____9____33632, ____9____33633,
       ____9____33636, ____9____33637, ____9____33638, ____9____33639;
  wire ____9____33640, ____9____33641, ____9____33642, ____9____33645,
       ____9____33646, ____9____33647, ____9____33648, ____9____33649;
  wire ____9____33650, ____9____33651, ____9____33652, ____9____33655,
       ____9____33656, ____9____33657, ____9____33658, ____9____33659;
  wire ____9____33660, ____9____33661, ____9____33662, ____9____34518,
       ____9____34519, ____090__28225, ____090__29166, ____090__30084;
  wire ____090__30988, ____090__31890, ____090__32840, ____090__33759,
       ____090__34618, ____90, ____90__19196, ____90__19292;
  wire ____90__19390, ____90__19487, ____90__19582, ____90__19677,
       ____90__19937, ____90__20031, ____90__20126, ____90__20217;
  wire ____90__20314, ____90__20410, ____90__20500, ____90__20595,
       ____90__20876, ____90__20972, ____90__21066, ____90__21156;
  wire ____90__21250, ____90__21345, ____90__21438, ____90__21533,
       ____90__21801, ____90__21895, ____90__22071, ____90__22346;
  wire ____90__22436, ____90__22709, ____90__22798, ____90__22885,
       ____90__22981, ____90__23074, ____90__23162, ____90__23250;
  wire ____90__23336, ____90__23609, ____90__23704, ____90__23792,
       ____90__23877, ____90__23965, ____90__24053, ____90__24235;
  wire ____90__24508, ____90__24598, ____90__24693, ____90__24782,
       ____90__24877, ____90__24974, ____90__25071, ____90__25165;
  wire ____90__25455, ____90__25549, ____90__25645, ____90__25741,
       ____90__25840, ____90__25939, ____90__26037, ____90__26137;
  wire ____90___28993, ____90___28994, ____90___28995, ____90___28996,
       ____90___28997, ____90___28998, ____90___28999, ____90___29000;
  wire ____90___29902, ____90___29903, ____90___29904, ____90___29905,
       ____90___29906, ____90___29907, ____90___29908, ____90___29909;
  wire ____90___30821, ____90___30822, ____90___30823, ____90___30824,
       ____90___30825, ____90___30826, ____90___31725, ____90___31726;
  wire ____90___31727, ____90___31728, ____90___31729, ____90___31730,
       ____90___31731, ____90___32657, ____90___32658, ____90___32659;
  wire ____90___32660, ____90___32661, ____90___32662, ____90___32663,
       ____90___33579, ____90___33580, ____90___33581, ____90___33582;
  wire ____90___33583, ____90___33584, ____90___33585, ____099__28234,
       ____099__29175, ____099__30093, ____099__30996, ____099__31899;
  wire ____099__32848, ____099__33768, ____099__34627, ____99,
       ____99__19113, ____99__19204, ____99__19301, ____99__19398;
  wire ____99__19591, ____99__19685, ____99__19946, ____99__20039,
       ____99__20135, ____99__20225, ____99__20323, ____99__20419;
  wire ____99__20509, ____99__20604, ____99__20885, ____99__20981,
       ____99__21074, ____99__21165, ____99__21259, ____99__21354;
  wire ____99__21445, ____99__21542, ____99__21810, ____99__21903,
       ____99__22080, ____99__22171, ____99__22260, ____99__22355;
  wire ____99__22445, ____99__22717, ____99__22806, ____99__22894,
       ____99__23083, ____99__23170, ____99__23258, ____99__23345;
  wire ____99__23617, ____99__23711, ____99__23801, ____99__23886,
       ____99__24062, ____99__24517, ____99__24607, ____99__24700;
  wire ____99__24791, ____99__24983, ____99__25079, ____99__25173,
       ____99__25463, ____99__25557, ____99__25654, ____99__25750;
  wire ____99__25849, ____99__25947, ____99__26046, ____99__26146,
       ____99___29074, ____99___29075, ____99___29076, ____99___29077;
  wire ____99___29078, ____99___29079, ____99___29080, ____99___29081,
       ____99___29991, ____99___29992, ____99___29993, ____99___29994;
  wire ____99___29995, ____99___29996, ____99___29997, ____99___29998,
       ____99___30898, ____99___30899, ____99___30900, ____99___30901;
  wire ____99___30902, ____99___30903, ____99___30904, ____99___31802,
       ____99___31803, ____99___31804, ____99___31805, ____99___31806;
  wire ____99___32744, ____99___32745, ____99___32746, ____99___32747,
       ____99___32748, ____99___32749, ____99___33665, ____99___33666;
  wire ____99___33667, ____99___33668, ____99___33669, ____99___33670,
       ____99___33671, ____99___33672, ____99___34522, ____99___34523;
  wire ____99___34524, ____99___34525, ____99___34526, ____99___34527,
       ____99___34528, ____99___34529, ____99___35108, ____900__28992;
  wire ____900__29901, ____900__30820, ____900__31724, ____900__32656,
       ____909__29001, ____909__29910, ____909__30827, ____909__31732;
  wire ____909__32664, ____909__33586, ____990__29073, ____990__29990,
       ____990__32743, ____990__33664, ____990__34521, ____999__29082;
  wire ____999__29999, ____999__30905, ____999__31807, ____999__32750,
       ____999__33673, ____999__34530, _____, _____0;
  wire _____00__28235, _____00__28331, _____00__28425, _____00__28523,
       _____00__28616, _____00__28705, _____00__28800, _____00__28898;
  wire _____00__29176, _____00__29265, _____00__29356, _____00__29446,
       _____00__29532, _____00__29615, _____00__29710, _____00__29803;
  wire _____00__30094, _____00__30178, _____00__30274, _____00__30364,
       _____00__30456, _____00__30545, _____00__30632, _____00__30726;
  wire _____00__30997, _____00__31093, _____00__31183, _____00__31269,
       _____00__31354, _____00__31446, _____00__31536, _____00__31632;
  wire _____00__31900, _____00__31997, _____00__32096, _____00__32194,
       _____00__32292, _____00__32386, _____00__32569, _____00__32849;
  wire _____00__32936, _____00__33029, _____00__33127, _____00__33220,
       _____00__33310, _____00__33401, _____00__33488, _____00__33769;
  wire _____00__33865, _____00__33954, _____00__34045, _____00__34144,
       _____00__34238, _____00__34333, _____00__34421, _____00__34628;
  wire _____00__34728, _____00__34828, _____00__34928, _____00__35028,
       _____0__19068, _____0__19086, _____0__19096, _____0__19124;
  wire _____0__19134, _____0__19144, _____0__19153, _____0__19163,
       _____0__19170, _____0__19187, _____0__19215, _____0__19225;
  wire _____0__19234, _____0__19243, _____0__19252, _____0__19262,
       _____0__19272, _____0__19282, _____0__19312, _____0__19321;
  wire _____0__19331, _____0__19341, _____0__19351, _____0__19361,
       _____0__19371, _____0__19380, _____0__19409, _____0__19419;
  wire _____0__19429, _____0__19439, _____0__19449, _____0__19468,
       _____0__19477, _____0__19506, _____0__19516, _____0__19525;
  wire _____0__19534, _____0__19552, _____0__19562, _____0__19572,
       _____0__19602, _____0__19612, _____0__19622, _____0__19639;
  wire _____0__19649, _____0__19659, _____0__19669, _____0__19862,
       _____0__19872, _____0__19882, _____0__19892, _____0__19909;
  wire _____0__19918, _____0__19927, _____0__19956, _____0__19966,
       _____0__19975, _____0__19985, _____0__19992, _____0__20002;
  wire _____0__20012, _____0__20021, _____0__20049, _____0__20059,
       _____0__20069, _____0__20079, _____0__20088, _____0__20097;
  wire _____0__20107, _____0__20116, _____0__20146, _____0__20156,
       _____0__20181, _____0__20189, _____0__20198, _____0__20207;
  wire _____0__20245, _____0__20254, _____0__20264, _____0__20274,
       _____0__20284, _____0__20294, _____0__20304, _____0__20332;
  wire _____0__20342, _____0__20352, _____0__20362, _____0__20372,
       _____0__20382, _____0__20392, _____0__20402, _____0__20429;
  wire _____0__20439, _____0__20456, _____0__20465, _____0__20474,
       _____0__20484, _____0__20492, _____0__20520, _____0__20530;
  wire _____0__20540, _____0__20549, _____0__20558, _____0__20567,
       _____0__20576, _____0__20585, _____0__20799, _____0__20807;
  wire _____0__20817, _____0__20827, _____0__20837, _____0__20847,
       _____0__20857, _____0__20866, _____0__20895, _____0__20904;
  wire _____0__20913, _____0__20923, _____0__20933, _____0__20942,
       _____0__20952, _____0__20962, _____0__20991, _____0__21001;
  wire _____0__21010, _____0__21020, _____0__21030, _____0__21046,
       _____0__21056, _____0__21085, _____0__21103, _____0__21120;
  wire _____0__21130, _____0__21140, _____0__21147, _____0__21173,
       _____0__21183, _____0__21191, _____0__21200, _____0__21210;
  wire _____0__21220, _____0__21230, _____0__21240, _____0__21270,
       _____0__21279, _____0__21288, _____0__21298, _____0__21308;
  wire _____0__21317, _____0__21327, _____0__21335, _____0__21365,
       _____0__21374, _____0__21384, _____0__21393, _____0__21401;
  wire _____0__21410, _____0__21419, _____0__21429, _____0__21455,
       _____0__21465, _____0__21475, _____0__21485, _____0__21494;
  wire _____0__21504, _____0__21514, _____0__21523, _____0__21729,
       _____0__21739, _____0__21749, _____0__21757, _____0__21763;
  wire _____0__21773, _____0__21783, _____0__21821, _____0__21831,
       _____0__21840, _____0__21849, _____0__21859, _____0__21876;
  wire _____0__21885, _____0__21914, _____0__21924, _____0__21934,
       _____0__21940, _____0__21948, _____0__21962, _____0__21971;
  wire _____0__21995, _____0__22005, _____0__22014, _____0__22023,
       _____0__22033, _____0__22043, _____0__22053, _____0__22063;
  wire _____0__22089, _____0__22099, _____0__22108, _____0__22118,
       _____0__22128, _____0__22138, _____0__22148, _____0__22157;
  wire _____0__22182, _____0__22192, _____0__22200, _____0__22206,
       _____0__22216, _____0__22224, _____0__22234, _____0__22242;
  wire _____0__22271, _____0__22281, _____0__22291, _____0__22300,
       _____0__22310, _____0__22319, _____0__22327, _____0__22337;
  wire _____0__22366, _____0__22375, _____0__22384, _____0__22400,
       _____0__22417, _____0__22427, _____0__22635, _____0__22644;
  wire _____0__22653, _____0__22670, _____0__22680, _____0__22690,
       _____0__22700, _____0__22725, _____0__22734, _____0__22744;
  wire _____0__22754, _____0__22764, _____0__22772, _____0__22780,
       _____0__22790, _____0__22816, _____0__22826, _____0__22833;
  wire _____0__22848, _____0__22855, _____0__22865, _____0__22875,
       _____0__22905, _____0__22914, _____0__22924, _____0__22934;
  wire _____0__22952, _____0__22962, _____0__22999, _____0__23009,
       _____0__23018, _____0__23028, _____0__23038, _____0__23056;
  wire _____0__23065, _____0__23092, _____0__23108, _____0__23115,
       _____0__23125, _____0__23134, _____0__23143, _____0__23152;
  wire _____0__23181, _____0__23190, _____0__23199, _____0__23208,
       _____0__23215, _____0__23223, _____0__23231, _____0__23241;
  wire _____0__23268, _____0__23276, _____0__23286, _____0__23294,
       _____0__23303, _____0__23312, _____0__23317, _____0__23326;
  wire _____0__23536, _____0__23545, _____0__23555, _____0__23572,
       _____0__23582, _____0__23591, _____0__23601, _____0__23628;
  wire _____0__23638, _____0__23656, _____0__23666, _____0__23675,
       _____0__23685, _____0__23695, _____0__23720, _____0__23728;
  wire _____0__23737, _____0__23747, _____0__23756, _____0__23765,
       _____0__23775, _____0__23785, _____0__23811, _____0__23821;
  wire _____0__23828, _____0__23837, _____0__23850, _____0__23860,
       _____0__23897, _____0__23915, _____0__23925, _____0__23933;
  wire _____0__23942, _____0__23950, _____0__23958, _____0__23992,
       _____0__23999, _____0__24008, _____0__24018, _____0__24027;
  wire _____0__24035, _____0__24044, _____0__24072, _____0__24082,
       _____0__24092, _____0__24102, _____0__24120, _____0__24130;
  wire _____0__24140, _____0__24163, _____0__24173, _____0__24182,
       _____0__24190, _____0__24199, _____0__24209, _____0__24219;
  wire _____0__24227, _____0__24437, _____0__24447, _____0__24456,
       _____0__24465, _____0__24473, _____0__24481, _____0__24491;
  wire _____0__24499, _____0__24525, _____0__24534, _____0__24541,
       _____0__24551, _____0__24560, _____0__24570, _____0__24579;
  wire _____0__24588, _____0__24616, _____0__24626, _____0__24636,
       _____0__24646, _____0__24656, _____0__24666, _____0__24676;
  wire _____0__24684, _____0__24710, _____0__24720, _____0__24729,
       _____0__24739, _____0__24746, _____0__24756, _____0__24764;
  wire _____0__24772, _____0__24809, _____0__24819, _____0__24829,
       _____0__24848, _____0__24867, _____0__24896, _____0__24906;
  wire _____0__24916, _____0__24926, _____0__24936, _____0__24946,
       _____0__24956, _____0__24965, _____0__24993, _____0__25002;
  wire _____0__25012, _____0__25022, _____0__25032, _____0__25041,
       _____0__25051, _____0__25061, _____0__25090, _____0__25109;
  wire _____0__25119, _____0__25127, _____0__25136, _____0__25146,
       _____0__25156, _____0__25377, _____0__25387, _____0__25397;
  wire _____0__25406, _____0__25416, _____0__25426, _____0__25436,
       _____0__25446, _____0__25472, _____0__25482, _____0__25492;
  wire _____0__25501, _____0__25511, _____0__25520, _____0__25529,
       _____0__25539, _____0__25568, _____0__25578, _____0__25588;
  wire _____0__25597, _____0__25607, _____0__25616, _____0__25625,
       _____0__25635, _____0__25665, _____0__25675, _____0__25685;
  wire _____0__25694, _____0__25703, _____0__25712, _____0__25721,
       _____0__25731, _____0__25770, _____0__25780, _____0__25790;
  wire _____0__25800, _____0__25810, _____0__25820, _____0__25830,
       _____0__25860, _____0__25870, _____0__25880, _____0__25890;
  wire _____0__25899, _____0__25909, _____0__25919, _____0__25929,
       _____0__25957, _____0__25967, _____0__25977, _____0__25987;
  wire _____0__25997, _____0__26007, _____0__26017, _____0__26027,
       _____0__26057, _____0__26067, _____0__26077, _____0__26087;
  wire _____0__26097, _____0__26107, _____0__26117, _____0__26127,
       _____0___28236, _____0___28237, _____0___28238, _____0___28239;
  wire _____0___28240, _____0___28241, _____0___28242, _____0___28332,
       _____0___28333, _____0___28334, _____0___28335, _____0___28336;
  wire _____0___28337, _____0___28338, _____0___28426, _____0___28427,
       _____0___28428, _____0___28429, _____0___28430, _____0___28431;
  wire _____0___28432, _____0___28433, _____0___28524, _____0___28525,
       _____0___28526, _____0___28527, _____0___28528, _____0___28529;
  wire _____0___28530, _____0___28617, _____0___28618, _____0___28619,
       _____0___28620, _____0___28621, _____0___28622, _____0___28623;
  wire _____0___28706, _____0___28707, _____0___28708, _____0___28709,
       _____0___28710, _____0___28711, _____0___28712, _____0___28801;
  wire _____0___28802, _____0___28803, _____0___28804, _____0___28805,
       _____0___28806, _____0___28807, _____0___28808, _____0___28899;
  wire _____0___28900, _____0___28901, _____0___28902, _____0___28903,
       _____0___28904, _____0___28905, _____0___29177, _____0___29178;
  wire _____0___29179, _____0___29180, _____0___29181, _____0___29182,
       _____0___29183, _____0___29184, _____0___29266, _____0___29267;
  wire _____0___29268, _____0___29269, _____0___29270, _____0___29271,
       _____0___29272, _____0___29273, _____0___29357, _____0___29358;
  wire _____0___29359, _____0___29360, _____0___29361, _____0___29362,
       _____0___29363, _____0___29364, _____0___29447, _____0___29448;
  wire _____0___29449, _____0___29450, _____0___29451, _____0___29452,
       _____0___29453, _____0___29454, _____0___29533, _____0___29534;
  wire _____0___29535, _____0___29616, _____0___29617, _____0___29618,
       _____0___29619, _____0___29620, _____0___29621, _____0___29622;
  wire _____0___29711, _____0___29712, _____0___29713, _____0___29714,
       _____0___29715, _____0___29716, _____0___29717, _____0___29804;
  wire _____0___29805, _____0___29806, _____0___29807, _____0___29808,
       _____0___29809, _____0___29810, _____0___29811, _____0___30095;
  wire _____0___30096, _____0___30097, _____0___30098, _____0___30099,
       _____0___30100, _____0___30101, _____0___30179, _____0___30180;
  wire _____0___30181, _____0___30182, _____0___30183, _____0___30184,
       _____0___30185, _____0___30186, _____0___30275, _____0___30276;
  wire _____0___30277, _____0___30278, _____0___30279, _____0___30280,
       _____0___30281, _____0___30365, _____0___30366, _____0___30367;
  wire _____0___30368, _____0___30369, _____0___30370, _____0___30371,
       _____0___30457, _____0___30458, _____0___30459, _____0___30460;
  wire _____0___30461, _____0___30462, _____0___30463, _____0___30546,
       _____0___30547, _____0___30548, _____0___30549, _____0___30550;
  wire _____0___30551, _____0___30552, _____0___30553, _____0___30633,
       _____0___30634, _____0___30635, _____0___30636, _____0___30637;
  wire _____0___30638, _____0___30639, _____0___30640, _____0___30727,
       _____0___30728, _____0___30729, _____0___30730, _____0___30731;
  wire _____0___30732, _____0___30733, _____0___30734, _____0___30998,
       _____0___30999, _____0___31000, _____0___31001, _____0___31002;
  wire _____0___31003, _____0___31004, _____0___31005, _____0___31094,
       _____0___31095, _____0___31096, _____0___31097, _____0___31098;
  wire _____0___31099, _____0___31100, _____0___31184, _____0___31185,
       _____0___31186, _____0___31187, _____0___31188, _____0___31189;
  wire _____0___31190, _____0___31191, _____0___31270, _____0___31271,
       _____0___31272, _____0___31273, _____0___31274, _____0___31275;
  wire _____0___31276, _____0___31355, _____0___31356, _____0___31357,
       _____0___31358, _____0___31359, _____0___31447, _____0___31448;
  wire _____0___31449, _____0___31450, _____0___31451, _____0___31452,
       _____0___31453, _____0___31454, _____0___31537, _____0___31538;
  wire _____0___31539, _____0___31540, _____0___31541, _____0___31542,
       _____0___31633, _____0___31634, _____0___31635, _____0___31636;
  wire _____0___31637, _____0___31638, _____0___31639, _____0___31901,
       _____0___31902, _____0___31903, _____0___31904, _____0___31905;
  wire _____0___31906, _____0___31907, _____0___31908, _____0___31998,
       _____0___31999, _____0___32000, _____0___32001, _____0___32002;
  wire _____0___32003, _____0___32004, _____0___32097, _____0___32098,
       _____0___32099, _____0___32100, _____0___32101, _____0___32102;
  wire _____0___32103, _____0___32104, _____0___32195, _____0___32196,
       _____0___32197, _____0___32198, _____0___32199, _____0___32200;
  wire _____0___32201, _____0___32202, _____0___32293, _____0___32294,
       _____0___32295, _____0___32296, _____0___32297, _____0___32298;
  wire _____0___32299, _____0___32300, _____0___32387, _____0___32388,
       _____0___32389, _____0___32390, _____0___32391, _____0___32392;
  wire _____0___32393, _____0___32394, _____0___32477, _____0___32478,
       _____0___32479, _____0___32480, _____0___32481, _____0___32482;
  wire _____0___32483, _____0___32484, _____0___32570, _____0___32571,
       _____0___32572, _____0___32573, _____0___32574, _____0___32575;
  wire _____0___32850, _____0___32851, _____0___32852, _____0___32853,
       _____0___32854, _____0___32855, _____0___32937, _____0___32938;
  wire _____0___32939, _____0___32940, _____0___32941, _____0___32942,
       _____0___32943, _____0___33030, _____0___33031, _____0___33032;
  wire _____0___33033, _____0___33034, _____0___33035, _____0___33036,
       _____0___33037, _____0___33128, _____0___33129, _____0___33130;
  wire _____0___33131, _____0___33132, _____0___33133, _____0___33134,
       _____0___33221, _____0___33222, _____0___33223, _____0___33224;
  wire _____0___33225, _____0___33226, _____0___33227, _____0___33311,
       _____0___33312, _____0___33313, _____0___33314, _____0___33315;
  wire _____0___33316, _____0___33402, _____0___33403, _____0___33404,
       _____0___33405, _____0___33406, _____0___33407, _____0___33408;
  wire _____0___33489, _____0___33490, _____0___33491, _____0___33492,
       _____0___33493, _____0___33494, _____0___33495, _____0___33770;
  wire _____0___33771, _____0___33772, _____0___33773, _____0___33774,
       _____0___33775, _____0___33776, _____0___33777, _____0___33866;
  wire _____0___33867, _____0___33868, _____0___33869, _____0___33870,
       _____0___33871, _____0___33872, _____0___33955, _____0___33956;
  wire _____0___33957, _____0___33958, _____0___33959, _____0___33960,
       _____0___33961, _____0___34046, _____0___34047, _____0___34048;
  wire _____0___34049, _____0___34050, _____0___34051, _____0___34052,
       _____0___34053, _____0___34145, _____0___34146, _____0___34147;
  wire _____0___34148, _____0___34149, _____0___34150, _____0___34151,
       _____0___34152, _____0___34239, _____0___34240, _____0___34241;
  wire _____0___34242, _____0___34243, _____0___34244, _____0___34245,
       _____0___34246, _____0___34334, _____0___34335, _____0___34336;
  wire _____0___34337, _____0___34338, _____0___34339, _____0___34340,
       _____0___34422, _____0___34423, _____0___34424, _____0___34425;
  wire _____0___34426, _____0___34427, _____0___34428, _____0___34429,
       _____0___34629, _____0___34630, _____0___34631, _____0___34632;
  wire _____0___34633, _____0___34634, _____0___34635, _____0___34636,
       _____0___34729, _____0___34730, _____0___34731, _____0___34732;
  wire _____0___34733, _____0___34734, _____0___34735, _____0___34736,
       _____0___34829, _____0___34830, _____0___34831, _____0___34832;
  wire _____0___34833, _____0___34834, _____0___34835, _____0___34836,
       _____0___34929, _____0___34930, _____0___34931, _____0___34932;
  wire _____0___34933, _____0___34934, _____0___34935, _____0___34936,
       _____0___35029, _____0___35030, _____0___35031, _____0___35032;
  wire _____0___35033, _____0___35034, _____0___35035, _____0___35036,
       _____0___35109, _____09__28243, _____09__28339, _____09__28434;
  wire _____09__28531, _____09__28624, _____09__28713, _____09__28809,
       _____09__28906, _____09__29185, _____09__29274, _____09__29365;
  wire _____09__29455, _____09__29536, _____09__29623, _____09__29718,
       _____09__29812, _____09__30102, _____09__30187, _____09__30282;
  wire _____09__30372, _____09__30464, _____09__30554, _____09__30641,
       _____09__30735, _____09__31006, _____09__31192, _____09__31277;
  wire _____09__31455, _____09__31543, _____09__31640, _____09__31909,
       _____09__32005, _____09__32105, _____09__32301, _____09__32395;
  wire _____09__32485, _____09__32576, _____09__32856, _____09__32944,
       _____09__33038, _____09__33135, _____09__33228, _____09__33317;
  wire _____09__33409, _____09__33496, _____09__33778, _____09__33873,
       _____09__33962, _____09__34054, _____09__34153, _____09__34247;
  wire _____09__34341, _____09__34430, _____09__34637, _____09__34737,
       _____09__34837, _____09__34937, _____09__35037, _____9;
  wire _____9__19085, _____9__19095, _____9__19105, _____9__19133,
       _____9__19143, _____9__19152, _____9__19162, _____9__19169;
  wire _____9__19177, _____9__19186, _____9__19195, _____9__19224,
       _____9__19233, _____9__19242, _____9__19251, _____9__19261;
  wire _____9__19271, _____9__19281, _____9__19291, _____9__19320,
       _____9__19330, _____9__19340, _____9__19350, _____9__19360;
  wire _____9__19370, _____9__19379, _____9__19389, _____9__19418,
       _____9__19428, _____9__19438, _____9__19448, _____9__19458;
  wire _____9__19467, _____9__19476, _____9__19486, _____9__19515,
       _____9__19524, _____9__19533, _____9__19543, _____9__19551;
  wire _____9__19561, _____9__19571, _____9__19581, _____9__19611,
       _____9__19621, _____9__19630, _____9__19638, _____9__19648;
  wire _____9__19658, _____9__19668, _____9__19676, _____9__19871,
       _____9__19881, _____9__19891, _____9__19900, _____9__19908;
  wire _____9__19917, _____9__19926, _____9__19936, _____9__19965,
       _____9__19984, _____9__19991, _____9__20001, _____9__20011;
  wire _____9__20020, _____9__20030, _____9__20058, _____9__20068,
       _____9__20078, _____9__20087, _____9__20096, _____9__20106;
  wire _____9__20115, _____9__20125, _____9__20155, _____9__20164,
       _____9__20172, _____9__20180, _____9__20188, _____9__20197;
  wire _____9__20206, _____9__20216, _____9__20244, _____9__20263,
       _____9__20273, _____9__20283, _____9__20293, _____9__20303;
  wire _____9__20313, _____9__20341, _____9__20351, _____9__20361,
       _____9__20371, _____9__20381, _____9__20391, _____9__20401;
  wire _____9__20438, _____9__20448, _____9__20455, _____9__20464,
       _____9__20483, _____9__20491, _____9__20499, _____9__20529;
  wire _____9__20539, _____9__20548, _____9__20557, _____9__20575,
       _____9__20584, _____9__20594, _____9__20806, _____9__20816;
  wire _____9__20826, _____9__20836, _____9__20846, _____9__20856,
       _____9__20865, _____9__20875, _____9__20903, _____9__20912;
  wire _____9__20922, _____9__20932, _____9__20951, _____9__20961,
       _____9__20971, _____9__21000, _____9__21009, _____9__21019;
  wire _____9__21029, _____9__21038, _____9__21045, _____9__21055,
       _____9__21065, _____9__21093, _____9__21102, _____9__21112;
  wire _____9__21119, _____9__21129, _____9__21139, _____9__21146,
       _____9__21155, _____9__21182, _____9__21190, _____9__21199;
  wire _____9__21209, _____9__21219, _____9__21229, _____9__21239,
       _____9__21249, _____9__21278, _____9__21287, _____9__21297;
  wire _____9__21307, _____9__21316, _____9__21326, _____9__21334,
       _____9__21344, _____9__21383, _____9__21392, _____9__21400;
  wire _____9__21428, _____9__21437, _____9__21464, _____9__21474,
       _____9__21484, _____9__21493, _____9__21503, _____9__21513;
  wire _____9__21522, _____9__21532, _____9__21738, _____9__21748,
       _____9__21756, _____9__21772, _____9__21782, _____9__21792;
  wire _____9__21800, _____9__21830, _____9__21839, _____9__21858,
       _____9__21867, _____9__21875, _____9__21884, _____9__21894;
  wire _____9__21923, _____9__21933, _____9__21939, _____9__21947,
       _____9__21956, _____9__21961, _____9__21970, _____9__21979;
  wire _____9__22004, _____9__22013, _____9__22022, _____9__22032,
       _____9__22042, _____9__22052, _____9__22062, _____9__22070;
  wire _____9__22098, _____9__22107, _____9__22117, _____9__22127,
       _____9__22137, _____9__22147, _____9__22156, _____9__22191;
  wire _____9__22199, _____9__22215, _____9__22223, _____9__22233,
       _____9__22241, _____9__22251, _____9__22280, _____9__22290;
  wire _____9__22299, _____9__22309, _____9__22326, _____9__22336,
       _____9__22345, _____9__22374, _____9__22391, _____9__22399;
  wire _____9__22408, _____9__22416, _____9__22426, _____9__22435,
       _____9__22643, _____9__22652, _____9__22669, _____9__22679;
  wire _____9__22689, _____9__22699, _____9__22708, _____9__22733,
       _____9__22743, _____9__22753, _____9__22763, _____9__22771;
  wire _____9__22779, _____9__22789, _____9__22797, _____9__22825,
       _____9__22832, _____9__22838, _____9__22847, _____9__22854;
  wire _____9__22864, _____9__22874, _____9__22884, _____9__22923,
       _____9__22933, _____9__22942, _____9__22951, _____9__22961;
  wire _____9__22971, _____9__22980, _____9__23008, _____9__23017,
       _____9__23027, _____9__23037, _____9__23047, _____9__23055;
  wire _____9__23064, _____9__23073, _____9__23099, _____9__23107,
       _____9__23124, _____9__23133, _____9__23142, _____9__23151;
  wire _____9__23161, _____9__23189, _____9__23214, _____9__23230,
       _____9__23240, _____9__23275, _____9__23285, _____9__23293;
  wire _____9__23302, _____9__23311, _____9__23325, _____9__23335,
       _____9__23544, _____9__23554, _____9__23563, _____9__23571;
  wire _____9__23581, _____9__23590, _____9__23600, _____9__23608,
       _____9__23637, _____9__23646, _____9__23655, _____9__23665;
  wire _____9__23674, _____9__23684, _____9__23694, _____9__23703,
       _____9__23727, _____9__23736, _____9__23746, _____9__23755;
  wire _____9__23764, _____9__23774, _____9__23784, _____9__23791,
       _____9__23820, _____9__23827, _____9__23836, _____9__23843;
  wire _____9__23859, _____9__23868, _____9__23876, _____9__23914,
       _____9__23924, _____9__23941, _____9__23957, _____9__23964;
  wire _____9__23991, _____9__24007, _____9__24017, _____9__24026,
       _____9__24034, _____9__24043, _____9__24052, _____9__24081;
  wire _____9__24091, _____9__24101, _____9__24110, _____9__24119,
       _____9__24129, _____9__24139, _____9__24147, _____9__24172;
  wire _____9__24181, _____9__24198, _____9__24208, _____9__24218,
       _____9__24234, _____9__24446, _____9__24464, _____9__24472;
  wire _____9__24480, _____9__24490, _____9__24498, _____9__24507,
       _____9__24533, _____9__24550, _____9__24559, _____9__24569;
  wire _____9__24578, _____9__24587, _____9__24597, _____9__24625,
       _____9__24635, _____9__24645, _____9__24655, _____9__24665;
  wire _____9__24675, _____9__24719, _____9__24738, _____9__24745,
       _____9__24755, _____9__24771, _____9__24781, _____9__24808;
  wire _____9__24818, _____9__24828, _____9__24838, _____9__24847,
       _____9__24857, _____9__24866, _____9__24876, _____9__24905;
  wire _____9__24915, _____9__24925, _____9__24935, _____9__24945,
       _____9__24955, _____9__24964, _____9__24973, _____9__25001;
  wire _____9__25011, _____9__25021, _____9__25031, _____9__25040,
       _____9__25050, _____9__25060, _____9__25070, _____9__25099;
  wire _____9__25108, _____9__25118, _____9__25126, _____9__25135,
       _____9__25145, _____9__25155, _____9__25164, _____9__25386;
  wire _____9__25396, _____9__25405, _____9__25415, _____9__25425,
       _____9__25435, _____9__25445, _____9__25454, _____9__25481;
  wire _____9__25491, _____9__25500, _____9__25510, _____9__25519,
       _____9__25528, _____9__25538, _____9__25548, _____9__25577;
  wire _____9__25587, _____9__25596, _____9__25606, _____9__25615,
       _____9__25624, _____9__25634, _____9__25644, _____9__25674;
  wire _____9__25684, _____9__25693, _____9__25702, _____9__25711,
       _____9__25720, _____9__25730, _____9__25740, _____9__25769;
  wire _____9__25779, _____9__25789, _____9__25799, _____9__25809,
       _____9__25819, _____9__25829, _____9__25839, _____9__25869;
  wire _____9__25879, _____9__25889, _____9__25908, _____9__25918,
       _____9__25928, _____9__25938, _____9__25966, _____9__25976;
  wire _____9__25986, _____9__25996, _____9__26006, _____9__26016,
       _____9__26026, _____9__26036, _____9__26066, _____9__26076;
  wire _____9__26086, _____9__26096, _____9__26106, _____9__26116,
       _____9__26126, _____9__26136, _____9___28322, _____9___28323;
  wire _____9___28324, _____9___28325, _____9___28326, _____9___28327,
       _____9___28328, _____9___28329, _____9___28417, _____9___28418;
  wire _____9___28419, _____9___28420, _____9___28421, _____9___28422,
       _____9___28423, _____9___28514, _____9___28515, _____9___28516;
  wire _____9___28517, _____9___28518, _____9___28519, _____9___28520,
       _____9___28521, _____9___28607, _____9___28608, _____9___28609;
  wire _____9___28610, _____9___28611, _____9___28612, _____9___28613,
       _____9___28614, _____9___28697, _____9___28698, _____9___28699;
  wire _____9___28700, _____9___28701, _____9___28702, _____9___28703,
       _____9___28792, _____9___28793, _____9___28794, _____9___28795;
  wire _____9___28796, _____9___28797, _____9___28798, _____9___28889,
       _____9___28890, _____9___28891, _____9___28892, _____9___28893;
  wire _____9___28894, _____9___28895, _____9___28896, _____9___28984,
       _____9___28985, _____9___28986, _____9___28987, _____9___28988;
  wire _____9___28989, _____9___28990, _____9___29257, _____9___29258,
       _____9___29259, _____9___29260, _____9___29261, _____9___29262;
  wire _____9___29263, _____9___29350, _____9___29351, _____9___29352,
       _____9___29353, _____9___29354, _____9___29438, _____9___29439;
  wire _____9___29440, _____9___29441, _____9___29442, _____9___29443,
       _____9___29444, _____9___29523, _____9___29524, _____9___29525;
  wire _____9___29526, _____9___29527, _____9___29528, _____9___29529,
       _____9___29530, _____9___29607, _____9___29608, _____9___29609;
  wire _____9___29610, _____9___29611, _____9___29612, _____9___29613,
       _____9___29701, _____9___29702, _____9___29703, _____9___29704;
  wire _____9___29705, _____9___29706, _____9___29707, _____9___29708,
       _____9___29794, _____9___29795, _____9___29796, _____9___29797;
  wire _____9___29798, _____9___29799, _____9___29800, _____9___29801,
       _____9___29892, _____9___29893, _____9___29894, _____9___29895;
  wire _____9___29896, _____9___29897, _____9___29898, _____9___29899,
       _____9___30171, _____9___30172, _____9___30173, _____9___30174;
  wire _____9___30175, _____9___30176, _____9___30177, _____9___30265,
       _____9___30266, _____9___30267, _____9___30268, _____9___30269;
  wire _____9___30270, _____9___30271, _____9___30272, _____9___30355,
       _____9___30356, _____9___30357, _____9___30358, _____9___30359;
  wire _____9___30360, _____9___30361, _____9___30362, _____9___30448,
       _____9___30449, _____9___30450, _____9___30451, _____9___30452;
  wire _____9___30453, _____9___30454, _____9___30539, _____9___30540,
       _____9___30541, _____9___30542, _____9___30543, _____9___30624;
  wire _____9___30625, _____9___30626, _____9___30627, _____9___30628,
       _____9___30629, _____9___30630, _____9___30718, _____9___30719;
  wire _____9___30720, _____9___30721, _____9___30722, _____9___30723,
       _____9___30724, _____9___30725, _____9___30811, _____9___30812;
  wire _____9___30813, _____9___30814, _____9___30815, _____9___30816,
       _____9___30817, _____9___30818, _____9___31085, _____9___31086;
  wire _____9___31087, _____9___31088, _____9___31089, _____9___31090,
       _____9___31091, _____9___31175, _____9___31176, _____9___31177;
  wire _____9___31178, _____9___31179, _____9___31180, _____9___31181,
       _____9___31263, _____9___31264, _____9___31265, _____9___31266;
  wire _____9___31267, _____9___31345, _____9___31346, _____9___31347,
       _____9___31348, _____9___31349, _____9___31350, _____9___31351;
  wire _____9___31352, _____9___31437, _____9___31438, _____9___31439,
       _____9___31440, _____9___31441, _____9___31442, _____9___31443;
  wire _____9___31444, _____9___31527, _____9___31528, _____9___31529,
       _____9___31530, _____9___31531, _____9___31532, _____9___31533;
  wire _____9___31534, _____9___31623, _____9___31624, _____9___31625,
       _____9___31626, _____9___31627, _____9___31628, _____9___31629;
  wire _____9___31630, _____9___31716, _____9___31717, _____9___31718,
       _____9___31719, _____9___31720, _____9___31721, _____9___31722;
  wire _____9___31988, _____9___31989, _____9___31990, _____9___31991,
       _____9___31992, _____9___31993, _____9___31994, _____9___31995;
  wire _____9___32087, _____9___32088, _____9___32089, _____9___32090,
       _____9___32091, _____9___32092, _____9___32093, _____9___32094;
  wire _____9___32185, _____9___32186, _____9___32187, _____9___32188,
       _____9___32189, _____9___32190, _____9___32191, _____9___32192;
  wire _____9___32283, _____9___32284, _____9___32285, _____9___32286,
       _____9___32287, _____9___32288, _____9___32289, _____9___32290;
  wire _____9___32378, _____9___32379, _____9___32380, _____9___32381,
       _____9___32382, _____9___32383, _____9___32384, _____9___32469;
  wire _____9___32470, _____9___32471, _____9___32472, _____9___32473,
       _____9___32474, _____9___32475, _____9___32561, _____9___32562;
  wire _____9___32563, _____9___32564, _____9___32565, _____9___32566,
       _____9___32567, _____9___32568, _____9___32647, _____9___32648;
  wire _____9___32649, _____9___32650, _____9___32651, _____9___32652,
       _____9___32653, _____9___32654, _____9___32929, _____9___32930;
  wire _____9___32931, _____9___32932, _____9___32933, _____9___32934,
       _____9___33020, _____9___33021, _____9___33022, _____9___33023;
  wire _____9___33024, _____9___33025, _____9___33026, _____9___33027,
       _____9___33118, _____9___33119, _____9___33120, _____9___33121;
  wire _____9___33122, _____9___33123, _____9___33124, _____9___33125,
       _____9___33213, _____9___33214, _____9___33215, _____9___33216;
  wire _____9___33217, _____9___33218, _____9___33303, _____9___33304,
       _____9___33305, _____9___33306, _____9___33307, _____9___33308;
  wire _____9___33392, _____9___33393, _____9___33394, _____9___33395,
       _____9___33396, _____9___33397, _____9___33398, _____9___33399;
  wire _____9___33480, _____9___33481, _____9___33482, _____9___33483,
       _____9___33484, _____9___33485, _____9___33486, _____9___33570;
  wire _____9___33571, _____9___33572, _____9___33573, _____9___33574,
       _____9___33575, _____9___33576, _____9___33577, _____9___33857;
  wire _____9___33858, _____9___33859, _____9___33860, _____9___33861,
       _____9___33862, _____9___33863, _____9___33945, _____9___33946;
  wire _____9___33947, _____9___33948, _____9___33949, _____9___33950,
       _____9___33951, _____9___33952, _____9___34037, _____9___34038;
  wire _____9___34039, _____9___34040, _____9___34041, _____9___34042,
       _____9___34043, _____9___34135, _____9___34136, _____9___34137;
  wire _____9___34138, _____9___34139, _____9___34140, _____9___34141,
       _____9___34142, _____9___34229, _____9___34230, _____9___34231;
  wire _____9___34232, _____9___34233, _____9___34234, _____9___34235,
       _____9___34236, _____9___34325, _____9___34326, _____9___34327;
  wire _____9___34328, _____9___34329, _____9___34330, _____9___34331,
       _____9___34412, _____9___34413, _____9___34414, _____9___34415;
  wire _____9___34416, _____9___34417, _____9___34418, _____9___34419,
       _____9___34509, _____9___34510, _____9___34511, _____9___34512;
  wire _____9___34513, _____9___34514, _____9___34515, _____9___34516,
       _____9___34719, _____9___34720, _____9___34721, _____9___34722;
  wire _____9___34723, _____9___34724, _____9___34725, _____9___34726,
       _____9___34819, _____9___34820, _____9___34821, _____9___34822;
  wire _____9___34823, _____9___34824, _____9___34825, _____9___34826,
       _____9___34919, _____9___34920, _____9___34921, _____9___34922;
  wire _____9___34923, _____9___34924, _____9___34925, _____9___34926,
       _____9___35019, _____9___35020, _____9___35021, _____9___35022;
  wire _____9___35023, _____9___35024, _____9___35025, _____9___35026,
       _____90__28321, _____90__28416, _____90__28606, _____90__28696;
  wire _____90__28791, _____90__28888, _____90__28983, _____90__29256,
       _____90__29349, _____90__29437, _____90__29522, _____90__29606;
  wire _____90__29700, _____90__29793, _____90__29891, _____90__30170,
       _____90__30264, _____90__30354, _____90__30447, _____90__30538;
  wire _____90__30623, _____90__30717, _____90__30810, _____90__31084,
       _____90__31174, _____90__31344, _____90__31526, _____90__31622;
  wire _____90__31715, _____90__31987, _____90__32086, _____90__32184,
       _____90__32282, _____90__32377, _____90__32468, _____90__32560;
  wire _____90__32646, _____90__32928, _____90__33117, _____90__33212,
       _____90__33302, _____90__33391, _____90__33479, _____90__33569;
  wire _____90__33944, _____90__34036, _____90__34134, _____90__34228,
       _____90__34324, _____90__34411, _____90__34508, _____90__34718;
  wire _____90__34818, _____90__34918, _____90__35018, _____99__28330,
       _____99__28424, _____99__28522, _____99__28615, _____99__28704;
  wire _____99__28799, _____99__28897, _____99__28991, _____99__29264,
       _____99__29355, _____99__29445, _____99__29531, _____99__29614;
  wire _____99__29709, _____99__29802, _____99__29900, _____99__30273,
       _____99__30363, _____99__30455, _____99__30544, _____99__30631;
  wire _____99__30819, _____99__31092, _____99__31182, _____99__31268,
       _____99__31353, _____99__31445, _____99__31535, _____99__31631;
  wire _____99__31723, _____99__31996, _____99__32095, _____99__32193,
       _____99__32291, _____99__32385, _____99__32476, _____99__32655;
  wire _____99__32935, _____99__33028, _____99__33126, _____99__33219,
       _____99__33309, _____99__33400, _____99__33487, _____99__33578;
  wire _____99__33864, _____99__33953, _____99__34044, _____99__34143,
       _____99__34237, _____99__34332, _____99__34420, _____99__34517;
  wire _____99__34727, _____99__34827, _____99__34927, _____99__35027,
       _____18906, _____18907, _____18908, _____18909;
  wire _____18910, _____18911, ______, ______0__18842, ______0__18849,
       ______0__18857, ______0__18865, ______0__28244;
  wire ______0__28254, ______0__28263, ______0__28273, ______0__28283,
       ______0__28292, ______0__28302, ______0__28311, ______0__28348;
  wire ______0__28358, ______0__28376, ______0__28386, ______0__28396,
       ______0__28406, ______0__28435, ______0__28445, ______0__28455;
  wire ______0__28465, ______0__28475, ______0__28485, ______0__28494,
       ______0__28504, ______0__28532, ______0__28542, ______0__28551;
  wire ______0__28569, ______0__28579, ______0__28589, ______0__28597,
       ______0__28625, ______0__28634, ______0__28643, ______0__28659;
  wire ______0__28677, ______0__28686, ______0__28714, ______0__28723,
       ______0__28733, ______0__28751, ______0__28761, ______0__28771;
  wire ______0__28781, ______0__28810, ______0__28820, ______0__28830,
       ______0__28840, ______0__28850, ______0__28860, ______0__28869;
  wire ______0__28878, ______0__28907, ______0__28917, ______0__28925,
       ______0__28935, ______0__28945, ______0__28955, ______0__28965;
  wire ______0__28974, ______0__29186, ______0__29196, ______0__29203,
       ______0__29212, ______0__29221, ______0__29230, ______0__29239;
  wire ______0__29247, ______0__29275, ______0__29283, ______0__29293,
       ______0__29301, ______0__29310, ______0__29320, ______0__29329;
  wire ______0__29339, ______0__29375, ______0__29385, ______0__29394,
       ______0__29403, ______0__29420, ______0__29429, ______0__29456;
  wire ______0__29466, ______0__29476, ______0__29484, ______0__29502,
       ______0__29512, ______0__29537, ______0__29545, ______0__29562;
  wire ______0__29571, ______0__29580, ______0__29597, ______0__29624,
       ______0__29634, ______0__29652, ______0__29662, ______0__29671;
  wire ______0__29680, ______0__29690, ______0__29719, ______0__29729,
       ______0__29739, ______0__29757, ______0__29766, ______0__29776;
  wire ______0__29813, ______0__29823, ______0__29833, ______0__29841,
       ______0__29851, ______0__29861, ______0__29871, ______0__29881;
  wire ______0__30103, ______0__30112, ______0__30121, ______0__30136,
       ______0__30143, ______0__30152, ______0__30162, ______0__30188;
  wire ______0__30198, ______0__30208, ______0__30217, ______0__30227,
       ______0__30237, ______0__30246, ______0__30255, ______0__30283;
  wire ______0__30291, ______0__30299, ______0__30309, ______0__30318,
       ______0__30327, ______0__30335, ______0__30345, ______0__30373;
  wire ______0__30382, ______0__30391, ______0__30399, ______0__30409,
       ______0__30418, ______0__30427, ______0__30437, ______0__30465;
  wire ______0__30475, ______0__30485, ______0__30494, ______0__30500,
       ______0__30510, ______0__30520, ______0__30530, ______0__30555;
  wire ______0__30564, ______0__30574, ______0__30582, ______0__30591,
       ______0__30600, ______0__30607, ______0__30642, ______0__30652;
  wire ______0__30662, ______0__30671, ______0__30680, ______0__30689,
       ______0__30698, ______0__30708, ______0__30736, ______0__30745;
  wire ______0__30764, ______0__30774, ______0__30784, ______0__30791,
       ______0__31007, ______0__31016, ______0__31025, ______0__31035;
  wire ______0__31044, ______0__31054, ______0__31064, ______0__31074,
       ______0__31101, ______0__31111, ______0__31121, ______0__31130;
  wire ______0__31140, ______0__31149, ______0__31159, ______0__31167,
       ______0__31193, ______0__31201, ______0__31211, ______0__31229;
  wire ______0__31238, ______0__31247, ______0__31254, ______0__31278,
       ______0__31286, ______0__31293, ______0__31299, ______0__31309;
  wire ______0__31317, ______0__31325, ______0__31334, ______0__31360,
       ______0__31370, ______0__31380, ______0__31390, ______0__31400;
  wire ______0__31410, ______0__31419, ______0__31427, ______0__31456,
       ______0__31466, ______0__31474, ______0__31482, ______0__31491;
  wire ______0__31501, ______0__31511, ______0__31544, ______0__31554,
       ______0__31564, ______0__31574, ______0__31583, ______0__31593;
  wire ______0__31602, ______0__31612, ______0__31641, ______0__31650,
       ______0__31659, ______0__31669, ______0__31678, ______0__31686;
  wire ______0__31696, ______0__31706, ______0__31910, ______0__31919,
       ______0__31929, ______0__31938, ______0__31948, ______0__31958;
  wire ______0__31968, ______0__31977, ______0__32006, ______0__32016,
       ______0__32026, ______0__32036, ______0__32046, ______0__32056;
  wire ______0__32066, ______0__32076, ______0__32106, ______0__32116,
       ______0__32126, ______0__32135, ______0__32145, ______0__32155;
  wire ______0__32164, ______0__32174, ______0__32203, ______0__32213,
       ______0__32223, ______0__32233, ______0__32243, ______0__32252;
  wire ______0__32262, ______0__32272, ______0__32302, ______0__32311,
       ______0__32321, ______0__32331, ______0__32341, ______0__32351;
  wire ______0__32360, ______0__32370, ______0__32396, ______0__32406,
       ______0__32416, ______0__32426, ______0__32436, ______0__32445;
  wire ______0__32453, ______0__32461, ______0__32486, ______0__32496,
       ______0__32506, ______0__32515, ______0__32524, ______0__32541;
  wire ______0__32550, ______0__32586, ______0__32594, ______0__32602,
       ______0__32611, ______0__32621, ______0__32628, ______0__32637;
  wire ______0__32857, ______0__32863, ______0__32873, ______0__32881,
       ______0__32890, ______0__32899, ______0__32909, ______0__32918;
  wire ______0__32945, ______0__32954, ______0__32964, ______0__32974,
       ______0__32984, ______0__32992, ______0__33000, ______0__33010;
  wire ______0__33039, ______0__33048, ______0__33058, ______0__33067,
       ______0__33077, ______0__33087, ______0__33097, ______0__33107;
  wire ______0__33136, ______0__33146, ______0__33156, ______0__33166,
       ______0__33175, ______0__33184, ______0__33193, ______0__33203;
  wire ______0__33229, ______0__33239, ______0__33248, ______0__33258,
       ______0__33276, ______0__33284, ______0__33292, ______0__33318;
  wire ______0__33327, ______0__33336, ______0__33354, ______0__33363,
       ______0__33373, ______0__33383, ______0__33419, ______0__33429;
  wire ______0__33437, ______0__33446, ______0__33454, ______0__33464,
       ______0__33473, ______0__33497, ______0__33506, ______0__33524;
  wire ______0__33533, ______0__33543, ______0__33553, ______0__33561,
       ______0__33779, ______0__33789, ______0__33799, ______0__33809;
  wire ______0__33819, ______0__33829, ______0__33839, ______0__33874,
       ______0__33883, ______0__33893, ______0__33900, ______0__33909;
  wire ______0__33918, ______0__33935, ______0__33963, ______0__33973,
       ______0__33983, ______0__33991, ______0__33999, ______0__34008;
  wire ______0__34018, ______0__34027, ______0__34055, ______0__34065,
       ______0__34075, ______0__34085, ______0__34095, ______0__34104;
  wire ______0__34114, ______0__34124, ______0__34154, ______0__34164,
       ______0__34174, ______0__34183, ______0__34192, ______0__34201;
  wire ______0__34210, ______0__34218, ______0__34248, ______0__34257,
       ______0__34265, ______0__34274, ______0__34284, ______0__34294;
  wire ______0__34304, ______0__34314, ______0__34342, ______0__34352,
       ______0__34360, ______0__34370, ______0__34380, ______0__34388;
  wire ______0__34396, ______0__34406, ______0__34431, ______0__34441,
       ______0__34451, ______0__34461, ______0__34471, ______0__34481;
  wire ______0__34491, ______0__34499, ______0__34638, ______0__34648,
       ______0__34658, ______0__34668, ______0__34678, ______0__34688;
  wire ______0__34698, ______0__34708, ______0__34738, ______0__34748,
       ______0__34758, ______0__34768, ______0__34778, ______0__34788;
  wire ______0__34798, ______0__34808, ______0__34838, ______0__34848,
       ______0__34858, ______0__34868, ______0__34878, ______0__34888;
  wire ______0__34898, ______0__34908, ______0__34938, ______0__34948,
       ______0__34958, ______0__34968, ______0__34978, ______0__34988;
  wire ______0__34998, ______0__35008, ______0__35038, ______0__35048,
       ______0__35058, ______0__35068, ______0__35078, ______0__35088;
  wire ______0__35098, ______9__18848, ______9__28253, ______9__28262,
       ______9__28272, ______9__28282, ______9__28291, ______9__28301;
  wire ______9__28310, ______9__28320, ______9__28347, ______9__28357,
       ______9__28375, ______9__28385, ______9__28395, ______9__28405;
  wire ______9__28415, ______9__28444, ______9__28454, ______9__28464,
       ______9__28474, ______9__28484, ______9__28493, ______9__28503;
  wire ______9__28513, ______9__28541, ______9__28560, ______9__28568,
       ______9__28578, ______9__28588, ______9__28596, ______9__28605;
  wire ______9__28633, ______9__28642, ______9__28658, ______9__28668,
       ______9__28676, ______9__28685, ______9__28695, ______9__28722;
  wire ______9__28732, ______9__28741, ______9__28750, ______9__28760,
       ______9__28770, ______9__28780, ______9__28790, ______9__28819;
  wire ______9__28829, ______9__28839, ______9__28849, ______9__28859,
       ______9__28868, ______9__28877, ______9__28887, ______9__28916;
  wire ______9__28934, ______9__28944, ______9__28954, ______9__28964,
       ______9__28973, ______9__28982, ______9__29195, ______9__29202;
  wire ______9__29211, ______9__29220, ______9__29229, ______9__29238,
       ______9__29246, ______9__29255, ______9__29282, ______9__29292;
  wire ______9__29300, ______9__29309, ______9__29319, ______9__29338,
       ______9__29348, ______9__29374, ______9__29384, ______9__29402;
  wire ______9__29419, ______9__29428, ______9__29465, ______9__29475,
       ______9__29491, ______9__29501, ______9__29511, ______9__29521;
  wire ______9__29544, ______9__29553, ______9__29561, ______9__29570,
       ______9__29579, ______9__29588, ______9__29596, ______9__29605;
  wire ______9__29633, ______9__29643, ______9__29651, ______9__29661,
       ______9__29670, ______9__29679, ______9__29689, ______9__29699;
  wire ______9__29728, ______9__29738, ______9__29747, ______9__29756,
       ______9__29765, ______9__29775, ______9__29792, ______9__29822;
  wire ______9__29832, ______9__29850, ______9__29860, ______9__29870,
       ______9__29880, ______9__29890, ______9__30111, ______9__30127;
  wire ______9__30135, ______9__30142, ______9__30161, ______9__30169,
       ______9__30197, ______9__30207, ______9__30216, ______9__30226;
  wire ______9__30236, ______9__30245, ______9__30254, ______9__30290,
       ______9__30298, ______9__30308, ______9__30317, ______9__30326;
  wire ______9__30334, ______9__30344, ______9__30353, ______9__30381,
       ______9__30398, ______9__30408, ______9__30417, ______9__30426;
  wire ______9__30436, ______9__30446, ______9__30474, ______9__30484,
       ______9__30493, ______9__30509, ______9__30519, ______9__30529;
  wire ______9__30537, ______9__30573, ______9__30581, ______9__30590,
       ______9__30599, ______9__30606, ______9__30622, ______9__30651;
  wire ______9__30661, ______9__30670, ______9__30679, ______9__30697,
       ______9__30707, ______9__30716, ______9__30744, ______9__30754;
  wire ______9__30763, ______9__30773, ______9__30783, ______9__30800,
       ______9__30809, ______9__31015, ______9__31024, ______9__31034;
  wire ______9__31043, ______9__31053, ______9__31063, ______9__31073,
       ______9__31083, ______9__31110, ______9__31120, ______9__31129;
  wire ______9__31139, ______9__31148, ______9__31158, ______9__31166,
       ______9__31200, ______9__31210, ______9__31219, ______9__31228;
  wire ______9__31237, ______9__31246, ______9__31253, ______9__31262,
       ______9__31292, ______9__31298, ______9__31308, ______9__31316;
  wire ______9__31324, ______9__31333, ______9__31343, ______9__31369,
       ______9__31379, ______9__31389, ______9__31399, ______9__31409;
  wire ______9__31418, ______9__31426, ______9__31436, ______9__31465,
       ______9__31473, ______9__31481, ______9__31490, ______9__31500;
  wire ______9__31510, ______9__31525, ______9__31553, ______9__31563,
       ______9__31573, ______9__31582, ______9__31592, ______9__31601;
  wire ______9__31611, ______9__31621, ______9__31649, ______9__31658,
       ______9__31668, ______9__31677, ______9__31685, ______9__31695;
  wire ______9__31705, ______9__31714, ______9__31918, ______9__31928,
       ______9__31947, ______9__31957, ______9__31967, ______9__31976;
  wire ______9__31986, ______9__32015, ______9__32025, ______9__32035,
       ______9__32045, ______9__32055, ______9__32065, ______9__32075;
  wire ______9__32085, ______9__32115, ______9__32125, ______9__32134,
       ______9__32144, ______9__32154, ______9__32163, ______9__32173;
  wire ______9__32183, ______9__32212, ______9__32222, ______9__32232,
       ______9__32242, ______9__32251, ______9__32261, ______9__32271;
  wire ______9__32281, ______9__32310, ______9__32320, ______9__32330,
       ______9__32340, ______9__32350, ______9__32369, ______9__32405;
  wire ______9__32415, ______9__32425, ______9__32435, ______9__32444,
       ______9__32460, ______9__32495, ______9__32505, ______9__32514;
  wire ______9__32523, ______9__32532, ______9__32540, ______9__32549,
       ______9__32559, ______9__32585, ______9__32593, ______9__32601;
  wire ______9__32610, ______9__32620, ______9__32636, ______9__32872,
       ______9__32880, ______9__32889, ______9__32898, ______9__32908;
  wire ______9__32917, ______9__32927, ______9__32963, ______9__32973,
       ______9__32983, ______9__32991, ______9__33009, ______9__33019;
  wire ______9__33047, ______9__33057, ______9__33076, ______9__33086,
       ______9__33096, ______9__33106, ______9__33116, ______9__33145;
  wire ______9__33155, ______9__33165, ______9__33183, ______9__33192,
       ______9__33202, ______9__33238, ______9__33247, ______9__33257;
  wire ______9__33266, ______9__33275, ______9__33283, ______9__33291,
       ______9__33301, ______9__33326, ______9__33335, ______9__33344;
  wire ______9__33353, ______9__33372, ______9__33382, ______9__33390,
       ______9__33418, ______9__33428, ______9__33436, ______9__33453;
  wire ______9__33463, ______9__33472, ______9__33505, ______9__33514,
       ______9__33523, ______9__33532, ______9__33542, ______9__33552;
  wire ______9__33560, ______9__33568, ______9__33788, ______9__33798,
       ______9__33808, ______9__33818, ______9__33828, ______9__33838;
  wire ______9__33848, ______9__33856, ______9__33882, ______9__33892,
       ______9__33899, ______9__33908, ______9__33917, ______9__33926;
  wire ______9__33934, ______9__33943, ______9__33972, ______9__33982,
       ______9__33990, ______9__34007, ______9__34017, ______9__34026;
  wire ______9__34035, ______9__34064, ______9__34074, ______9__34084,
       ______9__34094, ______9__34103, ______9__34113, ______9__34123;
  wire ______9__34133, ______9__34163, ______9__34173, ______9__34182,
       ______9__34191, ______9__34200, ______9__34209, ______9__34217;
  wire ______9__34227, ______9__34256, ______9__34264, ______9__34273,
       ______9__34283, ______9__34293, ______9__34303, ______9__34313;
  wire ______9__34323, ______9__34351, ______9__34359, ______9__34369,
       ______9__34379, ______9__34395, ______9__34405, ______9__34410;
  wire ______9__34440, ______9__34450, ______9__34460, ______9__34470,
       ______9__34480, ______9__34490, ______9__34498, ______9__34507;
  wire ______9__34647, ______9__34657, ______9__34667, ______9__34677,
       ______9__34687, ______9__34697, ______9__34707, ______9__34717;
  wire ______9__34747, ______9__34757, ______9__34767, ______9__34777,
       ______9__34787, ______9__34797, ______9__34807, ______9__34817;
  wire ______9__34847, ______9__34857, ______9__34867, ______9__34877,
       ______9__34887, ______9__34897, ______9__34907, ______9__34917;
  wire ______9__34947, ______9__34957, ______9__34967, ______9__34977,
       ______9__34987, ______9__34997, ______9__35007, ______9__35017;
  wire ______9__35047, ______9__35057, ______9__35067, ______9__35077,
       ______9__35087, ______9__35097, ______18912, ______18913;
  wire ______18914, ______18916, ______18917, ______18918, ______18919,
       ______18920, ______18922, ______18923;
  wire ______18924, ______18925, ______18927, ______18928, ______18929,
       ______18932, ______18933, ______18936;
  wire ______18937, ______18938, ______18939, ______18940, ______18941,
       ______18944, ______18945, ______18946;
  wire ______18947, ______18948, _______18950, _______18951,
       _______18954, _______18956, _______18957, _______18958;
  wire _______18960, _______18961, _______18962, _______18963,
       _______18964, _______18965, _______18966, _______18968;
  wire _______18969, _______18970, _______18971, _______18972,
       _______18973, _______18974, _______18990, _______18991;
  wire _______18992, _______18993, _______18994, _______18995,
       _______18998, _______18999, _______19000, _______19001;
  wire _______19002, _______19003, _______19004, _______19005,
       _______19008, _______19009, _______19010, _______19011;
  wire _______19012, _______19013, _______19014, _______19017,
       _______19018, _______19019, _______19020, _______19021;
  wire _______19022, _______19023, _______19024, _______19025,
       _______19026, _______19027, _______19028, _______19029;
  wire _______19037, _______19038, _______19039, _______19040,
       _______19043, _______19044, _______19047, _______19048;
  wire _______19049, _______19050, _______19051, _______19052,
       ________18840, ________18841, ________19060, ________19061;
  wire ________19062, ________19063, ________19064, ________19065,
       ________19066, ________19067, ________19069, ________19070;
  wire ________19071, ________19072, ________19073, ________19074,
       ________19075, ________19076, ________19077, ________19078;
  wire ________19079, ________19080, ________19081, ________19082,
       ________19083, ________19084, ________19087, ________19088;
  wire ________19089, ________19090, ________19091, ________19092,
       ________19093, ________19094, ________19097, ________19098;
  wire ________19099, ________19100, ________19101, ________19102,
       ________19103, ________19104, ________19125, ________19126;
  wire ________19127, ________19128, ________19129, ________19130,
       ________19131, ________19132, ________19135, ________19136;
  wire ________19137, ________19138, ________19139, ________19140,
       ________19141, ________19142, ________19145, ________19146;
  wire ________19147, ________19148, ________19149, ________19150,
       ________19151, ________19154, ________19155, ________19156;
  wire ________19157, ________19158, ________19159, ________19160,
       ________19161, ________19164, ________19165, ________19166;
  wire ________19167, ________19168, ________19171, ________19172,
       ________19173, ________19174, ________19175, ________19176;
  wire ________19178, ________19179, ________19180, ________19181,
       ________19182, ________19183, ________19184, ________19185;
  wire ________19188, ________19189, ________19190, ________19191,
       ________19192, ________19193, ________19194, ________19216;
  wire ________19217, ________19218, ________19219, ________19220,
       ________19221, ________19222, ________19223, ________19226;
  wire ________19227, ________19228, ________19229, ________19230,
       ________19231, ________19232, ________19235, ________19236;
  wire ________19237, ________19238, ________19239, ________19240,
       ________19241, ________19244, ________19245, ________19246;
  wire ________19247, ________19248, ________19249, ________19250,
       ________19253, ________19254, ________19255, ________19256;
  wire ________19257, ________19258, ________19259, ________19260,
       ________19263, ________19264, ________19265, ________19266;
  wire ________19267, ________19268, ________19269, ________19270,
       ________19273, ________19274, ________19275, ________19276;
  wire ________19277, ________19278, ________19279, ________19280,
       ________19283, ________19284, ________19285, ________19286;
  wire ________19287, ________19288, ________19289, ________19290,
       ________19313, ________19314, ________19315, ________19316;
  wire ________19317, ________19318, ________19319, ________19322,
       ________19323, ________19324, ________19325, ________19326;
  wire ________19327, ________19328, ________19329, ________19332,
       ________19333, ________19334, ________19335, ________19336;
  wire ________19337, ________19338, ________19339, ________19342,
       ________19343, ________19344, ________19345, ________19346;
  wire ________19347, ________19348, ________19349, ________19352,
       ________19353, ________19354, ________19355, ________19356;
  wire ________19357, ________19358, ________19359, ________19362,
       ________19363, ________19364, ________19365, ________19366;
  wire ________19367, ________19368, ________19369, ________19372,
       ________19373, ________19374, ________19375, ________19376;
  wire ________19377, ________19378, ________19381, ________19382,
       ________19383, ________19384, ________19385, ________19386;
  wire ________19387, ________19388, ________19410, ________19411,
       ________19412, ________19413, ________19414, ________19415;
  wire ________19416, ________19417, ________19420, ________19421,
       ________19422, ________19423, ________19424, ________19425;
  wire ________19426, ________19427, ________19430, ________19431,
       ________19432, ________19433, ________19434, ________19435;
  wire ________19436, ________19437, ________19440, ________19441,
       ________19442, ________19443, ________19444, ________19445;
  wire ________19446, ________19447, ________19450, ________19451,
       ________19452, ________19453, ________19454, ________19455;
  wire ________19456, ________19457, ________19459, ________19460,
       ________19461, ________19462, ________19463, ________19464;
  wire ________19465, ________19466, ________19469, ________19470,
       ________19471, ________19472, ________19473, ________19474;
  wire ________19475, ________19478, ________19479, ________19480,
       ________19481, ________19482, ________19483, ________19484;
  wire ________19485, ________19507, ________19508, ________19509,
       ________19510, ________19511, ________19512, ________19513;
  wire ________19514, ________19517, ________19518, ________19519,
       ________19520, ________19521, ________19522, ________19523;
  wire ________19526, ________19527, ________19528, ________19529,
       ________19530, ________19531, ________19532, ________19535;
  wire ________19536, ________19537, ________19538, ________19539,
       ________19540, ________19541, ________19542, ________19544;
  wire ________19545, ________19546, ________19547, ________19548,
       ________19549, ________19550, ________19553, ________19554;
  wire ________19555, ________19556, ________19557, ________19558,
       ________19559, ________19560, ________19563, ________19564;
  wire ________19565, ________19566, ________19567, ________19568,
       ________19569, ________19570, ________19573, ________19574;
  wire ________19575, ________19576, ________19577, ________19578,
       ________19579, ________19580, ________19603, ________19604;
  wire ________19605, ________19606, ________19607, ________19608,
       ________19609, ________19610, ________19613, ________19614;
  wire ________19615, ________19616, ________19617, ________19618,
       ________19619, ________19620, ________19623, ________19624;
  wire ________19625, ________19626, ________19627, ________19628,
       ________19629, ________19631, ________19632, ________19633;
  wire ________19634, ________19635, ________19636, ________19637,
       ________19640, ________19641, ________19642, ________19643;
  wire ________19644, ________19645, ________19646, ________19647,
       ________19650, ________19651, ________19652, ________19653;
  wire ________19654, ________19655, ________19656, ________19657,
       ________19660, ________19661, ________19662, ________19663;
  wire ________19664, ________19665, ________19666, ________19667,
       ________19670, ________19671, ________19672, ________19673;
  wire ________19674, ________19675, ________19863, ________19864,
       ________19865, ________19866, ________19867, ________19868;
  wire ________19869, ________19870, ________19873, ________19874,
       ________19875, ________19876, ________19877, ________19878;
  wire ________19879, ________19880, ________19883, ________19884,
       ________19885, ________19886, ________19887, ________19888;
  wire ________19889, ________19890, ________19893, ________19894,
       ________19895, ________19896, ________19897, ________19898;
  wire ________19899, ________19901, ________19902, ________19903,
       ________19904, ________19905, ________19906, ________19907;
  wire ________19910, ________19911, ________19912, ________19913,
       ________19914, ________19915, ________19916, ________19919;
  wire ________19920, ________19921, ________19922, ________19923,
       ________19924, ________19925, ________19928, ________19929;
  wire ________19930, ________19931, ________19932, ________19933,
       ________19934, ________19935, ________19957, ________19958;
  wire ________19959, ________19960, ________19961, ________19962,
       ________19963, ________19964, ________19967, ________19968;
  wire ________19969, ________19970, ________19971, ________19972,
       ________19973, ________19974, ________19976, ________19977;
  wire ________19978, ________19979, ________19980, ________19981,
       ________19982, ________19983, ________19986, ________19987;
  wire ________19988, ________19989, ________19990, ________19993,
       ________19994, ________19995, ________19996, ________19997;
  wire ________19998, ________19999, ________20000, ________20003,
       ________20004, ________20005, ________20006, ________20007;
  wire ________20008, ________20009, ________20010, ________20013,
       ________20014, ________20015, ________20016, ________20017;
  wire ________20018, ________20019, ________20022, ________20023,
       ________20024, ________20025, ________20026, ________20027;
  wire ________20028, ________20029, ________20050, ________20051,
       ________20052, ________20053, ________20054, ________20055;
  wire ________20056, ________20057, ________20060, ________20061,
       ________20062, ________20063, ________20064, ________20065;
  wire ________20066, ________20067, ________20070, ________20071,
       ________20072, ________20073, ________20074, ________20075;
  wire ________20076, ________20077, ________20080, ________20081,
       ________20082, ________20083, ________20084, ________20085;
  wire ________20086, ________20089, ________20090, ________20091,
       ________20092, ________20093, ________20094, ________20095;
  wire ________20098, ________20099, ________20100, ________20101,
       ________20102, ________20103, ________20104, ________20105;
  wire ________20108, ________20109, ________20110, ________20111,
       ________20112, ________20113, ________20114, ________20117;
  wire ________20118, ________20119, ________20120, ________20121,
       ________20122, ________20123, ________20124, ________20147;
  wire ________20148, ________20149, ________20150, ________20151,
       ________20152, ________20153, ________20154, ________20157;
  wire ________20158, ________20159, ________20160, ________20161,
       ________20162, ________20163, ________20165, ________20166;
  wire ________20167, ________20168, ________20169, ________20170,
       ________20171, ________20173, ________20174, ________20175;
  wire ________20176, ________20177, ________20178, ________20179,
       ________20182, ________20183, ________20184, ________20185;
  wire ________20186, ________20187, ________20190, ________20191,
       ________20192, ________20193, ________20194, ________20195;
  wire ________20196, ________20199, ________20200, ________20201,
       ________20202, ________20203, ________20204, ________20205;
  wire ________20208, ________20209, ________20210, ________20211,
       ________20212, ________20213, ________20214, ________20215;
  wire ________20236, ________20237, ________20238, ________20239,
       ________20240, ________20241, ________20242, ________20243;
  wire ________20246, ________20247, ________20248, ________20249,
       ________20250, ________20251, ________20252, ________20253;
  wire ________20255, ________20256, ________20257, ________20258,
       ________20259, ________20260, ________20261, ________20262;
  wire ________20265, ________20266, ________20267, ________20268,
       ________20269, ________20270, ________20271, ________20272;
  wire ________20275, ________20276, ________20277, ________20278,
       ________20279, ________20280, ________20281, ________20282;
  wire ________20285, ________20286, ________20287, ________20288,
       ________20289, ________20290, ________20291, ________20292;
  wire ________20295, ________20296, ________20297, ________20298,
       ________20299, ________20300, ________20301, ________20302;
  wire ________20305, ________20306, ________20307, ________20308,
       ________20309, ________20310, ________20311, ________20312;
  wire ________20333, ________20334, ________20335, ________20336,
       ________20337, ________20338, ________20339, ________20340;
  wire ________20343, ________20344, ________20345, ________20346,
       ________20347, ________20348, ________20349, ________20350;
  wire ________20353, ________20354, ________20355, ________20356,
       ________20357, ________20358, ________20359, ________20360;
  wire ________20363, ________20364, ________20365, ________20366,
       ________20367, ________20368, ________20369, ________20370;
  wire ________20373, ________20374, ________20375, ________20376,
       ________20377, ________20378, ________20379, ________20380;
  wire ________20383, ________20384, ________20385, ________20386,
       ________20387, ________20388, ________20389, ________20390;
  wire ________20393, ________20394, ________20395, ________20396,
       ________20397, ________20398, ________20399, ________20400;
  wire ________20403, ________20404, ________20405, ________20406,
       ________20407, ________20408, ________20409, ________20430;
  wire ________20431, ________20432, ________20433, ________20434,
       ________20435, ________20436, ________20437, ________20440;
  wire ________20441, ________20442, ________20443, ________20444,
       ________20445, ________20446, ________20447, ________20449;
  wire ________20450, ________20451, ________20452, ________20453,
       ________20454, ________20457, ________20458, ________20459;
  wire ________20460, ________20461, ________20462, ________20463,
       ________20466, ________20467, ________20468, ________20469;
  wire ________20470, ________20471, ________20472, ________20473,
       ________20475, ________20476, ________20477, ________20478;
  wire ________20479, ________20480, ________20481, ________20482,
       ________20485, ________20486, ________20487, ________20488;
  wire ________20489, ________20490, ________20493, ________20494,
       ________20495, ________20496, ________20497, ________20498;
  wire ________20521, ________20522, ________20523, ________20524,
       ________20525, ________20526, ________20527, ________20528;
  wire ________20531, ________20532, ________20533, ________20534,
       ________20535, ________20536, ________20537, ________20538;
  wire ________20541, ________20542, ________20543, ________20544,
       ________20545, ________20546, ________20547, ________20550;
  wire ________20551, ________20552, ________20553, ________20554,
       ________20555, ________20556, ________20559, ________20560;
  wire ________20561, ________20562, ________20563, ________20564,
       ________20565, ________20566, ________20568, ________20569;
  wire ________20570, ________20571, ________20572, ________20573,
       ________20574, ________20577, ________20578, ________20579;
  wire ________20580, ________20581, ________20582, ________20583,
       ________20586, ________20587, ________20588, ________20589;
  wire ________20590, ________20591, ________20592, ________20593,
       ________20800, ________20801, ________20802, ________20803;
  wire ________20804, ________20805, ________20808, ________20809,
       ________20810, ________20811, ________20812, ________20813;
  wire ________20814, ________20815, ________20818, ________20819,
       ________20820, ________20821, ________20822, ________20823;
  wire ________20824, ________20825, ________20828, ________20829,
       ________20830, ________20831, ________20832, ________20833;
  wire ________20834, ________20835, ________20838, ________20839,
       ________20840, ________20841, ________20842, ________20843;
  wire ________20844, ________20845, ________20848, ________20849,
       ________20850, ________20851, ________20852, ________20853;
  wire ________20854, ________20855, ________20858, ________20859,
       ________20860, ________20861, ________20862, ________20863;
  wire ________20864, ________20867, ________20868, ________20869,
       ________20870, ________20871, ________20872, ________20873;
  wire ________20874, ________20896, ________20897, ________20898,
       ________20899, ________20900, ________20901, ________20902;
  wire ________20905, ________20906, ________20907, ________20908,
       ________20909, ________20910, ________20911, ________20914;
  wire ________20915, ________20916, ________20917, ________20918,
       ________20919, ________20920, ________20921, ________20924;
  wire ________20925, ________20926, ________20927, ________20928,
       ________20929, ________20930, ________20931, ________20934;
  wire ________20935, ________20936, ________20937, ________20938,
       ________20939, ________20940, ________20941, ________20943;
  wire ________20944, ________20945, ________20946, ________20947,
       ________20948, ________20949, ________20950, ________20953;
  wire ________20954, ________20955, ________20956, ________20957,
       ________20958, ________20959, ________20960, ________20963;
  wire ________20964, ________20965, ________20966, ________20967,
       ________20968, ________20969, ________20970, ________20992;
  wire ________20993, ________20994, ________20995, ________20996,
       ________20997, ________20998, ________20999, ________21002;
  wire ________21003, ________21004, ________21005, ________21006,
       ________21007, ________21008, ________21011, ________21012;
  wire ________21013, ________21014, ________21015, ________21016,
       ________21017, ________21018, ________21021, ________21022;
  wire ________21023, ________21024, ________21025, ________21026,
       ________21027, ________21028, ________21031, ________21032;
  wire ________21033, ________21034, ________21035, ________21036,
       ________21037, ________21039, ________21040, ________21041;
  wire ________21042, ________21043, ________21044, ________21047,
       ________21048, ________21049, ________21050, ________21051;
  wire ________21052, ________21053, ________21054, ________21057,
       ________21058, ________21059, ________21060, ________21061;
  wire ________21062, ________21063, ________21064, ________21086,
       ________21087, ________21088, ________21089, ________21090;
  wire ________21091, ________21092, ________21094, ________21095,
       ________21096, ________21097, ________21098, ________21099;
  wire ________21100, ________21101, ________21104, ________21105,
       ________21106, ________21107, ________21108, ________21109;
  wire ________21110, ________21111, ________21113, ________21114,
       ________21115, ________21116, ________21117, ________21118;
  wire ________21121, ________21122, ________21123, ________21124,
       ________21125, ________21126, ________21127, ________21128;
  wire ________21131, ________21132, ________21133, ________21134,
       ________21135, ________21136, ________21137, ________21138;
  wire ________21141, ________21142, ________21143, ________21144,
       ________21145, ________21148, ________21149, ________21150;
  wire ________21151, ________21152, ________21153, ________21154,
       ________21174, ________21175, ________21176, ________21177;
  wire ________21178, ________21179, ________21180, ________21181,
       ________21184, ________21185, ________21186, ________21187;
  wire ________21188, ________21189, ________21192, ________21193,
       ________21194, ________21195, ________21196, ________21197;
  wire ________21198, ________21201, ________21202, ________21203,
       ________21204, ________21205, ________21206, ________21207;
  wire ________21208, ________21211, ________21212, ________21213,
       ________21214, ________21215, ________21216, ________21217;
  wire ________21218, ________21221, ________21222, ________21223,
       ________21224, ________21225, ________21226, ________21227;
  wire ________21228, ________21231, ________21232, ________21233,
       ________21234, ________21235, ________21236, ________21237;
  wire ________21238, ________21241, ________21242, ________21243,
       ________21244, ________21245, ________21246, ________21247;
  wire ________21248, ________21271, ________21272, ________21273,
       ________21274, ________21275, ________21276, ________21277;
  wire ________21280, ________21281, ________21282, ________21283,
       ________21284, ________21285, ________21286, ________21289;
  wire ________21290, ________21291, ________21292, ________21293,
       ________21294, ________21295, ________21296, ________21299;
  wire ________21300, ________21301, ________21302, ________21303,
       ________21304, ________21305, ________21306, ________21309;
  wire ________21310, ________21311, ________21312, ________21313,
       ________21314, ________21315, ________21318, ________21319;
  wire ________21320, ________21321, ________21322, ________21323,
       ________21324, ________21325, ________21328, ________21329;
  wire ________21330, ________21331, ________21332, ________21333,
       ________21336, ________21337, ________21338, ________21339;
  wire ________21340, ________21341, ________21342, ________21343,
       ________21366, ________21367, ________21368, ________21369;
  wire ________21370, ________21371, ________21372, ________21373,
       ________21375, ________21376, ________21377, ________21378;
  wire ________21379, ________21380, ________21381, ________21382,
       ________21385, ________21386, ________21387, ________21388;
  wire ________21389, ________21390, ________21391, ________21394,
       ________21395, ________21396, ________21397, ________21398;
  wire ________21399, ________21402, ________21403, ________21404,
       ________21405, ________21406, ________21407, ________21408;
  wire ________21409, ________21411, ________21412, ________21413,
       ________21414, ________21415, ________21416, ________21417;
  wire ________21418, ________21420, ________21421, ________21422,
       ________21423, ________21424, ________21425, ________21426;
  wire ________21427, ________21430, ________21431, ________21432,
       ________21433, ________21434, ________21435, ________21436;
  wire ________21456, ________21457, ________21458, ________21459,
       ________21460, ________21461, ________21462, ________21463;
  wire ________21466, ________21467, ________21468, ________21469,
       ________21470, ________21471, ________21472, ________21473;
  wire ________21476, ________21477, ________21478, ________21479,
       ________21480, ________21481, ________21482, ________21483;
  wire ________21486, ________21487, ________21488, ________21489,
       ________21490, ________21491, ________21492, ________21495;
  wire ________21496, ________21497, ________21498, ________21499,
       ________21500, ________21501, ________21502, ________21505;
  wire ________21506, ________21507, ________21508, ________21509,
       ________21510, ________21511, ________21512, ________21515;
  wire ________21516, ________21517, ________21518, ________21519,
       ________21520, ________21521, ________21524, ________21525;
  wire ________21526, ________21527, ________21528, ________21529,
       ________21530, ________21531, ________21730, ________21731;
  wire ________21732, ________21733, ________21734, ________21735,
       ________21736, ________21737, ________21740, ________21741;
  wire ________21742, ________21743, ________21744, ________21745,
       ________21746, ________21747, ________21750, ________21751;
  wire ________21752, ________21753, ________21754, ________21755,
       ________21758, ________21759, ________21760, ________21761;
  wire ________21762, ________21764, ________21765, ________21766,
       ________21767, ________21768, ________21769, ________21770;
  wire ________21771, ________21774, ________21775, ________21776,
       ________21777, ________21778, ________21779, ________21780;
  wire ________21781, ________21784, ________21785, ________21786,
       ________21787, ________21788, ________21789, ________21790;
  wire ________21791, ________21793, ________21794, ________21795,
       ________21796, ________21797, ________21798, ________21799;
  wire ________21822, ________21823, ________21824, ________21825,
       ________21826, ________21827, ________21828, ________21829;
  wire ________21832, ________21833, ________21834, ________21835,
       ________21836, ________21837, ________21838, ________21841;
  wire ________21842, ________21843, ________21844, ________21845,
       ________21846, ________21847, ________21848, ________21850;
  wire ________21851, ________21852, ________21853, ________21854,
       ________21855, ________21856, ________21857, ________21860;
  wire ________21861, ________21862, ________21863, ________21864,
       ________21865, ________21866, ________21868, ________21869;
  wire ________21870, ________21871, ________21872, ________21873,
       ________21874, ________21877, ________21878, ________21879;
  wire ________21880, ________21881, ________21882, ________21883,
       ________21886, ________21887, ________21888, ________21889;
  wire ________21890, ________21891, ________21892, ________21893,
       ________21915, ________21916, ________21917, ________21918;
  wire ________21919, ________21920, ________21921, ________21922,
       ________21925, ________21926, ________21927, ________21928;
  wire ________21929, ________21930, ________21931, ________21932,
       ________21935, ________21936, ________21937, ________21938;
  wire ________21941, ________21942, ________21943, ________21944,
       ________21945, ________21946, ________21949, ________21950;
  wire ________21951, ________21952, ________21953, ________21954,
       ________21955, ________21957, ________21958, ________21959;
  wire ________21960, ________21963, ________21964, ________21965,
       ________21966, ________21967, ________21968, ________21969;
  wire ________21972, ________21973, ________21974, ________21975,
       ________21976, ________21977, ________21978, ________21996;
  wire ________21997, ________21998, ________21999, ________22000,
       ________22001, ________22002, ________22003, ________22006;
  wire ________22007, ________22008, ________22009, ________22010,
       ________22011, ________22012, ________22015, ________22016;
  wire ________22017, ________22018, ________22019, ________22020,
       ________22021, ________22024, ________22025, ________22026;
  wire ________22027, ________22028, ________22029, ________22030,
       ________22031, ________22034, ________22035, ________22036;
  wire ________22037, ________22038, ________22039, ________22040,
       ________22041, ________22044, ________22045, ________22046;
  wire ________22047, ________22048, ________22049, ________22050,
       ________22051, ________22054, ________22055, ________22056;
  wire ________22057, ________22058, ________22059, ________22060,
       ________22061, ________22064, ________22065, ________22066;
  wire ________22067, ________22068, ________22069, ________22090,
       ________22091, ________22092, ________22093, ________22094;
  wire ________22095, ________22096, ________22097, ________22100,
       ________22101, ________22102, ________22103, ________22104;
  wire ________22105, ________22106, ________22109, ________22110,
       ________22111, ________22112, ________22113, ________22114;
  wire ________22115, ________22116, ________22119, ________22120,
       ________22121, ________22122, ________22123, ________22124;
  wire ________22125, ________22126, ________22129, ________22130,
       ________22131, ________22132, ________22133, ________22134;
  wire ________22135, ________22136, ________22139, ________22140,
       ________22141, ________22142, ________22143, ________22144;
  wire ________22145, ________22146, ________22149, ________22150,
       ________22151, ________22152, ________22153, ________22154;
  wire ________22155, ________22158, ________22159, ________22160,
       ________22161, ________22162, ________22183, ________22184;
  wire ________22185, ________22186, ________22187, ________22188,
       ________22189, ________22190, ________22193, ________22194;
  wire ________22195, ________22196, ________22197, ________22198,
       ________22201, ________22202, ________22203, ________22204;
  wire ________22205, ________22207, ________22208, ________22209,
       ________22210, ________22211, ________22212, ________22213;
  wire ________22214, ________22217, ________22218, ________22219,
       ________22220, ________22221, ________22222, ________22225;
  wire ________22226, ________22227, ________22228, ________22229,
       ________22230, ________22231, ________22232, ________22235;
  wire ________22236, ________22237, ________22238, ________22239,
       ________22240, ________22243, ________22244, ________22245;
  wire ________22246, ________22247, ________22248, ________22249,
       ________22250, ________22272, ________22273, ________22274;
  wire ________22275, ________22276, ________22277, ________22278,
       ________22279, ________22282, ________22283, ________22284;
  wire ________22285, ________22286, ________22287, ________22288,
       ________22289, ________22292, ________22293, ________22294;
  wire ________22295, ________22296, ________22297, ________22298,
       ________22301, ________22302, ________22303, ________22304;
  wire ________22305, ________22306, ________22307, ________22308,
       ________22311, ________22312, ________22313, ________22314;
  wire ________22315, ________22316, ________22317, ________22318,
       ________22320, ________22321, ________22322, ________22323;
  wire ________22324, ________22325, ________22328, ________22329,
       ________22330, ________22331, ________22332, ________22333;
  wire ________22334, ________22335, ________22338, ________22339,
       ________22340, ________22341, ________22342, ________22343;
  wire ________22344, ________22367, ________22368, ________22369,
       ________22370, ________22371, ________22372, ________22373;
  wire ________22376, ________22377, ________22378, ________22379,
       ________22380, ________22381, ________22382, ________22383;
  wire ________22385, ________22386, ________22387, ________22388,
       ________22389, ________22390, ________22392, ________22393;
  wire ________22394, ________22395, ________22396, ________22397,
       ________22398, ________22401, ________22402, ________22403;
  wire ________22404, ________22405, ________22406, ________22407,
       ________22409, ________22410, ________22411, ________22412;
  wire ________22413, ________22414, ________22415, ________22418,
       ________22419, ________22420, ________22421, ________22422;
  wire ________22423, ________22424, ________22425, ________22428,
       ________22429, ________22430, ________22431, ________22432;
  wire ________22433, ________22434, ________22636, ________22637,
       ________22638, ________22639, ________22640, ________22641;
  wire ________22642, ________22645, ________22646, ________22647,
       ________22648, ________22649, ________22650, ________22651;
  wire ________22654, ________22655, ________22656, ________22657,
       ________22658, ________22659, ________22660, ________22661;
  wire ________22662, ________22663, ________22664, ________22665,
       ________22666, ________22667, ________22668, ________22671;
  wire ________22672, ________22673, ________22674, ________22675,
       ________22676, ________22677, ________22678, ________22681;
  wire ________22682, ________22683, ________22684, ________22685,
       ________22686, ________22687, ________22688, ________22691;
  wire ________22692, ________22693, ________22694, ________22695,
       ________22696, ________22697, ________22698, ________22701;
  wire ________22702, ________22703, ________22704, ________22705,
       ________22706, ________22707, ________22726, ________22727;
  wire ________22728, ________22729, ________22730, ________22731,
       ________22732, ________22735, ________22736, ________22737;
  wire ________22738, ________22739, ________22740, ________22741,
       ________22742, ________22745, ________22746, ________22747;
  wire ________22748, ________22749, ________22750, ________22751,
       ________22752, ________22755, ________22756, ________22757;
  wire ________22758, ________22759, ________22760, ________22761,
       ________22762, ________22765, ________22766, ________22767;
  wire ________22768, ________22769, ________22770, ________22773,
       ________22774, ________22775, ________22776, ________22777;
  wire ________22778, ________22781, ________22782, ________22783,
       ________22784, ________22785, ________22786, ________22787;
  wire ________22788, ________22791, ________22792, ________22793,
       ________22794, ________22795, ________22796, ________22817;
  wire ________22818, ________22819, ________22820, ________22821,
       ________22822, ________22823, ________22824, ________22827;
  wire ________22828, ________22829, ________22830, ________22831,
       ________22834, ________22835, ________22836, ________22837;
  wire ________22839, ________22840, ________22841, ________22842,
       ________22843, ________22844, ________22845, ________22846;
  wire ________22849, ________22850, ________22851, ________22852,
       ________22853, ________22856, ________22857, ________22858;
  wire ________22859, ________22860, ________22861, ________22862,
       ________22863, ________22866, ________22867, ________22868;
  wire ________22869, ________22870, ________22871, ________22872,
       ________22873, ________22876, ________22877, ________22878;
  wire ________22879, ________22880, ________22881, ________22882,
       ________22883, ________22906, ________22907, ________22908;
  wire ________22909, ________22910, ________22911, ________22912,
       ________22913, ________22915, ________22916, ________22917;
  wire ________22918, ________22919, ________22920, ________22921,
       ________22922, ________22925, ________22926, ________22927;
  wire ________22928, ________22929, ________22930, ________22931,
       ________22932, ________22935, ________22936, ________22937;
  wire ________22938, ________22939, ________22940, ________22941,
       ________22943, ________22944, ________22945, ________22946;
  wire ________22947, ________22948, ________22949, ________22950,
       ________22953, ________22954, ________22955, ________22956;
  wire ________22957, ________22958, ________22959, ________22960,
       ________22963, ________22964, ________22965, ________22966;
  wire ________22967, ________22968, ________22969, ________22970,
       ________22972, ________22973, ________22974, ________22975;
  wire ________22976, ________22977, ________22978, ________22979,
       ________23000, ________23001, ________23002, ________23003;
  wire ________23004, ________23005, ________23006, ________23007,
       ________23010, ________23011, ________23012, ________23013;
  wire ________23014, ________23015, ________23016, ________23019,
       ________23020, ________23021, ________23022, ________23023;
  wire ________23024, ________23025, ________23026, ________23029,
       ________23030, ________23031, ________23032, ________23033;
  wire ________23034, ________23035, ________23036, ________23039,
       ________23040, ________23041, ________23042, ________23043;
  wire ________23044, ________23045, ________23046, ________23048,
       ________23049, ________23050, ________23051, ________23052;
  wire ________23053, ________23054, ________23057, ________23058,
       ________23059, ________23060, ________23061, ________23062;
  wire ________23063, ________23066, ________23067, ________23068,
       ________23069, ________23070, ________23071, ________23072;
  wire ________23093, ________23094, ________23095, ________23096,
       ________23097, ________23098, ________23100, ________23101;
  wire ________23102, ________23103, ________23104, ________23105,
       ________23106, ________23109, ________23110, ________23111;
  wire ________23112, ________23113, ________23114, ________23116,
       ________23117, ________23118, ________23119, ________23120;
  wire ________23121, ________23122, ________23123, ________23126,
       ________23127, ________23128, ________23129, ________23130;
  wire ________23131, ________23132, ________23135, ________23136,
       ________23137, ________23138, ________23139, ________23140;
  wire ________23141, ________23144, ________23145, ________23146,
       ________23147, ________23148, ________23149, ________23150;
  wire ________23153, ________23154, ________23155, ________23156,
       ________23157, ________23158, ________23159, ________23160;
  wire ________23182, ________23183, ________23184, ________23185,
       ________23186, ________23187, ________23188, ________23191;
  wire ________23192, ________23193, ________23194, ________23195,
       ________23196, ________23197, ________23198, ________23200;
  wire ________23201, ________23202, ________23203, ________23204,
       ________23205, ________23206, ________23207, ________23209;
  wire ________23210, ________23211, ________23212, ________23213,
       ________23216, ________23217, ________23218, ________23219;
  wire ________23220, ________23221, ________23222, ________23224,
       ________23225, ________23226, ________23227, ________23228;
  wire ________23229, ________23232, ________23233, ________23234,
       ________23235, ________23236, ________23237, ________23238;
  wire ________23239, ________23242, ________23243, ________23244,
       ________23245, ________23246, ________23247, ________23248;
  wire ________23249, ________23269, ________23270, ________23271,
       ________23272, ________23273, ________23274, ________23277;
  wire ________23278, ________23279, ________23280, ________23281,
       ________23282, ________23283, ________23284, ________23287;
  wire ________23288, ________23289, ________23290, ________23291,
       ________23292, ________23295, ________23296, ________23297;
  wire ________23298, ________23299, ________23300, ________23301,
       ________23304, ________23305, ________23306, ________23307;
  wire ________23308, ________23309, ________23310, ________23313,
       ________23314, ________23315, ________23316, ________23318;
  wire ________23319, ________23320, ________23321, ________23322,
       ________23323, ________23324, ________23327, ________23328;
  wire ________23329, ________23330, ________23331, ________23332,
       ________23333, ________23334, ________23537, ________23538;
  wire ________23539, ________23540, ________23541, ________23542,
       ________23543, ________23546, ________23547, ________23548;
  wire ________23549, ________23550, ________23551, ________23552,
       ________23553, ________23556, ________23557, ________23558;
  wire ________23559, ________23560, ________23561, ________23562,
       ________23564, ________23565, ________23566, ________23567;
  wire ________23568, ________23569, ________23570, ________23573,
       ________23574, ________23575, ________23576, ________23577;
  wire ________23578, ________23579, ________23580, ________23583,
       ________23584, ________23585, ________23586, ________23587;
  wire ________23588, ________23589, ________23592, ________23593,
       ________23594, ________23595, ________23596, ________23597;
  wire ________23598, ________23599, ________23602, ________23603,
       ________23604, ________23605, ________23606, ________23607;
  wire ________23629, ________23630, ________23631, ________23632,
       ________23633, ________23634, ________23635, ________23636;
  wire ________23639, ________23640, ________23641, ________23642,
       ________23643, ________23644, ________23645, ________23647;
  wire ________23648, ________23649, ________23650, ________23651,
       ________23652, ________23653, ________23654, ________23657;
  wire ________23658, ________23659, ________23660, ________23661,
       ________23662, ________23663, ________23664, ________23667;
  wire ________23668, ________23669, ________23670, ________23671,
       ________23672, ________23673, ________23676, ________23677;
  wire ________23678, ________23679, ________23680, ________23681,
       ________23682, ________23683, ________23686, ________23687;
  wire ________23688, ________23689, ________23690, ________23691,
       ________23692, ________23693, ________23696, ________23697;
  wire ________23698, ________23699, ________23700, ________23701,
       ________23702, ________23721, ________23722, ________23723;
  wire ________23724, ________23725, ________23726, ________23729,
       ________23730, ________23731, ________23732, ________23733;
  wire ________23734, ________23735, ________23738, ________23739,
       ________23740, ________23741, ________23742, ________23743;
  wire ________23744, ________23745, ________23748, ________23749,
       ________23750, ________23751, ________23752, ________23753;
  wire ________23754, ________23757, ________23758, ________23759,
       ________23760, ________23761, ________23762, ________23763;
  wire ________23766, ________23767, ________23768, ________23769,
       ________23770, ________23771, ________23772, ________23773;
  wire ________23776, ________23777, ________23778, ________23779,
       ________23780, ________23781, ________23782, ________23783;
  wire ________23786, ________23787, ________23788, ________23789,
       ________23790, ________23812, ________23813, ________23814;
  wire ________23815, ________23816, ________23817, ________23818,
       ________23819, ________23822, ________23823, ________23824;
  wire ________23825, ________23826, ________23829, ________23830,
       ________23831, ________23832, ________23833, ________23834;
  wire ________23835, ________23838, ________23839, ________23840,
       ________23841, ________23842, ________23844, ________23845;
  wire ________23846, ________23847, ________23848, ________23849,
       ________23851, ________23852, ________23853, ________23854;
  wire ________23855, ________23856, ________23857, ________23858,
       ________23861, ________23862, ________23863, ________23864;
  wire ________23865, ________23866, ________23867, ________23869,
       ________23870, ________23871, ________23872, ________23873;
  wire ________23874, ________23875, ________23898, ________23899,
       ________23900, ________23901, ________23902, ________23903;
  wire ________23904, ________23905, ________23906, ________23907,
       ________23908, ________23909, ________23910, ________23911;
  wire ________23912, ________23913, ________23916, ________23917,
       ________23918, ________23919, ________23920, ________23921;
  wire ________23922, ________23923, ________23926, ________23927,
       ________23928, ________23929, ________23930, ________23931;
  wire ________23932, ________23934, ________23935, ________23936,
       ________23937, ________23938, ________23939, ________23940;
  wire ________23943, ________23944, ________23945, ________23946,
       ________23947, ________23948, ________23949, ________23951;
  wire ________23952, ________23953, ________23954, ________23955,
       ________23956, ________23959, ________23960, ________23961;
  wire ________23962, ________23963, ________23984, ________23985,
       ________23986, ________23987, ________23988, ________23989;
  wire ________23990, ________23993, ________23994, ________23995,
       ________23996, ________23997, ________23998, ________24000;
  wire ________24001, ________24002, ________24003, ________24004,
       ________24005, ________24006, ________24009, ________24010;
  wire ________24011, ________24012, ________24013, ________24014,
       ________24015, ________24016, ________24019, ________24020;
  wire ________24021, ________24022, ________24023, ________24024,
       ________24025, ________24028, ________24029, ________24030;
  wire ________24031, ________24032, ________24033, ________24036,
       ________24037, ________24038, ________24039, ________24040;
  wire ________24041, ________24042, ________24045, ________24046,
       ________24047, ________24048, ________24049, ________24050;
  wire ________24051, ________24073, ________24074, ________24075,
       ________24076, ________24077, ________24078, ________24079;
  wire ________24080, ________24083, ________24084, ________24085,
       ________24086, ________24087, ________24088, ________24089;
  wire ________24090, ________24093, ________24094, ________24095,
       ________24096, ________24097, ________24098, ________24099;
  wire ________24100, ________24103, ________24104, ________24105,
       ________24106, ________24107, ________24108, ________24109;
  wire ________24111, ________24112, ________24113, ________24114,
       ________24115, ________24116, ________24117, ________24118;
  wire ________24121, ________24122, ________24123, ________24124,
       ________24125, ________24126, ________24127, ________24128;
  wire ________24131, ________24132, ________24133, ________24134,
       ________24135, ________24136, ________24137, ________24138;
  wire ________24141, ________24142, ________24143, ________24144,
       ________24145, ________24146, ________24164, ________24165;
  wire ________24166, ________24167, ________24168, ________24169,
       ________24170, ________24171, ________24174, ________24175;
  wire ________24176, ________24177, ________24178, ________24179,
       ________24180, ________24183, ________24184, ________24185;
  wire ________24186, ________24187, ________24188, ________24189,
       ________24191, ________24192, ________24193, ________24194;
  wire ________24195, ________24196, ________24197, ________24200,
       ________24201, ________24202, ________24203, ________24204;
  wire ________24205, ________24206, ________24207, ________24210,
       ________24211, ________24212, ________24213, ________24214;
  wire ________24215, ________24216, ________24217, ________24220,
       ________24221, ________24222, ________24223, ________24224;
  wire ________24225, ________24226, ________24228, ________24229,
       ________24230, ________24231, ________24232, ________24233;
  wire ________24438, ________24439, ________24440, ________24441,
       ________24442, ________24443, ________24444, ________24445;
  wire ________24448, ________24449, ________24450, ________24451,
       ________24452, ________24453, ________24454, ________24455;
  wire ________24457, ________24458, ________24459, ________24460,
       ________24461, ________24462, ________24463, ________24466;
  wire ________24467, ________24468, ________24469, ________24470,
       ________24471, ________24474, ________24475, ________24476;
  wire ________24477, ________24478, ________24479, ________24482,
       ________24483, ________24484, ________24485, ________24486;
  wire ________24487, ________24488, ________24489, ________24492,
       ________24493, ________24494, ________24495, ________24496;
  wire ________24497, ________24500, ________24501, ________24502,
       ________24503, ________24504, ________24505, ________24506;
  wire ________24526, ________24527, ________24528, ________24529,
       ________24530, ________24531, ________24532, ________24535;
  wire ________24536, ________24537, ________24538, ________24539,
       ________24540, ________24542, ________24543, ________24544;
  wire ________24545, ________24546, ________24547, ________24548,
       ________24549, ________24552, ________24553, ________24554;
  wire ________24555, ________24556, ________24557, ________24558,
       ________24561, ________24562, ________24563, ________24564;
  wire ________24565, ________24566, ________24567, ________24568,
       ________24571, ________24572, ________24573, ________24574;
  wire ________24575, ________24576, ________24577, ________24580,
       ________24581, ________24582, ________24583, ________24584;
  wire ________24585, ________24586, ________24589, ________24590,
       ________24591, ________24592, ________24593, ________24594;
  wire ________24595, ________24596, ________24617, ________24618,
       ________24619, ________24620, ________24621, ________24622;
  wire ________24623, ________24624, ________24627, ________24628,
       ________24629, ________24630, ________24631, ________24632;
  wire ________24633, ________24634, ________24637, ________24638,
       ________24639, ________24640, ________24641, ________24642;
  wire ________24643, ________24644, ________24647, ________24648,
       ________24649, ________24650, ________24651, ________24652;
  wire ________24653, ________24654, ________24657, ________24658,
       ________24659, ________24660, ________24661, ________24662;
  wire ________24663, ________24664, ________24667, ________24668,
       ________24669, ________24670, ________24671, ________24672;
  wire ________24673, ________24674, ________24677, ________24678,
       ________24679, ________24680, ________24681, ________24682;
  wire ________24683, ________24685, ________24686, ________24687,
       ________24688, ________24689, ________24690, ________24691;
  wire ________24692, ________24711, ________24712, ________24713,
       ________24714, ________24715, ________24716, ________24717;
  wire ________24718, ________24721, ________24722, ________24723,
       ________24724, ________24725, ________24726, ________24727;
  wire ________24728, ________24730, ________24731, ________24732,
       ________24733, ________24734, ________24735, ________24736;
  wire ________24737, ________24740, ________24741, ________24742,
       ________24743, ________24744, ________24747, ________24748;
  wire ________24749, ________24750, ________24751, ________24752,
       ________24753, ________24754, ________24757, ________24758;
  wire ________24759, ________24760, ________24761, ________24762,
       ________24763, ________24765, ________24766, ________24767;
  wire ________24768, ________24769, ________24770, ________24773,
       ________24774, ________24775, ________24776, ________24777;
  wire ________24778, ________24779, ________24780, ________24802,
       ________24803, ________24804, ________24805, ________24806;
  wire ________24807, ________24810, ________24811, ________24812,
       ________24813, ________24814, ________24815, ________24816;
  wire ________24817, ________24820, ________24821, ________24822,
       ________24823, ________24824, ________24825, ________24826;
  wire ________24827, ________24830, ________24831, ________24832,
       ________24833, ________24834, ________24835, ________24836;
  wire ________24837, ________24839, ________24840, ________24841,
       ________24842, ________24843, ________24844, ________24845;
  wire ________24846, ________24849, ________24850, ________24851,
       ________24852, ________24853, ________24854, ________24855;
  wire ________24856, ________24858, ________24859, ________24860,
       ________24861, ________24862, ________24863, ________24864;
  wire ________24865, ________24868, ________24869, ________24870,
       ________24871, ________24872, ________24873, ________24874;
  wire ________24875, ________24897, ________24898, ________24899,
       ________24900, ________24901, ________24902, ________24903;
  wire ________24904, ________24907, ________24908, ________24909,
       ________24910, ________24911, ________24912, ________24913;
  wire ________24914, ________24917, ________24918, ________24919,
       ________24920, ________24921, ________24922, ________24923;
  wire ________24924, ________24927, ________24928, ________24929,
       ________24930, ________24931, ________24932, ________24933;
  wire ________24934, ________24937, ________24938, ________24939,
       ________24940, ________24941, ________24942, ________24943;
  wire ________24944, ________24947, ________24948, ________24949,
       ________24950, ________24951, ________24952, ________24953;
  wire ________24954, ________24957, ________24958, ________24959,
       ________24960, ________24961, ________24962, ________24963;
  wire ________24966, ________24967, ________24968, ________24969,
       ________24970, ________24971, ________24972, ________24994;
  wire ________24995, ________24996, ________24997, ________24998,
       ________24999, ________25000, ________25003, ________25004;
  wire ________25005, ________25006, ________25007, ________25008,
       ________25009, ________25010, ________25013, ________25014;
  wire ________25015, ________25016, ________25017, ________25018,
       ________25019, ________25020, ________25023, ________25024;
  wire ________25025, ________25026, ________25027, ________25028,
       ________25029, ________25030, ________25033, ________25034;
  wire ________25035, ________25036, ________25037, ________25038,
       ________25039, ________25042, ________25043, ________25044;
  wire ________25045, ________25046, ________25047, ________25048,
       ________25049, ________25052, ________25053, ________25054;
  wire ________25055, ________25056, ________25057, ________25058,
       ________25059, ________25062, ________25063, ________25064;
  wire ________25065, ________25066, ________25067, ________25068,
       ________25069, ________25091, ________25092, ________25093;
  wire ________25094, ________25095, ________25096, ________25097,
       ________25098, ________25100, ________25101, ________25102;
  wire ________25103, ________25104, ________25105, ________25106,
       ________25107, ________25110, ________25111, ________25112;
  wire ________25113, ________25114, ________25115, ________25116,
       ________25117, ________25120, ________25121, ________25122;
  wire ________25123, ________25124, ________25125, ________25128,
       ________25129, ________25130, ________25131, ________25132;
  wire ________25133, ________25134, ________25137, ________25138,
       ________25139, ________25140, ________25141, ________25142;
  wire ________25143, ________25144, ________25147, ________25148,
       ________25149, ________25150, ________25151, ________25152;
  wire ________25153, ________25154, ________25157, ________25158,
       ________25159, ________25160, ________25161, ________25162;
  wire ________25163, ________25378, ________25379, ________25380,
       ________25381, ________25382, ________25383, ________25384;
  wire ________25385, ________25388, ________25389, ________25390,
       ________25391, ________25392, ________25393, ________25394;
  wire ________25395, ________25398, ________25399, ________25400,
       ________25401, ________25402, ________25403, ________25404;
  wire ________25407, ________25408, ________25409, ________25410,
       ________25411, ________25412, ________25413, ________25414;
  wire ________25417, ________25418, ________25419, ________25420,
       ________25421, ________25422, ________25423, ________25424;
  wire ________25427, ________25428, ________25429, ________25430,
       ________25431, ________25432, ________25433, ________25434;
  wire ________25437, ________25438, ________25439, ________25440,
       ________25441, ________25442, ________25443, ________25444;
  wire ________25447, ________25448, ________25449, ________25450,
       ________25451, ________25452, ________25453, ________25473;
  wire ________25474, ________25475, ________25476, ________25477,
       ________25478, ________25479, ________25480, ________25483;
  wire ________25484, ________25485, ________25486, ________25487,
       ________25488, ________25489, ________25490, ________25493;
  wire ________25494, ________25495, ________25496, ________25497,
       ________25498, ________25499, ________25502, ________25503;
  wire ________25504, ________25505, ________25506, ________25507,
       ________25508, ________25509, ________25512, ________25513;
  wire ________25514, ________25515, ________25516, ________25517,
       ________25518, ________25521, ________25522, ________25523;
  wire ________25524, ________25525, ________25526, ________25527,
       ________25530, ________25531, ________25532, ________25533;
  wire ________25534, ________25535, ________25536, ________25537,
       ________25540, ________25541, ________25542, ________25543;
  wire ________25544, ________25545, ________25546, ________25547,
       ________25569, ________25570, ________25571, ________25572;
  wire ________25573, ________25574, ________25575, ________25576,
       ________25579, ________25580, ________25581, ________25582;
  wire ________25583, ________25584, ________25585, ________25586,
       ________25589, ________25590, ________25591, ________25592;
  wire ________25593, ________25594, ________25595, ________25598,
       ________25599, ________25600, ________25601, ________25602;
  wire ________25603, ________25604, ________25605, ________25608,
       ________25609, ________25610, ________25611, ________25612;
  wire ________25613, ________25614, ________25617, ________25618,
       ________25619, ________25620, ________25621, ________25622;
  wire ________25623, ________25626, ________25627, ________25628,
       ________25629, ________25630, ________25631, ________25632;
  wire ________25633, ________25636, ________25637, ________25638,
       ________25639, ________25640, ________25641, ________25642;
  wire ________25643, ________25666, ________25667, ________25668,
       ________25669, ________25670, ________25671, ________25672;
  wire ________25673, ________25676, ________25677, ________25678,
       ________25679, ________25680, ________25681, ________25682;
  wire ________25683, ________25686, ________25687, ________25688,
       ________25689, ________25690, ________25691, ________25692;
  wire ________25695, ________25696, ________25697, ________25698,
       ________25699, ________25700, ________25701, ________25704;
  wire ________25705, ________25706, ________25707, ________25708,
       ________25709, ________25710, ________25713, ________25714;
  wire ________25715, ________25716, ________25717, ________25718,
       ________25719, ________25722, ________25723, ________25724;
  wire ________25725, ________25726, ________25727, ________25728,
       ________25729, ________25732, ________25733, ________25734;
  wire ________25735, ________25736, ________25737, ________25738,
       ________25739, ________25761, ________25762, ________25763;
  wire ________25764, ________25765, ________25766, ________25767,
       ________25768, ________25771, ________25772, ________25773;
  wire ________25774, ________25775, ________25776, ________25777,
       ________25778, ________25781, ________25782, ________25783;
  wire ________25784, ________25785, ________25786, ________25787,
       ________25788, ________25791, ________25792, ________25793;
  wire ________25794, ________25795, ________25796, ________25797,
       ________25798, ________25801, ________25802, ________25803;
  wire ________25804, ________25805, ________25806, ________25807,
       ________25808, ________25811, ________25812, ________25813;
  wire ________25814, ________25815, ________25816, ________25817,
       ________25818, ________25821, ________25822, ________25823;
  wire ________25824, ________25825, ________25826, ________25827,
       ________25828, ________25831, ________25832, ________25833;
  wire ________25834, ________25835, ________25836, ________25837,
       ________25838, ________25861, ________25862, ________25863;
  wire ________25864, ________25865, ________25866, ________25867,
       ________25868, ________25871, ________25872, ________25873;
  wire ________25874, ________25875, ________25876, ________25877,
       ________25878, ________25881, ________25882, ________25883;
  wire ________25884, ________25885, ________25886, ________25887,
       ________25888, ________25891, ________25892, ________25893;
  wire ________25894, ________25895, ________25896, ________25897,
       ________25898, ________25900, ________25901, ________25902;
  wire ________25903, ________25904, ________25905, ________25906,
       ________25907, ________25910, ________25911, ________25912;
  wire ________25913, ________25914, ________25915, ________25916,
       ________25917, ________25920, ________25921, ________25922;
  wire ________25923, ________25924, ________25925, ________25926,
       ________25927, ________25930, ________25931, ________25932;
  wire ________25933, ________25934, ________25935, ________25936,
       ________25937, ________25958, ________25959, ________25960;
  wire ________25961, ________25962, ________25963, ________25964,
       ________25965, ________25968, ________25969, ________25970;
  wire ________25971, ________25972, ________25973, ________25974,
       ________25975, ________25978, ________25979, ________25980;
  wire ________25981, ________25982, ________25983, ________25984,
       ________25985, ________25988, ________25989, ________25990;
  wire ________25991, ________25992, ________25993, ________25994,
       ________25995, ________25998, ________25999, ________26000;
  wire ________26001, ________26002, ________26003, ________26004,
       ________26005, ________26008, ________26009, ________26010;
  wire ________26011, ________26012, ________26013, ________26014,
       ________26015, ________26018, ________26019, ________26020;
  wire ________26021, ________26022, ________26023, ________26024,
       ________26025, ________26028, ________26029, ________26030;
  wire ________26031, ________26032, ________26033, ________26034,
       ________26035, ________26058, ________26059, ________26060;
  wire ________26061, ________26062, ________26063, ________26064,
       ________26065, ________26068, ________26069, ________26070;
  wire ________26071, ________26072, ________26073, ________26074,
       ________26075, ________26078, ________26079, ________26080;
  wire ________26081, ________26082, ________26083, ________26084,
       ________26085, ________26088, ________26089, ________26090;
  wire ________26091, ________26092, ________26093, ________26094,
       ________26095, ________26098, ________26099, ________26100;
  wire ________26101, ________26102, ________26103, ________26104,
       ________26105, ________26108, ________26109, ________26110;
  wire ________26111, ________26112, ________26113, ________26114,
       ________26115, ________26118, ________26119, ________26120;
  wire ________26121, ________26122, ________26123, ________26124,
       ________26125, ________26128, ________26129, ________26130;
  wire ________26131, ________26132, ________26133, ________26134,
       ________26135, ________35107, _________0_, _________0___18904;
  wire _________9_, _________9__9_, _________9___0_,
       _________9___18903, _________9____, _________9_____,
       _________9______18799, _________9______18800;
  wire _________9______18801, _________9______18802,
       _________9______18803, _________9_______18804,
       _________9_______18805, _________9_______18806,
       _________9_______18807, _________9_______18808;
  wire _________9_______18809, _________9_______18810,
       _________9_______18811, _________9_______18812,
       _________9_______18813, _________9_______18814, _________18843,
       _________18844;
  wire _________18845, _________18846, _________18847, _________18850,
       _________18851, _________18852, _________18853, _________18854;
  wire _________18855, _________18856, _________18858, _________18859,
       _________18860, _________18861, _________18862, _________18863;
  wire _________18864, _________18866, _________28245, _________28246,
       _________28247, _________28248, _________28249, _________28250;
  wire _________28251, _________28252, _________28255, _________28256,
       _________28257, _________28258, _________28259, _________28260;
  wire _________28261, _________28264, _________28265, _________28266,
       _________28267, _________28268, _________28269, _________28270;
  wire _________28271, _________28274, _________28275, _________28276,
       _________28277, _________28278, _________28279, _________28280;
  wire _________28281, _________28284, _________28285, _________28286,
       _________28287, _________28288, _________28289, _________28290;
  wire _________28293, _________28294, _________28295, _________28296,
       _________28297, _________28298, _________28299, _________28300;
  wire _________28303, _________28304, _________28305, _________28306,
       _________28307, _________28308, _________28309, _________28312;
  wire _________28313, _________28314, _________28315, _________28316,
       _________28317, _________28318, _________28319, _________28340;
  wire _________28341, _________28342, _________28343, _________28344,
       _________28345, _________28346, _________28349, _________28350;
  wire _________28351, _________28352, _________28353, _________28354,
       _________28355, _________28356, _________28359, _________28360;
  wire _________28361, _________28362, _________28363, _________28364,
       _________28365, _________28366, _________28367, _________28368;
  wire _________28369, _________28370, _________28371, _________28372,
       _________28373, _________28374, _________28377, _________28378;
  wire _________28379, _________28380, _________28381, _________28382,
       _________28383, _________28384, _________28387, _________28388;
  wire _________28389, _________28390, _________28391, _________28392,
       _________28393, _________28394, _________28397, _________28398;
  wire _________28399, _________28400, _________28401, _________28402,
       _________28403, _________28404, _________28407, _________28408;
  wire _________28409, _________28410, _________28411, _________28412,
       _________28413, _________28414, _________28436, _________28437;
  wire _________28438, _________28439, _________28440, _________28441,
       _________28442, _________28443, _________28446, _________28447;
  wire _________28448, _________28449, _________28450, _________28451,
       _________28452, _________28453, _________28456, _________28457;
  wire _________28458, _________28459, _________28460, _________28461,
       _________28462, _________28463, _________28466, _________28467;
  wire _________28468, _________28469, _________28470, _________28471,
       _________28472, _________28473, _________28476, _________28477;
  wire _________28478, _________28479, _________28480, _________28481,
       _________28482, _________28483, _________28486, _________28487;
  wire _________28488, _________28489, _________28490, _________28491,
       _________28492, _________28495, _________28496, _________28497;
  wire _________28498, _________28499, _________28500, _________28501,
       _________28502, _________28505, _________28506, _________28507;
  wire _________28508, _________28509, _________28510, _________28511,
       _________28512, _________28533, _________28534, _________28535;
  wire _________28536, _________28537, _________28538, _________28539,
       _________28540, _________28543, _________28544, _________28545;
  wire _________28546, _________28547, _________28548, _________28549,
       _________28550, _________28552, _________28553, _________28554;
  wire _________28555, _________28556, _________28557, _________28558,
       _________28559, _________28561, _________28562, _________28563;
  wire _________28564, _________28565, _________28566, _________28567,
       _________28570, _________28571, _________28572, _________28573;
  wire _________28574, _________28575, _________28576, _________28577,
       _________28580, _________28581, _________28582, _________28583;
  wire _________28584, _________28585, _________28586, _________28587,
       _________28590, _________28591, _________28592, _________28593;
  wire _________28594, _________28595, _________28598, _________28599,
       _________28600, _________28601, _________28602, _________28603;
  wire _________28604, _________28626, _________28627, _________28628,
       _________28629, _________28630, _________28631, _________28632;
  wire _________28635, _________28636, _________28637, _________28638,
       _________28639, _________28640, _________28641, _________28644;
  wire _________28645, _________28646, _________28647, _________28648,
       _________28649, _________28650, _________28651, _________28652;
  wire _________28653, _________28654, _________28655, _________28656,
       _________28657, _________28660, _________28661, _________28662;
  wire _________28663, _________28664, _________28665, _________28666,
       _________28667, _________28669, _________28670, _________28671;
  wire _________28672, _________28673, _________28674, _________28675,
       _________28678, _________28679, _________28680, _________28681;
  wire _________28682, _________28683, _________28684, _________28687,
       _________28688, _________28689, _________28690, _________28691;
  wire _________28692, _________28693, _________28694, _________28715,
       _________28716, _________28717, _________28718, _________28719;
  wire _________28720, _________28721, _________28724, _________28725,
       _________28726, _________28727, _________28728, _________28729;
  wire _________28730, _________28731, _________28734, _________28735,
       _________28736, _________28737, _________28738, _________28739;
  wire _________28740, _________28742, _________28743, _________28744,
       _________28745, _________28746, _________28747, _________28748;
  wire _________28749, _________28752, _________28753, _________28754,
       _________28755, _________28756, _________28757, _________28758;
  wire _________28759, _________28762, _________28763, _________28764,
       _________28765, _________28766, _________28767, _________28768;
  wire _________28769, _________28772, _________28773, _________28774,
       _________28775, _________28776, _________28777, _________28778;
  wire _________28779, _________28782, _________28783, _________28784,
       _________28785, _________28786, _________28787, _________28788;
  wire _________28789, _________28811, _________28812, _________28813,
       _________28814, _________28815, _________28816, _________28817;
  wire _________28818, _________28821, _________28822, _________28823,
       _________28824, _________28825, _________28826, _________28827;
  wire _________28828, _________28831, _________28832, _________28833,
       _________28834, _________28835, _________28836, _________28837;
  wire _________28838, _________28841, _________28842, _________28843,
       _________28844, _________28845, _________28846, _________28847;
  wire _________28848, _________28851, _________28852, _________28853,
       _________28854, _________28855, _________28856, _________28857;
  wire _________28858, _________28861, _________28862, _________28863,
       _________28864, _________28865, _________28866, _________28867;
  wire _________28870, _________28871, _________28872, _________28873,
       _________28874, _________28875, _________28876, _________28879;
  wire _________28880, _________28881, _________28882, _________28883,
       _________28884, _________28885, _________28886, _________28908;
  wire _________28909, _________28910, _________28911, _________28912,
       _________28913, _________28914, _________28915, _________28918;
  wire _________28919, _________28920, _________28921, _________28922,
       _________28923, _________28924, _________28926, _________28927;
  wire _________28928, _________28929, _________28930, _________28931,
       _________28932, _________28933, _________28936, _________28937;
  wire _________28938, _________28939, _________28940, _________28941,
       _________28942, _________28943, _________28946, _________28947;
  wire _________28948, _________28949, _________28950, _________28951,
       _________28952, _________28953, _________28956, _________28957;
  wire _________28958, _________28959, _________28960, _________28961,
       _________28962, _________28963, _________28966, _________28967;
  wire _________28968, _________28969, _________28970, _________28971,
       _________28972, _________28975, _________28976, _________28977;
  wire _________28978, _________28979, _________28980, _________28981,
       _________29187, _________29188, _________29189, _________29190;
  wire _________29191, _________29192, _________29193, _________29194,
       _________29197, _________29198, _________29199, _________29200;
  wire _________29201, _________29204, _________29205, _________29206,
       _________29207, _________29208, _________29209, _________29210;
  wire _________29213, _________29214, _________29215, _________29216,
       _________29217, _________29218, _________29219, _________29222;
  wire _________29223, _________29224, _________29225, _________29226,
       _________29227, _________29228, _________29231, _________29232;
  wire _________29233, _________29234, _________29235, _________29236,
       _________29237, _________29240, _________29241, _________29242;
  wire _________29243, _________29244, _________29245, _________29248,
       _________29249, _________29250, _________29251, _________29252;
  wire _________29253, _________29254, _________29276, _________29277,
       _________29278, _________29279, _________29280, _________29281;
  wire _________29284, _________29285, _________29286, _________29287,
       _________29288, _________29289, _________29290, _________29291;
  wire _________29294, _________29295, _________29296, _________29297,
       _________29298, _________29299, _________29302, _________29303;
  wire _________29304, _________29305, _________29306, _________29307,
       _________29308, _________29311, _________29312, _________29313;
  wire _________29314, _________29315, _________29316, _________29317,
       _________29318, _________29321, _________29322, _________29323;
  wire _________29324, _________29325, _________29326, _________29327,
       _________29328, _________29330, _________29331, _________29332;
  wire _________29333, _________29334, _________29335, _________29336,
       _________29337, _________29340, _________29341, _________29342;
  wire _________29343, _________29344, _________29345, _________29346,
       _________29347, _________29366, _________29367, _________29368;
  wire _________29369, _________29370, _________29371, _________29372,
       _________29373, _________29376, _________29377, _________29378;
  wire _________29379, _________29380, _________29381, _________29382,
       _________29383, _________29386, _________29387, _________29388;
  wire _________29389, _________29390, _________29391, _________29392,
       _________29393, _________29395, _________29396, _________29397;
  wire _________29398, _________29399, _________29400, _________29401,
       _________29404, _________29405, _________29406, _________29407;
  wire _________29408, _________29409, _________29410, _________29411,
       _________29412, _________29413, _________29414, _________29415;
  wire _________29416, _________29417, _________29418, _________29421,
       _________29422, _________29423, _________29424, _________29425;
  wire _________29426, _________29427, _________29430, _________29431,
       _________29432, _________29433, _________29434, _________29435;
  wire _________29436, _________29457, _________29458, _________29459,
       _________29460, _________29461, _________29462, _________29463;
  wire _________29464, _________29467, _________29468, _________29469,
       _________29470, _________29471, _________29472, _________29473;
  wire _________29474, _________29477, _________29478, _________29479,
       _________29480, _________29481, _________29482, _________29483;
  wire _________29485, _________29486, _________29487, _________29488,
       _________29489, _________29490, _________29492, _________29493;
  wire _________29494, _________29495, _________29496, _________29497,
       _________29498, _________29499, _________29500, _________29503;
  wire _________29504, _________29505, _________29506, _________29507,
       _________29508, _________29509, _________29510, _________29513;
  wire _________29514, _________29515, _________29516, _________29517,
       _________29518, _________29519, _________29520, _________29538;
  wire _________29539, _________29540, _________29541, _________29542,
       _________29543, _________29546, _________29547, _________29548;
  wire _________29549, _________29550, _________29551, _________29552,
       _________29554, _________29555, _________29556, _________29557;
  wire _________29558, _________29559, _________29560, _________29563,
       _________29564, _________29565, _________29566, _________29567;
  wire _________29568, _________29569, _________29572, _________29573,
       _________29574, _________29575, _________29576, _________29577;
  wire _________29578, _________29581, _________29582, _________29583,
       _________29584, _________29585, _________29586, _________29587;
  wire _________29589, _________29590, _________29591, _________29592,
       _________29593, _________29594, _________29595, _________29598;
  wire _________29599, _________29600, _________29601, _________29602,
       _________29603, _________29604, _________29625, _________29626;
  wire _________29627, _________29628, _________29629, _________29630,
       _________29631, _________29632, _________29635, _________29636;
  wire _________29637, _________29638, _________29639, _________29640,
       _________29641, _________29642, _________29644, _________29645;
  wire _________29646, _________29647, _________29648, _________29649,
       _________29650, _________29653, _________29654, _________29655;
  wire _________29656, _________29657, _________29658, _________29659,
       _________29660, _________29663, _________29664, _________29665;
  wire _________29666, _________29667, _________29668, _________29669,
       _________29672, _________29673, _________29674, _________29675;
  wire _________29676, _________29677, _________29678, _________29681,
       _________29682, _________29683, _________29684, _________29685;
  wire _________29686, _________29687, _________29688, _________29691,
       _________29692, _________29693, _________29694, _________29695;
  wire _________29696, _________29697, _________29698, _________29720,
       _________29721, _________29722, _________29723, _________29724;
  wire _________29725, _________29726, _________29727, _________29730,
       _________29731, _________29732, _________29733, _________29734;
  wire _________29735, _________29736, _________29737, _________29740,
       _________29741, _________29742, _________29743, _________29744;
  wire _________29745, _________29746, _________29748, _________29749,
       _________29750, _________29751, _________29752, _________29753;
  wire _________29754, _________29755, _________29758, _________29759,
       _________29760, _________29761, _________29762, _________29763;
  wire _________29764, _________29767, _________29768, _________29769,
       _________29770, _________29771, _________29772, _________29773;
  wire _________29774, _________29777, _________29778, _________29779,
       _________29780, _________29781, _________29782, _________29783;
  wire _________29784, _________29785, _________29786, _________29787,
       _________29788, _________29789, _________29790, _________29791;
  wire _________29814, _________29815, _________29816, _________29817,
       _________29818, _________29819, _________29820, _________29821;
  wire _________29824, _________29825, _________29826, _________29827,
       _________29828, _________29829, _________29830, _________29831;
  wire _________29834, _________29835, _________29836, _________29837,
       _________29838, _________29839, _________29840, _________29842;
  wire _________29843, _________29844, _________29845, _________29846,
       _________29847, _________29848, _________29849, _________29852;
  wire _________29853, _________29854, _________29855, _________29856,
       _________29857, _________29858, _________29859, _________29862;
  wire _________29863, _________29864, _________29865, _________29866,
       _________29867, _________29868, _________29869, _________29872;
  wire _________29873, _________29874, _________29875, _________29876,
       _________29877, _________29878, _________29879, _________29882;
  wire _________29883, _________29884, _________29885, _________29886,
       _________29887, _________29888, _________29889, _________30104;
  wire _________30105, _________30106, _________30107, _________30108,
       _________30109, _________30110, _________30113, _________30114;
  wire _________30115, _________30116, _________30117, _________30118,
       _________30119, _________30120, _________30122, _________30123;
  wire _________30124, _________30125, _________30126, _________30128,
       _________30129, _________30130, _________30131, _________30132;
  wire _________30133, _________30134, _________30137, _________30138,
       _________30139, _________30140, _________30141, _________30144;
  wire _________30145, _________30146, _________30147, _________30148,
       _________30149, _________30150, _________30151, _________30153;
  wire _________30154, _________30155, _________30156, _________30157,
       _________30158, _________30159, _________30160, _________30163;
  wire _________30164, _________30165, _________30166, _________30167,
       _________30168, _________30189, _________30190, _________30191;
  wire _________30192, _________30193, _________30194, _________30195,
       _________30196, _________30199, _________30200, _________30201;
  wire _________30202, _________30203, _________30204, _________30205,
       _________30206, _________30209, _________30210, _________30211;
  wire _________30212, _________30213, _________30214, _________30215,
       _________30218, _________30219, _________30220, _________30221;
  wire _________30222, _________30223, _________30224, _________30225,
       _________30228, _________30229, _________30230, _________30231;
  wire _________30232, _________30233, _________30234, _________30235,
       _________30238, _________30239, _________30240, _________30241;
  wire _________30242, _________30243, _________30244, _________30247,
       _________30248, _________30249, _________30250, _________30251;
  wire _________30252, _________30253, _________30256, _________30257,
       _________30258, _________30259, _________30260, _________30261;
  wire _________30262, _________30263, _________30284, _________30285,
       _________30286, _________30287, _________30288, _________30289;
  wire _________30292, _________30293, _________30294, _________30295,
       _________30296, _________30297, _________30300, _________30301;
  wire _________30302, _________30303, _________30304, _________30305,
       _________30306, _________30307, _________30310, _________30311;
  wire _________30312, _________30313, _________30314, _________30315,
       _________30316, _________30319, _________30320, _________30321;
  wire _________30322, _________30323, _________30324, _________30325,
       _________30328, _________30329, _________30330, _________30331;
  wire _________30332, _________30333, _________30336, _________30337,
       _________30338, _________30339, _________30340, _________30341;
  wire _________30342, _________30343, _________30346, _________30347,
       _________30348, _________30349, _________30350, _________30351;
  wire _________30352, _________30374, _________30375, _________30376,
       _________30377, _________30378, _________30379, _________30380;
  wire _________30383, _________30384, _________30385, _________30386,
       _________30387, _________30388, _________30389, _________30390;
  wire _________30392, _________30393, _________30394, _________30395,
       _________30396, _________30397, _________30400, _________30401;
  wire _________30402, _________30403, _________30404, _________30405,
       _________30406, _________30407, _________30410, _________30411;
  wire _________30412, _________30413, _________30414, _________30415,
       _________30416, _________30419, _________30420, _________30421;
  wire _________30422, _________30423, _________30424, _________30425,
       _________30428, _________30429, _________30430, _________30431;
  wire _________30432, _________30433, _________30434, _________30435,
       _________30438, _________30439, _________30440, _________30441;
  wire _________30442, _________30443, _________30444, _________30445,
       _________30466, _________30467, _________30468, _________30469;
  wire _________30470, _________30471, _________30472, _________30473,
       _________30476, _________30477, _________30478, _________30479;
  wire _________30480, _________30481, _________30482, _________30483,
       _________30486, _________30487, _________30488, _________30489;
  wire _________30490, _________30491, _________30492, _________30495,
       _________30496, _________30497, _________30498, _________30499;
  wire _________30501, _________30502, _________30503, _________30504,
       _________30505, _________30506, _________30507, _________30508;
  wire _________30511, _________30512, _________30513, _________30514,
       _________30515, _________30516, _________30517, _________30518;
  wire _________30521, _________30522, _________30523, _________30524,
       _________30525, _________30526, _________30527, _________30528;
  wire _________30531, _________30532, _________30533, _________30534,
       _________30535, _________30536, _________30556, _________30557;
  wire _________30558, _________30559, _________30560, _________30561,
       _________30562, _________30563, _________30565, _________30566;
  wire _________30567, _________30568, _________30569, _________30570,
       _________30571, _________30572, _________30575, _________30576;
  wire _________30577, _________30578, _________30579, _________30580,
       _________30583, _________30584, _________30585, _________30586;
  wire _________30587, _________30588, _________30589, _________30592,
       _________30593, _________30594, _________30595, _________30596;
  wire _________30597, _________30598, _________30601, _________30602,
       _________30603, _________30604, _________30605, _________30608;
  wire _________30609, _________30610, _________30611, _________30612,
       _________30613, _________30614, _________30615, _________30616;
  wire _________30617, _________30618, _________30619, _________30620,
       _________30621, _________30643, _________30644, _________30645;
  wire _________30646, _________30647, _________30648, _________30649,
       _________30650, _________30653, _________30654, _________30655;
  wire _________30656, _________30657, _________30658, _________30659,
       _________30660, _________30663, _________30664, _________30665;
  wire _________30666, _________30667, _________30668, _________30669,
       _________30672, _________30673, _________30674, _________30675;
  wire _________30676, _________30677, _________30678, _________30681,
       _________30682, _________30683, _________30684, _________30685;
  wire _________30686, _________30687, _________30688, _________30690,
       _________30691, _________30692, _________30693, _________30694;
  wire _________30695, _________30696, _________30699, _________30700,
       _________30701, _________30702, _________30703, _________30704;
  wire _________30705, _________30706, _________30709, _________30710,
       _________30711, _________30712, _________30713, _________30714;
  wire _________30715, _________30737, _________30738, _________30739,
       _________30740, _________30741, _________30742, _________30743;
  wire _________30746, _________30747, _________30748, _________30749,
       _________30750, _________30751, _________30752, _________30753;
  wire _________30755, _________30756, _________30757, _________30758,
       _________30759, _________30760, _________30761, _________30762;
  wire _________30765, _________30766, _________30767, _________30768,
       _________30769, _________30770, _________30771, _________30772;
  wire _________30775, _________30776, _________30777, _________30778,
       _________30779, _________30780, _________30781, _________30782;
  wire _________30785, _________30786, _________30787, _________30788,
       _________30789, _________30790, _________30792, _________30793;
  wire _________30794, _________30795, _________30796, _________30797,
       _________30798, _________30799, _________30801, _________30802;
  wire _________30803, _________30804, _________30805, _________30806,
       _________30807, _________30808, _________31008, _________31009;
  wire _________31010, _________31011, _________31012, _________31013,
       _________31014, _________31017, _________31018, _________31019;
  wire _________31020, _________31021, _________31022, _________31023,
       _________31026, _________31027, _________31028, _________31029;
  wire _________31030, _________31031, _________31032, _________31033,
       _________31036, _________31037, _________31038, _________31039;
  wire _________31040, _________31041, _________31042, _________31045,
       _________31046, _________31047, _________31048, _________31049;
  wire _________31050, _________31051, _________31052, _________31055,
       _________31056, _________31057, _________31058, _________31059;
  wire _________31060, _________31061, _________31062, _________31065,
       _________31066, _________31067, _________31068, _________31069;
  wire _________31070, _________31071, _________31072, _________31075,
       _________31076, _________31077, _________31078, _________31079;
  wire _________31080, _________31081, _________31082, _________31102,
       _________31103, _________31104, _________31105, _________31106;
  wire _________31107, _________31108, _________31109, _________31112,
       _________31113, _________31114, _________31115, _________31116;
  wire _________31117, _________31118, _________31119, _________31122,
       _________31123, _________31124, _________31125, _________31126;
  wire _________31127, _________31128, _________31131, _________31132,
       _________31133, _________31134, _________31135, _________31136;
  wire _________31137, _________31138, _________31141, _________31142,
       _________31143, _________31144, _________31145, _________31146;
  wire _________31147, _________31150, _________31151, _________31152,
       _________31153, _________31154, _________31155, _________31156;
  wire _________31157, _________31160, _________31161, _________31162,
       _________31163, _________31164, _________31165, _________31168;
  wire _________31169, _________31170, _________31171, _________31172,
       _________31173, _________31194, _________31195, _________31196;
  wire _________31197, _________31198, _________31199, _________31202,
       _________31203, _________31204, _________31205, _________31206;
  wire _________31207, _________31208, _________31209, _________31212,
       _________31213, _________31214, _________31215, _________31216;
  wire _________31217, _________31218, _________31220, _________31221,
       _________31222, _________31223, _________31224, _________31225;
  wire _________31226, _________31227, _________31230, _________31231,
       _________31232, _________31233, _________31234, _________31235;
  wire _________31236, _________31239, _________31240, _________31241,
       _________31242, _________31243, _________31244, _________31245;
  wire _________31248, _________31249, _________31250, _________31251,
       _________31252, _________31255, _________31256, _________31257;
  wire _________31258, _________31259, _________31260, _________31261,
       _________31279, _________31280, _________31281, _________31282;
  wire _________31283, _________31284, _________31285, _________31287,
       _________31288, _________31289, _________31290, _________31291;
  wire _________31294, _________31295, _________31296, _________31297,
       _________31300, _________31301, _________31302, _________31303;
  wire _________31304, _________31305, _________31306, _________31307,
       _________31310, _________31311, _________31312, _________31313;
  wire _________31314, _________31315, _________31318, _________31319,
       _________31320, _________31321, _________31322, _________31323;
  wire _________31326, _________31327, _________31328, _________31329,
       _________31330, _________31331, _________31332, _________31335;
  wire _________31336, _________31337, _________31338, _________31339,
       _________31340, _________31341, _________31342, _________31361;
  wire _________31362, _________31363, _________31364, _________31365,
       _________31366, _________31367, _________31368, _________31371;
  wire _________31372, _________31373, _________31374, _________31375,
       _________31376, _________31377, _________31378, _________31381;
  wire _________31382, _________31383, _________31384, _________31385,
       _________31386, _________31387, _________31388, _________31391;
  wire _________31392, _________31393, _________31394, _________31395,
       _________31396, _________31397, _________31398, _________31401;
  wire _________31402, _________31403, _________31404, _________31405,
       _________31406, _________31407, _________31408, _________31411;
  wire _________31412, _________31413, _________31414, _________31415,
       _________31416, _________31417, _________31420, _________31421;
  wire _________31422, _________31423, _________31424, _________31425,
       _________31428, _________31429, _________31430, _________31431;
  wire _________31432, _________31433, _________31434, _________31435,
       _________31457, _________31458, _________31459, _________31460;
  wire _________31461, _________31462, _________31463, _________31464,
       _________31467, _________31468, _________31469, _________31470;
  wire _________31471, _________31472, _________31475, _________31476,
       _________31477, _________31478, _________31479, _________31480;
  wire _________31483, _________31484, _________31485, _________31486,
       _________31487, _________31488, _________31489, _________31492;
  wire _________31493, _________31494, _________31495, _________31496,
       _________31497, _________31498, _________31499, _________31502;
  wire _________31503, _________31504, _________31505, _________31506,
       _________31507, _________31508, _________31509, _________31512;
  wire _________31513, _________31514, _________31515, _________31516,
       _________31517, _________31518, _________31519, _________31520;
  wire _________31521, _________31522, _________31523, _________31524,
       _________31545, _________31546, _________31547, _________31548;
  wire _________31549, _________31550, _________31551, _________31552,
       _________31555, _________31556, _________31557, _________31558;
  wire _________31559, _________31560, _________31561, _________31562,
       _________31565, _________31566, _________31567, _________31568;
  wire _________31569, _________31570, _________31571, _________31572,
       _________31575, _________31576, _________31577, _________31578;
  wire _________31579, _________31580, _________31581, _________31584,
       _________31585, _________31586, _________31587, _________31588;
  wire _________31589, _________31590, _________31591, _________31594,
       _________31595, _________31596, _________31597, _________31598;
  wire _________31599, _________31600, _________31603, _________31604,
       _________31605, _________31606, _________31607, _________31608;
  wire _________31609, _________31610, _________31613, _________31614,
       _________31615, _________31616, _________31617, _________31618;
  wire _________31619, _________31620, _________31642, _________31643,
       _________31644, _________31645, _________31646, _________31647;
  wire _________31648, _________31651, _________31652, _________31653,
       _________31654, _________31655, _________31656, _________31657;
  wire _________31660, _________31661, _________31662, _________31663,
       _________31664, _________31665, _________31666, _________31667;
  wire _________31670, _________31671, _________31672, _________31673,
       _________31674, _________31675, _________31676, _________31679;
  wire _________31680, _________31681, _________31682, _________31683,
       _________31684, _________31687, _________31688, _________31689;
  wire _________31690, _________31691, _________31692, _________31693,
       _________31694, _________31697, _________31698, _________31699;
  wire _________31700, _________31701, _________31702, _________31703,
       _________31704, _________31707, _________31708, _________31709;
  wire _________31710, _________31711, _________31712, _________31713,
       _________31911, _________31912, _________31913, _________31914;
  wire _________31915, _________31916, _________31917, _________31920,
       _________31921, _________31922, _________31923, _________31924;
  wire _________31925, _________31926, _________31927, _________31930,
       _________31931, _________31932, _________31933, _________31934;
  wire _________31935, _________31936, _________31937, _________31939,
       _________31940, _________31941, _________31942, _________31943;
  wire _________31944, _________31945, _________31946, _________31949,
       _________31950, _________31951, _________31952, _________31953;
  wire _________31954, _________31955, _________31956, _________31959,
       _________31960, _________31961, _________31962, _________31963;
  wire _________31964, _________31965, _________31966, _________31969,
       _________31970, _________31971, _________31972, _________31973;
  wire _________31974, _________31975, _________31978, _________31979,
       _________31980, _________31981, _________31982, _________31983;
  wire _________31984, _________31985, _________32007, _________32008,
       _________32009, _________32010, _________32011, _________32012;
  wire _________32013, _________32014, _________32017, _________32018,
       _________32019, _________32020, _________32021, _________32022;
  wire _________32023, _________32024, _________32027, _________32028,
       _________32029, _________32030, _________32031, _________32032;
  wire _________32033, _________32034, _________32037, _________32038,
       _________32039, _________32040, _________32041, _________32042;
  wire _________32043, _________32044, _________32047, _________32048,
       _________32049, _________32050, _________32051, _________32052;
  wire _________32053, _________32054, _________32057, _________32058,
       _________32059, _________32060, _________32061, _________32062;
  wire _________32063, _________32064, _________32067, _________32068,
       _________32069, _________32070, _________32071, _________32072;
  wire _________32073, _________32074, _________32077, _________32078,
       _________32079, _________32080, _________32081, _________32082;
  wire _________32083, _________32084, _________32107, _________32108,
       _________32109, _________32110, _________32111, _________32112;
  wire _________32113, _________32114, _________32117, _________32118,
       _________32119, _________32120, _________32121, _________32122;
  wire _________32123, _________32124, _________32127, _________32128,
       _________32129, _________32130, _________32131, _________32132;
  wire _________32133, _________32136, _________32137, _________32138,
       _________32139, _________32140, _________32141, _________32142;
  wire _________32143, _________32146, _________32147, _________32148,
       _________32149, _________32150, _________32151, _________32152;
  wire _________32153, _________32156, _________32157, _________32158,
       _________32159, _________32160, _________32161, _________32162;
  wire _________32165, _________32166, _________32167, _________32168,
       _________32169, _________32170, _________32171, _________32172;
  wire _________32175, _________32176, _________32177, _________32178,
       _________32179, _________32180, _________32181, _________32182;
  wire _________32204, _________32205, _________32206, _________32207,
       _________32208, _________32209, _________32210, _________32211;
  wire _________32214, _________32215, _________32216, _________32217,
       _________32218, _________32219, _________32220, _________32221;
  wire _________32224, _________32225, _________32226, _________32227,
       _________32228, _________32229, _________32230, _________32231;
  wire _________32234, _________32235, _________32236, _________32237,
       _________32238, _________32239, _________32240, _________32241;
  wire _________32244, _________32245, _________32246, _________32247,
       _________32248, _________32249, _________32250, _________32253;
  wire _________32254, _________32255, _________32256, _________32257,
       _________32258, _________32259, _________32260, _________32263;
  wire _________32264, _________32265, _________32266, _________32267,
       _________32268, _________32269, _________32270, _________32273;
  wire _________32274, _________32275, _________32276, _________32277,
       _________32278, _________32279, _________32280, _________32303;
  wire _________32304, _________32305, _________32306, _________32307,
       _________32308, _________32309, _________32312, _________32313;
  wire _________32314, _________32315, _________32316, _________32317,
       _________32318, _________32319, _________32322, _________32323;
  wire _________32324, _________32325, _________32326, _________32327,
       _________32328, _________32329, _________32332, _________32333;
  wire _________32334, _________32335, _________32336, _________32337,
       _________32338, _________32339, _________32342, _________32343;
  wire _________32344, _________32345, _________32346, _________32347,
       _________32348, _________32349, _________32352, _________32353;
  wire _________32354, _________32355, _________32356, _________32357,
       _________32358, _________32359, _________32361, _________32362;
  wire _________32363, _________32364, _________32365, _________32366,
       _________32367, _________32368, _________32371, _________32372;
  wire _________32373, _________32374, _________32375, _________32376,
       _________32397, _________32398, _________32399, _________32400;
  wire _________32401, _________32402, _________32403, _________32404,
       _________32407, _________32408, _________32409, _________32410;
  wire _________32411, _________32412, _________32413, _________32414,
       _________32417, _________32418, _________32419, _________32420;
  wire _________32421, _________32422, _________32423, _________32424,
       _________32427, _________32428, _________32429, _________32430;
  wire _________32431, _________32432, _________32433, _________32434,
       _________32437, _________32438, _________32439, _________32440;
  wire _________32441, _________32442, _________32443, _________32446,
       _________32447, _________32448, _________32449, _________32450;
  wire _________32451, _________32452, _________32454, _________32455,
       _________32456, _________32457, _________32458, _________32459;
  wire _________32462, _________32463, _________32464, _________32465,
       _________32466, _________32467, _________32487, _________32488;
  wire _________32489, _________32490, _________32491, _________32492,
       _________32493, _________32494, _________32497, _________32498;
  wire _________32499, _________32500, _________32501, _________32502,
       _________32503, _________32504, _________32507, _________32508;
  wire _________32509, _________32510, _________32511, _________32512,
       _________32513, _________32516, _________32517, _________32518;
  wire _________32519, _________32520, _________32521, _________32522,
       _________32525, _________32526, _________32527, _________32528;
  wire _________32529, _________32530, _________32531, _________32533,
       _________32534, _________32535, _________32536, _________32537;
  wire _________32538, _________32539, _________32542, _________32543,
       _________32544, _________32545, _________32546, _________32547;
  wire _________32548, _________32551, _________32552, _________32553,
       _________32554, _________32555, _________32556, _________32557;
  wire _________32558, _________32577, _________32578, _________32579,
       _________32580, _________32581, _________32582, _________32583;
  wire _________32584, _________32587, _________32588, _________32589,
       _________32590, _________32591, _________32592, _________32595;
  wire _________32596, _________32597, _________32598, _________32599,
       _________32600, _________32603, _________32604, _________32605;
  wire _________32606, _________32607, _________32608, _________32609,
       _________32612, _________32613, _________32614, _________32615;
  wire _________32616, _________32617, _________32618, _________32619,
       _________32622, _________32623, _________32624, _________32625;
  wire _________32626, _________32627, _________32629, _________32630,
       _________32631, _________32632, _________32633, _________32634;
  wire _________32635, _________32638, _________32639, _________32640,
       _________32641, _________32642, _________32643, _________32644;
  wire _________32645, _________32858, _________32859, _________32860,
       _________32861, _________32862, _________32864, _________32865;
  wire _________32866, _________32867, _________32868, _________32869,
       _________32870, _________32871, _________32874, _________32875;
  wire _________32876, _________32877, _________32878, _________32879,
       _________32882, _________32883, _________32884, _________32885;
  wire _________32886, _________32887, _________32888, _________32891,
       _________32892, _________32893, _________32894, _________32895;
  wire _________32896, _________32897, _________32900, _________32901,
       _________32902, _________32903, _________32904, _________32905;
  wire _________32906, _________32907, _________32910, _________32911,
       _________32912, _________32913, _________32914, _________32915;
  wire _________32916, _________32919, _________32920, _________32921,
       _________32922, _________32923, _________32924, _________32925;
  wire _________32926, _________32946, _________32947, _________32948,
       _________32949, _________32950, _________32951, _________32952;
  wire _________32953, _________32955, _________32956, _________32957,
       _________32958, _________32959, _________32960, _________32961;
  wire _________32962, _________32965, _________32966, _________32967,
       _________32968, _________32969, _________32970, _________32971;
  wire _________32972, _________32975, _________32976, _________32977,
       _________32978, _________32979, _________32980, _________32981;
  wire _________32982, _________32985, _________32986, _________32987,
       _________32988, _________32989, _________32990, _________32993;
  wire _________32994, _________32995, _________32996, _________32997,
       _________32998, _________32999, _________33001, _________33002;
  wire _________33003, _________33004, _________33005, _________33006,
       _________33007, _________33008, _________33011, _________33012;
  wire _________33013, _________33014, _________33015, _________33016,
       _________33017, _________33018, _________33040, _________33041;
  wire _________33042, _________33043, _________33044, _________33045,
       _________33046, _________33049, _________33050, _________33051;
  wire _________33052, _________33053, _________33054, _________33055,
       _________33056, _________33059, _________33060, _________33061;
  wire _________33062, _________33063, _________33064, _________33065,
       _________33066, _________33068, _________33069, _________33070;
  wire _________33071, _________33072, _________33073, _________33074,
       _________33075, _________33078, _________33079, _________33080;
  wire _________33081, _________33082, _________33083, _________33084,
       _________33085, _________33088, _________33089, _________33090;
  wire _________33091, _________33092, _________33093, _________33094,
       _________33095, _________33098, _________33099, _________33100;
  wire _________33101, _________33102, _________33103, _________33104,
       _________33105, _________33108, _________33109, _________33110;
  wire _________33111, _________33112, _________33113, _________33114,
       _________33115, _________33137, _________33138, _________33139;
  wire _________33140, _________33141, _________33142, _________33143,
       _________33144, _________33147, _________33148, _________33149;
  wire _________33150, _________33151, _________33152, _________33153,
       _________33154, _________33157, _________33158, _________33159;
  wire _________33160, _________33161, _________33162, _________33163,
       _________33164, _________33167, _________33168, _________33169;
  wire _________33170, _________33171, _________33172, _________33173,
       _________33174, _________33176, _________33177, _________33178;
  wire _________33179, _________33180, _________33181, _________33182,
       _________33185, _________33186, _________33187, _________33188;
  wire _________33189, _________33190, _________33191, _________33194,
       _________33195, _________33196, _________33197, _________33198;
  wire _________33199, _________33200, _________33201, _________33204,
       _________33205, _________33206, _________33207, _________33208;
  wire _________33209, _________33210, _________33211, _________33230,
       _________33231, _________33232, _________33233, _________33234;
  wire _________33235, _________33236, _________33237, _________33240,
       _________33241, _________33242, _________33243, _________33244;
  wire _________33245, _________33246, _________33249, _________33250,
       _________33251, _________33252, _________33253, _________33254;
  wire _________33255, _________33256, _________33259, _________33260,
       _________33261, _________33262, _________33263, _________33264;
  wire _________33265, _________33267, _________33268, _________33269,
       _________33270, _________33271, _________33272, _________33273;
  wire _________33274, _________33277, _________33278, _________33279,
       _________33280, _________33281, _________33282, _________33285;
  wire _________33286, _________33287, _________33288, _________33289,
       _________33290, _________33293, _________33294, _________33295;
  wire _________33296, _________33297, _________33298, _________33299,
       _________33300, _________33319, _________33320, _________33321;
  wire _________33322, _________33323, _________33324, _________33325,
       _________33328, _________33329, _________33330, _________33331;
  wire _________33332, _________33333, _________33334, _________33337,
       _________33338, _________33339, _________33340, _________33341;
  wire _________33342, _________33343, _________33345, _________33346,
       _________33347, _________33348, _________33349, _________33350;
  wire _________33351, _________33352, _________33355, _________33356,
       _________33357, _________33358, _________33359, _________33360;
  wire _________33361, _________33362, _________33364, _________33365,
       _________33366, _________33367, _________33368, _________33369;
  wire _________33370, _________33371, _________33374, _________33375,
       _________33376, _________33377, _________33378, _________33379;
  wire _________33380, _________33381, _________33384, _________33385,
       _________33386, _________33387, _________33388, _________33389;
  wire _________33410, _________33411, _________33412, _________33413,
       _________33414, _________33415, _________33416, _________33417;
  wire _________33420, _________33421, _________33422, _________33423,
       _________33424, _________33425, _________33426, _________33427;
  wire _________33430, _________33431, _________33432, _________33433,
       _________33434, _________33435, _________33438, _________33439;
  wire _________33440, _________33441, _________33442, _________33443,
       _________33444, _________33445, _________33447, _________33448;
  wire _________33449, _________33450, _________33451, _________33452,
       _________33455, _________33456, _________33457, _________33458;
  wire _________33459, _________33460, _________33461, _________33462,
       _________33465, _________33466, _________33467, _________33468;
  wire _________33469, _________33470, _________33471, _________33474,
       _________33475, _________33476, _________33477, _________33478;
  wire _________33498, _________33499, _________33500, _________33501,
       _________33502, _________33503, _________33504, _________33507;
  wire _________33508, _________33509, _________33510, _________33511,
       _________33512, _________33513, _________33515, _________33516;
  wire _________33517, _________33518, _________33519, _________33520,
       _________33521, _________33522, _________33525, _________33526;
  wire _________33527, _________33528, _________33529, _________33530,
       _________33531, _________33534, _________33535, _________33536;
  wire _________33537, _________33538, _________33539, _________33540,
       _________33541, _________33544, _________33545, _________33546;
  wire _________33547, _________33548, _________33549, _________33550,
       _________33551, _________33554, _________33555, _________33556;
  wire _________33557, _________33558, _________33559, _________33562,
       _________33563, _________33564, _________33565, _________33566;
  wire _________33567, _________33780, _________33781, _________33782,
       _________33783, _________33784, _________33785, _________33786;
  wire _________33787, _________33790, _________33791, _________33792,
       _________33793, _________33794, _________33795, _________33796;
  wire _________33797, _________33800, _________33801, _________33802,
       _________33803, _________33804, _________33805, _________33806;
  wire _________33807, _________33810, _________33811, _________33812,
       _________33813, _________33814, _________33815, _________33816;
  wire _________33817, _________33820, _________33821, _________33822,
       _________33823, _________33824, _________33825, _________33826;
  wire _________33827, _________33830, _________33831, _________33832,
       _________33833, _________33834, _________33835, _________33836;
  wire _________33837, _________33840, _________33841, _________33842,
       _________33843, _________33844, _________33845, _________33846;
  wire _________33847, _________33849, _________33850, _________33851,
       _________33852, _________33853, _________33854, _________33855;
  wire _________33875, _________33876, _________33877, _________33878,
       _________33879, _________33880, _________33881, _________33884;
  wire _________33885, _________33886, _________33887, _________33888,
       _________33889, _________33890, _________33891, _________33894;
  wire _________33895, _________33896, _________33897, _________33898,
       _________33901, _________33902, _________33903, _________33904;
  wire _________33905, _________33906, _________33907, _________33910,
       _________33911, _________33912, _________33913, _________33914;
  wire _________33915, _________33916, _________33919, _________33920,
       _________33921, _________33922, _________33923, _________33924;
  wire _________33925, _________33927, _________33928, _________33929,
       _________33930, _________33931, _________33932, _________33933;
  wire _________33936, _________33937, _________33938, _________33939,
       _________33940, _________33941, _________33942, _________33964;
  wire _________33965, _________33966, _________33967, _________33968,
       _________33969, _________33970, _________33971, _________33974;
  wire _________33975, _________33976, _________33977, _________33978,
       _________33979, _________33980, _________33981, _________33984;
  wire _________33985, _________33986, _________33987, _________33988,
       _________33989, _________33992, _________33993, _________33994;
  wire _________33995, _________33996, _________33997, _________33998,
       _________34000, _________34001, _________34002, _________34003;
  wire _________34004, _________34005, _________34006, _________34009,
       _________34010, _________34011, _________34012, _________34013;
  wire _________34014, _________34015, _________34016, _________34019,
       _________34020, _________34021, _________34022, _________34023;
  wire _________34024, _________34025, _________34028, _________34029,
       _________34030, _________34031, _________34032, _________34033;
  wire _________34034, _________34056, _________34057, _________34058,
       _________34059, _________34060, _________34061, _________34062;
  wire _________34063, _________34066, _________34067, _________34068,
       _________34069, _________34070, _________34071, _________34072;
  wire _________34073, _________34076, _________34077, _________34078,
       _________34079, _________34080, _________34081, _________34082;
  wire _________34083, _________34086, _________34087, _________34088,
       _________34089, _________34090, _________34091, _________34092;
  wire _________34093, _________34096, _________34097, _________34098,
       _________34099, _________34100, _________34101, _________34102;
  wire _________34105, _________34106, _________34107, _________34108,
       _________34109, _________34110, _________34111, _________34112;
  wire _________34115, _________34116, _________34117, _________34118,
       _________34119, _________34120, _________34121, _________34122;
  wire _________34125, _________34126, _________34127, _________34128,
       _________34129, _________34130, _________34131, _________34132;
  wire _________34155, _________34156, _________34157, _________34158,
       _________34159, _________34160, _________34161, _________34162;
  wire _________34165, _________34166, _________34167, _________34168,
       _________34169, _________34170, _________34171, _________34172;
  wire _________34175, _________34176, _________34177, _________34178,
       _________34179, _________34180, _________34181, _________34184;
  wire _________34185, _________34186, _________34187, _________34188,
       _________34189, _________34190, _________34193, _________34194;
  wire _________34195, _________34196, _________34197, _________34198,
       _________34199, _________34202, _________34203, _________34204;
  wire _________34205, _________34206, _________34207, _________34208,
       _________34211, _________34212, _________34213, _________34214;
  wire _________34215, _________34216, _________34219, _________34220,
       _________34221, _________34222, _________34223, _________34224;
  wire _________34225, _________34226, _________34249, _________34250,
       _________34251, _________34252, _________34253, _________34254;
  wire _________34255, _________34258, _________34259, _________34260,
       _________34261, _________34262, _________34263, _________34266;
  wire _________34267, _________34268, _________34269, _________34270,
       _________34271, _________34272, _________34275, _________34276;
  wire _________34277, _________34278, _________34279, _________34280,
       _________34281, _________34282, _________34285, _________34286;
  wire _________34287, _________34288, _________34289, _________34290,
       _________34291, _________34292, _________34295, _________34296;
  wire _________34297, _________34298, _________34299, _________34300,
       _________34301, _________34302, _________34305, _________34306;
  wire _________34307, _________34308, _________34309, _________34310,
       _________34311, _________34312, _________34315, _________34316;
  wire _________34317, _________34318, _________34319, _________34320,
       _________34321, _________34322, _________34343, _________34344;
  wire _________34345, _________34346, _________34347, _________34348,
       _________34349, _________34350, _________34353, _________34354;
  wire _________34355, _________34356, _________34357, _________34358,
       _________34361, _________34362, _________34363, _________34364;
  wire _________34365, _________34366, _________34367, _________34368,
       _________34371, _________34372, _________34373, _________34374;
  wire _________34375, _________34376, _________34377, _________34378,
       _________34381, _________34382, _________34383, _________34384;
  wire _________34385, _________34386, _________34387, _________34389,
       _________34390, _________34391, _________34392, _________34393;
  wire _________34394, _________34397, _________34398, _________34399,
       _________34400, _________34401, _________34402, _________34403;
  wire _________34404, _________34407, _________34408, _________34409,
       _________34432, _________34433, _________34434, _________34435;
  wire _________34436, _________34437, _________34438, _________34439,
       _________34442, _________34443, _________34444, _________34445;
  wire _________34446, _________34447, _________34448, _________34449,
       _________34452, _________34453, _________34454, _________34455;
  wire _________34456, _________34457, _________34458, _________34459,
       _________34462, _________34463, _________34464, _________34465;
  wire _________34466, _________34467, _________34468, _________34469,
       _________34472, _________34473, _________34474, _________34475;
  wire _________34476, _________34477, _________34478, _________34479,
       _________34482, _________34483, _________34484, _________34485;
  wire _________34486, _________34487, _________34488, _________34489,
       _________34492, _________34493, _________34494, _________34495;
  wire _________34496, _________34497, _________34500, _________34501,
       _________34502, _________34503, _________34504, _________34505;
  wire _________34506, _________34639, _________34640, _________34641,
       _________34642, _________34643, _________34644, _________34645;
  wire _________34646, _________34649, _________34650, _________34651,
       _________34652, _________34653, _________34654, _________34655;
  wire _________34656, _________34659, _________34660, _________34661,
       _________34662, _________34663, _________34664, _________34665;
  wire _________34666, _________34669, _________34670, _________34671,
       _________34672, _________34673, _________34674, _________34675;
  wire _________34676, _________34679, _________34680, _________34681,
       _________34682, _________34683, _________34684, _________34685;
  wire _________34686, _________34689, _________34690, _________34691,
       _________34692, _________34693, _________34694, _________34695;
  wire _________34696, _________34699, _________34700, _________34701,
       _________34702, _________34703, _________34704, _________34705;
  wire _________34706, _________34709, _________34710, _________34711,
       _________34712, _________34713, _________34714, _________34715;
  wire _________34716, _________34739, _________34740, _________34741,
       _________34742, _________34743, _________34744, _________34745;
  wire _________34746, _________34749, _________34750, _________34751,
       _________34752, _________34753, _________34754, _________34755;
  wire _________34756, _________34759, _________34760, _________34761,
       _________34762, _________34763, _________34764, _________34765;
  wire _________34766, _________34769, _________34770, _________34771,
       _________34772, _________34773, _________34774, _________34775;
  wire _________34776, _________34779, _________34780, _________34781,
       _________34782, _________34783, _________34784, _________34785;
  wire _________34786, _________34789, _________34790, _________34791,
       _________34792, _________34793, _________34794, _________34795;
  wire _________34796, _________34799, _________34800, _________34801,
       _________34802, _________34803, _________34804, _________34805;
  wire _________34806, _________34809, _________34810, _________34811,
       _________34812, _________34813, _________34814, _________34815;
  wire _________34816, _________34839, _________34840, _________34841,
       _________34842, _________34843, _________34844, _________34845;
  wire _________34846, _________34849, _________34850, _________34851,
       _________34852, _________34853, _________34854, _________34855;
  wire _________34856, _________34859, _________34860, _________34861,
       _________34862, _________34863, _________34864, _________34865;
  wire _________34866, _________34869, _________34870, _________34871,
       _________34872, _________34873, _________34874, _________34875;
  wire _________34876, _________34879, _________34880, _________34881,
       _________34882, _________34883, _________34884, _________34885;
  wire _________34886, _________34889, _________34890, _________34891,
       _________34892, _________34893, _________34894, _________34895;
  wire _________34896, _________34899, _________34900, _________34901,
       _________34902, _________34903, _________34904, _________34905;
  wire _________34906, _________34909, _________34910, _________34911,
       _________34912, _________34913, _________34914, _________34915;
  wire _________34916, _________34939, _________34940, _________34941,
       _________34942, _________34943, _________34944, _________34945;
  wire _________34946, _________34949, _________34950, _________34951,
       _________34952, _________34953, _________34954, _________34955;
  wire _________34956, _________34959, _________34960, _________34961,
       _________34962, _________34963, _________34964, _________34965;
  wire _________34966, _________34969, _________34970, _________34971,
       _________34972, _________34973, _________34974, _________34975;
  wire _________34976, _________34979, _________34980, _________34981,
       _________34982, _________34983, _________34984, _________34985;
  wire _________34986, _________34989, _________34990, _________34991,
       _________34992, _________34993, _________34994, _________34995;
  wire _________34996, _________34999, _________35000, _________35001,
       _________35002, _________35003, _________35004, _________35005;
  wire _________35006, _________35009, _________35010, _________35011,
       _________35012, _________35013, _________35014, _________35015;
  wire _________35016, _________35039, _________35040, _________35041,
       _________35042, _________35043, _________35044, _________35045;
  wire _________35046, _________35049, _________35050, _________35051,
       _________35052, _________35053, _________35054, _________35055;
  wire _________35056, _________35059, _________35060, _________35061,
       _________35062, _________35063, _________35064, _________35065;
  wire _________35066, _________35069, _________35070, _________35071,
       _________35072, _________35073, _________35074, _________35075;
  wire _________35076, _________35079, _________35080, _________35081,
       _________35082, _________35083, _________35084, _________35085;
  wire _________35086, _________35089, _________35090, _________35091,
       _________35092, _________35093, _________35094, _________35095;
  wire _________35096, _________35099, _________35100, _________35101,
       _________35102, _________35103, _________35104, _________35105;
  wire _________35106, _________35110, _________35111, __________,
       __________0__0_, __________0__9_, __________0___0_,
       __________0___0___18817;
  wire __________0___0___18823, __________0___9_, __________0_____,
       __________0_______18815, __________0_______18816,
       __________0_______18818, __________0_______18819,
       __________0_______18820;
  wire __________0_______18821, __________0_______18822, __________9_,
       ___________, ___________0___18872, ___________0___18877,
       ___________0___18883, ____________;
  wire ____________0_, ____________0___18686, ____________0___18704,
       ____________0___18753, ____________0___18769,
       ____________0___18786, ____________9_, ____________9___18692;
  wire ____________9___18707, ____________9___18758,
       ____________9___18773, ____________9___18791, ____________18893,
       _____________0___18679, _____________0___18684,
       _____________0___18697;
  wire _____________0___18708, _____________0___18715,
       _____________0___18729, _____________0___18740,
       _____________0___18759, _____________0___18764,
       _____________0___18779, _____________0___18784;
  wire _____________0___18798, _____________9___18703,
       _____________9___18714, _____________9___18719,
       _____________9___18751, _____________9___18767,
       _____________9___18778, _____________18894;
  wire _____________18895, _____________18896, _____________18897,
       _____________18898, _____________18899, _____________18900,
       _____________18901, _____________18902;
  wire _____________18905, ______________0___________________,
       ______________0___________________0,
       ______________0___________________9,
       ______________0___________________9__18827,
       ______________0____________________,
       ______________0______________________18824,
       ______________0______________________18825;
  wire ______________0______________________18826,
       ______________0______________________18828, ______________18867,
       ______________18868, ______________18869, ______________18870,
       ______________18871, _______________0__________________;
  wire _______________0__________________0,
       _______________0___________________,
       _______________0____________________18829,
       _______________0_____________________18830,
       _______________0_____________________18831,
       _______________0_____________________18832,
       _______________0_____________________18833,
       _______________0_____________________18834;
  wire _______________18873, _______________18874,
       _______________18875, _______________18876,
       _______________18878, _______________18879,
       _______________18880, _______________18881;
  wire _______________18882, _______________18884,
       ________________18673, ________________18674,
       ________________18675, ________________18676,
       ________________18677, ________________18678;
  wire ________________18687, ________________18688,
       ________________18689, ________________18690,
       ________________18691, ________________18705,
       ________________18706, ________________18721;
  wire ________________18722, ________________18723,
       ________________18724, ________________18735,
       ________________18736, ________________18737,
       ________________18738, ________________18739;
  wire ________________18754, ________________18755,
       ________________18756, ________________18757,
       ________________18770, ________________18771,
       ________________18772, ________________18787;
  wire ________________18788, ________________18789,
       ________________18790, _________________0___18597,
       _________________0___18607, _________________0___18618,
       _________________0___18633, _________________0___18660;
  wire _________________9___18606, _________________9___18616,
       _________________9___18627, _________________9___18642,
       _________________9___18669, _________________18680,
       _________________18681, _________________18682;
  wire _________________18683, _________________18685,
       _________________18693, _________________18694,
       _________________18695, _________________18696,
       _________________18698, _________________18699;
  wire _________________18700, _________________18701,
       _________________18702, _________________18709,
       _________________18710, _________________18711,
       _________________18712, _________________18713;
  wire _________________18716, _________________18717,
       _________________18718, _________________18720,
       _________________18725, _________________18726,
       _________________18727, _________________18728;
  wire _________________18730, _________________18731,
       _________________18732, _________________18733,
       _________________18734, _________________18741,
       _________________18742, _________________18743;
  wire _________________18744, _________________18745,
       _________________18746, _________________18747,
       _________________18748, _________________18749,
       _________________18750, _________________18752;
  wire _________________18760, _________________18761,
       _________________18762, _________________18763,
       _________________18765, _________________18766,
       _________________18768, _________________18774;
  wire _________________18775, _________________18776,
       _________________18777, _________________18780,
       _________________18781, _________________18782,
       _________________18783, _________________18785;
  wire _________________18792, _________________18793,
       _________________18794, _________________18795,
       _________________18796, _________________18797,
       __________________0_, __________________0___18628;
  wire __________________0___18643, __________________0___18670,
       ____________________, _____________________18598,
       _____________________18599, _____________________18600,
       _____________________18601, _____________________18602;
  wire _____________________18603, _____________________18604,
       _____________________18605, _____________________18608,
       _____________________18609, _____________________18610,
       _____________________18611, _____________________18612;
  wire _____________________18613, _____________________18614,
       _____________________18615, _____________________18619,
       _____________________18620, _____________________18621,
       _____________________18622, _____________________18623;
  wire _____________________18624, _____________________18625,
       _____________________18626, _____________________18634,
       _____________________18635, _____________________18636,
       _____________________18637, _____________________18638;
  wire _____________________18639, _____________________18640,
       _____________________18641, _____________________18661,
       _____________________18662, _____________________18663,
       _____________________18664, _____________________18665;
  wire _____________________18666, _____________________18667,
       _____________________18668, ______________________18617,
       ______________________18629, ______________________18630,
       ______________________18631, ______________________18632;
  wire ______________________18644, ______________________18671,
       ______________________18672, __________________________________,
       __________________________________0,
       __________________________________9,
       ___________________________________,
       ____________________________________18835;
  wire ____________________________________18836,
       _____________________________________18837,
       _____________________________________18838,
       _____________________________________18839,
       ______________________________________0__________0,
       ______________________________________0__________0__18892,
       ______________________________________0___________,
       ______________________________________0_____________18885;
  wire ______________________________________0_____________18886,
       ______________________________________0_____________18887,
       ______________________________________0_____________18888,
       ______________________________________0_____________18889,
       ______________________________________0_____________18890,
       ______________________________________0_____________18891;
  dffacs1 ________________(.CLRB (reset), .CLK (clk), .DIN
       (_________34408), .QN (_____________18905));
  nnd2s1 ____________0(.DIN1 (_________34407), .DIN2 (______9__30590),
       .Q (_________34408));
  nnd2s1 ___________9_(.DIN1 (___9____19692), .DIN2 (______9__34410),
       .Q (_________34407));
  dffacs1 ______________0_____(.CLRB (reset), .CLK (clk), .DIN
       (______0__34406), .QN (______9__34410));
  nnd2s1 ______0______(.DIN1 (______9__34405), .DIN2 (_________34393),
       .Q (______0__34406));
  xor2s1 _____________(.DIN1 (_________34383), .DIN2 (_________34404),
       .Q (______9__34405));
  xor2s1 _____________436009(.DIN1 (_________34402), .DIN2
       (_________33541), .Q (_________34404));
  dffacs1 ______________9_(.CLRB (reset), .CLK (clk), .DIN
       (_________34403), .QN (_________9___18903));
  or2s1 _________9___(.DIN1 (________20000), .DIN2 (_________34401), .Q
       (_________34403));
  xor2s1 _____________436010(.DIN1 (_________34399), .DIN2
       (_________33925), .Q (_________34402));
  dffacs1 ______________0___0_(.CLRB (reset), .CLK (clk), .DIN
       (_________34400), .Q (__________0___0___18823));
  nor2s1 ______9____09(.DIN1 (_____90__34411), .DIN2 (________19962),
       .Q (_________34401));
  nor2s1 _____________436011(.DIN1 (_________________0___18660), .DIN2
       (_________34397), .Q (_________34400));
  dffacs1 ________________436012(.CLRB (reset), .CLK (clk), .DIN
       (_________34398), .QN (_____________18902));
  nnd2s1 __________900(.DIN1 (______0__34396), .DIN2 (______9__34379),
       .Q (_________34399));
  dffacs1 ______________0___9_(.CLRB (reset), .CLK (clk), .DIN
       (_________34394), .Q (_____90__34411));
  nnd2s1 ___________9_436013(.DIN1 (_________34392), .DIN2
       (________19366), .Q (_________34398));
  xor2s1 _____________436014(.DIN1 (______0__34380), .DIN2
       (______9__34395), .Q (_________34397));
  or2s1 _____________436015(.DIN1 (_________34374), .DIN2
       (______9__34395), .Q (______0__34396));
  nnd2s1 _____________436016(.DIN1 (_________34391), .DIN2
       (_________34393), .Q (_________34394));
  nnd2s1 _____________436017(.DIN1 (___9____19692), .DIN2
       (__________0_______18822), .Q (_________34392));
  nor2s1 ______0___9__(.DIN1 (_________34353), .DIN2 (_________34390),
       .Q (______9__34395));
  dffacs1 ______________0_____436018(.CLRB (reset), .CLK (clk), .DIN
       (______0__34388), .Q (__________0_______18822));
  xor2s1 ______9____0_(.DIN1 (_________34361), .DIN2 (____0____34558),
       .Q (_________34391));
  dffacs1 ________________436019(.CLRB (reset), .CLK (clk), .DIN
       (_________34389), .QN (outData[27]));
  and2s1 _____________436020(.DIN1 (____0____34558), .DIN2
       (______9__34351), .Q (_________34390));
  nnd2s1 _____________436021(.DIN1 (_________34387), .DIN2
       (___9____21587), .Q (_________34389));
  nor2s1 ____________436022(.DIN1 (_________________0___18660), .DIN2
       (_________34386), .Q (______0__34388));
  nnd2s1 ___________0_(.DIN1 (___9____19692), .DIN2 (______0__34499),
       .Q (_________34387));
  xor2s1 ___________9_436023(.DIN1 (_________34385), .DIN2
       (_________34371), .Q (_________34386));
  dffacs1 ________________436024(.CLRB (reset), .CLK (clk), .DIN
       (_________34384), .QN (_____________18901));
  dffacs1 ______________0_____436025(.CLRB (reset), .CLK (clk), .DIN
       (_________34382), .Q (______0__34499));
  nnd2s1 ______0_____0(.DIN1 (_________34381), .DIN2 (________20100),
       .Q (_________34384));
  xor2s1 __________0_9(.DIN1 (_________34376), .DIN2 (_________34307),
       .Q (_________34383));
  xor2s1 _____________436026(.DIN1 (_________34377), .DIN2
       (_________34362), .Q (_________34385));
  nnd2s1 _________990_(.DIN1 (_________34378), .DIN2 (_________34365),
       .Q (_________34382));
  nnd2s1 ____________436027(.DIN1 (___9____19692), .DIN2
       (_____9___34412), .Q (_________34381));
  nnd2s1 ___________9_436028(.DIN1 (______9__34379), .DIN2
       (_________34375), .Q (______0__34380));
  xor2s1 _____________436029(.DIN1 (_________34363), .DIN2
       (_________34372), .Q (_________34378));
  nor2s1 _____________436030(.DIN1 (_________34347), .DIN2
       (_________34373), .Q (_________34377));
  xor2s1 _____________436031(.DIN1 (_________34367), .DIN2
       (_________34069), .Q (_________34376));
  dffacs1 ______________0_____436032(.CLRB (reset), .CLK (clk), .DIN
       (_________34366), .QN (_____9___34412));
  hi1s1 _____90(.DIN (_________34374), .Q (_________34375));
  dffacs1 ________________436033(.CLRB (reset), .CLK (clk), .DIN
       (_________34364), .QN (_____________18900));
  nor2s1 _________9___436034(.DIN1 (_________34348), .DIN2
       (_________34372), .Q (_________34373));
  nnd2s1 _____________436035(.DIN1 (______0__34370), .DIN2
       (_________34354), .Q (_________34371));
  nor2s1 _____9_____09(.DIN1 (_________34368), .DIN2 (______9__34369),
       .Q (_________34374));
  nnd2s1 _____9_______(.DIN1 (______9__34369), .DIN2 (_________34368),
       .Q (______9__34379));
  nnd2s1 _____00___900(.DIN1 (______0__34360), .DIN2 (_________34280),
       .Q (_________34367));
  nnd2s1 ______9____9_(.DIN1 (_________34357), .DIN2 (_________34365),
       .Q (_________34366));
  or2s1 ______0______436036(.DIN1 (_____9__21155), .DIN2
       (_________34358), .Q (_________34364));
  xor2s1 _____________436037(.DIN1 (_________34349), .DIN2
       (_________28828), .Q (_________34363));
  xor2s1 _____0_______(.DIN1 (______0__34294), .DIN2 (______9__34359),
       .Q (_________34368));
  nor2s1 ______9______(.DIN1 (_____9___34325), .DIN2 (_________34356),
       .Q (_________34372));
  xor2s1 _____9____9__(.DIN1 (_________34346), .DIN2 (_________34362),
       .Q (______0__34370));
  xor2s1 _____0_____0_(.DIN1 (______0__34352), .DIN2 (_________32215),
       .Q (_________34361));
  or2s1 _____________436038(.DIN1 (_________34279), .DIN2
       (______9__34359), .Q (______0__34360));
  nor2s1 _____________436039(.DIN1 (__________0_______18821), .DIN2
       (________19962), .Q (_________34358));
  xor2s1 _____9______0(.DIN1 (_____9___34327), .DIN2 (_________34355),
       .Q (_________34357));
  dffacs1 ________________436040(.CLRB (reset), .CLK (clk), .DIN
       (_________34343), .QN (_____________18899));
  nor2s1 _____99___0__(.DIN1 (_____9___34326), .DIN2 (_________34355),
       .Q (_________34356));
  and2s1 _____09____0_(.DIN1 (_________34350), .DIN2 (______0__34352),
       .Q (_________34353));
  or2s1 ______0____9_(.DIN1 (______0__34352), .DIN2 (_________34350),
       .Q (______9__34351));
  nor2s1 _____9_______436041(.DIN1 (_________34348), .DIN2
       (_________34347), .Q (_________34349));
  nor2s1 _____0______0(.DIN1 (_________34344), .DIN2 (_________34345),
       .Q (_________34346));
  nnd2s1 __________0_436042(.DIN1 (_________34345), .DIN2
       (_________34344), .Q (_________34354));
  nnd2s1 _____________436043(.DIN1 (_____0___34339), .DIN2
       (________20103), .Q (_________34343));
  dffacs1 ______________0_____436044(.CLRB (reset), .CLK (clk), .DIN
       (______0__34342), .QN (__________0_______18821));
  nor2s1 _________990_436045(.DIN1 (_____0___34242), .DIN2
       (_____09__34341), .Q (______9__34359));
  nor2s1 _____0______436046(.DIN1 (_________34320), .DIN2
       (_____0___34337), .Q (_________34355));
  xor2s1 ___________9_436047(.DIN1 (_____0___34335), .DIN2
       (_________________0___18618), .Q (_________34347));
  xor2s1 ______0______436048(.DIN1 (_________34252), .DIN2
       (_____0___34340), .Q (______0__34352));
  dffacs1 ________________436049(.CLRB (reset), .CLK (clk), .DIN
       (_____0___34338), .QN (outData[23]));
  nor2s1 _____0_______436050(.DIN1 (_________________0___18660), .DIN2
       (_____0___34336), .Q (______0__34342));
  xor2s1 ______9______436051(.DIN1 (_____9___34331), .DIN2
       (_________9_______18813), .Q (_________34344));
  nor2s1 _________9___436052(.DIN1 (_____0___34246), .DIN2
       (_____0___34340), .Q (_____09__34341));
  nnd2s1 _____9_______436053(.DIN1 (___9____19692), .DIN2
       (__________0_______18820), .Q (_____0___34339));
  nnd2s1 _____0_____09(.DIN1 (_____99__34332), .DIN2 (_________34295),
       .Q (_____0___34338));
  xor2s1 _____________436054(.DIN1 (_____9___34329), .DIN2
       (____0____32777), .Q (_____0___34337));
  dffacs1 ______________0_____436055(.CLRB (reset), .CLK (clk), .DIN
       (_____9___34330), .Q (__________0_______18820));
  xor2s1 __________436056(.DIN1 (_________34321), .DIN2
       (_____9___34328), .Q (_____0___34336));
  nnd2s1 ___________9_436057(.DIN1 (_____00__34333), .DIN2
       (_____0___34334), .Q (_____0___34335));
  nor2s1 _____________436058(.DIN1 (______9__34217), .DIN2
       (_____90__34324), .Q (_____0___34340));
  nor2s1 _____________436059(.DIN1 (_____0___34334), .DIN2
       (_____00__34333), .Q (_________34348));
  nor2s1 _____________436060(.DIN1 (_________34322), .DIN2
       (_____9__20273), .Q (_____99__34332));
  xor2s1 _____________436061(.DIN1 (______9__34323), .DIN2
       (_____________________________________18839), .Q
       (_____9___34331));
  nor2s1 __________9__(.DIN1 (_________________0___18660), .DIN2
       (_________34319), .Q (_____9___34330));
  xor2s1 ______9____0_436062(.DIN1 (_________34316), .DIN2
       (_____________________________________18839), .Q
       (_____0___34334));
  nnd2s1 ______0______436063(.DIN1 (_________34318), .DIN2
       (_____9___34328), .Q (_____9___34329));
  or2s1 _____________436064(.DIN1 (_____9___34326), .DIN2
       (_____9___34325), .Q (_____9___34327));
  nor2s1 ____________436065(.DIN1 (_________34214), .DIN2
       (______9__34323), .Q (_____90__34324));
  nor2s1 __________0__(.DIN1 (__________0_______18819), .DIN2
       (________19962), .Q (_________34322));
  or2s1 ___________0_436066(.DIN1 (_________34320), .DIN2
       (_________34317), .Q (_________34321));
  xor2s1 ___________9_436067(.DIN1 (_________34312), .DIN2
       (_________34272), .Q (_________34319));
  hi1s1 _______(.DIN (_________34317), .Q (_________34318));
  xor2s1 _____________436068(.DIN1 (_________34311), .DIN2
       (_____9___33022), .Q (_____9___34325));
  nor2s1 ______9_____0(.DIN1 (_______18956), .DIN2 (_________34315), .Q
       (______9__34323));
  dffacs1 ______________0_____436069(.CLRB (reset), .CLK (clk), .DIN
       (______9__34313), .Q (__________0_______18819));
  xor2s1 __________0_436070(.DIN1 (_________9_______18812), .DIN2
       (______0__34314), .Q (_________34316));
  xor2s1 _____________436071(.DIN1 (_________34308), .DIN2
       (_____9___33026), .Q (_________34317));
  nor2s1 _________990_436072(.DIN1 (______18948), .DIN2
       (______0__34314), .Q (_________34315));
  nor2s1 ____________436073(.DIN1 (_________________0___18660), .DIN2
       (_________34306), .Q (______9__34313));
  xor2s1 ___________9_436074(.DIN1 (_________34305), .DIN2
       (____00___31810), .Q (_________34312));
  nnd2s1 _____________436075(.DIN1 (_________34309), .DIN2
       (_________34310), .Q (_________34311));
  nor2s1 _____________436076(.DIN1 (_________34310), .DIN2
       (_________34309), .Q (_____9___34326));
  nor2s1 _____________436077(.DIN1 (______0__34304), .DIN2
       (_________34299), .Q (_________34308));
  xor2s1 _________9___436078(.DIN1 (_____99__34420), .DIN2
       (_________9_______18814), .Q (_________34307));
  nor2s1 ______9______436079(.DIN1 (________19446), .DIN2
       (______9__34303), .Q (______0__34314));
  xor2s1 ______0____09(.DIN1 (_________34275), .DIN2 (_________34297),
       .Q (_________34306));
  nnd2s1 _____________436080(.DIN1 (_________34301), .DIN2
       (_________34271), .Q (_____9___34328));
  xor2s1 __________436081(.DIN1 (_________34302), .DIN2
       (___99___19767), .Q (_________34310));
  xor2s1 ___________9_436082(.DIN1 (_________34300), .DIN2
       (_____00__30545), .Q (_________34305));
  dffacs1 ________________436083(.CLRB (reset), .CLK (clk), .DIN
       (_________34296), .QN (outData[22]));
  xor2s1 _____________436084(.DIN1 (_________34298), .DIN2
       (_________31578), .Q (______0__34304));
  nor2s1 _____________436085(.DIN1 (________19447), .DIN2
       (_________34302), .Q (______9__34303));
  or2s1 _____________436086(.DIN1 (_________34266), .DIN2
       (_________34300), .Q (_________34301));
  dffacs1 _____________9_____(.CLRB (reset), .CLK (clk), .DIN
       (______9__34293), .Q (_________9_______18814));
  and2s1 _____________436087(.DIN1 (_________34299), .DIN2
       (_________34298), .Q (_________34320));
  xor2s1 __________9__436088(.DIN1 (_________34289), .DIN2
       (____9_9__33643), .Q (_________34297));
  nnd2s1 ___________0_436089(.DIN1 (_________34292), .DIN2
       (_________34295), .Q (_________34296));
  xor2s1 _____________436090(.DIN1 (_________34290), .DIN2
       (______9__32232), .Q (_________34302));
  xor2s1 _____________436091(.DIN1 (______0__34284), .DIN2
       (__________________________________), .Q (______0__34294));
  nnd2s1 ____________436092(.DIN1 (_________34287), .DIN2
       (_________34288), .Q (_________34300));
  nor2s1 __________0__436093(.DIN1 (_________________0___18660), .DIN2
       (_________34291), .Q (______9__34293));
  xor2s1 ___________0_436094(.DIN1 (______9__34283), .DIN2
       (_________31290), .Q (_________34298));
  nor2s1 ______9____9_436095(.DIN1 (_________34285), .DIN2
       (___99___21627), .Q (_________34292));
  nor2s1 ______0______436096(.DIN1 (_________34277), .DIN2
       (_________34278), .Q (_________34291));
  nor2s1 ____________436097(.DIN1 (___9____24289), .DIN2
       (_________34282), .Q (_________34290));
  and2s1 __________0_436098(.DIN1 (_________34286), .DIN2
       (_________34288), .Q (_________34289));
  nnd2s1 _____________436099(.DIN1 (______0__34274), .DIN2
       (_________34286), .Q (_________34287));
  nor2s1 _________990_436100(.DIN1 (__________0_______18818), .DIN2
       (________19962), .Q (_________34285));
  xor2s1 ____________436101(.DIN1 (_____99__34420), .DIN2
       (_____0___33866), .Q (______0__34284));
  xnr2s1 ___________9_436102(.DIN1 (_________9_______18811), .DIN2
       (_________34281), .Q (______9__34283));
  nor2s1 _____________436103(.DIN1 (___9____24274), .DIN2
       (_________34281), .Q (_________34282));
  nnd2s1 _____________436104(.DIN1 (______9__31228), .DIN2
       (_________34276), .Q (_________34286));
  nnd2s1 ______9______436105(.DIN1 (_____99__34420), .DIN2
       (__________________________________), .Q (_________34280));
  nor2s1 ______0__9___(.DIN1 (__________________________________),
       .DIN2 (_____99__34420), .Q (_________34279));
  nnd2s1 _____________436106(.DIN1 (______9__34273), .DIN2
       (_________34251), .Q (_________34278));
  dffacs1 ______________0_____436107(.CLRB (reset), .CLK (clk), .DIN
       (_________34270), .Q (__________0_______18818));
  nor2s1 ___________09(.DIN1 (_________34269), .DIN2 (_________34216),
       .Q (_________34277));
  xor2s1 _____________436108(.DIN1 (_________34268), .DIN2
       (____0_0__30932), .Q (_________34276));
  xor2s1 __________436109(.DIN1 (______0__34274), .DIN2
       (_________31153), .Q (_________34275));
  nnd2s1 ___________9_436110(.DIN1 (_________34263), .DIN2
       (_________34260), .Q (_________34281));
  nnd2s1 _____________436111(.DIN1 (______9__34264), .DIN2
       (_______________18884), .Q (______9__34273));
  nnd2s1 _____90______(.DIN1 (______0__34265), .DIN2 (_________34271),
       .Q (_________34272));
  dffacs1 _____________9___0_(.CLRB (reset), .CLK (clk), .DIN
       (_________34267), .QN (_____99__34420));
  nor2s1 _____________436112(.DIN1 (_________________0___18660), .DIN2
       (_________34262), .Q (_________34270));
  nor2s1 _____________436113(.DIN1 (_________34255), .DIN2
       (_________34261), .Q (_________34269));
  nnd2s1 __________9__436114(.DIN1 (_________31226), .DIN2
       (_________34268), .Q (_________34288));
  nnd2s1 _____9_____0_(.DIN1 (______0__34257), .DIN2 (_________34365),
       .Q (_________34267));
  hi1s1 _____9_(.DIN (______0__34265), .Q (_________34266));
  nnd2s1 _____9_______436115(.DIN1 (____0_0__34560), .DIN2
       (______9__34256), .Q (______9__34264));
  nnd2s1 _____99______(.DIN1 (_________34259), .DIN2 (_____0___31184),
       .Q (_________34263));
  nnd2s1 _____00_____0(.DIN1 (_____9___31347), .DIN2 (_________34258),
       .Q (_________34271));
  xor2s1 ______9___0__(.DIN1 (_________34250), .DIN2 (_____0___33866),
       .Q (_________34262));
  nnd2s1 ___________0_436116(.DIN1 (_____0___34240), .DIN2
       (_________34253), .Q (______0__34274));
  nor2s1 _____9_____9_(.DIN1 (_________34254), .DIN2
       (_______________18884), .Q (_________34261));
  xor2s1 _____9_______436117(.DIN1 (_________34249), .DIN2
       (_________31431), .Q (_________34268));
  nnd2s1 _____0______436118(.DIN1 (_____90__31344), .DIN2
       (____0____34555), .Q (______0__34265));
  nnd2s1 _____0____0_9(.DIN1 (_____0___34245), .DIN2 (______9__34123),
       .Q (_________34260));
  nnd2s1 _____0_______436119(.DIN1 (_____0___34243), .DIN2
       (____0___19213), .Q (_________34259));
  hi1s1 _____09(.DIN (____0____34555), .Q (_________34258));
  xor2s1 ______0__990_(.DIN1 (_____00__34238), .DIN2 (______0__35078),
       .Q (______0__34257));
  nnd2s1 ____________436120(.DIN1 (_____09__34247), .DIN2
       (_____________0___18798), .Q (______9__34256));
  dffacs1 ______________0_(.CLRB (reset), .CLK (clk), .DIN
       (______0__34248), .QN (_________0_));
  nor2s1 _____0_____9_(.DIN1 (_____________0___18798), .DIN2
       (_____00__34421), .Q (_________34255));
  nnd2s1 _____0_______436121(.DIN1 (_____00__34421), .DIN2
       (_____________0___18798), .Q (_________34254));
  nnd2s1 _____9_______436122(.DIN1 (_____0___34239), .DIN2
       (____9____29986), .Q (_________34253));
  xor2s1 _________9___436123(.DIN1 (_________34221), .DIN2
       (__________________________________), .Q (_________34252));
  or2s1 _____________436124(.DIN1 (_____00__34421), .DIN2
       (_________34225), .Q (_________34251));
  dffacs1 ________________436125(.CLRB (reset), .CLK (clk), .DIN
       (_____0___34241), .QN (_____________18898));
  xor2s1 _____________436126(.DIN1 (_____9___34231), .DIN2
       (_____9___34235), .Q (_________34250));
  xor2s1 __________436127(.DIN1 (_____9___34230), .DIN2
       (_________33895), .Q (_________34249));
  nnd2s1 _____9_____9_436128(.DIN1 (_____99__34237), .DIN2
       (_____0__20264), .Q (______0__34248));
  hi1s1 _______436129(.DIN (_____00__34421), .Q (_____09__34247));
  and2s1 _____________436130(.DIN1 (_________9_______18813), .DIN2
       (__________________________________), .Q (_____0___34246));
  nor2s1 ______0______436131(.DIN1 (____9___19495), .DIN2
       (_____0___34244), .Q (_____0___34245));
  nnd2s1 ______9______436132(.DIN1 (_____0___34244), .DIN2
       (____09__19214), .Q (_____0___34243));
  nor2s1 _____________436133(.DIN1
       (__________________________________), .DIN2
       (_________9_______18813), .Q (_____0___34242));
  or2s1 _____0____9__(.DIN1 (________20900), .DIN2 (_____9___34233), .Q
       (_____0___34241));
  nnd2s1 _____0_____0_436134(.DIN1 (_____9___34234), .DIN2
       (___0_09__27568), .Q (_____0___34240));
  nnd2s1 _____________436135(.DIN1 (_____9___34236), .DIN2
       (_________34219), .Q (_____0___34239));
  xor2s1 _____________436136(.DIN1 (_________34226), .DIN2
       (_____________0___18798), .Q (_____00__34238));
  dffacs1 ___________________(.CLRB (reset), .CLK (clk), .DIN
       (_____9___34232), .Q (_____00__34421));
  nnd2s1 _____0______436137(.DIN1 (___9____19692), .DIN2
       (__________0___0___18817), .Q (_____99__34237));
  nor2s1 __________0__436138(.DIN1 (________22296), .DIN2
       (_____9___34229), .Q (_____0___34244));
  dffacs1 _____________9___9_(.CLRB (reset), .CLK (clk), .DIN
       (______9__34227), .Q (__________________________________));
  nnd2s1 ___________0_436139(.DIN1 (_____9___34235), .DIN2
       (_________34208), .Q (_____9___34236));
  nor2s1 ___________9_436140(.DIN1 (_____9___34235), .DIN2
       (_________34223), .Q (_____9___34234));
  nor2s1 _____________436141(.DIN1 (_____9___34413), .DIN2
       (________19962), .Q (_____9___34233));
  nnd2s1 ____________436142(.DIN1 (_________34222), .DIN2
       (_________34393), .Q (_____9___34232));
  nor2s1 ______0___0_9(.DIN1 (_________34220), .DIN2 (_________34224),
       .Q (_____9___34231));
  xnr2s1 _____________436143(.DIN1 (_____90__34228), .DIN2
       (________22297), .Q (_____9___34230));
  dffacs1 ______________0___0_436144(.CLRB (reset), .CLK (clk), .DIN
       (______0__34218), .Q (__________0___0___18817));
  and2s1 _________990_436145(.DIN1 (_____90__34228), .DIN2
       (________19248), .Q (_____9___34229));
  nnd2s1 ____________436146(.DIN1 (_________34213), .DIN2
       (_________34393), .Q (______9__34227));
  and2s1 ___________9_436147(.DIN1 (_________34215), .DIN2
       (_________34225), .Q (_________34226));
  dffacs1 ______________0_____436148(.CLRB (reset), .CLK (clk), .DIN
       (_________34212), .Q (_____9___34413));
  xor2s1 _____________436149(.DIN1 (______0__34210), .DIN2
       (_________31479), .Q (_____9___34235));
  nor2s1 _____________436150(.DIN1 (_________33268), .DIN2
       (_________34223), .Q (_________34224));
  xor2s1 _____________436151(.DIN1 (_________34206), .DIN2
       (_____9___34137), .Q (_________34222));
  xor2s1 ______0__9___436152(.DIN1 (_________9_______18813), .DIN2
       (_________34077), .Q (_________34221));
  nor2s1 _____________436153(.DIN1 (______9__33247), .DIN2
       (_________34219), .Q (_________34220));
  nor2s1 ___________436154(.DIN1 (_________34187), .DIN2
       (______9__34209), .Q (______0__34218));
  and2s1 _____________436155(.DIN1 (_________9_______18813), .DIN2
       (_____________________________________18839), .Q
       (______9__34217));
  nor2s1 __________436156(.DIN1 (_________34199), .DIN2
       (_________34211), .Q (_____90__34228));
  or2s1 _____________436157(.DIN1 (_________31290), .DIN2
       (_________34216), .Q (_________34215));
  nor2s1 _____________436158(.DIN1 (_________9_______18813), .DIN2
       (_____________________________________18839), .Q
       (_________34214));
  xor2s1 _____________436159(.DIN1 (_________34203), .DIN2
       (____9____31787), .Q (_________34213));
  nnd2s1 ______0______436160(.DIN1 (_________34204), .DIN2
       (_________34393), .Q (_________34212));
  xor2s1 __________9__436161(.DIN1 (_________31161), .DIN2
       (_________34207), .Q (_________34223));
  nor2s1 ___________0_436162(.DIN1 (_________29736), .DIN2
       (______9__34200), .Q (_________34211));
  nnd2s1 ______9______436163(.DIN1 (_________34202), .DIN2
       (_________34176), .Q (______0__34210));
  xor2s1 _____________436164(.DIN1 (_________34195), .DIN2
       (_________34181), .Q (______9__34209));
  or2s1 ____________436165(.DIN1 (_________34207), .DIN2
       (_________34205), .Q (_________34208));
  xor2s1 ______9___0__436166(.DIN1 (_________34194), .DIN2
       (_____90__32282), .Q (_________34206));
  nnd2s1 ___________0_436167(.DIN1 (_________34205), .DIN2
       (_________34207), .Q (_________34219));
  nnd2s1 ___________9_436168(.DIN1 (_________34225), .DIN2
       (____99___34522), .Q (_________34216));
  dffacs1 _____________9_____436169(.CLRB (reset), .CLK (clk), .DIN
       (_________34198), .Q (_________9_______18813));
  xor2s1 _____________436170(.DIN1 (_________34177), .DIN2
       (______0__34201), .Q (_________34204));
  and2s1 ____________436171(.DIN1 (_________34197), .DIN2
       (____99___34522), .Q (_________34203));
  or2s1 __________0_436172(.DIN1 (_________34169), .DIN2
       (______0__34201), .Q (_________34202));
  nor2s1 _____________436173(.DIN1 (________19451), .DIN2
       (______0__34192), .Q (______9__34200));
  nor2s1 _________990_436174(.DIN1 (____0____32807), .DIN2
       (_________34196), .Q (_________34199));
  nnd2s1 ____________436175(.DIN1 (_________34190), .DIN2
       (___0____24415), .Q (_________34198));
  nnd2s1 ______9____9_436176(.DIN1 (_________34197), .DIN2
       (_________31290), .Q (_________34225));
  nnd2s1 _____________436177(.DIN1 (_________34196), .DIN2
       (_________34193), .Q (_________34207));
  xor2s1 ______0______436178(.DIN1 (_________34184), .DIN2
       (______9__33828), .Q (_________34195));
  dffacs1 ______________9_436179(.CLRB (reset), .CLK (clk), .DIN
       (_________34186), .QN (_________9_));
  xor2s1 _____________436180(.DIN1 (_________34179), .DIN2
       (______9__33856), .Q (_________34194));
  dffacs1 _________________0_(.CLRB (reset), .CLK (clk), .DIN
       (_________34188), .Q (_____________0___18798));
  or2s1 ______9______436181(.DIN1 (_________34189), .DIN2
       (______9__34191), .Q (_________34193));
  nor2s1 ______0____436182(.DIN1 (________19450), .DIN2
       (______9__34191), .Q (______0__34192));
  nor2s1 _____________436183(.DIN1 (______0__34183), .DIN2
       (______9__34182), .Q (______0__34201));
  nnd2s1 __________436184(.DIN1 (_________34178), .DIN2
       (_________34159), .Q (_________34190));
  nnd2s1 ___________9_436185(.DIN1 (______9__34191), .DIN2
       (_________34189), .Q (_________34196));
  nnd2s1 _____________436186(.DIN1 (_________34185), .DIN2
       (_____0___34422), .Q (_________34197));
  nor2s1 ______0______436187(.DIN1 (_________34187), .DIN2
       (______9__34173), .Q (_________34188));
  dffacs1 _____________9_____436188(.CLRB (reset), .CLK (clk), .DIN
       (_________34175), .Q
       (_____________________________________18839));
  nnd2s1 _____________436189(.DIN1 (______0__34174), .DIN2
       (___99___20697), .Q (_________34186));
  nor2s1 _____________436190(.DIN1 (______0__34183), .DIN2
       (_________34180), .Q (_________34184));
  nor2s1 __________9__436191(.DIN1 (_________34181), .DIN2
       (_________34180), .Q (______9__34182));
  nor2s1 ___________0_436192(.DIN1 (_________34156), .DIN2
       (_________34171), .Q (______9__34191));
  dffacs1 _____________9_____436193(.CLRB (reset), .CLK (clk), .DIN
       (_________34172), .Q (_________9_______18812));
  nor2s1 ____90_______(.DIN1 (_________34096), .DIN2 (_________34166),
       .Q (_________34179));
  xor2s1 _____9_______436194(.DIN1 (______0__34164), .DIN2
       (_________34167), .Q (_________34178));
  nnd2s1 ____________436195(.DIN1 (_________34176), .DIN2
       (_________34170), .Q (_________34177));
  nor2s1 ____90____0__(.DIN1 (______9__34163), .DIN2 (_________34168),
       .Q (_________34185));
  nnd2s1 _____90____0_(.DIN1 (_________34160), .DIN2 (________22248),
       .Q (_________34175));
  nnd2s1 _____9_____9_436196(.DIN1 (___9____19692), .DIN2
       (__________0___9_), .Q (______0__34174));
  xor2s1 _____9_______436197(.DIN1 (_________34098), .DIN2
       (_________34165), .Q (______9__34173));
  dffacs1 _________________9_(.CLRB (reset), .CLK (clk), .DIN
       (_________34161), .QN (_____0___34422));
  nnd2s1 _____9______436198(.DIN1 (_________34155), .DIN2
       (_____0__22865), .Q (_________34172));
  nor2s1 _____9____0_9(.DIN1 (_________30595), .DIN2 (_________34157),
       .Q (_________34171));
  xor2s1 ______9______436199(.DIN1 (_____0___34149), .DIN2
       (____0_0__31861), .Q (_________34180));
  hi1s1 _____9_436200(.DIN (_________34169), .Q (_________34170));
  nor2s1 ____9____990_(.DIN1 (_________34162), .DIN2 (_________34167),
       .Q (_________34168));
  nor2s1 ____9_______0(.DIN1 (_________34097), .DIN2 (_________34165),
       .Q (_________34166));
  nor2s1 ____9_9____9_(.DIN1 (______9__34163), .DIN2 (_________34162),
       .Q (______0__34164));
  nnd2s1 ____9________(.DIN1 (_____0___34150), .DIN2 (_________34393),
       .Q (_________34161));
  dffacs1 _____________9_____436201(.CLRB (reset), .CLK (clk), .DIN
       (_____0___34152), .Q (_________9_______18809));
  dffacs1 ________________436202(.CLRB (reset), .CLK (clk), .DIN
       (______0__34154), .QN (_____________18897));
  dffacs1 ______________0___9_436203(.CLRB (reset), .CLK (clk), .DIN
       (_____09__34153), .Q (__________0___9_));
  nnd2s1 ____9________436204(.DIN1 (_____0___34151), .DIN2
       (_________34159), .Q (_________34160));
  nor2s1 _____99______436205(.DIN1 (_________34158), .DIN2
       (____0____30985), .Q (_________34169));
  nnd2s1 ____900__9___(.DIN1 (____0____30986), .DIN2 (_________34158),
       .Q (_________34176));
  nor2s1 ____9________436206(.DIN1 (_________32149), .DIN2
       (_____9___34139), .Q (_________34167));
  nor2s1 ____9_0____09(.DIN1 (_________34131), .DIN2 (_____9___34140),
       .Q (_________34165));
  dffacs1 ________________436207(.CLRB (reset), .CLK (clk), .DIN
       (_____00__34144), .QN (outData[17]));
  nor2s1 ____90_______436208(.DIN1 (_________33992), .DIN2
       (_____0___34146), .Q (_________34157));
  nor2s1 ____90____900(.DIN1 (_________32081), .DIN2 (_____99__34143),
       .Q (_________34156));
  nnd2s1 ____9______9_(.DIN1 (_____9___34141), .DIN2 (_________34159),
       .Q (_________34155));
  nnd2s1 ____9_0______(.DIN1 (_____9___34135), .DIN2 (________21272),
       .Q (______0__34154));
  nor2s1 ____9________436209(.DIN1 (_________________0___18660), .DIN2
       (_____90__34134), .Q (_____09__34153));
  nor2s1 ____9________436210(.DIN1 (_____0___34147), .DIN2
       (_____0___34148), .Q (______0__34183));
  xor2s1 ____9________436211(.DIN1 (_____0___34145), .DIN2
       (_____9___34142), .Q (_________34158));
  nnd2s1 ____90____9__(.DIN1 (______0__33991), .DIN2 (_____9___34136),
       .Q (_____0___34152));
  xor2s1 ____9______0_(.DIN1 (_________32151), .DIN2 (_____9___34138),
       .Q (_____0___34151));
  nor2s1 ____9________436212(.DIN1 (_________34122), .DIN2
       (_________34132), .Q (_____0___34150));
  nnd2s1 ____9________436213(.DIN1 (_____0___34148), .DIN2
       (_____0___34147), .Q (_____0___34149));
  nor2s1 ____9_0_____0(.DIN1 (______9__34133), .DIN2 (_____0___35109),
       .Q (_________34162));
  nor2s1 ____9_____0__(.DIN1 (_________33993), .DIN2 (_____0___34145),
       .Q (_____0___34146));
  nnd2s1 ____9______0_436214(.DIN1 (_________34129), .DIN2
       (______9__34084), .Q (_____00__34144));
  nnd2s1 ____9_9____9_436215(.DIN1 (_____0___34145), .DIN2
       (_____9___34142), .Q (_____99__34143));
  xor2s1 ____9________436216(.DIN1 (_________34125), .DIN2
       (_________________18796), .Q (_____9___34141));
  xor2s1 ____9_9_____0(.DIN1 (_________34130), .DIN2 (_________32554),
       .Q (_____9___34140));
  nor2s1 ____9_____0_9(.DIN1 (_________32150), .DIN2 (_____9___34138),
       .Q (_____9___34139));
  xor2s1 ____9________436217(.DIN1 (______0__34124), .DIN2
       (_________________18785), .Q (_____9___34137));
  nnd2s1 ____9____990_436218(.DIN1 (_________34128), .DIN2
       (_________34110), .Q (_________34181));
  nor2s1 ____9_______436219(.DIN1 (_____0___34423), .DIN2
       (_______________18884), .Q (______9__34163));
  nnd2s1 ____9______9_436220(.DIN1 (_________34126), .DIN2
       (inData[14]), .Q (_____9___34136));
  nnd2s1 ____9________436221(.DIN1 (_________34116), .DIN2
       (_____9___34414), .Q (_____9___34135));
  xor2s1 ____9________436222(.DIN1 (_________34120), .DIN2
       (______0__34114), .Q (_____0___34147));
  xor2s1 ____9________436223(.DIN1 (_________34112), .DIN2
       (_________34127), .Q (_____90__34134));
  hi1s1 ____9__(.DIN (_____0___34423), .Q (______9__34133));
  nor2s1 ____9____9___(.DIN1 (_________34131), .DIN2 (_________34130),
       .Q (_________34132));
  nor2s1 ____9________436224(.DIN1 (________21877), .DIN2
       (_________34117), .Q (_________34129));
  dffacs1 ___________________436225(.CLRB (reset), .CLK (clk), .DIN
       (_________34107), .QN (_____0___34423));
  nnd2s1 ____9______09(.DIN1 (_________34115), .DIN2 (_________34119),
       .Q (_____0___34145));
  nnd2s1 ____9________436226(.DIN1 (_________34127), .DIN2
       (_________34111), .Q (_________34128));
  nor2s1 ____9_____900(.DIN1 (_____9___34039), .DIN2 (_________34109),
       .Q (_____9___34138));
  dffacs1 _____________9_____436227(.CLRB (reset), .CLK (clk), .DIN
       (_________34118), .Q (_________9_______18810));
  nor2s1 ____9______9_436228(.DIN1 (_________34106), .DIN2
       (______9__33899), .Q (_________34126));
  dffacs1 ______________0_____436229(.CLRB (reset), .CLK (clk), .DIN
       (_________34105), .QN (_____9___34414));
  xor2s1 ____9________436230(.DIN1 (_________34108), .DIN2
       (_____9___34038), .Q (_________34125));
  xor2s1 ____9_9______(.DIN1 (_________34099), .DIN2 (______9__34123),
       .Q (______0__34124));
  nor2s1 ____9________436231(.DIN1 (_________34078), .DIN2
       (_________34121), .Q (_________34122));
  nnd2s1 ____9________436232(.DIN1 (_________34121), .DIN2
       (_________34063), .Q (_________34130));
  dffacs1 ___________________436233(.CLRB (reset), .CLK (clk), .DIN
       (______0__34104), .QN (_________________18797));
  nnd2s1 ____9_9___9__(.DIN1 (______9__34113), .DIN2 (_________34119),
       .Q (_________34120));
  nnd2s1 ____9______0_436234(.DIN1 (______9__34103), .DIN2
       (___99___22530), .Q (_________34118));
  and2s1 ____9________436235(.DIN1 (_________34116), .DIN2
       (__________0_______18816), .Q (_________34117));
  nnd2s1 ____9_0______436236(.DIN1 (______0__34114), .DIN2
       (______9__34113), .Q (_________34115));
  and2s1 ____9_______436237(.DIN1 (_________34111), .DIN2
       (_________34110), .Q (_________34112));
  and2s1 ____9_____0__436238(.DIN1 (_________34108), .DIN2
       (_____9___34037), .Q (_________34109));
  nnd2s1 ____9_9____0_(.DIN1 (_________34100), .DIN2 (_________34365),
       .Q (_________34107));
  nnd2s1 ____9______9_436239(.DIN1 (_________34102), .DIN2
       (_________34080), .Q (_________34127));
  dffacs1 _____________9_____436240(.CLRB (reset), .CLK (clk), .DIN
       (_________34101), .Q (_________9_______18811));
  xor2s1 ____9________436241(.DIN1 (_________34088), .DIN2
       (______9__33982), .Q (_________34106));
  nnd2s1 ____9_______436242(.DIN1 (_________34093), .DIN2
       (_________34365), .Q (_________34105));
  nnd2s1 ____9_0___0_9(.DIN1 (_________34092), .DIN2 (________20524),
       .Q (______0__34104));
  nnd2s1 ____9________436243(.DIN1 (_________34091), .DIN2
       (____99___34524), .Q (_________34121));
  dffacs1 _____________9____(.CLRB (reset), .CLK (clk), .DIN
       (_________34089), .Q (_________18851));
  dffacs1 ______________0_____436244(.CLRB (reset), .CLK (clk), .DIN
       (_________34086), .QN (__________0_______18816));
  nnd2s1 ____9____990_436245(.DIN1 (_________34087), .DIN2
       (_________34159), .Q (______9__34103));
  nnd2s1 ____9_______436246(.DIN1 (_________34083), .DIN2
       (_____9___34042), .Q (_________34102));
  nnd2s1 ____9_9____9_436247(.DIN1 (_________34081), .DIN2
       (____00__23084), .Q (_________34101));
  nnd2s1 ____9________436248(.DIN1 (______9__34094), .DIN2
       (______0__34095), .Q (_________34111));
  xnr2s1 ____9________436249(.DIN1 (________19986), .DIN2
       (______0__34075), .Q (______9__34113));
  xor2s1 ____9________436250(.DIN1 (_________34090), .DIN2
       (_________33995), .Q (_________34100));
  xor2s1 ____00___9___(.DIN1 (_________34070), .DIN2 (outData[31]), .Q
       (_________34099));
  nor2s1 ____99_______(.DIN1 (_________34097), .DIN2 (_________34096),
       .Q (_________34098));
  xor2s1 ____9______436251(.DIN1 (_________34076), .DIN2
       (____9____30874), .Q (_________34108));
  or2s1 ____9________436252(.DIN1 (______0__34095), .DIN2
       (______9__34094), .Q (_________34110));
  dffacs1 ________________436253(.CLRB (reset), .CLK (clk), .DIN
       (______0__34085), .QN (outData[16]));
  xor2s1 ____9_____436254(.DIN1 (_________34082), .DIN2
       (_____9___34043), .Q (_________34093));
  nnd2s1 ____9______9_436255(.DIN1 (_________34068), .DIN2
       (_________34071), .Q (_________34092));
  or2s1 ____990______(.DIN1 (_________33977), .DIN2 (_________34090),
       .Q (_________34091));
  nnd2s1 ____99_______436256(.DIN1 (_____0___29271), .DIN2
       (_________34072), .Q (_________34089));
  nnd2s1 ____99_______436257(.DIN1 (______9__34074), .DIN2
       (_________33910), .Q (______0__34114));
  xor2s1 ____9_0______436258(.DIN1
       (____________________________________18836), .DIN2
       (__________________________________0), .Q (_________34088));
  xor2s1 ____9_____9__(.DIN1 (_________34062), .DIN2 (______0__34988),
       .Q (_________34087));
  nor2s1 ____9______0_436259(.DIN1 (_________34187), .DIN2
       (_________34067), .Q (_________34086));
  nnd2s1 ____9________436260(.DIN1 (_________34066), .DIN2
       (______9__34084), .Q (______0__34085));
  or2s1 ____9________436261(.DIN1 (_________34079), .DIN2
       (_________34082), .Q (_________34083));
  nnd2s1 ____99______0(.DIN1 (______0__34065), .DIN2 (_________34159),
       .Q (_________34081));
  nnd2s1 ____9_9___0__(.DIN1 (_________34082), .DIN2 (_________34079),
       .Q (_________34080));
  nor2s1 ____0______0_(.DIN1 (______9__34064), .DIN2 (_________34131),
       .Q (_________34078));
  xor2s1 ____0______9_(.DIN1 (_________34057), .DIN2 (_________34077),
       .Q (_________34096));
  xor2s1 ____99_______436262(.DIN1 (_________33912), .DIN2
       (_________34073), .Q (______0__34095));
  nnd2s1 ____999_____0(.DIN1 (_________34061), .DIN2 (_________32077),
       .Q (_________34076));
  and2s1 ____9_____0_436263(.DIN1
       (______________________________________0_____________18885),
       .DIN2 (__________________________________0), .Q
       (______0__34075));
  nnd2s1 ____00_______(.DIN1 (_________34073), .DIN2 (_________33911),
       .Q (______9__34074));
  or2s1 ____9____990_436264(.DIN1
       (__________________________________0), .DIN2
       (______________________________________0_____________18885), .Q
       (_________34119));
  or2s1 ____00______0(.DIN1 (_________34071), .DIN2 (_________34058),
       .Q (_________34072));
  xor2s1 ____0______9_436265(.DIN1 (_____0___34048), .DIN2
       (_________34069), .Q (_________34070));
  xor2s1 ____00_______436266(.DIN1 (_________34012), .DIN2
       (_____0___34051), .Q (_________34068));
  xor2s1 ____00_______436267(.DIN1 (_____0___34050), .DIN2
       (________35107), .Q (_________34090));
  dffacs1 ________________436268(.CLRB (reset), .CLK (clk), .DIN
       (_________34059), .QN (_____________18896));
  xor2s1 ____99_______436269(.DIN1 (_____0___34047), .DIN2
       (_____0___34052), .Q (_________34067));
  nor2s1 ____99___9___(.DIN1 (_____9__21738), .DIN2 (_____09__34054),
       .Q (_________34066));
  xor2s1 ____00_______436270(.DIN1 (_____90__32086), .DIN2
       (_________34060), .Q (______0__34065));
  hi1s1 ____0__(.DIN (_________34063), .Q (______9__34064));
  nnd2s1 ____00_____09(.DIN1 (_____0___34053), .DIN2 (_____0___34046),
       .Q (_________34082));
  xor2s1 ____00_______436271(.DIN1 (______0__32026), .DIN2
       (_________34033), .Q (_________34062));
  or2s1 ____009___900(.DIN1 (______9__32075), .DIN2 (_________34060),
       .Q (_________34061));
  nnd2s1 ____99_____9_(.DIN1 (_____00__34045), .DIN2 (____0___20137),
       .Q (_________34059));
  dffacs1 _____________9___0_436272(.CLRB (reset), .CLK (clk), .DIN
       (_____99__34044), .Q (__________________________________0));
  nor2s1 ____0________(.DIN1 (_____9___34040), .DIN2 (_____0__20362),
       .Q (_________34058));
  nnd2s1 ____0________436273(.DIN1 (______0__34055), .DIN2
       (_________34056), .Q (_________34057));
  nor2s1 ____0________436274(.DIN1 (_________34024), .DIN2
       (_____9___34041), .Q (_________34073));
  nor2s1 ____0________436275(.DIN1 (_________34056), .DIN2
       (______0__34055), .Q (_________34097));
  nnd2s1 ____0_0___9__(.DIN1 (______9__34026), .DIN2 (____99___34523),
       .Q (_________34063));
  and2s1 ____0______0_436276(.DIN1 (_________34116), .DIN2
       (__________0_______18815), .Q (_____09__34054));
  or2s1 ____0________436277(.DIN1 (______9__34035), .DIN2
       (_____0___34052), .Q (_____0___34053));
  nor2s1 ____0________436278(.DIN1 (_________34028), .DIN2
       (_____0___34049), .Q (_____0___34051));
  or2s1 ____0_______0(.DIN1 (_____0___34049), .DIN2 (_________34029),
       .Q (_____0___34050));
  xor2s1 ____0_____0__(.DIN1 (_____________0___18784), .DIN2
       (______0__34027), .Q (_____0___34048));
  nnd2s1 ____0______0_436279(.DIN1 (_________34034), .DIN2
       (_____0___34046), .Q (_____0___34047));
  nnd2s1 ____0______9_436280(.DIN1 (_________34116), .DIN2
       (_____9___34415), .Q (_____00__34045));
  or2s1 ____0_0______(.DIN1 (_________33989), .DIN2 (_________34031),
       .Q (_____99__34044));
  xnr2s1 ____0_______436281(.DIN1 (_________34079), .DIN2
       (_____9___34042), .Q (_____9___34043));
  nnd2s1 ____0_____0_9(.DIN1 (_________34032), .DIN2 (_____9___31990),
       .Q (_________34060));
  nor2s1 ____0________436282(.DIN1 (_________34023), .DIN2
       (_________34030), .Q (_____9___34041));
  xnr2s1 ____0____990_(.DIN1 (___00___19775), .DIN2
       (_________________18796), .Q (_____9___34040));
  nor2s1 ____0_9_____0(.DIN1 (_____90__34036), .DIN2 (_____9___34038),
       .Q (_____9___34039));
  nnd2s1 ____0_9______(.DIN1 (_____9___34038), .DIN2 (_____90__34036),
       .Q (_____9___34037));
  xor2s1 ____0________436283(.DIN1 (_________34021), .DIN2
       (_________31290), .Q (_________34056));
  dffacs1 ______________0_____436284(.CLRB (reset), .CLK (clk), .DIN
       (_________34025), .QN (__________0_______18815));
  hi1s1 ____0__436285(.DIN (_________34034), .Q (______9__34035));
  xnr2s1 ____0_0______436286(.DIN1 (_________________18795), .DIN2
       (____0____34562), .Q (_________34033));
  xor2s1 ____0____9___(.DIN1 (_________34011), .DIN2 (___0____21656),
       .Q (_____0___34049));
  nnd2s1 ____0________436287(.DIN1 (____0____34562), .DIN2
       (_________32011), .Q (_________34032));
  nnd2s1 ____0______09(.DIN1 (_________33890), .DIN2 (______0__34018),
       .Q (_________34031));
  dffacs1 ______________0_____436288(.CLRB (reset), .CLK (clk), .DIN
       (_________34019), .QN (_____9___34415));
  nor2s1 ____0________436289(.DIN1 (____99__19301), .DIN2
       (_________34015), .Q (_________34030));
  nnd2s1 ____0_____900(.DIN1 (_________30596), .DIN2 (______9__34017),
       .Q (_________34034));
  nor2s1 ____0______9_436290(.DIN1 (_________34028), .DIN2
       (_________34013), .Q (_________34029));
  nor2s1 ____0________436291(.DIN1 (_________33785), .DIN2
       (_________34010), .Q (______0__34027));
  dffacs1 ___________________436292(.CLRB (reset), .CLK (clk), .DIN
       (______0__34008), .QN (_________18850));
  hi1s1 ____0__436293(.DIN (_________________18796), .Q
       (_____90__34036));
  nor2s1 ____0_9______436294(.DIN1 (_________34022), .DIN2
       (______9__34026), .Q (_________34131));
  dffacs1 ________________436295(.CLRB (reset), .CLK (clk), .DIN
       (_________34020), .QN (_____________18895));
  nor2s1 ____0________436296(.DIN1 (_________34187), .DIN2
       (_________34003), .Q (_________34025));
  and2s1 ____0________436297(.DIN1 (_________34005), .DIN2
       (_________34023), .Q (_________34024));
  nnd2s1 ____0_9___9__(.DIN1 (_________30535), .DIN2 (_________34016),
       .Q (_____0___34046));
  xnr2s1 ____09_____0_(.DIN1 (_____________0___18784), .DIN2
       (_________34009), .Q (_________34021));
  xor2s1 ____0________436298(.DIN1 (_________34014), .DIN2
       (_________34004), .Q (_________34079));
  dffacs1 ___________________436299(.CLRB (reset), .CLK (clk), .DIN
       (_________34002), .QN (_________________18796));
  nnd2s1 ____0________436300(.DIN1 (_________34000), .DIN2
       (_____9__20903), .Q (_________34020));
  nnd2s1 ____0_______436301(.DIN1 (_________34001), .DIN2
       (_________34393), .Q (_________34019));
  nnd2s1 ____0_9___0__(.DIN1 (_________33797), .DIN2 (______0__33999),
       .Q (______0__34018));
  hi1s1 ____0__436302(.DIN (_________34016), .Q (______9__34017));
  nor2s1 ____0______0_436303(.DIN1 (____9___19300), .DIN2
       (_________34014), .Q (_________34015));
  hi1s1 _____0_(.DIN (_________34012), .Q (_________34013));
  nnd2s1 ____0________436304(.DIN1 (_________34006), .DIN2
       (______9__34007), .Q (_________34011));
  nor2s1 _____0______436305(.DIN1 (_________33780), .DIN2
       (_________34009), .Q (_________34010));
  nnd2s1 ____0_____0_436306(.DIN1 (_________33994), .DIN2
       (_________33916), .Q (______0__34008));
  xor2s1 ____09_______(.DIN1 (_________33987), .DIN2 (_____0___31191),
       .Q (_________34022));
  nor2s1 ____0____990_436307(.DIN1 (_____0___33957), .DIN2
       (_________33997), .Q (_____0___34052));
  nor2s1 ____0_______436308(.DIN1 (______9__34007), .DIN2
       (_________34006), .Q (_________34028));
  nor2s1 ____0______9_436309(.DIN1 (_________34004), .DIN2
       (_________33998), .Q (_________34005));
  xor2s1 ____0_0______436310(.DIN1 (_________33996), .DIN2
       (_____0___33958), .Q (_________34003));
  xor2s1 ____0________436311(.DIN1 (_________33985), .DIN2
       (_________31281), .Q (_________34016));
  nnd2s1 ____0________436312(.DIN1 (_________33988), .DIN2
       (________19990), .Q (_________34002));
  xor2s1 _________9___436313(.DIN1 (_________33981), .DIN2
       (_____0___33866), .Q (_________34012));
  dffacs1 _____________9_____436314(.CLRB (reset), .CLK (clk), .DIN
       (______9__33990), .Q
       (____________________________________18836));
  xor2s1 ____0________436315(.DIN1 (_________33970), .DIN2
       (______0__33963), .Q (_________34001));
  nnd2s1 ____0______436316(.DIN1 (_________34116), .DIN2
       (_____9___34416), .Q (_________34000));
  nnd2s1 ____0_0______436317(.DIN1 (_________33986), .DIN2 (inData[8]),
       .Q (______0__33999));
  hi1s1 ____0__436318(.DIN (_________33998), .Q (_________34014));
  and2s1 ____0______9_436319(.DIN1 (_________33996), .DIN2
       (_____9___33947), .Q (_________33997));
  nnd2s1 _____________436320(.DIN1 (_________33976), .DIN2
       (____99___34524), .Q (_________33995));
  nor2s1 _____00______(.DIN1 (________23574), .DIN2 (_________33978),
       .Q (_________33994));
  xor2s1 ____09_______436321(.DIN1 (_________33969), .DIN2
       (_____9___32930), .Q (______9__34007));
  nor2s1 _____________436322(.DIN1 (____09___33762), .DIN2
       (_________33980), .Q (_________34009));
  nor2s1 ____0_____9__(.DIN1 (_________33993), .DIN2 (_________33992),
       .Q (_____9___34142));
  nnd2s1 ____0______0_436323(.DIN1 (_________33974), .DIN2
       (_____00__33954), .Q (______0__33991));
  or2s1 ____0_9______436324(.DIN1 (_________33989), .DIN2
       (_________33971), .Q (______9__33990));
  nnd2s1 ____099______(.DIN1 (_________33968), .DIN2 (_________34071),
       .Q (_________33988));
  xor2s1 ____________436325(.DIN1 (_________33979), .DIN2
       (_________34435), .Q (_________33987));
  nnd2s1 ____0_0___0__(.DIN1 (______0__33973), .DIN2 (________19073),
       .Q (_________33998));
  dffacs1 ______________0_____436326(.CLRB (reset), .CLK (clk), .DIN
       (_________33967), .QN (_____9___34416));
  xor2s1 ____0______0_436327(.DIN1 (_________9_______18808), .DIN2
       (____________________________________18836), .Q
       (_________33986));
  xor2s1 ____0______9_436328(.DIN1 (_________9_______18806), .DIN2
       (______9__33972), .Q (_________33985));
  nnd2s1 ____0_____0_436329(.DIN1 (_________33975), .DIN2
       (_________9_______18809), .Q (______9__33982));
  nor2s1 _____________436330(.DIN1 (_____0___33961), .DIN2
       (_____9___33949), .Q (_________33981));
  nor2s1 _________990_436331(.DIN1 (____09___33760), .DIN2
       (_________33979), .Q (_________33980));
  nor2s1 ____________436332(.DIN1 (______0__33918), .DIN2
       (_____0___33959), .Q (_________33978));
  hi1s1 _______436333(.DIN (_________33976), .Q (_________33977));
  nor2s1 ____09_______436334(.DIN1 (_________33966), .DIN2
       (_________33964), .Q (_________33996));
  nor2s1 ____09_______436335(.DIN1 (_________33975), .DIN2
       (_________31940), .Q (_________33992));
  xor2s1 ____0_9______436336(.DIN1 (_________32014), .DIN2
       (_____09__33962), .Q (_________33974));
  nnd2s1 ____0____9___436337(.DIN1 (______9__33972), .DIN2
       (________19093), .Q (______0__33973));
  nnd2s1 ____0________436338(.DIN1 (_____0___33955), .DIN2
       (____99__21259), .Q (_________33971));
  nnd2s1 ____09_____09(.DIN1 (_________33940), .DIN2 (_________33965),
       .Q (_________33970));
  xor2s1 _____________436339(.DIN1 (_____9___33952), .DIN2
       (_________28828), .Q (_________33969));
  xor2s1 __________436340(.DIN1 (_____9___33951), .DIN2
       (_____0___33960), .Q (_________33968));
  nnd2s1 ___________9_436341(.DIN1 (_____0___32202), .DIN2
       (_____0___33956), .Q (_________33976));
  nor2s1 ____09_______436342(.DIN1 (_________9_______18808), .DIN2
       (_______________18881), .Q (_________33993));
  nnd2s1 ____090______(.DIN1 (_____99__33953), .DIN2 (_________34365),
       .Q (_________33967));
  hi1s1 _____0_436343(.DIN (_________33965), .Q (_________33966));
  nor2s1 _____0_______436344(.DIN1 (______0__33963), .DIN2
       (_________33941), .Q (_________33964));
  hi1s1 ____09_(.DIN (_________9_______18808), .Q (_________33975));
  nnd2s1 _____0_______436345(.DIN1 (_____9___31988), .DIN2
       (_____09__33962), .Q (_________33984));
  nor2s1 __________9__436346(.DIN1 (_____9___33950), .DIN2
       (_____0___33960), .Q (_____0___33961));
  xor2s1 ___________0_436347(.DIN1 (_________33939), .DIN2
       (____0____34568), .Q (_____0___33959));
  nor2s1 ______0______436348(.DIN1 (_____0___33957), .DIN2
       (_____9___33948), .Q (_____0___33958));
  nnd2s1 _____________436349(.DIN1 (_____9___33946), .DIN2
       (______0__31238), .Q (_________33979));
  nnd2s1 _____0______436350(.DIN1 (_________33942), .DIN2
       (_____00__33954), .Q (_____0___33955));
  dffacs1 _____________9_____436351(.CLRB (reset), .CLK (clk), .DIN
       (_____90__33944), .QN (_________9_______18808));
  nnd2s1 _____09___0__(.DIN1 (_________30473), .DIN2 (______9__33943),
       .Q (_________33965));
  xor2s1 ___________0_436352(.DIN1 (_________33931), .DIN2
       (____9____32728), .Q (______9__33972));
  xor2s1 ___________9_436353(.DIN1 (_________31240), .DIN2
       (_____9___33945), .Q (_____0___33956));
  xor2s1 _____0_______436354(.DIN1 (______9__33926), .DIN2
       (____9____31798), .Q (_____99__33953));
  nnd2s1 ____________436355(.DIN1 (____0____34566), .DIN2
       (____0____34564), .Q (______0__33963));
  nnd2s1 __________0_436356(.DIN1 (______0__33935), .DIN2
       (_____09__31909), .Q (_____09__33962));
  dffacs1 ___________________436357(.CLRB (reset), .CLK (clk), .DIN
       (_________33932), .Q (_________________18795));
  xor2s1 _____________436358(.DIN1 (_________33927), .DIN2
       (____9_0__33587), .Q (_____9___33952));
  or2s1 _________990_436359(.DIN1 (_____9___33950), .DIN2
       (_____9___33949), .Q (_____9___33951));
  hi1s1 ______9(.DIN (_____9___33947), .Q (_____9___33948));
  nnd2s1 ______0_____436360(.DIN1 (_____9___33945), .DIN2
       (_________31239), .Q (_____9___33946));
  nor2s1 ___________9_436361(.DIN1 (_________33930), .DIN2
       (_________33938), .Q (_____0___33960));
  nnd2s1 _____________436362(.DIN1 (_________33928), .DIN2
       (____9___21161), .Q (_____90__33944));
  xor2s1 ______0______436363(.DIN1 (_________33933), .DIN2
       (____0____31872), .Q (______9__33943));
  xor2s1 _____________436364(.DIN1 (______0__31929), .DIN2
       (______9__33934), .Q (_________33942));
  hi1s1 _______436365(.DIN (_________33940), .Q (_________33941));
  or2s1 ______9__9___(.DIN1 (_________33929), .DIN2 (_________33938),
       .Q (_________33939));
  nor2s1 _____________436366(.DIN1 (_________33936), .DIN2
       (_________33937), .Q (_____0___33957));
  nnd2s1 ___________436367(.DIN1 (_________33937), .DIN2
       (_________33936), .Q (_____9___33947));
  or2s1 ______9___900(.DIN1 (______9__33934), .DIN2 (______9__31928),
       .Q (______0__33935));
  nnd2s1 ___________9_436368(.DIN1 (______9__30474), .DIN2
       (_________33933), .Q (_________33940));
  dffacs1 ___________________436369(.CLRB (reset), .CLK (clk), .DIN
       (______9__33917), .QN (_____0___34424));
  or2s1 _____________436370(.DIN1 (________23668), .DIN2
       (_________33919), .Q (_________33932));
  nor2s1 _____________436371(.DIN1 (______0__33799), .DIN2
       (_________33924), .Q (_________33931));
  nor2s1 _____________436372(.DIN1 (____0____34568), .DIN2
       (_________33929), .Q (_________33930));
  xor2s1 ______0______436373(.DIN1 (_________33913), .DIN2
       (____0____32762), .Q (_____9___33949));
  nor2s1 ______9___9__(.DIN1 (______9__31110), .DIN2 (_________33921),
       .Q (_____9___33945));
  nnd2s1 ___________0_436374(.DIN1 (_________33914), .DIN2
       (_____00__33954), .Q (_________33928));
  xor2s1 ______9______436375(.DIN1 (_________33800), .DIN2
       (_________33923), .Q (_________33936));
  dffacs1 _____________9_____436376(.CLRB (reset), .CLK (clk), .DIN
       (_________33915), .QN (_________9_______18807));
  xnr2s1 _____________436377(.DIN1 (_________________18782), .DIN2
       (_________33920), .Q (_________33927));
  xor2s1 ______0___0__(.DIN1 (_________33922), .DIN2 (______9__33882),
       .Q (______9__33926));
  xor2s1 ___________0_436378(.DIN1 (_________33905), .DIN2
       (_________33925), .Q (_________33938));
  and2s1 ___________9_436379(.DIN1 (_________33923), .DIN2
       (______9__33788), .Q (_________33924));
  xor2s1 ____________436380(.DIN1 (_________33897), .DIN2
       (_______________18878), .Q (_________33933));
  nor2s1 __________0_436381(.DIN1 (_________31711), .DIN2
       (_________33907), .Q (______9__33934));
  nor2s1 _____________436382(.DIN1 (_________31125), .DIN2
       (_________33920), .Q (_________33921));
  nor2s1 _________990_436383(.DIN1 (______0__33918), .DIN2
       (_________33904), .Q (_________33919));
  nnd2s1 ____________436384(.DIN1 (_________33903), .DIN2
       (_________33916), .Q (______9__33917));
  nnd2s1 _____________436385(.DIN1 (_________33791), .DIN2
       (______0__33900), .Q (_________33915));
  xor2s1 _____________436386(.DIN1 (_________31712), .DIN2
       (_________33906), .Q (_________33914));
  nor2s1 _____________436387(.DIN1 (_________33902), .DIN2
       (_____0___31999), .Q (_________33929));
  nnd2s1 _____90__9___(.DIN1 (______9__33908), .DIN2 (______0__33909),
       .Q (_________33913));
  and2s1 ___________436388(.DIN1 (_________33911), .DIN2
       (_________33910), .Q (_________33912));
  nor2s1 _____9_______436389(.DIN1 (______0__33909), .DIN2
       (______9__33908), .Q (_____9___33950));
  and2s1 __________436390(.DIN1 (_________33906), .DIN2
       (_________31693), .Q (_________33907));
  nor2s1 _____09____9_(.DIN1 (_________33901), .DIN2 (_____0___32000),
       .Q (_________33905));
  nor2s1 _____________436391(.DIN1 (_________33896), .DIN2
       (_________33889), .Q (_________33923));
  dffacs1 ________________436392(.CLRB (reset), .CLK (clk), .DIN
       (_________33886), .QN (outData[13]));
  xor2s1 _____9_______436393(.DIN1 (_________33885), .DIN2
       (_____9___30624), .Q (_________33904));
  nor2s1 _____________436394(.DIN1 (___9_0__23386), .DIN2
       (_________33887), .Q (_________33903));
  nnd2s1 _____0____9__436395(.DIN1 (______9__33892), .DIN2
       (______0__31044), .Q (_________33920));
  nnd2s1 ___________0_436396(.DIN1 (_________33898), .DIN2
       (_________33881), .Q (_________33922));
  hi1s1 ______0(.DIN (_________33901), .Q (_________33902));
  or2s1 _____________436397(.DIN1 (_________33884), .DIN2
       (______9__33899), .Q (______0__33900));
  xor2s1 _____________436398(.DIN1 (_________31045), .DIN2
       (_________33891), .Q (______0__33909));
  nor2s1 ____________436399(.DIN1 (_________33888), .DIN2
       (_________33896), .Q (_________33897));
  xor2s1 __________0__436400(.DIN1 (_________33875), .DIN2
       (_________33895), .Q (_________33911));
  or2s1 _____________436401(.DIN1 (____0____30970), .DIN2
       (_________33891), .Q (______9__33892));
  nnd2s1 ______9_____436402(.DIN1 (_________33876), .DIN2
       (_____00__33954), .Q (_________33890));
  xor2s1 __________0_436403(.DIN1 (______0__33874), .DIN2
       (___9____24307), .Q (_________33901));
  nor2s1 ______0______436404(.DIN1 (_________31058), .DIN2
       (_________33888), .Q (_________33889));
  nor2s1 ______9__990_(.DIN1 (______0__33918), .DIN2 (_________33880),
       .Q (_________33887));
  nnd2s1 ____________436405(.DIN1 (_________33879), .DIN2
       (______9__34084), .Q (_________33886));
  xnr2s1 ___________9_436406(.DIN1 (_________33895), .DIN2
       (____0_0__34570), .Q (_________33906));
  nnd2s1 _____________436407(.DIN1 (_____0___33872), .DIN2
       (_________33877), .Q (_________33898));
  xor2s1 _____________436408(.DIN1 (_____0___33869), .DIN2
       (_________33878), .Q (_________33885));
  xor2s1 _____________436409(.DIN1
       (_____________________________________18838), .DIN2
       (____0____33753), .Q (_________33884));
  and2s1 _____9___9___(.DIN1 (______9__33882), .DIN2 (_________33881),
       .Q (______0__33883));
  nor2s1 _____00______436410(.DIN1 (_________9_______18805), .DIN2
       (_____0___33871), .Q (_________33896));
  xor2s1 _____0_____436411(.DIN1 (_____9___33863), .DIN2
       (_________33832), .Q (_________33880));
  nor2s1 _____________436412(.DIN1 (________21869), .DIN2
       (_____00__33865), .Q (_________33879));
  xor2s1 __________436413(.DIN1 (_____9___33862), .DIN2
       (_________28828), .Q (_________33891));
  and2s1 ___________9_436414(.DIN1 (_________33878), .DIN2
       (_____0___33868), .Q (______0__33893));
  xor2s1 _____9_______436415(.DIN1 (_____09__33873), .DIN2
       (_________33385), .Q (_________33877));
  xor2s1 _____________436416(.DIN1 (_____99__33864), .DIN2
       (_________30166), .Q (_________33876));
  nor2s1 _____99______436417(.DIN1
       (_____________________________________18838), .DIN2
       (______________________________________0_____________18886), .Q
       (_________33875));
  nnd2s1 _____9_______436418(.DIN1
       (______________________________________0_____________18886),
       .DIN2 (_____________________________________18838), .Q
       (_________33910));
  nor2s1 _____9____9__436419(.DIN1 (____99___33668), .DIN2
       (_____0___33870), .Q (_________33888));
  xor2s1 ______9____0_436420(.DIN1 (_____9___33859), .DIN2
       (_________33852), .Q (______0__33874));
  or2s1 ______0______436421(.DIN1 (_____09__33873), .DIN2
       (_____0___33872), .Q (_________33881));
  hi1s1 _____0_436422(.DIN (_____0___33870), .Q (_____0___33871));
  and2s1 ____________436423(.DIN1 (_____0___33868), .DIN2
       (_____0___33867), .Q (_____0___33869));
  xor2s1 __________0__436424(.DIN1 (_________33854), .DIN2
       (_____0___33866), .Q (_____0___33870));
  nnd2s1 ___________0_436425(.DIN1 (_____9___33860), .DIN2
       (_________33842), .Q (_________33878));
  and2s1 ___________9_436426(.DIN1 (_________34116), .DIN2
       (______9__34498), .Q (_____00__33865));
  dffacs1 _____________9___9_436427(.CLRB (reset), .CLK (clk), .DIN
       (_____9___33861), .QN
       (_____________________________________18838));
  dffacs1 ________________436428(.CLRB (reset), .CLK (clk), .DIN
       (_____9___33857), .QN (_____________18894));
  xor2s1 _____________436429(.DIN1 (______9__33848), .DIN2
       (_________31697), .Q (_____99__33864));
  xor2s1 __________0_436430(.DIN1 (_________33841), .DIN2
       (_________33845), .Q (_____9___33863));
  nor2s1 _____________436431(.DIN1 (_____9___33858), .DIN2
       (_________33853), .Q (_____9___33862));
  xor2s1 _________990_436432(.DIN1 (_________33847), .DIN2
       (_________33835), .Q (_____09__33873));
  or2s1 ____________436433(.DIN1 (_________33989), .DIN2
       (_________33849), .Q (_____9___33861));
  or2s1 ___________9_436434(.DIN1 (_________33840), .DIN2
       (_________33831), .Q (_____9___33860));
  nnd2s1 _____________436435(.DIN1 (____0____31868), .DIN2
       (_________33844), .Q (_____0___33867));
  nor2s1 ______9______436436(.DIN1 (_____9___33858), .DIN2
       (______9__33838), .Q (_____9___33859));
  dffacs1 ______________0_____436437(.CLRB (reset), .CLK (clk), .DIN
       (_________33851), .Q (______9__34498));
  nnd2s1 _____0_______436438(.DIN1 (_________33850), .DIN2
       (________20121), .Q (_____9___33857));
  nor2s1 ___________436439(.DIN1 (_________33846), .DIN2
       (_________33836), .Q (_________33854));
  and2s1 _____________436440(.DIN1 (_________33837), .DIN2
       (_________33852), .Q (_________33853));
  nnd2s1 __________436441(.DIN1 (____0____31869), .DIN2
       (_________33843), .Q (_____0___33868));
  dffacs1 ___________________436442(.CLRB (reset), .CLK (clk), .DIN
       (_________33834), .Q (_________________18794));
  nnd2s1 ___________9_436443(.DIN1 (______0__33829), .DIN2
       (_________34393), .Q (_________33851));
  nnd2s1 _____________436444(.DIN1 (_________33817), .DIN2
       (__________0_____), .Q (_________33850));
  nnd2s1 _____________436445(.DIN1 (_________33824), .DIN2
       (______9__33798), .Q (_________33849));
  xor2s1 _____________436446(.DIN1 (_________33833), .DIN2
       (_____0___34426), .Q (______9__33848));
  or2s1 _____________436447(.DIN1 (_________33846), .DIN2
       (_________33826), .Q (_________33847));
  xor2s1 __________9__436448(.DIN1 (_________33823), .DIN2
       (_________33444), .Q (_________33845));
  hi1s1 _______436449(.DIN (_________33843), .Q (_________33844));
  nnd2s1 ___________0_436450(.DIN1 (_________33841), .DIN2
       (______0__33839), .Q (_________33842));
  nor2s1 _____________436451(.DIN1 (______0__33839), .DIN2
       (_________33841), .Q (_________33840));
  hi1s1 ______436452(.DIN (_________33837), .Q (______9__33838));
  dffacs1 ________________436453(.CLRB (reset), .CLK (clk), .DIN
       (_________33827), .QN (___________));
  and2s1 _____________436454(.DIN1 (_________33825), .DIN2
       (_________33835), .Q (_________33836));
  nnd2s1 ____________436455(.DIN1 (_________33821), .DIN2
       (___9_9__23365), .Q (_________33834));
  nnd2s1 __________0__436456(.DIN1 (_________31605), .DIN2
       (_________33833), .Q (_________33855));
  nnd2s1 ______9____0_436457(.DIN1 (_________33822), .DIN2
       (_________33794), .Q (______9__33882));
  xor2s1 ______0____9_436458(.DIN1 (_________33831), .DIN2
       (_________31951), .Q (_________33832));
  xor2s1 _____________436459(.DIN1 (_________33814), .DIN2
       (_________________18781), .Q (_________33843));
  nnd2s1 ____________436460(.DIN1 (_________33830), .DIN2
       (_______________0_____________________18834), .Q
       (_________33837));
  nor2s1 __________0_436461(.DIN1
       (_______________0_____________________18834), .DIN2
       (_________33830), .Q (_____9___33858));
  dffacs1 ______________0_____436462(.CLRB (reset), .CLK (clk), .DIN
       (______0__33819), .Q (__________0_____));
  xor2s1 _____________436463(.DIN1 (_________33813), .DIN2
       (______9__33828), .Q (______0__33829));
  nnd2s1 ______0__990_436464(.DIN1 (______9__33818), .DIN2
       (____99__20323), .Q (_________33827));
  hi1s1 _______436465(.DIN (_________33825), .Q (_________33826));
  nnd2s1 ____________436466(.DIN1 (_________33816), .DIN2
       (_____00__33954), .Q (_________33824));
  hi1s1 _______436467(.DIN (_________33823), .Q (______0__33839));
  dffacs1 ___________________436468(.CLRB (reset), .CLK (clk), .DIN
       (_________33815), .Q (_____0___34425));
  xor2s1 ___________9_436469(.DIN1 (_________33806), .DIN2
       (____99___35108), .Q (_________33822));
  or2s1 _____________436470(.DIN1 (______0__33918), .DIN2
       (_________33810), .Q (_________33821));
  nor2s1 _____________436471(.DIN1 (_________9_______18804), .DIN2
       (_________33820), .Q (_________33846));
  xor2s1 _____9_______436472(.DIN1 (_________33801), .DIN2
       (_________________0___18618), .Q (_________33823));
  nnd2s1 _________9___436473(.DIN1 (_________33812), .DIN2
       (_________31462), .Q (_________33833));
  nnd2s1 _____________436474(.DIN1 (_________33820), .DIN2
       (_________9_______18804), .Q (_________33825));
  nnd2s1 _____9_____436475(.DIN1 (______0__33809), .DIN2
       (____9____33591), .Q (_________33830));
  nor2s1 _____________436476(.DIN1 (_________________0___18660), .DIN2
       (_________33807), .Q (______0__33819));
  nnd2s1 __________436477(.DIN1 (_________33817), .DIN2
       (_____9___34417), .Q (______9__33818));
  xor2s1 ______9____9_436478(.DIN1 (_________31503), .DIN2
       (_________33811), .Q (_________33816));
  nnd2s1 _____________436479(.DIN1 (_________33802), .DIN2
       (_________33916), .Q (_________33815));
  xor2s1 _____0_______436480(.DIN1 (______9__33808), .DIN2
       (____9____33600), .Q (_________33814));
  nor2s1 ______9______436481(.DIN1 (____09___33761), .DIN2
       (_________33804), .Q (_________33831));
  xor2s1 _____________436482(.DIN1 (_________33795), .DIN2
       (_________33805), .Q (_________33813));
  nnd2s1 __________9__436483(.DIN1 (_________33811), .DIN2
       (_________31488), .Q (_________33812));
  xor2s1 ___________0_436484(.DIN1 (_____0___33771), .DIN2
       (_________33803), .Q (_________33810));
  nnd2s1 _____09______(.DIN1 (______9__33808), .DIN2 (____9____33601),
       .Q (______0__33809));
  xor2s1 _____________436485(.DIN1 (_________33793), .DIN2
       (_____0___33866), .Q (_________33820));
  xor2s1 ______0_____436486(.DIN1 (_________33790), .DIN2
       (____0_9__33749), .Q (_________33807));
  dffacs1 ______________0_____436487(.CLRB (reset), .CLK (clk), .DIN
       (_________33796), .QN (_____9___34417));
  nor2s1 __________0__436488(.DIN1 (_____0___33773), .DIN2
       (_________33805), .Q (_________33806));
  nor2s1 ___________0_436489(.DIN1 (____09___33766), .DIN2
       (_________33803), .Q (_________33804));
  nor2s1 _____9_____9_436490(.DIN1 (________23560), .DIN2
       (_________33792), .Q (_________33802));
  xor2s1 _____________436491(.DIN1 (_________33783), .DIN2
       (_________________18780), .Q (_________33801));
  xor2s1 _____9______436492(.DIN1 (_____0___33774), .DIN2
       (_________33384), .Q (_________33811));
  nnd2s1 ______9___0_9(.DIN1 (_________33786), .DIN2 (_________33781),
       .Q (______9__33808));
  dffacs1 ___________________436493(.CLRB (reset), .CLK (clk), .DIN
       (_________33784), .Q (_________________18785));
  dffacs1 ______________0_436494(.CLRB (reset), .CLK (clk), .DIN
       (______0__33789), .QN (outData[10]));
  nor2s1 ______9______436495(.DIN1 (______0__33799), .DIN2
       (_________33787), .Q (_________33800));
  nnd2s1 _________990_436496(.DIN1 (_________33797), .DIN2
       (_____0___33776), .Q (______9__33798));
  nnd2s1 ____________436497(.DIN1 (______0__33779), .DIN2
       (_________34365), .Q (_________33796));
  nor2s1 _____9_____9_436498(.DIN1 (____0____33748), .DIN2
       (_____09__33778), .Q (_________33805));
  nnd2s1 _____0_______436499(.DIN1 (_____0___33772), .DIN2
       (_________33794), .Q (_________33795));
  nnd2s1 _____9_______436500(.DIN1 (_____0___33775), .DIN2
       (____0____33757), .Q (_________33793));
  nor2s1 _____________436501(.DIN1 (______0__33918), .DIN2
       (_____0___33770), .Q (_________33792));
  xor2s1 _____0___9___(.DIN1 (____09___33763), .DIN2 (_________31431),
       .Q (_________33803));
  nnd2s1 _____9_______436502(.DIN1 (____09___33767), .DIN2
       (_____00__33954), .Q (_________33791));
  xor2s1 _____90____09(.DIN1 (_____0___33777), .DIN2 (______0__31325),
       .Q (_________33790));
  nnd2s1 _____________436503(.DIN1 (_____00__33769), .DIN2
       (_________34295), .Q (______0__33789));
  hi1s1 _____0_436504(.DIN (_________33787), .Q (______9__33788));
  nnd2s1 __________436505(.DIN1 (_________33782), .DIN2
       (_________________18780), .Q (_________33786));
  nor2s1 ___________9_436506(.DIN1 (_____________0___18784), .DIN2
       (_______________18884), .Q (_________33785));
  nor2s1 _____________436507(.DIN1 (_________________0___18660), .DIN2
       (____0_9__33758), .Q (_________33784));
  and2s1 _____________436508(.DIN1 (_________33782), .DIN2
       (_________33781), .Q (_________33783));
  and2s1 _____________436509(.DIN1 (_________35111), .DIN2
       (_____________0___18784), .Q (_________33780));
  dffacs1 _____________9_____436510(.CLRB (reset), .CLK (clk), .DIN
       (____099__33768), .Q (_________9_______18806));
  xor2s1 _____0_______436511(.DIN1 (____0____33736), .DIN2
       (____0____33720), .Q (______0__33779));
  nor2s1 _____0____9__436512(.DIN1 (____0____34574), .DIN2
       (_____0___33777), .Q (_____09__33778));
  nnd2s1 _____9_____0_436513(.DIN1 (____0____33754), .DIN2 (inData[0]),
       .Q (_____0___33776));
  nnd2s1 _____________436514(.DIN1 (____0____34572), .DIN2
       (_________34077), .Q (_____0___33775));
  xor2s1 _____0_______436515(.DIN1 (____0____33745), .DIN2
       (________19986), .Q (_________33787));
  nnd2s1 ____________436516(.DIN1 (____0____33756), .DIN2
       (_________31392), .Q (_____0___33774));
  hi1s1 _______436517(.DIN (_____0___33772), .Q (_____0___33773));
  xor2s1 ______0___0__436518(.DIN1 (____09___33764), .DIN2
       (____09___33765), .Q (_____0___33771));
  xor2s1 ___________0_436519(.DIN1 (____0____33738), .DIN2
       (____0_0__33741), .Q (_____0___33770));
  nnd2s1 ______0____9_436520(.DIN1 (____9____29932), .DIN2
       (____0____33751), .Q (_________33794));
  dffacs1 _________________0_436521(.CLRB (reset), .CLK (clk), .DIN
       (____0____33752), .Q (_____0___34426));
  nor2s1 _____0_______436522(.DIN1 (____9___20879), .DIN2
       (____0____33744), .Q (_____00__33769));
  nnd2s1 ______0_____436523(.DIN1 (____0____33747), .DIN2
       (________19628), .Q (____099__33768));
  xor2s1 __________0_436524(.DIN1 (______9__31436), .DIN2
       (____0____33755), .Q (____09___33767));
  nor2s1 _____________436525(.DIN1 (____09___33765), .DIN2
       (____09___33764), .Q (____09___33766));
  nnd2s1 _________990_436526(.DIN1 (____0____33739), .DIN2
       (____0_9__33740), .Q (____09___33763));
  nnd2s1 ______9_____436527(.DIN1 (____9____29933), .DIN2
       (____0____33750), .Q (_____0___33772));
  and2s1 _____9_____9_436528(.DIN1 (____090__33759), .DIN2
       (_________34435), .Q (____09___33762));
  and2s1 _____________436529(.DIN1 (____09___33764), .DIN2
       (____09___33765), .Q (____09___33761));
  nor2s1 _____9_______436530(.DIN1 (_________34435), .DIN2
       (____090__33759), .Q (____09___33760));
  xor2s1 _____9_______436531(.DIN1 (________24540), .DIN2
       (____0____33730), .Q (____0_9__33758));
  nnd2s1 _________9___436532(.DIN1 (____0____33743), .DIN2
       (_____0___30733), .Q (_________33782));
  dffacs1 _________________0_436533(.CLRB (reset), .CLK (clk), .DIN
       (____0____33737), .QN (_____________0___18784));
  dffacs1 _____________9_(.CLRB (reset), .CLK (clk), .DIN
       (____0____33746), .QN (outData[9]));
  or2s1 _____________436534(.DIN1 (_________34077), .DIN2
       (____0_9__33731), .Q (____0____33757));
  nnd2s1 ___________436535(.DIN1 (______9__31399), .DIN2
       (____0____33755), .Q (____0____33756));
  xor2s1 _____________436536(.DIN1 (____0____33753), .DIN2
       (____________________________________18835), .Q
       (____0____33754));
  nnd2s1 __________436537(.DIN1 (____0____33733), .DIN2
       (____0____33735), .Q (_____0___33777));
  nnd2s1 ___________9_436538(.DIN1 (____0____33729), .DIN2
       (_________33916), .Q (____0____33752));
  hi1s1 _______436539(.DIN (____0____33750), .Q (____0____33751));
  nnd2s1 _____________436540(.DIN1 (____0____33742), .DIN2
       (_____9___33396), .Q (_________33781));
  nor2s1 _____________436541(.DIN1 (____0____34574), .DIN2
       (____0____33748), .Q (____0_9__33749));
  nnd2s1 _____________436542(.DIN1 (____0____33727), .DIN2
       (____0_9__33692), .Q (____0____33747));
  nnd2s1 __________9__436543(.DIN1 (____0____33728), .DIN2
       (_________34295), .Q (____0____33746));
  and2s1 ___________0_436544(.DIN1 (_______________18879), .DIN2
       (____________________________________18835), .Q
       (____0____33745));
  and2s1 _____________436545(.DIN1 (_________33817), .DIN2
       (__________0___0_), .Q (____0____33744));
  nor2s1 _____________436546(.DIN1
       (____________________________________18835), .DIN2
       (_______________18879), .Q (______0__33799));
  xor2s1 ____________436547(.DIN1 (________20296), .DIN2
       (____0____33734), .Q (____0____33750));
  hi1s1 _______436548(.DIN (____0____33742), .Q (____0____33743));
  nnd2s1 ______9___0__436549(.DIN1 (____0____33725), .DIN2
       (____0_9__33740), .Q (____0_0__33741));
  or2s1 ___________0_436550(.DIN1 (____0____33726), .DIN2
       (____0____33738), .Q (____0____33739));
  nor2s1 _____00____9_(.DIN1 (_________34187), .DIN2 (____0____33723),
       .Q (____0____33737));
  nnd2s1 ______9______436551(.DIN1 (____0____33735), .DIN2
       (____0_0__33732), .Q (____0____33736));
  xor2s1 ______9_____436552(.DIN1 (____0_9__33711), .DIN2
       (____0____33715), .Q (____09___33765));
  dffacs1 _________________9_436553(.CLRB (reset), .CLK (clk), .DIN
       (____0____33724), .Q (_________34435));
  nnd2s1 _____________436554(.DIN1 (____0____33719), .DIN2
       (____0_0__33732), .Q (____0____33733));
  nnd2s1 _________990_436555(.DIN1 (____0____33734), .DIN2
       (________20295), .Q (____0_9__33731));
  nor2s1 ______9_____436556(.DIN1 (_________31197), .DIN2
       (____0____33718), .Q (____0____33755));
  nor2s1 ___________9_436557(.DIN1 (_________33518), .DIN2
       (____0____33714), .Q (____0____33730));
  nor2s1 _____________436558(.DIN1 (________23673), .DIN2
       (____0_0__33712), .Q (____0____33729));
  nnd2s1 _____________436559(.DIN1 (____0____33716), .DIN2
       (____0____33710), .Q (____0____33742));
  dffacs1 _____________9_____436560(.CLRB (reset), .CLK (clk), .DIN
       (____0_0__33722), .Q (_________9_______18804));
  dffacs1 _______________(.CLRB (reset), .CLK (clk), .DIN
       (____0_9__33721), .QN (outData[8]));
  nor2s1 _____________436561(.DIN1 (___099__20789), .DIN2
       (____0____33706), .Q (____0____33728));
  dffacs1 ______________0___0_436562(.CLRB (reset), .CLK (clk), .DIN
       (____0____33707), .QN (__________0___0_));
  xor2s1 _________9___436563(.DIN1 (_________31280), .DIN2
       (____0____33717), .Q (____0____33727));
  nnd2s1 ______9______436564(.DIN1 (_________29865), .DIN2
       (____0____33705), .Q (____0____33735));
  xor2s1 ______0____436565(.DIN1 (____0____33696), .DIN2
       (_________32901), .Q (____0____33748));
  dffacs1 _____________9_____436566(.CLRB (reset), .CLK (clk), .DIN
       (____0____33708), .Q
       (____________________________________18835));
  hi1s1 _____436567(.DIN (____0____33725), .Q (____0____33726));
  nnd2s1 _____________436568(.DIN1 (____0_9__33701), .DIN2
       (_________34365), .Q (____0____33724));
  xor2s1 __________436569(.DIN1 (_________33519), .DIN2
       (____0____33713), .Q (____0____33723));
  xor2s1 ___________9_436570(.DIN1 (____0____33695), .DIN2
       (_________33204), .Q (____0____33738));
  nnd2s1 _____9_______436571(.DIN1 (_________31555), .DIN2
       (____0____33703), .Q (____0_9__33740));
  dffacs1 _________________9_436572(.CLRB (reset), .CLK (clk), .DIN
       (____0____33700), .QN (_____0___34427));
  or2s1 _____________436573(.DIN1 (____99___33669), .DIN2
       (____0____33697), .Q (____0_0__33722));
  nnd2s1 _____________436574(.DIN1 (____0____33699), .DIN2
       (_________34295), .Q (____0_9__33721));
  xnr2s1 _____________436575(.DIN1 (_________31431), .DIN2
       (____0____33719), .Q (____0____33720));
  nor2s1 __________9__436576(.DIN1 (_____9___31177), .DIN2
       (____0____33717), .Q (____0____33718));
  nnd2s1 ___________0_436577(.DIN1 (_________29866), .DIN2
       (____0____33704), .Q (____0_0__33732));
  nnd2s1 _____0_______436578(.DIN1 (____0____33709), .DIN2
       (____0____33715), .Q (____0____33716));
  nor2s1 _____________436579(.DIN1 (_________33517), .DIN2
       (____0____33713), .Q (____0____33714));
  nor2s1 _____9______436580(.DIN1 (______0__33918), .DIN2
       (____0____33698), .Q (____0_0__33712));
  and2s1 _____0____0__(.DIN1 (____0____33710), .DIN2 (____0____33709),
       .Q (____0_9__33711));
  nnd2s1 _____9_____0_436581(.DIN1 (_________31556), .DIN2
       (____0_0__33702), .Q (____0____33725));
  xor2s1 ______0____9_436582(.DIN1 (____0____33690), .DIN2
       (____0____32823), .Q (____0____33734));
  nnd2s1 _____________436583(.DIN1 (____0_0__33693), .DIN2
       (___0____20774), .Q (____0____33708));
  nor2s1 ____________436584(.DIN1 (_________________0___18660), .DIN2
       (____0____33691), .Q (____0____33707));
  and2s1 __________0_436585(.DIN1 (_________33817), .DIN2
       (__________0__9_), .Q (____0____33706));
  hi1s1 _______436586(.DIN (____0____33704), .Q (____0____33705));
  hi1s1 _____436587(.DIN (____0_0__33702), .Q (____0____33703));
  xor2s1 _____________436588(.DIN1 (____00___33682), .DIN2
       (_________29500), .Q (____0_9__33701));
  nnd2s1 _________990_436589(.DIN1 (____0____33688), .DIN2
       (____9____33613), .Q (____0____33700));
  dffacs1 ________________0_(.CLRB (reset), .CLK (clk), .DIN
       (____0____33687), .QN (____________0___18769));
  nor2s1 ___________9_436590(.DIN1 (________20943), .DIN2
       (____0_0__33684), .Q (____0____33699));
  xor2s1 _____________436591(.DIN1 (____99___33666), .DIN2
       (____00___33680), .Q (____0____33698));
  nnd2s1 _____________436592(.DIN1 (____9_9__33596), .DIN2
       (____0____33686), .Q (____0____33697));
  nor2s1 _____9_______436593(.DIN1 (____0____33689), .DIN2
       (_________29840), .Q (____0____33696));
  nor2s1 _________9___436594(.DIN1 (____9____33655), .DIN2
       (____0____33685), .Q (____0____33717));
  xor2s1 _____________436595(.DIN1 (____99___33672), .DIN2
       (_________35050), .Q (____0____33704));
  nor2s1 ___________436596(.DIN1 (____99___33665), .DIN2
       (____00___33681), .Q (____0____33695));
  xor2s1 _____________436597(.DIN1 (____990__33664), .DIN2
       (______0__34988), .Q (____0_0__33702));
  nnd2s1 __________436598(.DIN1 (____0____33694), .DIN2
       (_______________0_____________________18830), .Q
       (____0____33709));
  or2s1 ___________9_436599(.DIN1
       (_______________0_____________________18830), .DIN2
       (____0____33694), .Q (____0____33710));
  nor2s1 ______0______436600(.DIN1 (____00___33679), .DIN2
       (____9____33661), .Q (____0____33713));
  dffacs1 ___________________436601(.CLRB (reset), .CLK (clk), .DIN
       (____009__33683), .Q (_________________18780));
  nnd2s1 _____________436602(.DIN1 (____00___33675), .DIN2
       (____0_9__33692), .Q (____0_0__33693));
  xor2s1 _____________436603(.DIN1 (____9____33658), .DIN2
       (____999__33673), .Q (____0____33691));
  dffacs1 ______________0__9_(.CLRB (reset), .CLK (clk), .DIN
       (____00___33676), .QN (__________0__9_));
  nnd2s1 _____99______436604(.DIN1 (____000__33674), .DIN2
       (____9____33618), .Q (____0____33719));
  nnd2s1 __________9__436605(.DIN1 (____99___33671), .DIN2
       (________25636), .Q (____0____33690));
  nor2s1 _____0_____0_436606(.DIN1 (_________34894), .DIN2
       (____99___33667), .Q (____0____33688));
  nnd2s1 _____________436607(.DIN1 (______9__28982), .DIN2
       (____9_9__33663), .Q (____0____33687));
  dffacs1 ________________0_436608(.CLRB (reset), .CLK (clk), .DIN
       (____9____33662), .Q (____________0___18786));
  nnd2s1 _____0_______436609(.DIN1 (____9___19587), .DIN2
       (____9____33657), .Q (____0____33686));
  and2s1 _____0______436610(.DIN1 (_________31230), .DIN2
       (____9____33660), .Q (____0____33685));
  and2s1 __________0__436611(.DIN1 (_________33817), .DIN2
       (_________34505), .Q (____0_0__33684));
  xnr2s1 ______0____0_(.DIN1 (____99___33670), .DIN2 (________25637),
       .Q (____0____33689));
  nnd2s1 ___________9_436612(.DIN1 (_________33339), .DIN2
       (____9____33656), .Q (____009__33683));
  nnd2s1 _____________436613(.DIN1 (____00___33678), .DIN2
       (____9____33645), .Q (____00___33682));
  and2s1 ____________436614(.DIN1 (____00___33680), .DIN2
       (____9____33651), .Q (____00___33681));
  nor2s1 __________0_436615(.DIN1 (____00___33677), .DIN2
       (____00___33678), .Q (____00___33679));
  xor2s1 _____________436616(.DIN1 (____9____33650), .DIN2
       (____00___33677), .Q (____0____33694));
  nor2s1 _________990_436617(.DIN1 (_________________0___18660), .DIN2
       (____9_0__33654), .Q (____00___33676));
  xor2s1 ____________436618(.DIN1 (______0__31229), .DIN2
       (____9____33659), .Q (____00___33675));
  nnd2s1 ___________9_436619(.DIN1 (____999__33673), .DIN2
       (____9_9__33625), .Q (____000__33674));
  xor2s1 ______9______436620(.DIN1 (____9____33640), .DIN2
       (_____0___30458), .Q (____99___33672));
  or2s1 _____________436621(.DIN1 (________25106), .DIN2
       (____99___33670), .Q (____99___33671));
  nor2s1 _____________436622(.DIN1 (____99___33668), .DIN2
       (________20019), .Q (____99___33669));
  nor2s1 ______9__9___436623(.DIN1 (____9_0__33597), .DIN2
       (____9_9__33653), .Q (____99___33667));
  nor2s1 ______9______436624(.DIN1 (____9____33652), .DIN2
       (____99___33665), .Q (____99___33666));
  xor2s1 ______9____436625(.DIN1 (____9____33636), .DIN2
       (_________30569), .Q (____990__33664));
  nnd2s1 _____________436626(.DIN1 (____9____33649), .DIN2
       (inData[10]), .Q (____9_9__33663));
  nnd2s1 __________436627(.DIN1 (____00___29088), .DIN2
       (____9____33648), .Q (____9____33662));
  and2s1 ___________9_436628(.DIN1 (____9____33646), .DIN2
       (____00___33677), .Q (____9____33661));
  or2s1 _____________436629(.DIN1 (_____0___34429), .DIN2
       (____9____33659), .Q (____9____33660));
  xor2s1 _____________436630(.DIN1 (____9____33624), .DIN2
       (____9_0__33635), .Q (____9____33658));
  dffacs1 ______________0____(.CLRB (reset), .CLK (clk), .DIN
       (____9____33642), .Q (_________34505));
  nor2s1 _____________436631(.DIN1 (_________9_______18805), .DIN2
       (________19283), .Q (____9____33657));
  nnd2s1 _____99______436632(.DIN1 (____9____33647), .DIN2
       (____9____33637), .Q (____9____33656));
  and2s1 __________9__436633(.DIN1 (____9____33659), .DIN2
       (_____0___34429), .Q (____9____33655));
  nnd2s1 ___________0_436634(.DIN1 (____90___33585), .DIN2
       (____9____33639), .Q (____00___33678));
  nnd2s1 _____________436635(.DIN1 (____9_0__33644), .DIN2
       (_________33567), .Q (____00___33680));
  dffacs1 _______________436636(.CLRB (reset), .CLK (clk), .DIN
       (____9____33641), .QN (____________18893));
  xor2s1 _____________436637(.DIN1 (____9____33621), .DIN2
       (____9____33592), .Q (____9_0__33654));
  xor2s1 ____________436638(.DIN1 (____9____33607), .DIN2
       (____9_0__33616), .Q (____9_9__33653));
  hi1s1 _______436639(.DIN (_________9_______18805), .Q
       (____99___33668));
  nnd2s1 ______0___0__436640(.DIN1 (____9_9__33634), .DIN2
       (_________33535), .Q (____99___33670));
  xor2s1 ___________0_436641(.DIN1 (____9____33611), .DIN2
       (____90___33582), .Q (____999__33673));
  hi1s1 _______436642(.DIN (____9____33651), .Q (____9____33652));
  nnd2s1 ______9____9_436643(.DIN1 (____9____33632), .DIN2
       (_________30570), .Q (____9____33650));
  nnd2s1 _____9_______436644(.DIN1 (____9____33628), .DIN2
       (____9____33603), .Q (____9____33649));
  nnd2s1 _____0______436645(.DIN1 (____9____33647), .DIN2
       (____9____33631), .Q (____9____33648));
  nnd2s1 _____0____0_436646(.DIN1 (____9____33630), .DIN2
       (____9_0__33626), .Q (____9____33646));
  nnd2s1 _____09______436647(.DIN1 (____9____33629), .DIN2
       (____9____33638), .Q (____9____33645));
  xnr2s1 _________990_436648(.DIN1 (____9_9__33643), .DIN2
       (____9_0__33606), .Q (____9_0__33644));
  nnd2s1 ______0_____436649(.DIN1 (____9____33622), .DIN2
       (_________34393), .Q (____9____33642));
  nnd2s1 ___________9_436650(.DIN1 (____9____33617), .DIN2
       (________21186), .Q (____9____33641));
  xor2s1 ______0______436651(.DIN1
       (__________________________________9), .DIN2 (____9____33633),
       .Q (____9____33640));
  xnr2s1 _____________436652(.DIN1 (_________35050), .DIN2
       (____0____34576), .Q (____9____33659));
  dffacs1 ___________________436653(.CLRB (reset), .CLK (clk), .DIN
       (____9____33614), .QN (_____0___34428));
  dffacs1 _____________9_____436654(.CLRB (reset), .CLK (clk), .DIN
       (____9____33620), .Q (_________9_______18805));
  hi1s1 _______436655(.DIN (____9____33638), .Q (____9____33639));
  nnd2s1 _____________436656(.DIN1 (____9____33609), .DIN2
       (____9____33590), .Q (____9____33637));
  xor2s1 _________9___436657(.DIN1 (_________34436), .DIN2
       (____0____34578), .Q (____9____33636));
  nnd2s1 ______9______436658(.DIN1 (______9__31473), .DIN2
       (____9____33612), .Q (____9____33651));
  dffacs1 _____________9___0_436659(.CLRB (reset), .CLK (clk), .DIN
       (____9____33619), .QN (_________9___0_));
  dffacs1 ___________________436660(.CLRB (reset), .CLK (clk), .DIN
       (____9____33610), .Q (_________________18783));
  dffacs1 ___________________436661(.CLRB (reset), .CLK (clk), .DIN
       (____9_9__33615), .QN (_________________18793));
  xor2s1 ___________436662(.DIN1 (____9____33623), .DIN2
       (______0__35008), .Q (____9_0__33635));
  nnd2s1 _____________436663(.DIN1 (____9____33633), .DIN2
       (_________33534), .Q (____9_9__33634));
  nnd2s1 _____9____900(.DIN1 (____0____34578), .DIN2 (_____0___30553),
       .Q (____9____33632));
  xor2s1 ______0____9_436664(.DIN1 (_________________18780), .DIN2
       (____9____33608), .Q (____9____33631));
  nnd2s1 _____________436665(.DIN1 (____9____33629), .DIN2
       (____9____33627), .Q (____9____33630));
  nnd2s1 _____________436666(.DIN1 (____9____33602), .DIN2
       (_________33530), .Q (____9____33628));
  nnd2s1 _____________436667(.DIN1 (____9____33627), .DIN2
       (____9_0__33626), .Q (____9____33638));
  nnd2s1 _____________436668(.DIN1 (____9____33624), .DIN2
       (____9____33623), .Q (____9_9__33625));
  xor2s1 __________9__436669(.DIN1 (_________33540), .DIN2
       (____90___33583), .Q (____9____33622));
  xor2s1 ___________0_436670(.DIN1 (____90___33584), .DIN2
       (_____9___33572), .Q (____9____33621));
  nnd2s1 _____________436671(.DIN1 (____9____33594), .DIN2
       (_________35100), .Q (____9____33620));
  nnd2s1 _____________436672(.DIN1 (______0__33318), .DIN2
       (____9____33595), .Q (____9____33619));
  or2s1 ____________436673(.DIN1 (____9____33623), .DIN2
       (____9____33624), .Q (____9____33618));
  nnd2s1 __________0__436674(.DIN1 (_________33817), .DIN2
       (_____9___34418), .Q (____9____33617));
  xnr2s1 _____9_____0_436675(.DIN1 (_________31486), .DIN2
       (____9_9__33605), .Q (____9_0__33616));
  nnd2s1 ___________9_436676(.DIN1 (____9____33598), .DIN2
       (________23855), .Q (____9_9__33615));
  nnd2s1 _____________436677(.DIN1 (____909__33586), .DIN2
       (____9____33613), .Q (____9____33614));
  xor2s1 ____________436678(.DIN1 (____9____33604), .DIN2
       (_________33007), .Q (____9____33612));
  nnd2s1 __________0_436679(.DIN1 (____9____33593), .DIN2
       (_____9___33574), .Q (____9____33611));
  nor2s1 _____________436680(.DIN1 (_________34187), .DIN2
       (____9____33588), .Q (____9____33610));
  nnd2s1 _________990_436681(.DIN1 (____9____33608), .DIN2
       (_________________18780), .Q (____9____33609));
  dffacs1 ___________________436682(.CLRB (reset), .CLK (clk), .DIN
       (____9____33589), .QN (_________________18768));
  xor2s1 ______9_____436683(.DIN1 (______9__33568), .DIN2
       (_________33333), .Q (____9____33607));
  nnd2s1 _____0_____9_436684(.DIN1 (____9_9__33605), .DIN2
       (_________33566), .Q (____9_0__33606));
  nor2s1 _____________436685(.DIN1 (____9____33604), .DIN2
       (______0__31474), .Q (____99___33665));
  nnd2s1 _____________436686(.DIN1 (____90___33581), .DIN2
       (___00____27248), .Q (____9____33633));
  nnd2s1 _________9___436687(.DIN1 (_________33522), .DIN2
       (_____________9___18767), .Q (____9____33603));
  nor2s1 _____________436688(.DIN1 (_____________9___18767), .DIN2
       (_________33511), .Q (____9____33602));
  nnd2s1 ___________436689(.DIN1 (____9____33600), .DIN2
       (____90___33579), .Q (____9____33601));
  nnd2s1 _____________436690(.DIN1 (____9____33599), .DIN2
       (_____________9___18767), .Q (____9____33627));
  or2s1 __________436691(.DIN1 (_____________9___18767), .DIN2
       (____9____33599), .Q (____9_0__33626));
  or2s1 _____00______436692(.DIN1 (____9_0__33597), .DIN2
       (_____90__33569), .Q (____9____33598));
  nnd2s1 _____________436693(.DIN1 (_____9___33577), .DIN2
       (____0_9__33692), .Q (____9_9__33596));
  nnd2s1 _____________436694(.DIN1 (______9__33436), .DIN2
       (_____9___33576), .Q (____9____33595));
  nor2s1 _____________436695(.DIN1 (_____9__20020), .DIN2
       (_____9___33575), .Q (____9____33594));
  nnd2s1 __________9__436696(.DIN1 (____9____33592), .DIN2
       (_____9___33571), .Q (____9____33593));
  dffacs1 ______________0____436697(.CLRB (reset), .CLK (clk), .DIN
       (_____99__33578), .QN (_____9___34418));
  xor2s1 _____9_____0_436698(.DIN1 (___0__0__27599), .DIN2
       (____90___33580), .Q (____9____33623));
  nnd2s1 _____________436699(.DIN1 (_____0___33226), .DIN2
       (_________________18781), .Q (____9____33591));
  nnd2s1 _____________436700(.DIN1 (_________33527), .DIN2
       (_________________18781), .Q (____9____33590));
  nnd2s1 ____________436701(.DIN1 (_________33544), .DIN2
       (_________33565), .Q (____9____33589));
  xor2s1 __________0__436702(.DIN1 (_________33557), .DIN2
       (____9_0__33587), .Q (____9____33588));
  nor2s1 _____0_____0_436703(.DIN1 (________23595), .DIN2
       (_____9___33570), .Q (____909__33586));
  nor2s1 ___________9_436704(.DIN1 (_________33509), .DIN2
       (_________________18781), .Q (____9____33608));
  hi1s1 _______436705(.DIN (____90___33585), .Q (____9____33629));
  xor2s1 _____9______436706(.DIN1 (_____9___33573), .DIN2
       (_________35094), .Q (____90___33584));
  xor2s1 _____90___0_9(.DIN1 (_________33551), .DIN2 (____90___33582),
       .Q (____90___33583));
  nnd2s1 _____9_______436707(.DIN1 (____90___33580), .DIN2
       (___0_____27449), .Q (____90___33581));
  nnd2s1 ______0__990_436708(.DIN1 (_________33562), .DIN2
       (_________33441), .Q (____9_9__33605));
  hi1s1 _______436709(.DIN (_________________18781), .Q
       (____90___33579));
  nor2s1 ___________9_436710(.DIN1 (_________33556), .DIN2
       (_________33558), .Q (____90___33585));
  xor2s1 _____________436711(.DIN1 (_________30306), .DIN2
       (_________33547), .Q (____9____33604));
  dffacs1 _________________9_436712(.CLRB (reset), .CLK (clk), .DIN
       (______9__33560), .Q (_____________9___18767));
  nnd2s1 _____________436713(.DIN1 (_________33548), .DIN2
       (_________34365), .Q (_____99__33578));
  xor2s1 _____________436714(.DIN1 (_________33538), .DIN2
       (_________32606), .Q (_____9___33577));
  and2s1 _____9___9___436715(.DIN1 (______0__33553), .DIN2
       (inData[22]), .Q (_____9___33576));
  and2s1 _____0_______436716(.DIN1 (_________33554), .DIN2
       (____0_9__33692), .Q (_____9___33575));
  or2s1 _____0_____436717(.DIN1 (_____9___33573), .DIN2
       (_____9___33572), .Q (_____9___33574));
  nnd2s1 _____0_______436718(.DIN1 (_____9___33572), .DIN2
       (_____9___33573), .Q (_____9___33571));
  nor2s1 __________436719(.DIN1 (____9_0__33597), .DIN2
       (______0__33543), .Q (_____9___33570));
  xor2s1 ___________9_436720(.DIN1 (______9__33472), .DIN2
       (______0__33561), .Q (_____90__33569));
  and2s1 _____________436721(.DIN1 (_________33567), .DIN2
       (_________33566), .Q (______9__33568));
  nnd2s1 _____________436722(.DIN1 (______9__33542), .DIN2
       (inData[20]), .Q (_________33565));
  nor2s1 _____________436723(.DIN1 (_________33550), .DIN2
       (______9__33552), .Q (____9____33592));
  dffacs1 ___________________436724(.CLRB (reset), .CLK (clk), .DIN
       (_________33545), .Q (_________________18782));
  dffacs1 ___________________436725(.CLRB (reset), .CLK (clk), .DIN
       (_________33546), .Q (_________________18781));
  nnd2s1 ___________0_436726(.DIN1 (______0__33561), .DIN2
       (_________33451), .Q (_________33562));
  nnd2s1 ______9______436727(.DIN1 (_________33537), .DIN2
       (_________33332), .Q (____90___33580));
  nnd2s1 ______9______436728(.DIN1 (______9__33532), .DIN2
       (_________33531), .Q (______9__33560));
  nor2s1 _____00____0_(.DIN1 (____9_0__33587), .DIN2 (_________33555),
       .Q (_________33558));
  or2s1 _____0_____9_436729(.DIN1 (_________33556), .DIN2
       (_________33555), .Q (_________33557));
  xor2s1 _____________436730(.DIN1 (______0__33533), .DIN2
       (____9____30879), .Q (_________33554));
  xor2s1 ______9_____436731(.DIN1
       (__________________________________9), .DIN2 (_________9__9_),
       .Q (______0__33553));
  nor2s1 __________0_436732(.DIN1 (_________33539), .DIN2
       (_________33549), .Q (______9__33552));
  nor2s1 _____________436733(.DIN1 (_________33550), .DIN2
       (_________33549), .Q (_________33551));
  xor2s1 _____0___990_(.DIN1 (____99___34525), .DIN2 (_____9___33482),
       .Q (_________33548));
  xor2s1 ____________436734(.DIN1 (_________33361), .DIN2
       (_________33536), .Q (_____9___33573));
  dffacs1 _____________9_____436735(.CLRB (reset), .CLK (clk), .DIN
       (_________33526), .Q (_________9_____));
  xnr2s1 ___________9_436736(.DIN1 (_____________0___18779), .DIN2
       (____0_0__34580), .Q (_________33547));
  nnd2s1 _____________436737(.DIN1 (_________33470), .DIN2
       (______0__33524), .Q (_________33546));
  nnd2s1 _____________436738(.DIN1 (_________33520), .DIN2
       (____0___21077), .Q (_________33545));
  nnd2s1 ______9______436739(.DIN1 (_________33528), .DIN2
       (_________33279), .Q (_________33544));
  xor2s1 _________9___436740(.DIN1 (_________33516), .DIN2
       (_________35104), .Q (______0__33543));
  nnd2s1 _____0_______436741(.DIN1 (_________33525), .DIN2
       (_________33512), .Q (______9__33542));
  xor2s1 ___________436742(.DIN1 (_________33507), .DIN2
       (_________33541), .Q (_________33567));
  dffacs1 ___________________436743(.CLRB (reset), .CLK (clk), .DIN
       (______9__33523), .Q
       (_______________0_____________________18831));
  xor2s1 ______0______436744(.DIN1 (_________33539), .DIN2
       (____009__31815), .Q (_________33540));
  xor2s1 __________436745(.DIN1 (_________33504), .DIN2
       (____0____30918), .Q (_________33538));
  nnd2s1 ______0____9_436746(.DIN1 (_________33536), .DIN2
       (______0__33327), .Q (_________33537));
  or2s1 ______0______436747(.DIN1
       (__________________________________9), .DIN2 (_________34409),
       .Q (_________33535));
  nnd2s1 ______9______436748(.DIN1 (_________34409), .DIN2
       (__________________________________9), .Q (_________33534));
  nor2s1 _____________436749(.DIN1 (____9____30873), .DIN2
       (______0__33533), .Q (_________33563));
  nor2s1 _____0_______436750(.DIN1 (_________33508), .DIN2
       (_________33371), .Q (______9__33532));
  nnd2s1 __________9__436751(.DIN1 (_________33510), .DIN2
       (_________33530), .Q (_________33531));
  nnd2s1 ___________0_436752(.DIN1 (______9__33514), .DIN2
       (_________33515), .Q (______0__33561));
  nor2s1 _____________436753(.DIN1 (_________30336), .DIN2
       (____0_0__34580), .Q (_________33559));
  and2s1 ______0______436754(.DIN1 (_________33529), .DIN2
       (_________18859), .Q (_________33556));
  nor2s1 ____________436755(.DIN1 (_________18859), .DIN2
       (_________33529), .Q (_________33555));
  xor2s1 _____9____0__(.DIN1 (_____0___33490), .DIN2 (________22792),
       .Q (_________33528));
  nnd2s1 ___________0_436756(.DIN1
       (_______________0_____________________18834), .DIN2
       (_________________18780), .Q (_________33527));
  nnd2s1 ___________9_436757(.DIN1 (_________33503), .DIN2
       (________19347), .Q (_________33526));
  or2s1 _____________436758(.DIN1 (____________0___18769), .DIN2
       (_________33521), .Q (_________33525));
  xor2s1 ____________436759(.DIN1 (_____0___33493), .DIN2
       (_________31983), .Q (_________33549));
  nnd2s1 __________0_436760(.DIN1 (____9____33647), .DIN2
       (_______________0_____________________18834), .Q
       (______0__33524));
  nnd2s1 _____________436761(.DIN1 (_________33502), .DIN2
       (____90___32662), .Q (______9__33523));
  nnd2s1 _________990_436762(.DIN1 (_________33521), .DIN2
       (___0____19820), .Q (_________33522));
  nnd2s1 ______0_____436763(.DIN1 (_________33501), .DIN2
       (_________32639), .Q (_________33520));
  or2s1 ___________9_436764(.DIN1 (_________33518), .DIN2
       (_________33517), .Q (_________33519));
  and2s1 _____9_______436765(.DIN1 (_________33513), .DIN2
       (_________33515), .Q (_________33516));
  nnd2s1 ______9______436766(.DIN1 (_________35104), .DIN2
       (_________33513), .Q (______9__33514));
  nor2s1 _________9___436767(.DIN1 (______9__30783), .DIN2
       (______0__33497), .Q (______0__33533));
  nnd2s1 ______0______436768(.DIN1 (_____9___33481), .DIN2
       (_____0___33494), .Q (_________33536));
  dffacs1 _____________9_____436769(.CLRB (reset), .CLK (clk), .DIN
       (_________33498), .QN (__________________________________9));
  dffacs1 ___________________436770(.CLRB (reset), .CLK (clk), .DIN
       (_____0___33495), .QN (_____0___34429));
  or2s1 ______9____436771(.DIN1 (___0__0__27481), .DIN2
       (_________33511), .Q (_________33512));
  hi1s1 ______436772(.DIN (_________33521), .Q (_________33510));
  hi1s1 _______436773(.DIN
       (_______________0_____________________18834), .Q
       (_________33509));
  nor2s1 _____________436774(.DIN1 (_________33530), .DIN2
       (_________33511), .Q (_________33508));
  nor2s1 _____9____436775(.DIN1 (______9__33505), .DIN2
       (______0__33506), .Q (_________33507));
  nor2s1 ___________9_436776(.DIN1 (____0____30960), .DIN2
       (_____0___33492), .Q (_________33529));
  nnd2s1 _____9_______436777(.DIN1 (______0__33506), .DIN2
       (______9__33505), .Q (_________33566));
  xor2s1 _____________436778(.DIN1 (_____09__33496), .DIN2
       (______0__18849), .Q (_________33504));
  nnd2s1 ______0______436779(.DIN1 (_____00__33488), .DIN2
       (____0_9__33692), .Q (_________33503));
  nor2s1 __________9__436780(.DIN1 (____9___21541), .DIN2
       (_____9___33486), .Q (_________33502));
  nor2s1 ___________0_436781(.DIN1 (_________33499), .DIN2
       (_____9___33483), .Q (_________33539));
  xor2s1 _____________436782(.DIN1 (_____0___33491), .DIN2
       (____0____30968), .Q (_________33501));
  nor2s1 _____________436783(.DIN1 (_________33500), .DIN2
       (_____0___31191), .Q (_________33517));
  nnd2s1 ____________436784(.DIN1 (_____0___33489), .DIN2
       (_________33500), .Q (_________33521));
  dffacs1 ___________________436785(.CLRB (reset), .CLK (clk), .DIN
       (_____99__33487), .QN
       (_______________0_____________________18834));
  nnd2s1 ______0___0__436786(.DIN1 (_________33374), .DIN2
       (_____90__33479), .Q (_________33498));
  and2s1 ___________0_436787(.DIN1 (_____09__33496), .DIN2
       (______0__30784), .Q (______0__33497));
  nnd2s1 ___________9_436788(.DIN1 (_____9___33484), .DIN2
       (____9____33613), .Q (_____0___33495));
  nnd2s1 _____90______436789(.DIN1 (_____9___33485), .DIN2
       (___0_____27896), .Q (_____0___33494));
  nor2s1 _____9______436790(.DIN1 (_____9___33480), .DIN2
       (_________29541), .Q (_____0___33493));
  nor2s1 ______9___0_436791(.DIN1 (____0____30959), .DIN2
       (_____0___33491), .Q (_____0___33492));
  xor2s1 _____________436792(.DIN1 (_________33469), .DIN2
       (_________________18752), .Q (_____0___33490));
  xor2s1 ____________436793(.DIN1 (_________33471), .DIN2
       (_________33206), .Q (______9__33505));
  xor2s1 ______9____9_436794(.DIN1 (_________33475), .DIN2
       (_________33564), .Q (_________33513));
  nor2s1 _____________436795(.DIN1 (_________34438), .DIN2
       (____090__33759), .Q (_________33518));
  nnd2s1 ______0______436796(.DIN1 (_____0___33489), .DIN2
       (_________34438), .Q (_________33511));
  xor2s1 _____9_______436797(.DIN1 (_________33455), .DIN2
       (______9__18848), .Q (_____00__33488));
  nor2s1 _____9___9___436798(.DIN1 (____99___34527), .DIN2
       (_________29539), .Q (_________33550));
  xor2s1 _____________436799(.DIN1 (_________33465), .DIN2
       (_________33894), .Q (_________33499));
  dffacs1 _____________9_____436800(.CLRB (reset), .CLK (clk), .DIN
       (_________33477), .Q (_________18852));
  nnd2s1 ___________436801(.DIN1 (_________33468), .DIN2
       (_________33350), .Q (_____99__33487));
  nor2s1 _____________436802(.DIN1 (_________31648), .DIN2
       (_________33467), .Q (_____9___33486));
  hi1s1 _______436803(.DIN (_________34438), .Q (_________33500));
  nnd2s1 _____0_____9_436804(.DIN1 (_________33461), .DIN2
       (_____9___33214), .Q (_____9___33485));
  nor2s1 _____99______436805(.DIN1 (_____0__23666), .DIN2
       (_________33452), .Q (_____9___33484));
  nor2s1 _____9_______436806(.DIN1 (_________33476), .DIN2
       (_____9___33482), .Q (_____9___33483));
  nnd2s1 _____0_______436807(.DIN1 (______0__33464), .DIN2
       (______0__34988), .Q (_____9___33481));
  hi1s1 ______436808(.DIN (____99___34527), .Q (_____9___33480));
  dffacs1 ___________________436809(.CLRB (reset), .CLK (clk), .DIN
       (_________33466), .QN (_____09__34430));
  nnd2s1 _____________436810(.DIN1 (______0__33373), .DIN2
       (_________33462), .Q (_____90__33479));
  nor2s1 _____00______436811(.DIN1 (_____9___30818), .DIN2
       (_________33458), .Q (_____0___33491));
  nnd2s1 _____________436812(.DIN1 (_________33456), .DIN2
       (______9__33453), .Q (_____09__33496));
  dffacs1 _________________0_436813(.CLRB (reset), .CLK (clk), .DIN
       (_________33449), .QN (_________34438));
  nnd2s1 ____________436814(.DIN1 (_________33447), .DIN2
       (________21271), .Q (_________33477));
  nor2s1 __________0__436815(.DIN1 (______0__33473), .DIN2
       (_________33474), .Q (_________33475));
  nnd2s1 ___________9_436816(.DIN1 (_________33474), .DIN2
       (______0__33473), .Q (_________33515));
  xor2s1 ____________436817(.DIN1 (_________33450), .DIN2
       (_________33440), .Q (______9__33472));
  xor2s1 ______9___0_436818(.DIN1 (_________33448), .DIN2
       (_____________9___18778), .Q (_________33471));
  nnd2s1 _____________436819(.DIN1 (_________33445), .DIN2
       (_________33442), .Q (_________33470));
  xor2s1 _____9___990_(.DIN1 (_________33433), .DIN2 (_________35111),
       .Q (_________33469));
  nor2s1 _____9______436820(.DIN1 (___9_9__22490), .DIN2
       (_________33443), .Q (_________33468));
  xor2s1 _____0_____9_436821(.DIN1 (_________33457), .DIN2
       (____9____30836), .Q (_________33467));
  nnd2s1 _____________436822(.DIN1 (_________33439), .DIN2
       (_________33379), .Q (_________33466));
  nnd2s1 _____________436823(.DIN1 (_________33459), .DIN2
       (_________33460), .Q (_________33465));
  nor2s1 _____________436824(.DIN1 (_____0___33223), .DIN2
       (______9__33463), .Q (______0__33464));
  nnd2s1 _________9___436825(.DIN1 (______0__33437), .DIN2
       (inData[28]), .Q (_________33462));
  nnd2s1 _____________436826(.DIN1 (______9__33463), .DIN2
       (_____9___33213), .Q (_________33461));
  nor2s1 ___________436827(.DIN1 (_________33460), .DIN2
       (_________33459), .Q (_________33476));
  dffacs2 _____________________0_(.CLRB (reset), .CLK (clk), .DIN
       (_________33438), .Q (_________________0___18618));
  nor2s1 _____________436828(.DIN1 (_____99__30819), .DIN2
       (_________33457), .Q (_________33458));
  nnd2s1 __________436829(.DIN1 (______0__33454), .DIN2
       (______9__18848), .Q (_________33456));
  and2s1 ___________9_436830(.DIN1 (______0__33454), .DIN2
       (______9__33453), .Q (_________33455));
  nor2s1 ______9______436831(.DIN1 (____9_0__33597), .DIN2
       (_________33435), .Q (_________33452));
  nnd2s1 _____________436832(.DIN1 (______9__31292), .DIN2
       (_________33450), .Q (_________33451));
  nnd2s1 _____0_______436833(.DIN1 (_________33434), .DIN2
       (_________34295), .Q (_________33449));
  nnd2s1 _____________436834(.DIN1 (_________33448), .DIN2
       (_________33207), .Q (_________33478));
  nnd2s1 __________9__436835(.DIN1 (____0____34582), .DIN2
       (____0_9__33692), .Q (_________33447));
  xor2s1 _____0_______436836(.DIN1 (______0__33419), .DIN2
       (_________33444), .Q (_________33445));
  and2s1 ______9_____436837(.DIN1 (_________33431), .DIN2
       (_________33442), .Q (_________33443));
  nnd2s1 __________0__436838(.DIN1 (_________33440), .DIN2
       (_________33432), .Q (_________33441));
  xor2s1 _____9_____0_436839(.DIN1 (_________33421), .DIN2
       (_________32442), .Q (______0__33473));
  and2s1 ___________9_436840(.DIN1 (_________33426), .DIN2
       (_________33430), .Q (_________33439));
  nnd2s1 _____________436841(.DIN1 (__9_____26378), .DIN2
       (______0__33429), .Q (_________33438));
  and2s1 ____________436842(.DIN1 (______9__33436), .DIN2
       (_________33424), .Q (______0__33437));
  xor2s1 ______0___0_436843(.DIN1 (_____9___33398), .DIN2
       (____0____34584), .Q (_________33435));
  xor2s1 _____________436844(.DIN1 (_________33416), .DIN2
       (_______________18874), .Q (_________33460));
  nnd2s1 _________990_436845(.DIN1 (_________33425), .DIN2
       (_________33414), .Q (______9__33463));
  nor2s1 ____________436846(.DIN1 (____9___20032), .DIN2
       (_________33420), .Q (_________33434));
  xor2s1 ___________9_436847(.DIN1 (_________32048), .DIN2
       (_________33412), .Q (_________33433));
  hi1s1 _____0_436848(.DIN (_________33432), .Q (_________33450));
  nnd2s1 _____________436849(.DIN1 (______9__33428), .DIN2
       (_________30604), .Q (______0__33454));
  nnd2s1 _____99______436850(.DIN1 (_________33423), .DIN2
       (_________30195), .Q (_________33448));
  nor2s1 _____________436851(.DIN1 (_________33249), .DIN2
       (______9__33418), .Q (_________33457));
  nnd2s1 _____________436852(.DIN1 (_________33427), .DIN2
       (_________30611), .Q (______9__33453));
  xor2s1 ___________436853(.DIN1 (_________33251), .DIN2
       (_________33417), .Q (_________33431));
  xor2s1 ______0______436854(.DIN1 (_________30196), .DIN2
       (_________33422), .Q (_________33432));
  nnd2s1 ______9___436855(.DIN1 (____0____34584), .DIN2
       (_____9___33393), .Q (______0__33446));
  nnd2s1 ___________9_436856(.DIN1 (______0__33336), .DIN2
       (_____09__33409), .Q (_________33430));
  or2s1 _____________436857(.DIN1 (_________33411), .DIN2
       (___0_9__22581), .Q (______0__33429));
  hi1s1 _______436858(.DIN (_________33427), .Q (______9__33428));
  nor2s1 _____________436859(.DIN1 (_____0___33408), .DIN2
       (_____9___33308), .Q (_________33426));
  nnd2s1 _____________436860(.DIN1 (_________33415), .DIN2
       (_____0___33407), .Q (_________33425));
  dffacs1 ___________________436861(.CLRB (reset), .CLK (clk), .DIN
       (_____0___33406), .QN (_________________18792));
  xor2s1 _____________436862(.DIN1 (_________33413), .DIN2
       (______9__33326), .Q (_________33424));
  or2s1 ______0___9__436863(.DIN1 (_________30163), .DIN2
       (_________33422), .Q (_________33423));
  xor2s1 ___________0_436864(.DIN1 (_____99__33400), .DIN2
       (_________33388), .Q (_________33421));
  nor2s1 ______0______436865(.DIN1 (_________33370), .DIN2
       (_____0___33405), .Q (_________33420));
  xor2s1 _____________436866(.DIN1 (_____9___33397), .DIN2
       (_________________18766), .Q (______0__33419));
  nor2s1 ____________436867(.DIN1 (_________33250), .DIN2
       (_________33417), .Q (______9__33418));
  xor2s1 _____9____0__436868(.DIN1 (_________33415), .DIN2
       (_________9______18803), .Q (_________33416));
  nnd2s1 ______0____0_436869(.DIN1 (_____0___33404), .DIN2
       (______0__30437), .Q (_________33427));
  nnd2s1 _____0_____9_436870(.DIN1 (_______________18874), .DIN2
       (_________33413), .Q (_________33414));
  nor2s1 _____________436871(.DIN1 (_________32130), .DIN2
       (_____0___33402), .Q (_________33412));
  nnd2s1 _____9____0_436872(.DIN1 (___9____26209), .DIN2
       (_________9______18803), .Q (_________33411));
  xor2s1 _____90______436873(.DIN1 (_____0___33403), .DIN2
       (___0____21656), .Q (_________33410));
  nor2s1 _____9___990_436874(.DIN1 (______9__18848), .DIN2
       (________23232), .Q (_____09__33409));
  and2s1 _____9______436875(.DIN1 (_________33241), .DIN2
       (______9__18848), .Q (_____0___33408));
  dffacs1 ___________________436876(.CLRB (reset), .CLK (clk), .DIN
       (_____9___33395), .Q (______0__18849));
  nnd2s1 _____0_____9_436877(.DIN1 (____0____30075), .DIN2
       (_________9______18803), .Q (_____0___33407));
  nnd2s1 _____0_______436878(.DIN1 (_____9___33394), .DIN2
       (____0___24156), .Q (_____0___33406));
  xor2s1 _____________436879(.DIN1 (______0__32135), .DIN2
       (_____00__33401), .Q (_____0___33405));
  nor2s1 _____________436880(.DIN1 (_____9___33399), .DIN2
       (_________33389), .Q (_________33422));
  nor2s1 _________9___436881(.DIN1 (_________30715), .DIN2
       (_________33387), .Q (_________33417));
  or2s1 _____9_______436882(.DIN1 (______9__30436), .DIN2
       (_____0___33403), .Q (_____0___33404));
  hi1s1 _______436883(.DIN (_________9______18803), .Q
       (_________33413));
  nor2s1 _____________436884(.DIN1 (_________32127), .DIN2
       (_____00__33401), .Q (_____0___33402));
  nor2s1 __________436885(.DIN1 (_____9___33399), .DIN2
       (______9__33382), .Q (_____99__33400));
  xor2s1 ___________9_436886(.DIN1 (_____90__33391), .DIN2
       (_____9___33392), .Q (_____9___33398));
  xor2s1 _____________436887(.DIN1 (_________33386), .DIN2
       (_____9___33396), .Q (_____9___33397));
  nnd2s1 _____________436888(.DIN1 (_________33377), .DIN2
       (____9____33613), .Q (_____9___33395));
  or2s1 _____________436889(.DIN1 (____9_0__33597), .DIN2
       (_________33376), .Q (_____9___33394));
  dffacs1 _____________9____436890(.CLRB (reset), .CLK (clk), .DIN
       (_________33378), .Q (_________9______18803));
  dffacs1 ___________________436891(.CLRB (reset), .CLK (clk), .DIN
       (_________33380), .QN (______9__18848));
  or2s1 _____________436892(.DIN1 (_____9___33392), .DIN2
       (_____90__33391), .Q (_____9___33393));
  and2s1 __________9__436893(.DIN1 (_____90__33391), .DIN2
       (_____9___33392), .Q (______9__33390));
  and2s1 ___________0_436894(.DIN1 (_________33381), .DIN2
       (_________33388), .Q (_________33389));
  and2s1 _____________436895(.DIN1 (_________33386), .DIN2
       (_____9___30721), .Q (_________33387));
  xor2s1 ____________436896(.DIN1 (_________33366), .DIN2
       (_________33384), .Q (_____0___33403));
  dffacs1 ___________________436897(.CLRB (reset), .CLK (clk), .DIN
       (_________33369), .Q (_________18859));
  hi1s1 _______436898(.DIN (_________33381), .Q (______9__33382));
  xor2s1 ___________0_436899(.DIN1 (_________33367), .DIN2
       (_________________0___18607), .Q (_____00__33401));
  nnd2s1 ___________9_436900(.DIN1 (_________33365), .DIN2
       (_________33379), .Q (_________33380));
  nnd2s1 _____________436901(.DIN1 (_________33139), .DIN2
       (_________33368), .Q (_________33378));
  nor2s1 ____________436902(.DIN1 (________23639), .DIN2
       (_________33364), .Q (_________33377));
  dffacs1 ___________________436903(.CLRB (reset), .CLK (clk), .DIN
       (______0__33363), .QN (_________34439));
  xor2s1 __________0_436904(.DIN1 (_____90__33302), .DIN2
       (______9__33372), .Q (_________33376));
  nnd2s1 _____________436905(.DIN1 (_________33375), .DIN2
       (_________________18776), .Q (_________33381));
  nor2s1 _________990_436906(.DIN1 (_________________18776), .DIN2
       (_________33375), .Q (_____9___33399));
  xnr2s1 ____________436907(.DIN1 (____0____31820), .DIN2
       (____0____34586), .Q (_________33386));
  xor2s1 ___________9_436908(.DIN1 (_________33359), .DIN2
       (_________28828), .Q (_____9___33392));
  or2s1 _____________436909(.DIN1 (______0__33373), .DIN2
       (_________33362), .Q (_________33374));
  or2s1 ______9______436910(.DIN1 (_________33290), .DIN2
       (______9__33372), .Q (______0__33383));
  nor2s1 _____________436911(.DIN1 (_________33370), .DIN2
       (_________33358), .Q (_________33371));
  nnd2s1 ______9__9___436912(.DIN1 (_________33360), .DIN2
       (_________34295), .Q (_________33369));
  nnd2s1 _____________436913(.DIN1 (_________33348), .DIN2
       (inData[16]), .Q (_________33368));
  nnd2s1 _____0_____436914(.DIN1 (______0__33354), .DIN2
       (_________32117), .Q (_________33367));
  dffacs1 ___________________436915(.CLRB (reset), .CLK (clk), .DIN
       (_________33351), .Q
       (_______________0_____________________18830));
  dffacs1 ___________________436916(.CLRB (reset), .CLK (clk), .DIN
       (_________33357), .QN (______0__34431));
  nor2s1 _____________436917(.DIN1 (_________30380), .DIN2
       (_________33356), .Q (_________33366));
  and2s1 ______0___900(.DIN1 (_________33352), .DIN2 (___9____23357),
       .Q (_________33365));
  nor2s1 ______9____9_436918(.DIN1 (____9_0__33597), .DIN2
       (_________33349), .Q (_________33364));
  nnd2s1 _____________436919(.DIN1 (_________33347), .DIN2
       (_________34295), .Q (______0__33363));
  xor2s1 _____________436920(.DIN1 (_________33346), .DIN2
       (_________33385), .Q (_________33375));
  xor2s1 _____________436921(.DIN1 (_________30392), .DIN2
       (_________33355), .Q (_________33362));
  xor2s1 ______0___9__436922(.DIN1 (_______________18875), .DIN2
       (_________33334), .Q (_________33361));
  nor2s1 _____9_____0_436923(.DIN1 (_________33280), .DIN2
       (_________33345), .Q (_________33360));
  xor2s1 _____________436924(.DIN1 (_________33342), .DIN2
       (_________33330), .Q (_________33359));
  xor2s1 _____9_______436925(.DIN1 (_________32119), .DIN2
       (______9__33353), .Q (_________33358));
  nor2s1 ____________436926(.DIN1 (_________33282), .DIN2
       (______9__33344), .Q (______9__33372));
  nnd2s1 __________0__436927(.DIN1 (_________33338), .DIN2
       (_________33379), .Q (_________33357));
  nor2s1 ___________0_436928(.DIN1 (______0__30373), .DIN2
       (_________33355), .Q (_________33356));
  nnd2s1 _____09____9_436929(.DIN1 (______9__33353), .DIN2
       (_________32118), .Q (______0__33354));
  nor2s1 _____________436930(.DIN1 (____9___23882), .DIN2
       (_________33337), .Q (_________33352));
  nnd2s1 _____90_____0(.DIN1 (_________33340), .DIN2 (_________33350),
       .Q (_________33351));
  xor2s1 ______0___0_436931(.DIN1 (______9__33283), .DIN2
       (_________33343), .Q (_________33349));
  and2s1 ______9______436932(.DIN1 (______9__33436), .DIN2
       (______9__33335), .Q (_________33348));
  nor2s1 _____9___990_436933(.DIN1 (________20582), .DIN2
       (_________33341), .Q (_________33347));
  nor2s1 _____00_____436934(.DIN1 (____99___34526), .DIN2
       (_________33331), .Q (_________33346));
  nor2s1 _____0_____9_436935(.DIN1 (_________33370), .DIN2
       (_________33328), .Q (_________33345));
  nor2s1 _____________436936(.DIN1 (_________33281), .DIN2
       (_________33343), .Q (______9__33344));
  nor2s1 _____________436937(.DIN1 (____99___34526), .DIN2
       (_________33329), .Q (_________33342));
  nor2s1 _____0___9___436938(.DIN1 (_________33370), .DIN2
       (_________33323), .Q (_________33341));
  and2s1 _____0_______436939(.DIN1 (_________33322), .DIN2
       (_________33237), .Q (_________33340));
  nnd2s1 ___________436940(.DIN1 (_____09__33317), .DIN2
       (_________33442), .Q (_________33339));
  nor2s1 _____________436941(.DIN1 (_____0___31998), .DIN2
       (_________33321), .Q (______9__33353));
  nor2s1 __________436942(.DIN1 (____99__23617), .DIN2
       (_____0___33316), .Q (_________33338));
  nor2s1 ______0____9_436943(.DIN1 (______0__33336), .DIN2
       (_________33319), .Q (_________33337));
  xnr2s1 _____________436944(.DIN1 (_________9__9_), .DIN2
       (_________9___0_), .Q (______9__33335));
  xnr2s1 _____________436945(.DIN1 (_________9__9_), .DIN2
       (_________33333), .Q (_________33334));
  nnd2s1 _____________436946(.DIN1 (_____0___33315), .DIN2
       (_______________18875), .Q (_________33332));
  xnr2s1 _____________436947(.DIN1 (____000__32751), .DIN2
       (_____0___33314), .Q (_________33355));
  nor2s1 __________9__436948(.DIN1 (_________33330), .DIN2
       (_________33329), .Q (_________33331));
  xor2s1 ___________0_436949(.DIN1 (_________32009), .DIN2
       (_________33320), .Q (_________33328));
  nnd2s1 _____________436950(.DIN1 (____09___30086), .DIN2
       (_________9__9_), .Q (______0__33327));
  nnd2s1 ______0_____436951(.DIN1 (_________9__9_), .DIN2
       (___00____27191), .Q (______9__33326));
  nor2s1 _______436952(.DIN1 (_________33176), .DIN2 (_____0___33313),
       .Q (_________33343));
  xor2s1 _______436953(.DIN1 (_____9___33304), .DIN2 (______9__33856),
       .Q (_________33323));
  nnd2s1 _______436954(.DIN1 (_____99__33309), .DIN2 (_________33442),
       .Q (_________33322));
  nor2s1 ______436955(.DIN1 (_____9___31995), .DIN2 (_________33320),
       .Q (_________33321));
  xor2s1 _______436956(.DIN1 (______9__33192), .DIN2 (_____0___33312),
       .Q (_________33319));
  or2s1 _______436957(.DIN1 (______0__33373), .DIN2 (_____9___33307),
       .Q (______0__33318));
  xor2s1 _______436958(.DIN1 (_________30526), .DIN2 (____0_0__34588),
       .Q (_____09__33317));
  nor2s1 _______436959(.DIN1 (______0__33336), .DIN2 (_____0___33311),
       .Q (_____0___33316));
  hi1s1 ______436960(.DIN (_________9__9_), .Q (_____0___33315));
  nor2s1 _______436961(.DIN1 (_________________18775), .DIN2
       (_____00__33310), .Q (_________33329));
  or2s1 _______436962(.DIN1 (_____0___30459), .DIN2 (____0_0__34588),
       .Q (_________33324));
  nor2s1 _____9_436963(.DIN1 (_________30235), .DIN2 (_____9___33306),
       .Q (_____0___33314));
  nor2s1 _____9_436964(.DIN1 (_________33185), .DIN2 (_____0___33312),
       .Q (_____0___33313));
  dffacs1 _____________9__9_(.CLRB (reset), .CLK (clk), .DIN
       (_____9___33305), .Q (_________9__9_));
  xor2s1 _____99(.DIN1 (_________33296), .DIN2 (_________33144), .Q
       (_____0___33311));
  xor2s1 _______436965(.DIN1 (_________33294), .DIN2 (_________28737),
       .Q (_____99__33309));
  nor2s1 _____9_436966(.DIN1 (______0__33336), .DIN2 (_____9___33303),
       .Q (_____9___33308));
  xor2s1 _____9_436967(.DIN1 (______9__30308), .DIN2 (____0____34590),
       .Q (_____9___33307));
  nor2s1 _______436968(.DIN1 (_________32911), .DIN2 (_________33300),
       .Q (_________33320));
  dffacs1 ___________________436969(.CLRB (reset), .CLK (clk), .DIN
       (______9__33301), .QN (______9__34440));
  nor2s1 _____0_436970(.DIN1 (______9__30236), .DIN2 (____0____34590),
       .Q (_____9___33306));
  nnd2s1 _____0_436971(.DIN1 (_________33295), .DIN2 (___9____19741),
       .Q (_____9___33305));
  nor2s1 _______436972(.DIN1 (_________33199), .DIN2 (_________33298),
       .Q (_____0___33312));
  xor2s1 _______436973(.DIN1 (_________32913), .DIN2 (_________33299),
       .Q (_____9___33304));
  xor2s1 ______436974(.DIN1 (_________33288), .DIN2
       (_________________0___18618), .Q (_____00__33310));
  xor2s1 ______436975(.DIN1 (_____9___33218), .DIN2 (_________33297),
       .Q (_____9___33303));
  xor2s1 ______436976(.DIN1 (______0__33292), .DIN2 (______9__33291),
       .Q (_____90__33302));
  nnd2s1 _______436977(.DIN1 (_________33287), .DIN2 (_____0___31454),
       .Q (______9__33301));
  nor2s1 _______436978(.DIN1 (_________32912), .DIN2 (_________33299),
       .Q (_________33300));
  dffacs1 ___________________436979(.CLRB (reset), .CLK (clk), .DIN
       (_________33286), .Q (_________34436));
  dffacs1 __________________(.CLRB (reset), .CLK (clk), .DIN
       (_________33289), .Q (_________34432));
  nor2s1 _______436980(.DIN1 (_________33198), .DIN2 (_________33297),
       .Q (_________33298));
  xor2s1 _______436981(.DIN1 (_________33260), .DIN2 (_________33274),
       .Q (_________33296));
  or2s1 _______436982(.DIN1 (______0__33373), .DIN2 (______0__33284),
       .Q (_________33295));
  xor2s1 _______436983(.DIN1 (_________33270), .DIN2
       (_________________18765), .Q (_________33294));
  and2s1 _______436984(.DIN1 (______0__33292), .DIN2 (______9__33291),
       .Q (_________33293));
  nor2s1 _______436985(.DIN1 (______9__33291), .DIN2 (______0__33292),
       .Q (_________33290));
  dffacs1 __________________436986(.CLRB (reset), .CLK (clk), .DIN
       (_________33285), .QN (________________18788));
  nnd2s1 _______436987(.DIN1 (_________33272), .DIN2 (_________33379),
       .Q (_________33289));
  nor2s1 ______436988(.DIN1 (_________29831), .DIN2 (______0__33276),
       .Q (_________33288));
  and2s1 _______436989(.DIN1 (_________33271), .DIN2 (________20909),
       .Q (_________33287));
  nnd2s1 _______436990(.DIN1 (_________33267), .DIN2 (_________33350),
       .Q (_________33286));
  nor2s1 _______436991(.DIN1 (______0__33248), .DIN2 (_________33269),
       .Q (_________33299));
  or2s1 ______436992(.DIN1 (______9__33266), .DIN2 (_________32968), .Q
       (_________33285));
  xor2s1 _______436993(.DIN1 (______0__33239), .DIN2 (_________33256),
       .Q (______0__33284));
  nor2s1 _______436994(.DIN1 (_________33273), .DIN2 (_________33261),
       .Q (_________33297));
  dffacs1 _________________0_436995(.CLRB (reset), .CLK (clk), .DIN
       (_________33265), .QN (_________18847));
  or2s1 _______436996(.DIN1 (_________33282), .DIN2 (_________33281),
       .Q (______9__33283));
  nor2s1 _______436997(.DIN1 (_________33262), .DIN2 (_________33279),
       .Q (_________33280));
  xor2s1 ______436998(.DIN1 (______9__29850), .DIN2 (______9__33275),
       .Q (______9__33291));
  nor2s1 _______436999(.DIN1 (_________29830), .DIN2 (______9__33275),
       .Q (______0__33276));
  nor2s1 _______437000(.DIN1 (_________33273), .DIN2 (_________33255),
       .Q (_________33274));
  nor2s1 _______437001(.DIN1 (_________33253), .DIN2 (_____0___33130),
       .Q (_________33272));
  nnd2s1 _____9_437002(.DIN1 (_________33244), .DIN2 (_________33186),
       .Q (_________33271));
  xor2s1 _____9_437003(.DIN1 (______9__33257), .DIN2 (_________30507),
       .Q (_________33270));
  nor2s1 _____9_437004(.DIN1 (_________33268), .DIN2 (_________33245),
       .Q (_________33269));
  nor2s1 _____9_437005(.DIN1 (________22409), .DIN2 (_________33246),
       .Q (_________33267));
  dffacs1 _________________0_437006(.CLRB (reset), .CLK (clk), .DIN
       (_________33252), .Q (_____________0___18779));
  nor2s1 _______437007(.DIN1 (____99___34528), .DIN2 (________23662),
       .Q (______9__33266));
  nnd2s1 _______437008(.DIN1 (_________33242), .DIN2 (_________33379),
       .Q (_________33265));
  nor2s1 ______437009(.DIN1 (_________32437), .DIN2 (______9__33238),
       .Q (_________33262));
  and2s1 ______437010(.DIN1 (_________33254), .DIN2 (_________33260),
       .Q (_________33261));
  and2s1 ______437011(.DIN1 (______0__33258), .DIN2 (_________33259),
       .Q (_________33282));
  nor2s1 _____437012(.DIN1 (_________33259), .DIN2 (______0__33258), .Q
       (_________33281));
  nor2s1 ____90_(.DIN1 (_________30489), .DIN2 (______9__33257), .Q
       (_________33277));
  nor2s1 _______437013(.DIN1 (_________33240), .DIN2 (_________33232),
       .Q (_________33256));
  hi1s1 _______437014(.DIN (_________33254), .Q (_________33255));
  nor2s1 ______437015(.DIN1 (_________33230), .DIN2 (_________33180),
       .Q (_________33253));
  nnd2s1 _______437016(.DIN1 (_________33233), .DIN2 (___9____24254),
       .Q (_________33252));
  nor2s1 _____9_437017(.DIN1 (_________33250), .DIN2 (_________33249),
       .Q (_________33251));
  nor2s1 ____90_437018(.DIN1 (______9__33247), .DIN2 (_________33243),
       .Q (______0__33248));
  nor2s1 ____90_437019(.DIN1 (_________33236), .DIN2 (_____0___33227),
       .Q (_________33246));
  nor2s1 ____9__437020(.DIN1 (_________32916), .DIN2 (_____09__33228),
       .Q (_________33245));
  nnd2s1 ____909(.DIN1 (_________33243), .DIN2 (_____9___33216), .Q
       (_________33244));
  nor2s1 _____437021(.DIN1 (_____00__33220), .DIN2 (______0__33229), .Q
       (______9__33275));
  nor2s1 _______437022(.DIN1 (_________33241), .DIN2 (_____0___33224),
       .Q (_________33242));
  nor2s1 _______437023(.DIN1 (_________33234), .DIN2 (_________33235),
       .Q (_________33273));
  nor2s1 _______437024(.DIN1 (_________33240), .DIN2 (______0__33239),
       .Q (_________33263));
  xor2s1 _____9_437025(.DIN1 (_________18858), .DIN2 (_____0__20962),
       .Q (______9__33238));
  nnd2s1 _______437026(.DIN1 (_________33236), .DIN2 (_____9___33217),
       .Q (_________33237));
  nor2s1 ____90_437027(.DIN1 (_________33208), .DIN2 (_____0___33221),
       .Q (_________33259));
  nor2s1 ____9__437028(.DIN1 (_________30332), .DIN2 (_____9___33215),
       .Q (______9__33257));
  nnd2s1 ______437029(.DIN1 (_________33235), .DIN2 (_________33234),
       .Q (_________33254));
  nnd2s1 ____90_437030(.DIN1 (_____90__33212), .DIN2 (_________33153),
       .Q (_________33233));
  hi1s1 _______437031(.DIN (_________33231), .Q (_________33232));
  xor2s1 _______437032(.DIN1 (_______19026), .DIN2
       (____________9___18791), .Q (_________33230));
  xor2s1 ____9_0(.DIN1 (_____99__33219), .DIN2 (_____99__29264), .Q
       (______0__33229));
  nor2s1 ____9__437033(.DIN1 (____999__34530), .DIN2 (_____0___33225),
       .Q (_____09__33228));
  xor2s1 ____9__437034(.DIN1 (_____9___30357), .DIN2 (____0____34592),
       .Q (_____0___33227));
  nor2s1 ____9__437035(.DIN1 (_________18858), .DIN2 (_____0___33226),
       .Q (_________33249));
  nnd2s1 ____9_9(.DIN1 (_____0___33225), .DIN2 (_________32922), .Q
       (_________33243));
  and2s1 ____9__437036(.DIN1 (_____0___33226), .DIN2 (_________18858),
       .Q (_________33250));
  or2s1 _______437037(.DIN1 (___0_0__23509), .DIN2 (_________33209), .Q
       (_____0___33224));
  nor2s1 _______437038(.DIN1 (____________9___18791), .DIN2
       (_____0___33222), .Q (_________33240));
  nnd2s1 _______437039(.DIN1 (_____0___33222), .DIN2
       (____________9___18791), .Q (_________33231));
  xor2s1 ______437040(.DIN1 (______0__33203), .DIN2 (____9___19200), .Q
       (_________33235));
  nor2s1 ____9__437041(.DIN1 (_____00__33220), .DIN2 (_____99__33219),
       .Q (_____0___33221));
  xor2s1 ____9__437042(.DIN1 (_________33200), .DIN2 (_________31326),
       .Q (_____9___33218));
  nnd2s1 ____90_437043(.DIN1 (_________33210), .DIN2 (inData[28]), .Q
       (_____9___33217));
  nnd2s1 ____9__437044(.DIN1 (_________33211), .DIN2 (_________32923),
       .Q (_____9___33216));
  nor2s1 ____9__437045(.DIN1 (_________30337), .DIN2 (____0____34592),
       .Q (_____9___33215));
  nnd2s1 ____90_437046(.DIN1 (_____9___33214), .DIN2 (_____9___33213),
       .Q (_____0___33223));
  dffacs1 ___________________437047(.CLRB (reset), .CLK (clk), .DIN
       (______9__33202), .Q (_________18858));
  xor2s1 ____9__437048(.DIN1 (_________33191), .DIN2 (_________31431),
       .Q (_____90__33212));
  hi1s1 ____9__437049(.DIN (_________33211), .Q (_____0___33225));
  dffacs1 ___________________437050(.CLRB (reset), .CLK (clk), .DIN
       (_________33197), .QN (_________________18774));
  xor2s1 ____9__437051(.DIN1 (_____________0___18779), .DIN2
       (_____________9___18778), .Q (_________33210));
  nor2s1 _____9_437052(.DIN1 (______0__33336), .DIN2 (_________33194),
       .Q (_________33209));
  nor2s1 ____9__437053(.DIN1 (_____0___29807), .DIN2 (_________33205),
       .Q (_________33208));
  dffacs1 ________________9_(.CLRB (reset), .CLK (clk), .DIN
       (_________33195), .Q (____________9___18791));
  nnd2s1 ____9_437054(.DIN1 (_________33206), .DIN2 (_________33196),
       .Q (_________33207));
  nnd2s1 ____9__437055(.DIN1 (_________33205), .DIN2 (_________29759),
       .Q (_____99__33219));
  xor2s1 ____9__437056(.DIN1 (_________33182), .DIN2 (_________33204),
       .Q (_________33211));
  dffacs1 ___________________437057(.CLRB (reset), .CLK (clk), .DIN
       (______0__33193), .Q (_________________18777));
  nor2s1 ____9__437058(.DIN1 (______9__33096), .DIN2 (_________33189),
       .Q (______0__33203));
  nnd2s1 ____9__437059(.DIN1 (_________33187), .DIN2 (________22059),
       .Q (______9__33202));
  nnd2s1 ____9_437060(.DIN1
       (______________________________________0_____________18890),
       .DIN2 (_________33190), .Q (_____9___33214));
  nnd2s1 ____9_437061(.DIN1 (______9__30135), .DIN2
       (_____________9___18778), .Q (_________33201));
  nor2s1 ____9__437062(.DIN1 (_________33199), .DIN2 (_________33198),
       .Q (_________33200));
  nnd2s1 ____9__437063(.DIN1 (_________32986), .DIN2 (______9__33183),
       .Q (_________33197));
  hi1s1 ____9__437064(.DIN (_____________9___18778), .Q
       (_________33196));
  nnd2s1 ____90_437065(.DIN1 (_________33181), .DIN2 (________23899),
       .Q (_________33195));
  xor2s1 ____9__437066(.DIN1 (_________33105), .DIN2 (_________33188),
       .Q (_________33194));
  nnd2s1 ____9__437067(.DIN1 (_________33078), .DIN2 (_________33178),
       .Q (______0__33193));
  nnd2s1 ____9_437068(.DIN1 (_________30104), .DIN2
       (_____________________________________18837), .Q
       (_____9___33213));
  xor2s1 ____9__437069(.DIN1 (______0__33175), .DIN2 (______0__33184),
       .Q (______9__33192));
  xor2s1 ____9__437070(.DIN1 (_________33167), .DIN2
       (_____________0___18764), .Q (_________33191));
  xnr2s1 ____9__437071(.DIN1 (_________32644), .DIN2 (_________33168),
       .Q (_________33205));
  dffacs1 ___________________437072(.CLRB (reset), .CLK (clk), .DIN
       (_________33179), .Q (_________________18765));
  hi1s1 ____9_437073(.DIN (_____________________________________18837),
       .Q (_________33190));
  nor2s1 ____9__437074(.DIN1 (_________33094), .DIN2 (_________33188),
       .Q (_________33189));
  nnd2s1 ____9__437075(.DIN1 (_________33171), .DIN2 (_________33186),
       .Q (_________33187));
  dffacs1 _________________9_437076(.CLRB (reset), .CLK (clk), .DIN
       (_________33172), .Q (_____________9___18778));
  nor2s1 ____9__437077(.DIN1 (______0__33184), .DIN2 (______9__30581),
       .Q (_________33185));
  nnd2s1 ____9_437078(.DIN1 (_________33177), .DIN2 (_________33169),
       .Q (______9__33183));
  nnd2s1 ____9_437079(.DIN1 (_________33170), .DIN2 (_____09__33135),
       .Q (_________33182));
  xor2s1 ____9__437080(.DIN1 (_________33161), .DIN2 (_________33384),
       .Q (_________33198));
  nnd2s1 ____9__437081(.DIN1 (_________33163), .DIN2 (_________33180),
       .Q (_________33181));
  nnd2s1 ____9__437082(.DIN1 (_________33059), .DIN2 (______9__33165),
       .Q (_________33179));
  dffacs1 _____________9____437083(.CLRB (reset), .CLK (clk), .DIN
       (_________33164), .QN
       (_____________________________________18837));
  nnd2s1 ____9_437084(.DIN1 (_________33177), .DIN2 (_________33162),
       .Q (_________33178));
  nor2s1 ____9__437085(.DIN1 (______0__33166), .DIN2 (______0__33175),
       .Q (_________33176));
  nnd2s1 ____9__437086(.DIN1 (_________33154), .DIN2 (________23569),
       .Q (_________33172));
  xor2s1 ____9__437087(.DIN1 (______9__33145), .DIN2 (_________32902),
       .Q (_________33171));
  nor2s1 ____9__437088(.DIN1 (_________33071), .DIN2 (_________33157),
       .Q (_________33188));
  nnd2s1 ____9_437089(.DIN1 (_________30107), .DIN2 (______9__33155),
       .Q (______0__33239));
  nor2s1 ____9__437090(.DIN1 (_________33148), .DIN2 (_________32895),
       .Q (_________33170));
  nnd2s1 ____9__437091(.DIN1 (_________33150), .DIN2 (______0__33136),
       .Q (_________33169));
  nnd2s1 ____9__437092(.DIN1 (_________33152), .DIN2 (_________29751),
       .Q (_________33168));
  xor2s1 ____9__437093(.DIN1 (_________33158), .DIN2 (_________33206),
       .Q (_________33167));
  hi1s1 ____9_437094(.DIN (______0__33166), .Q (______0__33184));
  nnd2s1 ____9__437095(.DIN1 (_____0___33034), .DIN2 (_________33143),
       .Q (______9__33165));
  nnd2s1 ____9__437096(.DIN1 (_________33147), .DIN2 (_________34393),
       .Q (_________33164));
  xor2s1 ____9__437097(.DIN1 (______0__33156), .DIN2 (_________33091),
       .Q (_________33163));
  xor2s1 ____9__437098(.DIN1 (_________________18774), .DIN2
       (_________33149), .Q (_________33162));
  nnd2s1 ____9__437099(.DIN1 (_________33159), .DIN2 (_________33160),
       .Q (_________33161));
  xor2s1 ____9__437100(.DIN1 (_________29752), .DIN2 (_________33151),
       .Q (______0__33166));
  nor2s1 ____9__437101(.DIN1 (_________33160), .DIN2 (_________33159),
       .Q (_________33199));
  nor2s1 ____999(.DIN1 (_____99__33028), .DIN2 (_________33158), .Q
       (_________33173));
  dffacs1 ___________________437102(.CLRB (reset), .CLK (clk), .DIN
       (______0__33146), .Q (_________________18766));
  and2s1 ____9__437103(.DIN1 (______0__33156), .DIN2 (_________33073),
       .Q (_________33157));
  nor2s1 ____9_437104(.DIN1 (____0____30034), .DIN2 (_________33142),
       .Q (______9__33155));
  nnd2s1 ____9__437105(.DIN1 (_________33140), .DIN2 (_________33153),
       .Q (_________33154));
  nnd2s1 ____9__437106(.DIN1 (_________33151), .DIN2 (_________29750),
       .Q (_________33152));
  or2s1 ____9_437107(.DIN1 (_________________18774), .DIN2
       (_________33149), .Q (_________33150));
  nor2s1 ____99_(.DIN1 (_________33138), .DIN2 (_________32871), .Q
       (_________33148));
  xor2s1 ____9__437108(.DIN1 (_________33141), .DIN2 (_________30106),
       .Q (_________33147));
  nnd2s1 ____990(.DIN1 (_____0___33133), .DIN2 (____9___23610), .Q
       (______0__33146));
  dffacs1 ___________________437109(.CLRB (reset), .CLK (clk), .DIN
       (_____0___33134), .QN (______0__34441));
  xor2s1 ____99_437110(.DIN1 (_________33137), .DIN2 (_________33144),
       .Q (______9__33145));
  xor2s1 ____99_437111(.DIN1 (_____9___33124), .DIN2 (_____9___33020),
       .Q (_________33143));
  nor2s1 ___90__(.DIN1 (_________33113), .DIN2 (_____0___33132), .Q
       (_________33158));
  xor2s1 ____99_437112(.DIN1 (_____00__33127), .DIN2 (_________31020),
       .Q (_________33160));
  nor2s1 ____9__437113(.DIN1 (_________33141), .DIN2 (____0_0__30056),
       .Q (_________33142));
  xor2s1 ____99_437114(.DIN1 (_____9___33120), .DIN2 (_____0___33131),
       .Q (_________33140));
  or2s1 ____9__437115(.DIN1 (______0__33373), .DIN2 (_____0___33129),
       .Q (_________33139));
  xor2s1 ____9__437116(.DIN1 (_____9___33123), .DIN2 (_____0___32570),
       .Q (______0__33156));
  nor2s1 ___900_(.DIN1 (_____9___31529), .DIN2 (_________33137), .Q
       (_________33138));
  nnd2s1 ___900_437117(.DIN1 (_________33082), .DIN2
       (_________________18775), .Q (______0__33136));
  nnd2s1 ___900_437118(.DIN1 (_________33137), .DIN2 (______9__32872),
       .Q (_____09__33135));
  nnd2s1 ___900_437119(.DIN1 (_____0___33128), .DIN2 (_____9___33125),
       .Q (_________33151));
  or2s1 ___90__437120(.DIN1 (_________________18775), .DIN2
       (_________________18776), .Q (_________33149));
  or2s1 ___900_437121(.DIN1 (_________31569), .DIN2 (_____9___33122),
       .Q (_____0___33134));
  nnd2s1 ___900_437122(.DIN1 (_____9___33121), .DIN2 (_________33103),
       .Q (_____0___33133));
  nor2s1 ___90__437123(.DIN1 (_____9___33119), .DIN2 (_____0___33131),
       .Q (_____0___33132));
  nor2s1 ____99_437124(.DIN1 (______0__33336), .DIN2 (______9__33116),
       .Q (_____0___33130));
  xor2s1 ____9_437125(.DIN1 (______9__33106), .DIN2 (_________33114),
       .Q (_____0___33129));
  nnd2s1 ___90__437126(.DIN1 (_____99__33126), .DIN2 (_________29508),
       .Q (_____0___33128));
  nnd2s1 ___9000(.DIN1 (_________33115), .DIN2 (______0__33097), .Q
       (_________33141));
  and2s1 ___90__437127(.DIN1 (_____99__33126), .DIN2 (_____9___33125),
       .Q (_____00__33127));
  xor2s1 ___90__437128(.DIN1 (_____9___33118), .DIN2 (_________34442),
       .Q (_____9___33124));
  nor2s1 ___90_9(.DIN1 (_________31616), .DIN2 (_________33112), .Q
       (_________33137));
  dffacs1 ___________________437129(.CLRB (reset), .CLK (clk), .DIN
       (_________33110), .Q (_________________18775));
  nor2s1 ____99_437130(.DIN1 (_________33101), .DIN2 (_________33108),
       .Q (_____9___33123));
  nnd2s1 ___90__437131(.DIN1 (_________33104), .DIN2 (_________31619),
       .Q (_____9___33122));
  xor2s1 ___90__437132(.DIN1 (_________31617), .DIN2 (_________33111),
       .Q (_____9___33121));
  xor2s1 ___90__437133(.DIN1 (_________18844), .DIN2 (_____90__33117),
       .Q (_____9___33120));
  nor2s1 ___90__437134(.DIN1 (_____9___33118), .DIN2 (_____90__33117),
       .Q (_____9___33119));
  nor2s1 ___9009(.DIN1 (______0__33087), .DIN2 (_________33102), .Q
       (______9__33116));
  or2s1 ___900_437135(.DIN1 (_________33099), .DIN2 (_________33114),
       .Q (_________33115));
  nor2s1 ___90__437136(.DIN1 (_________18844), .DIN2 (____0____30070),
       .Q (_________33113));
  xor2s1 ___90__437137(.DIN1 (_________33089), .DIN2 (____0____32835),
       .Q (_________33260));
  and2s1 ___90_0(.DIN1 (_________33111), .DIN2 (_________31597), .Q
       (_________33112));
  nnd2s1 ___90_437138(.DIN1 (______9__33047), .DIN2 (_________33092),
       .Q (_________33110));
  nnd2s1 ___90__437139(.DIN1 (_________33109), .DIN2
       (_______________0___________________), .Q (_____99__33126));
  or2s1 ___90__437140(.DIN1 (_______________0___________________),
       .DIN2 (_________33109), .Q (_____9___33125));
  xnr2s1 ___90_437141(.DIN1 (_________33204), .DIN2 (_________33088),
       .Q (_____0___33131));
  xor2s1 ___900_437142(.DIN1 (_________33100), .DIN2 (______0__33107),
       .Q (_________33108));
  xor2s1 ___90_437143(.DIN1 (_________33098), .DIN2
       (________________18790), .Q (______9__33106));
  xor2s1 ___90__437144(.DIN1 (_________30242), .DIN2 (_________33095),
       .Q (_________33105));
  nnd2s1 ___90__437145(.DIN1 (_________33090), .DIN2 (_________33103),
       .Q (_________33104));
  hi1s1 ___90__437146(.DIN (_________18844), .Q (_____9___33118));
  nor2s1 ___90__437147(.DIN1 (_________33101), .DIN2 (_________33100),
       .Q (_________33102));
  nor2s1 ___90__437148(.DIN1 (________________18790), .DIN2
       (_________33098), .Q (_________33099));
  nnd2s1 ___90__437149(.DIN1 (_________33098), .DIN2
       (________________18790), .Q (______0__33097));
  nor2s1 ___90__437150(.DIN1 (_________33095), .DIN2 (_________33093),
       .Q (______9__33096));
  and2s1 ___90__437151(.DIN1 (_________33093), .DIN2 (_________33095),
       .Q (_________33094));
  nnd2s1 ___90__437152(.DIN1 (_________33079), .DIN2 (inData[28]), .Q
       (_________33092));
  xor2s1 ___90_437153(.DIN1 (______0__33077), .DIN2 (_________32624),
       .Q (_________33091));
  nor2s1 ___90__437154(.DIN1 (_________31548), .DIN2 (_________33084),
       .Q (_________33111));
  nor2s1 ___90__437155(.DIN1 (____0____32834), .DIN2 (_________33081),
       .Q (_________33109));
  dffacs1 _________________9_437156(.CLRB (reset), .CLK (clk), .DIN
       (_________33085), .Q (_________18844));
  xor2s1 ___90__437157(.DIN1 (_________31550), .DIN2 (_________33083),
       .Q (_________33090));
  xor2s1 ___90_437158(.DIN1 (____09___32842), .DIN2 (_________33080),
       .Q (_________33089));
  nnd2s1 ___90_437159(.DIN1 (______9__33076), .DIN2 (_________33066),
       .Q (_________33088));
  nor2s1 ___90__437160(.DIN1 (_________33054), .DIN2 (______9__33086),
       .Q (______0__33087));
  nnd2s1 ___90__437161(.DIN1 (______9__33086), .DIN2 (_________33017),
       .Q (_________33100));
  xor2s1 ___90__437162(.DIN1 (_________33068), .DIN2 (_________31956),
       .Q (_________33095));
  dffacs1 __________________437163(.CLRB (reset), .CLK (clk), .DIN
       (_________33074), .Q (________________18790));
  or2s1 ___90__437164(.DIN1 (_____0___33037), .DIN2 (_________33075),
       .Q (_________33085));
  nor2s1 ___90__437165(.DIN1 (_________31549), .DIN2 (_________33083),
       .Q (_________33084));
  or2s1 ___90__437166(.DIN1 (_________________18776), .DIN2
       (_________________18774), .Q (_________33082));
  nor2s1 ___90__437167(.DIN1 (____0____32836), .DIN2 (_________33080),
       .Q (_________33081));
  nor2s1 ___90__437168(.DIN1 (_________________18776), .DIN2
       (_____0__23837), .Q (_________33079));
  nnd2s1 ___90__437169(.DIN1 (_________33069), .DIN2 (_________33153),
       .Q (_________33078));
  xor2s1 ___90_437170(.DIN1 (____0____30045), .DIN2 (_________33072),
       .Q (______0__33077));
  nor2s1 ___90__437171(.DIN1 (______0__33010), .DIN2 (______0__33067),
       .Q (______9__33076));
  nnd2s1 ___90__437172(.DIN1 (_________32971), .DIN2 (_________33064),
       .Q (_________33075));
  nor2s1 ___90__437173(.DIN1 (_________________0___18660), .DIN2
       (_________33062), .Q (_________33074));
  nor2s1 ___90__437174(.DIN1 (_____0___29363), .DIN2 (______9__33057),
       .Q (_________33080));
  xor2s1 ___90_437175(.DIN1 (_________33055), .DIN2 (_________32410),
       .Q (______9__33086));
  nnd2s1 ___90_437176(.DIN1 (_________33070), .DIN2 (_________33072),
       .Q (_________33073));
  nor2s1 ___90_437177(.DIN1 (_________33072), .DIN2 (_________33070),
       .Q (_________33071));
  nnd2s1 ___90__437178(.DIN1 (_________33060), .DIN2 (____9____32737),
       .Q (_________33083));
  dffacs1 ___________________437179(.CLRB (reset), .CLK (clk), .DIN
       (_________33063), .QN (_________________18763));
  dffacs1 ___________________437180(.CLRB (reset), .CLK (clk), .DIN
       (_________33061), .QN (_________________18776));
  xor2s1 ___90__437181(.DIN1 (_________33049), .DIN2 (_________33053),
       .Q (_________33069));
  xor2s1 ___90__437182(.DIN1 (_____0___29364), .DIN2 (_________33056),
       .Q (_________33068));
  nor2s1 ___90_437183(.DIN1 (_________31431), .DIN2 (_________33065),
       .Q (______0__33067));
  nnd2s1 ___90__437184(.DIN1 (_________33065), .DIN2 (_________35110),
       .Q (_________33066));
  nnd2s1 ___90__437185(.DIN1 (______0__33058), .DIN2 (_________33052),
       .Q (_________33064));
  nnd2s1 ___90__437186(.DIN1 (_________32888), .DIN2 (_________33051),
       .Q (_________33063));
  xor2s1 ___90__437187(.DIN1 (_________33046), .DIN2 (____0____34594),
       .Q (_________33062));
  nnd2s1 ___90__437188(.DIN1 (_________33050), .DIN2 (________23603),
       .Q (_________33061));
  xor2s1 ___90__437189(.DIN1 (_________33040), .DIN2 (_________35066),
       .Q (_________33060));
  or2s1 ___90_437190(.DIN1 (______0__33058), .DIN2 (______0__33048), .Q
       (_________33059));
  nor2s1 ___90__437191(.DIN1 (_________29345), .DIN2 (_________33056),
       .Q (______9__33057));
  xor2s1 ___90__437192(.DIN1 (_________33042), .DIN2 (_____0___33031),
       .Q (_________33072));
  nor2s1 ___90__437193(.DIN1 (_________33045), .DIN2 (_________33044),
       .Q (_________33055));
  nor2s1 ___90__437194(.DIN1 (_________33018), .DIN2 (_________33101),
       .Q (_________33054));
  nor2s1 ___909_(.DIN1 (_________33014), .DIN2 (_________33053), .Q
       (_________33065));
  dffacs1 ___________________437195(.CLRB (reset), .CLK (clk), .DIN
       (_____09__33038), .Q (_________34442));
  nnd2s1 ___90__437196(.DIN1 (_____0___33033), .DIN2 (inData[22]), .Q
       (_________33052));
  nnd2s1 ___90__437197(.DIN1 (_____0___33035), .DIN2 (inData[18]), .Q
       (_________33051));
  nnd2s1 ___90_437198(.DIN1 (_____00__33029), .DIN2 (_________33153),
       .Q (_________33050));
  xor2s1 ___909_437199(.DIN1 (____99___34529), .DIN2 (_________33388),
       .Q (_________33049));
  xor2s1 ___909_437200(.DIN1 (____9____32739), .DIN2 (______0__33039),
       .Q (______0__33048));
  nor2s1 ___909_437201(.DIN1 (_________33041), .DIN2 (_____0___33032),
       .Q (_________33056));
  dffacs1 __________________437202(.CLRB (reset), .CLK (clk), .DIN
       (_____0___33036), .Q (________________18789));
  nnd2s1 ___90__437203(.DIN1 (_____9___33027), .DIN2 (_________33153),
       .Q (______9__33047));
  nor2s1 ___90__437204(.DIN1 (_________33045), .DIN2 (_________33043),
       .Q (_________33046));
  nor2s1 ___90__437205(.DIN1 (_________33043), .DIN2 (____0____34594),
       .Q (_________33044));
  xor2s1 ___909_437206(.DIN1 (_________33015), .DIN2 (_____0___33866),
       .Q (_________33101));
  nor2s1 ___9_0_(.DIN1 (_____0___33030), .DIN2 (_________33041), .Q
       (_________33042));
  and2s1 ___9_00(.DIN1 (____9____32738), .DIN2 (______0__33039), .Q
       (_________33040));
  or2s1 ___9099(.DIN1 (_____0___33037), .DIN2 (_____9___33023), .Q
       (_____09__33038));
  nor2s1 ___9_0_437207(.DIN1 (____90___29905), .DIN2 (_____9___33025),
       .Q (_________33053));
  nnd2s1 ___90__437208(.DIN1 (______9__33019), .DIN2 (________24108),
       .Q (_____0___33036));
  and2s1 ___909_437209(.DIN1 (_____0___33034), .DIN2 (_________33016),
       .Q (_____0___33035));
  xnr2s1 ___9_0_437210(.DIN1 (_________34442), .DIN2
       (_____________0___18764), .Q (_____0___33033));
  nor2s1 ___9_0_437211(.DIN1 (_____0___33031), .DIN2 (_____0___33030),
       .Q (_____0___33032));
  xor2s1 ___9_0_437212(.DIN1 (____9____29924), .DIN2 (_____9___33024),
       .Q (_____00__33029));
  nor2s1 ___9_0_437213(.DIN1 (_____________0___18764), .DIN2
       (_________33206), .Q (_____99__33028));
  xor2s1 ___9_0_437214(.DIN1 (_________33002), .DIN2 (_____9___33026),
       .Q (_____9___33027));
  nor2s1 ___9__0(.DIN1 (_____9___29892), .DIN2 (_____9___33024), .Q
       (_____9___33025));
  nnd2s1 ___9_09(.DIN1 (_________33011), .DIN2 (___0____23470), .Q
       (_____9___33023));
  xor2s1 ___909_437215(.DIN1 (_________33006), .DIN2 (_____9___33022),
       .Q (_________33043));
  nnd2s1 ___9___(.DIN1 (_________33206), .DIN2
       (_____________0___18764), .Q (_____9___33021));
  nnd2s1 ___9___437216(.DIN1 (_____________0___18764), .DIN2
       (_________________18765), .Q (_____9___33020));
  nor2s1 ___9__9(.DIN1 (____________9___18773), .DIN2 (_________33013),
       .Q (_________33041));
  nnd2s1 ___9___437217(.DIN1 (______9__33009), .DIN2 (____0____32811),
       .Q (______0__33039));
  dffacs1 _________________0_437218(.CLRB (reset), .CLK (clk), .DIN
       (_________33008), .QN (_________34448));
  nnd2s1 ___9090(.DIN1 (_________33005), .DIN2 (_________32925), .Q
       (______9__33019));
  hi1s1 ___9___437219(.DIN (_________33017), .Q (_________33018));
  xor2s1 ___9___437220(.DIN1 (_________32960), .DIN2 (_________18843),
       .Q (_________33016));
  nnd2s1 ___9___437221(.DIN1 (____9____29962), .DIN2 (_________33001),
       .Q (_________33015));
  nor2s1 ___9__437222(.DIN1 (____9____32718), .DIN2 (_________33012),
       .Q (_____0___33030));
  and2s1 ___9___437223(.DIN1 (_________33388), .DIN2 (_________18843),
       .Q (_________33014));
  hi1s1 ___9___437224(.DIN (_________33012), .Q (_________33013));
  or2s1 ___9___437225(.DIN1 (______0__33058), .DIN2 (_________32998),
       .Q (_________33011));
  nnd2s1 ___9___437226(.DIN1 (____9____29963), .DIN2 (______0__33000),
       .Q (_________33017));
  nor2s1 ___9___437227(.DIN1 (_________18843), .DIN2 (_________33388),
       .Q (______0__33010));
  xor2s1 ___9___437228(.DIN1 (_________32994), .DIN2 (_________33385),
       .Q (______9__33009));
  or2s1 ___9__437229(.DIN1 (_________32919), .DIN2 (_________32997), .Q
       (_________33008));
  xor2s1 ___9___437230(.DIN1 (______0__32992), .DIN2 (_________33007),
       .Q (_____9___33024));
  dffacs1 _________________0_437231(.CLRB (reset), .CLK (clk), .DIN
       (_________32999), .Q (_____________0___18764));
  nnd2s1 ___9___437232(.DIN1 (_________33003), .DIN2 (_________33004),
       .Q (_________33006));
  xor2s1 ___9_0_437233(.DIN1 (______9__32991), .DIN2 (_________31154),
       .Q (_________33005));
  nor2s1 ___9___437234(.DIN1 (_________33004), .DIN2 (_________33003),
       .Q (_________33045));
  nnd2s1 ___9___437235(.DIN1 (_________32996), .DIN2 (____0____29130),
       .Q (_________33012));
  xor2s1 ___9___437236(.DIN1 (_________32988), .DIN2 (______0__32899),
       .Q (_________33002));
  hi1s1 ___9__437237(.DIN (______0__33000), .Q (_________33001));
  nnd2s1 ___9__437238(.DIN1 (_________32989), .DIN2 (_________34844),
       .Q (_________32999));
  xor2s1 ___9___437239(.DIN1 (____0____29141), .DIN2 (_________32995),
       .Q (______0__33000));
  xor2s1 ___9___437240(.DIN1 (____0____32812), .DIN2 (_________32993),
       .Q (_________32998));
  nnd2s1 ___9___437241(.DIN1 (_________32905), .DIN2 (_________32987),
       .Q (_________32997));
  dffacs1 ___________________437242(.CLRB (reset), .CLK (clk), .DIN
       (_________32990), .Q (_________18843));
  or2s1 ___9___437243(.DIN1 (____0____29129), .DIN2 (_________32995),
       .Q (_________32996));
  xor2s1 ___9___437244(.DIN1 (_________32982), .DIN2 (_____9___28896),
       .Q (_________33004));
  or2s1 ___9___437245(.DIN1 (_________32993), .DIN2 (____0_9__32809),
       .Q (_________32994));
  nnd2s1 ___9___437246(.DIN1 (______0__32984), .DIN2 (_________32900),
       .Q (______0__32992));
  xor2s1 ___9___437247(.DIN1 (_________32978), .DIN2 (_________32966),
       .Q (______9__32991));
  or2s1 ___9___437248(.DIN1 (_____0___33037), .DIN2 (_________32981),
       .Q (_________32990));
  or2s1 ___9__437249(.DIN1 (______0__33058), .DIN2 (_________32980), .Q
       (_________32989));
  xor2s1 ___9___437250(.DIN1 (_________34443), .DIN2 (______9__32983),
       .Q (_________32988));
  nnd2s1 ___9___437251(.DIN1 (______9__32927), .DIN2 (_________32979),
       .Q (_________32987));
  nnd2s1 ___9___437252(.DIN1 (_________32975), .DIN2 (_________33153),
       .Q (_________32986));
  nnd2s1 ___9__437253(.DIN1 (_________32887), .DIN2 (______9__32983),
       .Q (______0__32984));
  nor2s1 ___9___437254(.DIN1 (____00___32752), .DIN2 (_________32977),
       .Q (_________32995));
  nor2s1 ___9__437255(.DIN1 (____0____32796), .DIN2 (______0__32974),
       .Q (_________32993));
  xor2s1 ___9___437256(.DIN1 (_________32976), .DIN2
       (________________18772), .Q (_________32982));
  nnd2s1 ___9___437257(.DIN1 (_____9___32933), .DIN2 (_________32970),
       .Q (_________32981));
  xor2s1 ___9___437258(.DIN1 (____0____32804), .DIN2 (______9__32973),
       .Q (_________32980));
  nnd2s1 ___9___437259(.DIN1 (_________32969), .DIN2 (inData[2]), .Q
       (_________32979));
  xor2s1 ___9___437260(.DIN1 (_________32972), .DIN2 (_________32965),
       .Q (_________32978));
  and2s1 ___9___437261(.DIN1 (_________32976), .DIN2 (____999__32750),
       .Q (_________32977));
  xor2s1 ___9___437262(.DIN1 (_________32958), .DIN2 (_________32962),
       .Q (_________32975));
  and2s1 ___9__437263(.DIN1 (______9__32973), .DIN2 (____0____32792),
       .Q (______0__32974));
  and2s1 ___9___437264(.DIN1 (______0__32964), .DIN2 (_________32972),
       .Q (_________32985));
  nor2s1 ___9___437265(.DIN1 (_________32957), .DIN2 (______9__32963),
       .Q (______9__32983));
  or2s1 ___9___437266(.DIN1 (______0__33058), .DIN2 (_________32959),
       .Q (_________32971));
  nnd2s1 ___9___437267(.DIN1 (______0__33058), .DIN2 (_________32961),
       .Q (_________32970));
  xnr2s1 ___9__437268(.DIN1 (_________________18752), .DIN2
       (____99__21810), .Q (_________32969));
  nor2s1 ___9___437269(.DIN1 (____0____31829), .DIN2 (_________32955),
       .Q (_________32968));
  or2s1 ___9___437270(.DIN1 (_________32966), .DIN2 (_________32965),
       .Q (_________32967));
  nnd2s1 ___9___437271(.DIN1 (_________32965), .DIN2 (_________32966),
       .Q (______0__32964));
  nor2s1 ___9___437272(.DIN1 (_________32953), .DIN2 (_________32962),
       .Q (______9__32963));
  xor2s1 ___9___437273(.DIN1 (_________32951), .DIN2 (____9____31746),
       .Q (_________32976));
  nnd2s1 ___9__437274(.DIN1 (______0__32954), .DIN2 (_________31022),
       .Q (______9__32973));
  xor2s1 ___9___437275(.DIN1 (_________32960), .DIN2
       (_________________18762), .Q (_________32961));
  nnd2s1 ___9___437276(.DIN1 (_________32952), .DIN2 (_____0___32941),
       .Q (_________32972));
  xor2s1 ___9___437277(.DIN1 (_________31023), .DIN2 (____0____34596),
       .Q (_________32959));
  xor2s1 ___9___437278(.DIN1 (_________32956), .DIN2
       (_________________18762), .Q (_________32958));
  nor2s1 ___9___437279(.DIN1 (_________32950), .DIN2 (_________32956),
       .Q (_________32957));
  xor2s1 ___9___437280(.DIN1 (_____0___32942), .DIN2 (_____0___32939),
       .Q (_________32955));
  xor2s1 ___9___437281(.DIN1 (______0__32945), .DIN2 (_________32946),
       .Q (_________32966));
  or2s1 ___9___437282(.DIN1 (____0____30974), .DIN2 (____0____34596),
       .Q (______0__32954));
  nor2s1 ___9__437283(.DIN1 (_________________18762), .DIN2
       (_____9___29707), .Q (_________32953));
  dffacs1 ___________________437284(.CLRB (reset), .CLK (clk), .DIN
       (_________32949), .Q (_________________18752));
  xor2s1 ___9___437285(.DIN1 (_____0___32940), .DIN2 (____0____30981),
       .Q (_________32952));
  nor2s1 ___9_90(.DIN1 (_____09__32944), .DIN2 (_________32947), .Q
       (_________32951));
  hi1s1 ___9_9_(.DIN (_________________18762), .Q (_________32950));
  dffacs1 __________________437286(.CLRB (reset), .CLK (clk), .DIN
       (_________32948), .QN (_________34433));
  dffacs1 ___________________437287(.CLRB (reset), .CLK (clk), .DIN
       (_____0___32938), .Q (_________________18762));
  nnd2s1 ___9_437288(.DIN1 (_____0___32937), .DIN2 (_________34992), .Q
       (_________32949));
  or2s1 ___9___437289(.DIN1 (______9__30207), .DIN2 (_____00__32936),
       .Q (_________32948));
  nor2s1 ___9_9_437290(.DIN1 (_________32946), .DIN2 (_____0___32943),
       .Q (_________32947));
  nor2s1 ___9_9_437291(.DIN1 (_____09__32944), .DIN2 (_____0___32943),
       .Q (______0__32945));
  and2s1 ___9_9_437292(.DIN1 (_____99__32935), .DIN2 (_____0___32941),
       .Q (_____0___32942));
  nor2s1 ___9_9_437293(.DIN1 (_____0___32939), .DIN2 (_____9___32934),
       .Q (_____0___32940));
  nnd2s1 ___9_0_437294(.DIN1 (____0____32794), .DIN2 (_____9___32931),
       .Q (_____0___32938));
  nor2s1 ___9__437295(.DIN1 (________22240), .DIN2 (_____90__32928), .Q
       (_____0___32937));
  nnd2s1 ___9___437296(.DIN1 (_________32926), .DIN2 (________22976),
       .Q (_____00__32936));
  and2s1 ___9_0_437297(.DIN1 (_____9___32932), .DIN2
       (________________18771), .Q (_____09__32944));
  hi1s1 ___9_0_437298(.DIN (_____9___32934), .Q (_____99__32935));
  or2s1 ___9_0_437299(.DIN1 (______0__33058), .DIN2 (_________32924),
       .Q (_____9___32933));
  nor2s1 ___9_0_437300(.DIN1 (________________18771), .DIN2
       (_____9___32932), .Q (_____0___32943));
  nnd2s1 ___9_437301(.DIN1 (_________32921), .DIN2 (inData[20]), .Q
       (_____9___32931));
  xor2s1 ___9_0_437302(.DIN1 (_________32914), .DIN2 (_________33894),
       .Q (_____9___32934));
  nor2s1 ___9___437303(.DIN1 (______9__32927), .DIN2 (______0__32918),
       .Q (_____90__32928));
  dffacs1 ___________________437304(.CLRB (reset), .CLK (clk), .DIN
       (_________32920), .QN (_________34449));
  nnd2s1 ___9_9_437305(.DIN1 (_________32915), .DIN2 (_________32925),
       .Q (_________32926));
  xor2s1 ___9___437306(.DIN1 (____9_0__30854), .DIN2 (______9__32917),
       .Q (_________32924));
  hi1s1 ___9___437307(.DIN (_________32922), .Q (_________32923));
  xnr2s1 ___9___437308(.DIN1 (___0____21656), .DIN2 (_________32910),
       .Q (_____9___32932));
  or2s1 ___9___437309(.DIN1 (______9__32908), .DIN2 (_________32891),
       .Q (_________32921));
  or2s1 ___9__437310(.DIN1 (_________32919), .DIN2 (______0__32909), .Q
       (_________32920));
  nnd2s1 ___9___437311(.DIN1 (_________29575), .DIN2 (_________32907),
       .Q (_____0___32941));
  xor2s1 ___9___437312(.DIN1 (_________32434), .DIN2 (______9__32898),
       .Q (______0__32918));
  and2s1 ___9___437313(.DIN1 (______9__32917), .DIN2 (____0_0__34541),
       .Q (_____9___32929));
  nor2s1 ___9___437314(.DIN1 (____999__34530), .DIN2 (_________32916),
       .Q (_________32922));
  xor2s1 ___9_0_437315(.DIN1 (______0__32890), .DIN2 (_________32903),
       .Q (_________32915));
  nor2s1 ___9___437316(.DIN1 (______0__32881), .DIN2 (_________32904),
       .Q (_____0___32939));
  nnd2s1 ___9___437317(.DIN1 (_________29576), .DIN2 (_________32906),
       .Q (_________32914));
  nor2s1 ___9___437318(.DIN1 (_________32912), .DIN2 (_________32911),
       .Q (_________32913));
  nnd2s1 ___9___437319(.DIN1 (_________32893), .DIN2 (_________28848),
       .Q (_________32910));
  nnd2s1 ___9__437320(.DIN1 (____09___32847), .DIN2 (_________32892),
       .Q (______0__32909));
  and2s1 ___9__437321(.DIN1 (_________32897), .DIN2
       (_________________18763), .Q (______9__32908));
  hi1s1 ___9___437322(.DIN (_________32906), .Q (_________32907));
  or2s1 ___9__437323(.DIN1 (______9__32927), .DIN2 (_________32885), .Q
       (_________32905));
  xor2s1 ___9__437324(.DIN1 (_________32876), .DIN2 (_____9___33022),
       .Q (______9__32917));
  dffacs1 _________________0_437325(.CLRB (reset), .CLK (clk), .DIN
       (_________32896), .QN
       (_______________0_____________________18833));
  dffacs1 _________________9_437326(.CLRB (reset), .CLK (clk), .DIN
       (______9__32889), .QN (_____________9___18751));
  nor2s1 ___9__437327(.DIN1 (_________32884), .DIN2 (_________32903),
       .Q (_________32904));
  xor2s1 ___9___437328(.DIN1 (_________32894), .DIN2 (_________32901),
       .Q (_________32902));
  xnr2s1 ___9___437329(.DIN1 (____0_0__34598), .DIN2 (______9__28849),
       .Q (_________32906));
  nnd2s1 ___9___437330(.DIN1 (______0__32899), .DIN2 (______9__32880),
       .Q (_________32900));
  nor2s1 ___9__437331(.DIN1 (_________32419), .DIN2 (_________32878),
       .Q (______9__32898));
  nor2s1 ___9__437332(.DIN1 (_________32879), .DIN2 (_________31923),
       .Q (_________32912));
  nor2s1 ___9___437333(.DIN1 (_________32862), .DIN2 (_________32886),
       .Q (_________32916));
  and2s1 ___9___437334(.DIN1 (________22246), .DIN2 (_________34443),
       .Q (_________32897));
  nnd2s1 ___9___437335(.DIN1 (______0__32873), .DIN2 (_________32874),
       .Q (_________32896));
  and2s1 ___9___437336(.DIN1 (_________32894), .DIN2 (_____99__31353),
       .Q (_________32895));
  or2s1 ___9__437337(.DIN1 (_____9___28702), .DIN2 (____0_0__34598), .Q
       (_________32893));
  nnd2s1 ___9___437338(.DIN1 (______9__32927), .DIN2 (_________32870),
       .Q (_________32892));
  nor2s1 ___9___437339(.DIN1 (_________34443), .DIN2 (________22745),
       .Q (_________32891));
  xor2s1 ___9___437340(.DIN1 (_________32882), .DIN2 (_________32883),
       .Q (______0__32890));
  nnd2s1 ___9___437341(.DIN1 (_________32868), .DIN2 (________21870),
       .Q (______9__32889));
  or2s1 ___9___437342(.DIN1 (______0__33058), .DIN2 (_________32869),
       .Q (_________32888));
  nnd2s1 ___9___437343(.DIN1 (_________29854), .DIN2 (_________34443),
       .Q (_________32887));
  xor2s1 ___9___437344(.DIN1 (_________32423), .DIN2 (_________32877),
       .Q (_________32885));
  nor2s1 ___9___437345(.DIN1 (____0____34600), .DIN2 (_________31924),
       .Q (_________32911));
  nnd2s1 ___9___437346(.DIN1 (_________34443), .DIN2 (____90___29904),
       .Q (_________32960));
  dffacs1 ___________________437347(.CLRB (reset), .CLK (clk), .DIN
       (_________32875), .Q (_________18845));
  nor2s1 ___9___437348(.DIN1 (_________32883), .DIN2 (_________32882),
       .Q (_________32884));
  and2s1 ___9___437349(.DIN1 (_________32882), .DIN2 (_________32883),
       .Q (______0__32881));
  hi1s1 ___9___437350(.DIN (_________34443), .Q (______9__32880));
  hi1s1 ___9___437351(.DIN (____0____34600), .Q (_________32879));
  nor2s1 ___9__437352(.DIN1 (_________32421), .DIN2 (_________32877),
       .Q (_________32878));
  nnd2s1 ___9__437353(.DIN1 (_________32867), .DIN2 (____00___34532),
       .Q (_________32876));
  xor2s1 ___9___437354(.DIN1 (____000__34531), .DIN2 (________21041),
       .Q (_________32886));
  nnd2s1 ___9__437355(.DIN1 (_________32864), .DIN2 (_________32874),
       .Q (_________32875));
  nor2s1 ___9__437356(.DIN1 (______0__32863), .DIN2 (____9____32700),
       .Q (______0__32873));
  xnr2s1 ___9___437357(.DIN1 (______9__32872), .DIN2 (_________32871),
       .Q (_________32894));
  dffacs1 ___________________437358(.CLRB (reset), .CLK (clk), .DIN
       (_________32865), .QN (_________34443));
  xor2s1 ___9___437359(.DIN1 (_________32859), .DIN2 (____0_0__32830),
       .Q (_________32870));
  xor2s1 ___9___437360(.DIN1 (_________32588), .DIN2 (_________32866),
       .Q (_________32869));
  or2s1 ___9__437361(.DIN1 (______9__32927), .DIN2 (_________32860), .Q
       (_________32868));
  dffacs1 ___________________437362(.CLRB (reset), .CLK (clk), .DIN
       (_________32861), .QN (_________18856));
  xor2s1 ___9___437363(.DIN1 (_____0___32855), .DIN2 (____0____32837),
       .Q (_________32883));
  nnd2s1 ___9___437364(.DIN1 (_________32866), .DIN2 (_________32587),
       .Q (_________32867));
  nor2s1 ___9_9_437365(.DIN1 (_________32362), .DIN2 (_________32858),
       .Q (_________32877));
  nnd2s1 ___9___437366(.DIN1 (_____09__32856), .DIN2 (________22746),
       .Q (_________32865));
  and2s1 ___9___437367(.DIN1 (____099__32848), .DIN2 (_____0___32853),
       .Q (_________32864));
  nor2s1 ___9___437368(.DIN1 (_____0___32854), .DIN2 (____00___32758),
       .Q (______0__32863));
  nnd2s1 ___9___437369(.DIN1 (_____0___32852), .DIN2 (________22636),
       .Q (_________32861));
  xor2s1 ___9_9_437370(.DIN1 (_________32363), .DIN2 (______0__32857),
       .Q (_________32860));
  xor2s1 ___9___437371(.DIN1 (____090__32840), .DIN2 (____0____32826),
       .Q (_________32871));
  nnd2s1 ___9_9_437372(.DIN1 (____09___32845), .DIN2 (____0____32827),
       .Q (_________32862));
  xor2s1 ___9_9_437373(.DIN1 (_________18855), .DIN2 (______9__34450),
       .Q (_________32859));
  nor2s1 ___9_437374(.DIN1 (_________32361), .DIN2 (______0__32857), .Q
       (_________32858));
  nnd2s1 ___9_99(.DIN1 (____09___32846), .DIN2 (______9__32636), .Q
       (_________32866));
  nnd2s1 ___9___437375(.DIN1 (____09___32844), .DIN2 (____0____32793),
       .Q (_____09__32856));
  xor2s1 ___9___437376(.DIN1 (____0____32832), .DIN2 (____0____32816),
       .Q (_____0___32855));
  xor2s1 ___9___437377(.DIN1 (____0____32831), .DIN2 (____99___32748),
       .Q (_____0___32854));
  nnd2s1 ___9___437378(.DIN1 (____0_9__32819), .DIN2 (____09___32843),
       .Q (_____0___32853));
  or2s1 ___9_0_437379(.DIN1 (______9__32927), .DIN2 (____0____32838),
       .Q (_____0___32852));
  nor2s1 ___9___437380(.DIN1 (______9__34450), .DIN2 (____9_0__31767),
       .Q (_____00__32849));
  dffacs1 ___________________437381(.CLRB (reset), .CLK (clk), .DIN
       (____09___32841), .QN (_______________0__________________));
  nor2s1 ___9___437382(.DIN1 (____0____32833), .DIN2 (____0_0__32820),
       .Q (____099__32848));
  or2s1 ___9_0_437383(.DIN1 (______9__32927), .DIN2 (____0____32824),
       .Q (____09___32847));
  nnd2s1 ___9_0_437384(.DIN1 (____0_9__32829), .DIN2 (_________32625),
       .Q (____09___32846));
  nnd2s1 ___9___437385(.DIN1 (____0_9__32839), .DIN2 (____0____32825),
       .Q (____09___32845));
  nor2s1 ___9___437386(.DIN1 (_________32334), .DIN2 (____0____32822),
       .Q (______0__32857));
  xor2s1 ___9___437387(.DIN1 (____0____32828), .DIN2 (_________32635),
       .Q (____09___32844));
  nor2s1 ___9_0_437388(.DIN1 (____09___32842), .DIN2 (___0____22594),
       .Q (____09___32843));
  nnd2s1 ___9_9_437389(.DIN1 (____0____32818), .DIN2 (_________32874),
       .Q (____09___32841));
  xor2s1 ___9___437390(.DIN1 (_________________18750), .DIN2
       (____0_9__32839), .Q (____090__32840));
  xor2s1 ___9___437391(.DIN1 (_________32342), .DIN2 (____0____32821),
       .Q (____0____32838));
  and2s1 ___9___437392(.DIN1 (____0____32837), .DIN2 (____0____32817),
       .Q (_____0___32850));
  dffacs1 ___________________437393(.CLRB (reset), .CLK (clk), .DIN
       (____0____32815), .Q (______9__34450));
  dffacs1 ___________________437394(.CLRB (reset), .CLK (clk), .DIN
       (____0____32814), .QN (________18841));
  and2s1 ___9__437395(.DIN1 (____0____32835), .DIN2
       (_______________0_____________________18832), .Q
       (____0____32836));
  nor2s1 ___9_437396(.DIN1
       (_______________0_____________________18832), .DIN2
       (____0____32835), .Q (____0____32834));
  nor2s1 ___9_0_437397(.DIN1
       (_______________0_____________________18832), .DIN2
       (____0_0__32780), .Q (____0____32833));
  xor2s1 ___9___437398(.DIN1 (________________18770), .DIN2
       (_________31667), .Q (____0____32832));
  xor2s1 ___9___437399(.DIN1 (________________18770), .DIN2
       (____________9___18773), .Q (____0____32831));
  dffacs1 ___________________437400(.CLRB (reset), .CLK (clk), .DIN
       (____0_0__32810), .Q (______0__18842));
  nor2s1 ___9___437401(.DIN1 (_________31917), .DIN2
       (_________________18750), .Q (____0_0__32830));
  nnd2s1 ___9__437402(.DIN1 (____0____32828), .DIN2 (______0__32621),
       .Q (____0_9__32829));
  or2s1 ___9__437403(.DIN1 (_________________18750), .DIN2
       (____0____32826), .Q (____0____32827));
  nnd2s1 ___9___437404(.DIN1 (____0____32826), .DIN2
       (_________________18750), .Q (____0____32825));
  xor2s1 ___9___437405(.DIN1 (____0____32801), .DIN2 (____0____32823),
       .Q (____0____32824));
  nor2s1 ___9___437406(.DIN1 (_________32338), .DIN2 (____0____32821),
       .Q (____0____32822));
  nor2s1 ___9_0_437407(.DIN1 (____0_9__32819), .DIN2 (____0____32806),
       .Q (____0_0__32820));
  and2s1 ___9_0_437408(.DIN1 (____0____32805), .DIN2 (________22667),
       .Q (____0____32818));
  nnd2s1 ___9___437409(.DIN1 (____0____32816), .DIN2
       (________________18770), .Q (____0____32817));
  hi1s1 ___9__437410(.DIN (_______________0_____________________18832),
       .Q (____09___32842));
  nnd2s1 ___9__437411(.DIN1 (____0____32802), .DIN2 (_________32407),
       .Q (____0____32815));
  nnd2s1 ___9__437412(.DIN1 (____9_9__32704), .DIN2 (____0____32803),
       .Q (____0____32814));
  or2s1 ___9___437413(.DIN1 (________________18770), .DIN2
       (____0____32816), .Q (____0____32813));
  nnd2s1 ___9___437414(.DIN1 (____0____32808), .DIN2 (____0____32811),
       .Q (____0____32812));
  nnd2s1 ___9__437415(.DIN1 (____0_9__32799), .DIN2 (____9_0__32685),
       .Q (____0_0__32810));
  nor2s1 ___9___437416(.DIN1 (_________29724), .DIN2 (____0____32798),
       .Q (_________32962));
  dffacs1 ___________________437417(.CLRB (reset), .CLK (clk), .DIN
       (____0_0__32800), .Q
       (_______________0_____________________18832));
  hi1s1 ___9___437418(.DIN (____0____32808), .Q (____0_9__32809));
  nor2s1 ___9___437419(.DIN1 (_________32327), .DIN2 (____0_9__32789),
       .Q (____0____32821));
  xor2s1 ___9__437420(.DIN1 (____0____32782), .DIN2 (____0____32807),
       .Q (____0____32828));
  dffacs1 ___________________437421(.CLRB (reset), .CLK (clk), .DIN
       (____0_0__32790), .QN (_________________18750));
  xor2s1 ___9___437422(.DIN1 (____0____32797), .DIN2 (_________29725),
       .Q (____0____32806));
  nor2s1 ___9___437423(.DIN1 (________23246), .DIN2 (____0____32786),
       .Q (____0____32805));
  xor2s1 ___9___437424(.DIN1 (____0____32795), .DIN2 (____99___30900),
       .Q (____0____32804));
  dffacs1 __________________437425(.CLRB (reset), .CLK (clk), .DIN
       (____0____32785), .QN (________________18770));
  nnd2s1 ___9___437426(.DIN1 (____9____32723), .DIN2 (____0____32784),
       .Q (____0____32803));
  nor2s1 ___9___437427(.DIN1 (____99__20419), .DIN2 (____0____32783),
       .Q (____0____32802));
  xor2s1 ___9___437428(.DIN1 (_________32328), .DIN2 (____0____32788),
       .Q (____0____32801));
  xor2s1 ___9___437429(.DIN1 (____0____32776), .DIN2 (______0__34988),
       .Q (____0____32808));
  dffacs1 ___________________437430(.CLRB (reset), .CLK (clk), .DIN
       (____0____32787), .Q (_______________0___________________));
  nnd2s1 ___9___437431(.DIN1 (____0____32781), .DIN2 (_________32874),
       .Q (____0_0__32800));
  nor2s1 ___9___437432(.DIN1 (____9_0__32705), .DIN2 (____0_9__32779),
       .Q (____0_9__32799));
  and2s1 ___9___437433(.DIN1 (____0____32797), .DIN2 (_________29683),
       .Q (____0____32798));
  nor2s1 ___9___437434(.DIN1 (____0____32791), .DIN2 (____0____32795),
       .Q (____0____32796));
  nnd2s1 ___9___437435(.DIN1 (____0____32775), .DIN2 (____0____32793),
       .Q (____0____32794));
  nnd2s1 ___9___437436(.DIN1 (____0____32795), .DIN2 (____0____32791),
       .Q (____0____32792));
  nor2s1 ___9__437437(.DIN1 (_________33370), .DIN2 (____0____32778),
       .Q (____0_0__32790));
  nor2s1 ___9___437438(.DIN1 (_________32326), .DIN2 (____0____32788),
       .Q (____0_9__32789));
  nnd2s1 ___9___437439(.DIN1 (____0____32772), .DIN2 (_________32874),
       .Q (____0____32787));
  nor2s1 ___9___437440(.DIN1 (____0_9__32819), .DIN2 (____0____32771),
       .Q (____0____32786));
  nnd2s1 ___9___437441(.DIN1 (_________31614), .DIN2 (____0_0__32770),
       .Q (____0____32785));
  nnd2s1 ___9___437442(.DIN1 (____0_9__32769), .DIN2 (inData[26]), .Q
       (____0____32784));
  nor2s1 ___9__437443(.DIN1 (______9__32927), .DIN2 (____0____32767),
       .Q (____0____32783));
  nor2s1 ___9___437444(.DIN1 (_____9___32561), .DIN2 (____0____32768),
       .Q (____0____32782));
  and2s1 ___9___437445(.DIN1 (____0____32764), .DIN2 (____0_0__32780),
       .Q (____0____32781));
  and2s1 ___9__437446(.DIN1 (____0____32763), .DIN2 (____0____32793),
       .Q (____0_9__32779));
  xor2s1 ___9___437447(.DIN1 (____00___32754), .DIN2 (____0____32777),
       .Q (____0____32778));
  nnd2s1 ___9___437448(.DIN1 (____0____32766), .DIN2 (_________29492),
       .Q (____0____32797));
  or2s1 ___9___437449(.DIN1 (____0____32773), .DIN2 (____0____32774),
       .Q (____0____32776));
  xor2s1 ___9___437450(.DIN1 (_____9___32567), .DIN2 (____0____34602),
       .Q (____0____32775));
  nnd2s1 ___9___437451(.DIN1 (____0____32774), .DIN2 (____0____32773),
       .Q (____0____32811));
  nor2s1 ___9___437452(.DIN1 (______0__32302), .DIN2 (____0_0__32761),
       .Q (____0____32788));
  xor2s1 ___9___437453(.DIN1 (____00___32755), .DIN2 (____0____30938),
       .Q (____0____32795));
  and2s1 ___9___437454(.DIN1 (____00___32759), .DIN2 (________22726),
       .Q (____0____32772));
  xor2s1 ___9__437455(.DIN1 (_____9___29528), .DIN2 (____0____32765),
       .Q (____0____32771));
  nnd2s1 ___9__437456(.DIN1 (____9____32719), .DIN2 (____00___32757),
       .Q (____0_0__32770));
  nor2s1 ___9__437457(.DIN1 (____00___32756), .DIN2 (____9____32697),
       .Q (____0_9__32769));
  nor2s1 ___9__437458(.DIN1 (_____9___32566), .DIN2 (____0____34602),
       .Q (____0____32768));
  xor2s1 ___9___437459(.DIN1 (_________32308), .DIN2 (____009__32760),
       .Q (____0____32767));
  or2s1 ___9___437460(.DIN1 (_________29490), .DIN2 (____0____32765),
       .Q (____0____32766));
  and2s1 ___9___437461(.DIN1 (____00___32753), .DIN2 (________22752),
       .Q (____0____32764));
  xor2s1 ___9___437462(.DIN1 (____99___32745), .DIN2 (____0____32762),
       .Q (____0____32763));
  nor2s1 ___9___437463(.DIN1 (_____0___32298), .DIN2 (____009__32760),
       .Q (____0_0__32761));
  nnd2s1 ___9_437464(.DIN1 (____99___32747), .DIN2 (____0____30939), .Q
       (____0____32773));
  nnd2s1 ___9___437465(.DIN1 (____99___32746), .DIN2 (____00___32758),
       .Q (____00___32759));
  xor2s1 ___9___437466(.DIN1 (____________9___18773), .DIN2
       (________________18772), .Q (____00___32757));
  xor2s1 ___9_9_437467(.DIN1 (________18840), .DIN2 (____9____32691),
       .Q (____00___32756));
  xor2s1 ___9_9_437468(.DIN1 (________18840), .DIN2 (_________31978),
       .Q (____00___32755));
  xor2s1 ___9_9_437469(.DIN1 (______9__34460), .DIN2 (____9_9__32742),
       .Q (____00___32754));
  nnd2s1 ___9___437470(.DIN1 (____99___32744), .DIN2 (____00___32758),
       .Q (____00___32753));
  nor2s1 ___9__437471(.DIN1 (________________18772), .DIN2
       (____99___32749), .Q (____00___32752));
  xor2s1 ___9___437472(.DIN1 (____9____32736), .DIN2 (____000__32751),
       .Q (____0____32765));
  nnd2s1 ___9_9_437473(.DIN1 (____99___32749), .DIN2
       (________________18772), .Q (____999__32750));
  nor2s1 ___9_9_437474(.DIN1 (_____0___29362), .DIN2
       (________________18772), .Q (____99___32748));
  nnd2s1 ___9_0_437475(.DIN1 (_____0___31000), .DIN2 (________18840),
       .Q (____99___32747));
  nor2s1 ___9_437476(.DIN1 (____9____32740), .DIN2 (____990__32743), .Q
       (____009__32760));
  xor2s1 ___9___437477(.DIN1 (____9____32732), .DIN2 (_________32049),
       .Q (____99___32746));
  xor2s1 ___9_9_437478(.DIN1 (____9____32731), .DIN2 (_________32494),
       .Q (____99___32745));
  dffacs1 ___________________437479(.CLRB (reset), .CLK (clk), .DIN
       (____9____32735), .QN (_________________18749));
  xor2s1 ___9_9_437480(.DIN1 (____9_0__32725), .DIN2 (____99___35108),
       .Q (____99___32744));
  nor2s1 ___9_0_437481(.DIN1 (______9__34460), .DIN2 (____9____32741),
       .Q (____990__32743));
  dffacs1 __________________437482(.CLRB (reset), .CLK (clk), .DIN
       (____9____32733), .QN (________________18772));
  nor2s1 ___9_437483(.DIN1 (____9____32741), .DIN2 (____9____32740), .Q
       (____9_9__32742));
  nnd2s1 ___9___437484(.DIN1 (____9____32738), .DIN2 (____9____32737),
       .Q (____9____32739));
  dffacs1 _________________0_437485(.CLRB (reset), .CLK (clk), .DIN
       (____9____32730), .QN (________18840));
  nnd2s1 ___9_0_437486(.DIN1 (____9____32727), .DIN2 (_________29430),
       .Q (____9____32736));
  nnd2s1 ___9_0_437487(.DIN1 (____9_9__32724), .DIN2 (____0____29099),
       .Q (____9____32735));
  nnd2s1 ___9___437488(.DIN1 (_________32622), .DIN2 (____9____32720),
       .Q (____9____32733));
  xor2s1 ___9_0_437489(.DIN1 (_________29493), .DIN2 (____9____32726),
       .Q (____9____32732));
  xor2s1 ___9___437490(.DIN1 (_________30261), .DIN2 (____9____32722),
       .Q (____9____32731));
  dffacs1 ___________________437491(.CLRB (reset), .CLK (clk), .DIN
       (____9____32721), .QN (_________________18761));
  nnd2s1 ___9___437492(.DIN1 (_________32629), .DIN2 (____9____32717),
       .Q (____9____32730));
  nor2s1 ___9__437493(.DIN1 (____9____32729), .DIN2 (____0_9__32839),
       .Q (____9____32741));
  and2s1 ___9___437494(.DIN1 (____0_9__32839), .DIN2 (____9____32729),
       .Q (____9____32740));
  xor2s1 ___9___437495(.DIN1 (____9_9__32714), .DIN2 (____9____32728),
       .Q (____9____32738));
  nnd2s1 ___9_0_437496(.DIN1 (____9____32726), .DIN2 (_________29427),
       .Q (____9____32727));
  xor2s1 ___9___437497(.DIN1 (____9____32712), .DIN2 (____9____32693),
       .Q (____9_0__32725));
  or2s1 ___9___437498(.DIN1 (____9____32723), .DIN2 (____9____32716),
       .Q (____9_9__32724));
  nor2s1 ___9__437499(.DIN1 (_________32491), .DIN2 (____9____32722),
       .Q (____9_9__32734));
  dffacs1 ___________________437500(.CLRB (reset), .CLK (clk), .DIN
       (____9_0__32715), .QN (_________________18748));
  nnd2s1 ___9___437501(.DIN1 (____9____32713), .DIN2 (____0___22173),
       .Q (____9____32721));
  nnd2s1 ___9___437502(.DIN1 (____9____32719), .DIN2 (____9____32718),
       .Q (____9____32720));
  nnd2s1 ___9__437503(.DIN1 (____9____32723), .DIN2 (____9____32711),
       .Q (____9____32717));
  and2s1 ___9___437504(.DIN1 (____9____32710), .DIN2 (_________32238),
       .Q (____9____32729));
  nor2s1 ___9___437505(.DIN1 (____9_9__32694), .DIN2 (____9____32708),
       .Q (____9____32726));
  nor2s1 ___9___437506(.DIN1 (_________32525), .DIN2 (____9____32703),
       .Q (____9____32722));
  xor2s1 ___9___437507(.DIN1 (_________32240), .DIN2 (____9____32709),
       .Q (____9____32716));
  nnd2s1 ___9___437508(.DIN1 (____9____32671), .DIN2 (____9____32706),
       .Q (____9_0__32715));
  nnd2s1 ___9___437509(.DIN1 (______9__31409), .DIN2 (____9____32702),
       .Q (____9_9__32714));
  nnd2s1 ___9___437510(.DIN1 (____9____32699), .DIN2 (____0____32793),
       .Q (____9____32713));
  xor2s1 ___9__437511(.DIN1 (_________________18760), .DIN2
       (____9____32707), .Q (____9____32712));
  hi1s1 ___9__437512(.DIN (____________9___18773), .Q (____9____32718));
  nnd2s1 ___9___437513(.DIN1 (____9____32698), .DIN2 (inData[10]), .Q
       (____9____32711));
  nnd2s1 ___9___437514(.DIN1 (____9____32709), .DIN2 (_________32239),
       .Q (____9____32710));
  nnd2s1 ___9___437515(.DIN1 (______0__31410), .DIN2 (____9____32701),
       .Q (____9____32737));
  nor2s1 ___9___437516(.DIN1 (____9____32687), .DIN2 (____9____32707),
       .Q (____9____32708));
  nnd2s1 ___9__437517(.DIN1 (____0____29098), .DIN2 (____9____32692),
       .Q (____9____32706));
  nor2s1 ___9___437518(.DIN1 (____9____32696), .DIN2 (____0____32793),
       .Q (____9_0__32705));
  dffacs1 ________________9_437519(.CLRB (reset), .CLK (clk), .DIN
       (____9_0__32695), .QN (____________9___18773));
  or2s1 ___9__437520(.DIN1 (____9____32723), .DIN2 (____9____32690), .Q
       (____9_9__32704));
  nor2s1 ___9___437521(.DIN1 (_________________0___18633), .DIN2
       (____9____32689), .Q (____9____32703));
  hi1s1 ___9__437522(.DIN (____9____32701), .Q (____9____32702));
  xor2s1 ___9___437523(.DIN1 (____9____32678), .DIN2 (____9____32681),
       .Q (____0____32774));
  nor2s1 ___9___437524(.DIN1 (____0_9__32819), .DIN2 (____9_9__32684),
       .Q (____9____32700));
  xnr2s1 ___9___437525(.DIN1 (____9____32688), .DIN2 (____0____34610),
       .Q (____9____32699));
  nor2s1 ___9___437526(.DIN1 (______9__31379), .DIN2 (____9____32680),
       .Q (____9____32709));
  nor2s1 ___9___437527(.DIN1 (____9____32683), .DIN2 (____9____32697),
       .Q (____9____32698));
  nnd2s1 ___9___437528(.DIN1 (____9____32682), .DIN2 (____9____32677),
       .Q (____9____32701));
  dffacs1 ___________________437529(.CLRB (reset), .CLK (clk), .DIN
       (____9____32686), .QN (_________34444));
  xor2s1 ___9___437530(.DIN1 (_________________18760), .DIN2
       (________19636), .Q (____9____32696));
  nnd2s1 ___9___437531(.DIN1 (____9_9__32674), .DIN2 (___9____23364),
       .Q (____9_0__32695));
  nor2s1 ___9__437532(.DIN1 (____9_0__32675), .DIN2 (____9____32693),
       .Q (____9_9__32694));
  xnr2s1 ___9___437533(.DIN1 (________18841), .DIN2 (____9____32691),
       .Q (____9____32692));
  xor2s1 ___9___437534(.DIN1 (_________31406), .DIN2 (____9____32679),
       .Q (____9____32690));
  nnd2s1 ___9___437535(.DIN1 (____9____32688), .DIN2 (_________32508),
       .Q (____9____32689));
  nor2s1 ___9___437536(.DIN1 (_________29327), .DIN2 (____9____32673),
       .Q (____9____32707));
  nor2s1 ___9___437537(.DIN1 (_________________18760), .DIN2
       (_________30531), .Q (____9____32687));
  nnd2s1 ___9___437538(.DIN1 (____9____32669), .DIN2 (____9_0__32685),
       .Q (____9____32686));
  xor2s1 ___9___437539(.DIN1 (____9____32672), .DIN2 (_________29328),
       .Q (____9_9__32684));
  nnd2s1 ___9___437540(.DIN1 (____9____32691), .DIN2 (____9____32670),
       .Q (____9____32683));
  nnd2s1 ___9___437541(.DIN1 (____9____32676), .DIN2 (____9____32681),
       .Q (____9____32682));
  nor2s1 ___9___437542(.DIN1 (____9____32679), .DIN2 (_________31378),
       .Q (____9____32680));
  and2s1 ___9___437543(.DIN1 (____9____32677), .DIN2 (____9____32676),
       .Q (____9____32678));
  hi1s1 ___9___437544(.DIN (_________________18760), .Q
       (____9_0__32675));
  nnd2s1 ___9___437545(.DIN1 (____9____32667), .DIN2 (____00___32758),
       .Q (____9_9__32674));
  and2s1 ___9__437546(.DIN1 (______9__29300), .DIN2 (____9____32672),
       .Q (____9____32673));
  or2s1 ___9___437547(.DIN1 (____9____32723), .DIN2 (____9_0__32665),
       .Q (____9____32671));
  nnd2s1 ___9___437548(.DIN1 (____9____32666), .DIN2 (____90___32657),
       .Q (____9____32688));
  nnd2s1 ___9___437549(.DIN1 (_________________18748), .DIN2
       (_________________18747), .Q (____9____32670));
  nor2s1 ___9__437550(.DIN1 (________22843), .DIN2 (____90___32661), .Q
       (____9____32669));
  nnd2s1 ___9__437551(.DIN1 (____90___32660), .DIN2 (_________31311),
       .Q (____9____32679));
  dffacs1 ___________________437552(.CLRB (reset), .CLK (clk), .DIN
       (____909__32664), .Q (_________________18760));
  or2s1 ___9___437553(.DIN1 (_________________18747), .DIN2
       (____9____32668), .Q (____9____32677));
  nnd2s1 ___9___437554(.DIN1 (____9____32668), .DIN2
       (_________________18747), .Q (____9____32676));
  or2s1 ___9___437555(.DIN1 (_________________18747), .DIN2
       (_________________18748), .Q (____9____32691));
  dffacs1 __________________437556(.CLRB (reset), .CLK (clk), .DIN
       (____90___32663), .QN (_________18861));
  xor2s1 ___9___437557(.DIN1 (____9__19036), .DIN2 (_____9___32651), .Q
       (____9____32667));
  nnd2s1 ___9___437558(.DIN1 (____90___32658), .DIN2 (_____9___32648),
       .Q (____9____32672));
  nor2s1 ___9___437559(.DIN1 (____0____30053), .DIN2 (____900__32656),
       .Q (____9____32666));
  xor2s1 ___9___437560(.DIN1 (_________31319), .DIN2 (____90___32659),
       .Q (____9_0__32665));
  nnd2s1 ___9___437561(.DIN1 (_____9___32654), .DIN2 (____9___22802),
       .Q (____909__32664));
  nnd2s1 ___9__437562(.DIN1 (_____9___32653), .DIN2 (____90___32662),
       .Q (____90___32663));
  and2s1 ___9___437563(.DIN1 (_____9___32652), .DIN2 (____0____32793),
       .Q (____90___32661));
  nnd2s1 ___9_437564(.DIN1 (______0__31293), .DIN2 (____90___32659), .Q
       (____90___32660));
  dffacs1 ___________________437565(.CLRB (reset), .CLK (clk), .DIN
       (_____9___32649), .QN (_________________18747));
  or2s1 ___9__437566(.DIN1 (_____9___32650), .DIN2 (_____90__32646), .Q
       (____90___32658));
  nnd2s1 ___9_9_437567(.DIN1 (_____99__32655), .DIN2 (_________35110),
       .Q (____90___32657));
  nor2s1 ___9_9_437568(.DIN1 (_________31431), .DIN2 (_____99__32655),
       .Q (____900__32656));
  nnd2s1 ___9___437569(.DIN1 (_________32645), .DIN2 (____0____32793),
       .Q (_____9___32654));
  nor2s1 ___9_9_437570(.DIN1 (_________29876), .DIN2 (_________32643),
       .Q (_____9___32653));
  xor2s1 ___9_9_437571(.DIN1 (____0_9__30055), .DIN2 (____0____34604),
       .Q (_____9___32652));
  xor2s1 ___9_9_437572(.DIN1 (_____9___32647), .DIN2 (_____9___32650),
       .Q (_____9___32651));
  nnd2s1 ___9_9_437573(.DIN1 (_________32641), .DIN2 (_________35096),
       .Q (_____9___32649));
  nnd2s1 ___9_437574(.DIN1 (_________32642), .DIN2 (_________31198), .Q
       (____90___32659));
  or2s1 ___9_437575(.DIN1 (____________9___18758), .DIN2
       (_____9___32647), .Q (_____9___32648));
  and2s1 ___9_0_437576(.DIN1 (_____9___32647), .DIN2
       (____________9___18758), .Q (_____90__32646));
  nor2s1 ___9_0_437577(.DIN1 (____0____30054), .DIN2 (____0____34604),
       .Q (_____99__32655));
  xor2s1 ___9_9_437578(.DIN1 (_________32634), .DIN2 (_________32644),
       .Q (_________32645));
  nnd2s1 ___9_0_437579(.DIN1 (_________32640), .DIN2 (_________29786),
       .Q (_________32643));
  xor2s1 ___9_0_437580(.DIN1 (_________32633), .DIN2 (_________35105),
       .Q (_________32642));
  or2s1 ___9_437581(.DIN1 (____9____32723), .DIN2 (_________32638), .Q
       (_________32641));
  nor2s1 ___9_0_437582(.DIN1 (______0__32628), .DIN2 (______0__32637),
       .Q (_____9___32647));
  nnd2s1 ___9_0_437583(.DIN1 (_________32631), .DIN2 (_________32639),
       .Q (_________32640));
  xor2s1 ___9___437584(.DIN1 (_____9___34509), .DIN2 (_________32632),
       .Q (_________32638));
  dffacs1 _________________9_437585(.CLRB (reset), .CLK (clk), .DIN
       (_________32630), .QN (______0__34451));
  and2s1 ___9___437586(.DIN1 (_________32627), .DIN2 (____99___32749),
       .Q (______0__32637));
  or2s1 ___9_0_437587(.DIN1 (______9__32620), .DIN2 (_________32635),
       .Q (______9__32636));
  xor2s1 ___9__437588(.DIN1 (_________32618), .DIN2 (_________32446),
       .Q (_________32634));
  nor2s1 ___9___437589(.DIN1 (_________32632), .DIN2 (_________31173),
       .Q (_________32633));
  xor2s1 ___9__437590(.DIN1 (_____9___28986), .DIN2 (____0____34606),
       .Q (_________32631));
  nnd2s1 ___9___437591(.DIN1 (_________32619), .DIN2 (_____0___32574),
       .Q (_________32630));
  or2s1 ___9__437592(.DIN1 (____9____32723), .DIN2 (_________32616), .Q
       (_________32629));
  dffacs1 _________________0_437593(.CLRB (reset), .CLK (clk), .DIN
       (_________32617), .QN (_____________0___18759));
  nor2s1 ___9___437594(.DIN1 (_________32626), .DIN2 (____0____34606),
       .Q (______0__32628));
  nnd2s1 ___9___437595(.DIN1 (____0____34606), .DIN2 (_________32626),
       .Q (_________32627));
  nnd2s1 ___9__437596(.DIN1 (_________32615), .DIN2 (_________32625),
       .Q (_________32635));
  nnd2s1 ___9___437597(.DIN1 (_________32613), .DIN2 (_________31979),
       .Q (_________32632));
  nnd2s1 ___9___437598(.DIN1 (_________32609), .DIN2 (_________33103),
       .Q (_________32622));
  nnd2s1 ___9___437599(.DIN1 (_________32614), .DIN2 (______9__32620),
       .Q (______0__32621));
  dffacs1 __________________437600(.CLRB (reset), .CLK (clk), .DIN
       (______9__32610), .QN (_________34445));
  nor2s1 ___9___437601(.DIN1 (_____0___32571), .DIN2 (_________32607),
       .Q (_________32619));
  xor2s1 ___9___437602(.DIN1 (______0__32611), .DIN2 (______0__32445),
       .Q (_________32618));
  nnd2s1 ___9___437603(.DIN1 (_________32608), .DIN2 (_________32590),
       .Q (_________32617));
  xor2s1 ___9__437604(.DIN1 (____00___34535), .DIN2 (_________32612),
       .Q (_________32616));
  hi1s1 ___9___437605(.DIN (_________32614), .Q (_________32615));
  nnd2s1 ___9___437606(.DIN1 (_________32612), .DIN2 (______0__31977),
       .Q (_________32613));
  nor2s1 ___9___437607(.DIN1 (_________32447), .DIN2 (______0__32611),
       .Q (_________32623));
  nnd2s1 ___9___437608(.DIN1 (_________32605), .DIN2 (____0___23718),
       .Q (______9__32610));
  xor2s1 ___9___437609(.DIN1 (_________32599), .DIN2 (_____0___32851),
       .Q (_________32609));
  dffacs1 ________________9_437610(.CLRB (reset), .CLK (clk), .DIN
       (_________32603), .QN (____________9___18758));
  nnd2s1 ___9__437611(.DIN1 (______0__32602), .DIN2 (_________32604),
       .Q (_________32608));
  nor2s1 ___9___437612(.DIN1 (_____0___32572), .DIN2 (______9__32601),
       .Q (_________32607));
  xor2s1 ___9___437613(.DIN1 (_________32600), .DIN2 (_________32606),
       .Q (_________32614));
  nor2s1 ___9___437614(.DIN1 (_________32464), .DIN2 (_________32596),
       .Q (______0__32611));
  nor2s1 ___9___437615(.DIN1 (____99___30902), .DIN2 (_________32592),
       .Q (_________32612));
  nnd2s1 ___9___437616(.DIN1 (_________32591), .DIN2 (_________32604),
       .Q (_________32605));
  nnd2s1 ___9___437617(.DIN1 (_________32589), .DIN2 (________24577),
       .Q (_________32603));
  xor2s1 ___9___437618(.DIN1 (_________32467), .DIN2 (_________32595),
       .Q (______0__32602));
  xor2s1 ___9___437619(.DIN1 (____99___30904), .DIN2 (____0_0__34608),
       .Q (______9__32601));
  nor2s1 ___9__437620(.DIN1 (_________32597), .DIN2 (_________32598),
       .Q (_________32600));
  xor2s1 ___9__437621(.DIN1 (_________32584), .DIN2 (_________32946),
       .Q (_________32599));
  nnd2s1 ___9___437622(.DIN1 (_________32598), .DIN2 (_________32597),
       .Q (_________32625));
  nor2s1 ___9___437623(.DIN1 (_________32462), .DIN2 (_________32595),
       .Q (_________32596));
  nor2s1 ___9__437624(.DIN1 (____0_0__34608), .DIN2 (____99___30903),
       .Q (_________32592));
  xor2s1 ___9___437625(.DIN1 (_________32581), .DIN2 (____0____30044),
       .Q (_________32591));
  dffacs1 ___________________437626(.CLRB (reset), .CLK (clk), .DIN
       (_________32582), .QN (_________________18746));
  nnd2s1 ___9___437627(.DIN1 (_________31261), .DIN2 (______0__32586),
       .Q (_________32590));
  nnd2s1 ___9___437628(.DIN1 (______9__32585), .DIN2 (_________32604),
       .Q (_________32589));
  xor2s1 ___9__437629(.DIN1 (_____09__32576), .DIN2 (______9__32514),
       .Q (_________32598));
  nor2s1 ___9___437630(.DIN1 (_________32577), .DIN2 (_________32583),
       .Q (______9__32593));
  and2s1 ___9___437631(.DIN1 (_________32587), .DIN2 (____00___34532),
       .Q (_________32588));
  nor2s1 ___9___437632(.DIN1 (_____9___32470), .DIN2 (_________32580),
       .Q (_________32595));
  xor2s1 ___9___437633(.DIN1 (_________34445), .DIN2 (_________34446),
       .Q (______0__32586));
  dffacs1 ___________________437634(.CLRB (reset), .CLK (clk), .DIN
       (_____0___32575), .QN (_________34452));
  xor2s1 ___9___437635(.DIN1 (______9__34507), .DIN2 (_________32579),
       .Q (______9__32585));
  xor2s1 ___9___437636(.DIN1 (_________34446), .DIN2 (_________32583),
       .Q (_________32584));
  nnd2s1 ___9___437637(.DIN1 (_____0___32573), .DIN2 (________22294),
       .Q (_________32582));
  xor2s1 ___9___437638(.DIN1 (_____9___32564), .DIN2 (______0__32486),
       .Q (_________32581));
  nor2s1 ___9__437639(.DIN1 (_________32466), .DIN2 (_________32579),
       .Q (_________32580));
  nnd2s1 ___9___437640(.DIN1 (_________32946), .DIN2 (_________34446),
       .Q (_________32578));
  nor2s1 ___9___437641(.DIN1 (_________34446), .DIN2 (_________32946),
       .Q (_________32577));
  xor2s1 ___9___437642(.DIN1 (_________32555), .DIN2 (_____9___30449),
       .Q (_____09__32576));
  nnd2s1 ___9___437643(.DIN1 (_____9___32563), .DIN2 (_____0___32574),
       .Q (_____0___32575));
  or2s1 ___9__437644(.DIN1 (_____0___32572), .DIN2 (_____9___32562), .Q
       (_____0___32573));
  nnd2s1 ___9___437645(.DIN1 (_________30709), .DIN2 (_____9___32568),
       .Q (_________32587));
  and2s1 ___9__437646(.DIN1 (_____0___32572), .DIN2 (_________32556),
       .Q (_____0___32571));
  nnd2s1 ___9___437647(.DIN1 (_________32558), .DIN2 (_________32501),
       .Q (_________32579));
  dffacs1 __________________437648(.CLRB (reset), .CLK (clk), .DIN
       (______9__32559), .QN (_________34446));
  xor2s1 ___9___437649(.DIN1 (_____9___32565), .DIN2 (_____90__32560),
       .Q (_____9___32567));
  nor2s1 ___9___437650(.DIN1 (_____9___32565), .DIN2 (_________32552),
       .Q (_____9___32566));
  xor2s1 ___9___437651(.DIN1 (______9__32505), .DIN2 (_________32557),
       .Q (_____9___32564));
  nor2s1 ___9_437652(.DIN1 (________22794), .DIN2 (_________32551), .Q
       (_____9___32563));
  xor2s1 ___9_9_437653(.DIN1 (______0__30708), .DIN2 (_________32553),
       .Q (_____9___32562));
  nnd2s1 ___9_9_437654(.DIN1 (______0__32550), .DIN2 (_____9___30450),
       .Q (_____9___32568));
  nor2s1 ___9___437655(.DIN1 (_____09__30282), .DIN2 (_____90__32560),
       .Q (_____9___32561));
  nnd2s1 ___9_9_437656(.DIN1 (______9__32549), .DIN2 (_________34880),
       .Q (______9__32559));
  or2s1 ___9_9_437657(.DIN1 (______0__32506), .DIN2 (_________32557),
       .Q (_________32558));
  xor2s1 ___9_9_437658(.DIN1 (_________34452), .DIN2 (_________34453),
       .Q (_________32556));
  xor2s1 ___9_9_437659(.DIN1 (_________34453), .DIN2 (_________32554),
       .Q (_________32555));
  and2s1 ___9_437660(.DIN1 (_________30665), .DIN2 (_________32553), .Q
       (_____00__32569));
  hi1s1 ___9_9_437661(.DIN (_____90__32560), .Q (_________32552));
  nor2s1 ___9_0_437662(.DIN1 (_____0___32572), .DIN2 (_________32547),
       .Q (_________32551));
  or2s1 ___9_0_437663(.DIN1 (_________34453), .DIN2 (______9__30446),
       .Q (______0__32550));
  nnd2s1 ___9_0_437664(.DIN1 (_________32548), .DIN2 (_________32536),
       .Q (_________32597));
  xor2s1 ___9_437665(.DIN1 (_________32539), .DIN2 (_________32535), .Q
       (_____90__32560));
  dffacs1 ___________________437666(.CLRB (reset), .CLK (clk), .DIN
       (_________32543), .QN (_________________18744));
  nnd2s1 ___9_0_437667(.DIN1 (_________32545), .DIN2 (_________32604),
       .Q (______9__32549));
  nor2s1 ___9_0_437668(.DIN1 (______9__32540), .DIN2 (_________32546),
       .Q (_________32557));
  nnd2s1 ___9_437669(.DIN1 (_________32542), .DIN2 (_________30566), .Q
       (_________32553));
  dffacs1 ___________________437670(.CLRB (reset), .CLK (clk), .DIN
       (_________32537), .Q (_________34453));
  nnd2s1 ___9___437671(.DIN1 (_________32538), .DIN2 (_________32534),
       .Q (_________32548));
  xor2s1 ___9___437672(.DIN1 (_________30586), .DIN2 (______0__32541),
       .Q (_________32547));
  nor2s1 ___9_0_437673(.DIN1 (_________35106), .DIN2 (_________32544),
       .Q (_________32546));
  nnd2s1 ___9___437674(.DIN1 (_________32544), .DIN2 (_________32531),
       .Q (_________32545));
  nnd2s1 ___9___437675(.DIN1 (_____9___32474), .DIN2 (______9__32532),
       .Q (_________32543));
  or2s1 ___9__437676(.DIN1 (_________30565), .DIN2 (______0__32541), .Q
       (_________32542));
  nor2s1 ___9_0_437677(.DIN1 (_________________0___18633), .DIN2
       (_________32527), .Q (______9__32540));
  xor2s1 ___9___437678(.DIN1 (_________________18745), .DIN2
       (_________32538), .Q (_________32539));
  dffacs1 ___________________437679(.CLRB (reset), .CLK (clk), .DIN
       (_________32528), .QN (_________________18741));
  nnd2s1 ___9___437680(.DIN1 (_________32526), .DIN2 (_____0___32574),
       .Q (_________32537));
  nnd2s1 ___9___437681(.DIN1 (_________32535), .DIN2 (_________32533),
       .Q (_________32536));
  or2s1 ___9___437682(.DIN1 (_________32533), .DIN2 (_________32535),
       .Q (_________32534));
  or2s1 ___9___437683(.DIN1 (_________________18745), .DIN2
       (_________32487), .Q (______9__32532));
  nnd2s1 ___9___437684(.DIN1 (_________32529), .DIN2 (_________32530),
       .Q (_________32531));
  nnd2s1 ___9___437685(.DIN1 (____9____31799), .DIN2 (______0__32524),
       .Q (______0__32541));
  or2s1 ___9___437686(.DIN1 (_________32530), .DIN2 (_________32529),
       .Q (_________32544));
  nnd2s1 ___9__437687(.DIN1 (_________32422), .DIN2 (_________32522),
       .Q (_________32528));
  dffacs1 ___________________437688(.CLRB (reset), .CLK (clk), .DIN
       (_________32520), .QN (_________________18742));
  nor2s1 ___9___437689(.DIN1 (______9__32523), .DIN2 (_________32521),
       .Q (_________32527));
  nor2s1 ___9__437690(.DIN1 (________22651), .DIN2 (_________32519), .Q
       (_________32526));
  hi1s1 ___9___437691(.DIN (_________________18745), .Q
       (_________32533));
  dffacs1 ___________________437692(.CLRB (reset), .CLK (clk), .DIN
       (_________32518), .QN (_________________18745));
  nor2s1 ___9___437693(.DIN1 (_________32502), .DIN2 (______0__32515),
       .Q (______0__32524));
  or2s1 ___9___437694(.DIN1 (_________32517), .DIN2 (______9__32523),
       .Q (_________32529));
  nnd2s1 ___9__437695(.DIN1 (_________32513), .DIN2 (clk), .Q
       (_________32522));
  and2s1 ___9___437696(.DIN1 (_________32516), .DIN2 (_________32530),
       .Q (_________32521));
  nnd2s1 ___9___437697(.DIN1 (______0__32436), .DIN2 (_________32512),
       .Q (_________32520));
  nor2s1 ___9___437698(.DIN1 (_____0___32572), .DIN2 (_________32511),
       .Q (_________32519));
  nnd2s1 ___9___437699(.DIN1 (_________32489), .DIN2 (_________32507),
       .Q (_________32518));
  xor2s1 ___9___437700(.DIN1 (_________32498), .DIN2 (_________35105),
       .Q (_________32525));
  hi1s1 ___9__437701(.DIN (_________32516), .Q (_________32517));
  and2s1 ___9___437702(.DIN1 (______9__32514), .DIN2 (_________32504),
       .Q (______0__32515));
  nor2s1 ___9__437703(.DIN1 (_________32499), .DIN2 (_________32492),
       .Q (_________32513));
  nnd2s1 ___9___437704(.DIN1 (_________32509), .DIN2 (_________32510),
       .Q (_________32516));
  nnd2s1 ___9___437705(.DIN1 (_________32493), .DIN2 (inData[10]), .Q
       (_________32512));
  xor2s1 ___9__437706(.DIN1 (____99___31804), .DIN2 (_________32503),
       .Q (_________32511));
  nor2s1 ___9___437707(.DIN1 (_________32510), .DIN2 (_________32509),
       .Q (______9__32523));
  nnd2s1 ___9___437708(.DIN1 (_________32488), .DIN2 (inData[22]), .Q
       (_________32507));
  nor2s1 ___9__437709(.DIN1 (______9__32505), .DIN2 (_________32500),
       .Q (______0__32506));
  nnd2s1 ___9__437710(.DIN1 (_________32503), .DIN2 (____9____31762),
       .Q (_________32504));
  nor2s1 ___9___437711(.DIN1 (_________34462), .DIN2 (_________32503),
       .Q (_________32502));
  nnd2s1 ___9___437712(.DIN1 (_________32500), .DIN2 (______9__32505),
       .Q (_________32501));
  xor2s1 ___9___437713(.DIN1 (_____0___32481), .DIN2 (______0__32453),
       .Q (_________32499));
  or2s1 ___9___437714(.DIN1 (______0__32496), .DIN2 (_________32497),
       .Q (_________32498));
  nnd2s1 ___9__437715(.DIN1 (_________32497), .DIN2 (______0__32496),
       .Q (_________32508));
  xor2s1 ___9___437716(.DIN1 (_____0___32482), .DIN2 (____099__30093),
       .Q (_________32509));
  nnd2s1 ___9___437717(.DIN1 (_________32490), .DIN2 (_________32494),
       .Q (______9__32495));
  nor2s1 ___9___437718(.DIN1 (_____09__32485), .DIN2 (_________32492),
       .Q (_________32493));
  nor2s1 ___9___437719(.DIN1 (_________32494), .DIN2 (_________32490),
       .Q (_________32491));
  or2s1 ___9___437720(.DIN1 (_____0___32572), .DIN2 (_____0___32484),
       .Q (_________32489));
  nor2s1 ___9___437721(.DIN1 (_____0___32483), .DIN2 (_________32487),
       .Q (_________32488));
  hi1s1 ___9___437722(.DIN (______0__32486), .Q (_________32500));
  nnd2s1 ___9___437723(.DIN1 (_____0___32480), .DIN2 (_________30239),
       .Q (_________32503));
  and2s1 ___9___437724(.DIN1 (_____0___32478), .DIN2 (_____9___32472),
       .Q (_____09__32485));
  xor2s1 ___9___437725(.DIN1 (_____9___32473), .DIN2 (_________30122),
       .Q (_________32497));
  xor2s1 ___9__437726(.DIN1 (_____9___30266), .DIN2 (_____0___32479),
       .Q (_____0___32484));
  nnd2s1 ___9___437727(.DIN1 (_____99__32476), .DIN2 (_________29407),
       .Q (______0__32486));
  nnd2s1 ___9___437728(.DIN1 (_____9___32475), .DIN2 (_________30167),
       .Q (_________32494));
  xnr2s1 ___9__437729(.DIN1 (_____0___32477), .DIN2
       (_________________18742), .Q (_____0___32483));
  xor2s1 ___9___437730(.DIN1 (________________18739), .DIN2
       (_____9___29443), .Q (_____0___32482));
  xor2s1 ___9___437731(.DIN1 (________________18739), .DIN2
       (_____________0___18740), .Q (_____0___32481));
  or2s1 ___9___437732(.DIN1 (_________30240), .DIN2 (_____0___32479),
       .Q (_____0___32480));
  or2s1 ___9___437733(.DIN1 (_________________18742), .DIN2
       (_____0___32477), .Q (_____0___32478));
  or2s1 ___9___437734(.DIN1 (________________18739), .DIN2
       (_________29462), .Q (_____99__32476));
  nor2s1 ___9___437735(.DIN1 (______0__30162), .DIN2 (_____9___32471),
       .Q (_____9___32475));
  or2s1 ___9___437736(.DIN1 (_____0___32572), .DIN2 (_____9___32469),
       .Q (_____9___32474));
  xor2s1 ___9__437737(.DIN1 (_________________18743), .DIN2
       (______0__30121), .Q (_____9___32473));
  nor2s1 ___9___437738(.DIN1 (_____9___30171), .DIN2 (_____90__32468),
       .Q (_____0___32479));
  or2s1 ___9__437739(.DIN1 (_________________18743), .DIN2 (___9_), .Q
       (_____9___32472));
  nnd2s1 ___9___437740(.DIN1 (_________________18743), .DIN2
       (___0_9___27842), .Q (_____0___32477));
  dffacs1 __________________437741(.CLRB (reset), .CLK (clk), .DIN
       (_________32465), .QN (________________18739));
  nor2s1 ___9___437742(.DIN1 (_________________18743), .DIN2
       (_________30123), .Q (_____9___32471));
  xor2s1 ___9___437743(.DIN1 (_____0___30186), .DIN2 (____0____34612),
       .Q (_____9___32469));
  and2s1 ___9___437744(.DIN1 (____0____34612), .DIN2 (_____90__30170),
       .Q (_____90__32468));
  xor2s1 ___9_9_437745(.DIN1 (______0__32461), .DIN2 (_________32463),
       .Q (_________32467));
  dffacs1 ___________________437746(.CLRB (reset), .CLK (clk), .DIN
       (______9__32460), .QN (_________________18743));
  nnd2s1 ___9_9_437747(.DIN1 (_________31157), .DIN2 (_________32459),
       .Q (_________32465));
  nor2s1 ___9_9_437748(.DIN1 (_________32463), .DIN2 (_________32443),
       .Q (_________32464));
  nor2s1 ___9_9_437749(.DIN1 (_________32458), .DIN2 (______0__32461),
       .Q (_________32462));
  nnd2s1 ___9_9_437750(.DIN1 (_________32455), .DIN2 (____9___23082),
       .Q (______9__32460));
  nor2s1 ___9_9_437751(.DIN1 (_________32456), .DIN2 (_________32457),
       .Q (_________32466));
  or2s1 ___9_9_437752(.DIN1 (_________32454), .DIN2 (_________32492),
       .Q (_________32459));
  hi1s1 ___9_0_437753(.DIN (_________32458), .Q (_________32463));
  and2s1 ___9_437754(.DIN1 (_________32457), .DIN2 (_________32456), .Q
       (_____9___32470));
  nnd2s1 ___9_0_437755(.DIN1 (_________32451), .DIN2 (_________29558),
       .Q (_________32458));
  nnd2s1 ___9_0_437756(.DIN1 (_________32450), .DIN2 (_________32440),
       .Q (_________32455));
  xor2s1 ___9_0_437757(.DIN1 (_________34454), .DIN2
       (_____________0___18740), .Q (_________32454));
  xor2s1 ___9_0_437758(.DIN1 (_________29559), .DIN2 (_________34454),
       .Q (_________32457));
  nnd2s1 ___9_0_437759(.DIN1 (_________34454), .DIN2 (_________29696),
       .Q (______0__32453));
  nnd2s1 ___9_437760(.DIN1 (_____9___29530), .DIN2 (_________34454), .Q
       (_________32451));
  xor2s1 ___9__437761(.DIN1 (_________32449), .DIN2 (_________30153),
       .Q (_________32450));
  dffacs1 ________________9_437762(.CLRB (reset), .CLK (clk), .DIN
       (_________32448), .QN (_________34454));
  nnd2s1 ___9___437763(.DIN1 (_________30134), .DIN2 (_________32449),
       .Q (_________32452));
  nnd2s1 ___9___437764(.DIN1 (_________32418), .DIN2 (_________32441),
       .Q (_________32448));
  and2s1 ___9___437765(.DIN1 (_________32446), .DIN2 (______0__32445),
       .Q (_________32447));
  or2s1 ___9___437766(.DIN1 (______0__32445), .DIN2 (_________32446),
       .Q (______9__32444));
  xor2s1 ___9___437767(.DIN1 (_________32439), .DIN2 (_________31431),
       .Q (_________32449));
  hi1s1 ___9___437768(.DIN (_________32443), .Q (______0__32461));
  xor2s1 ___9___437769(.DIN1 (_________32433), .DIN2 (_________32442),
       .Q (_________32443));
  or2s1 ___9__437770(.DIN1 (_________32438), .DIN2 (_________32440), .Q
       (_________32441));
  nor2s1 ___9___437771(.DIN1 (_________32428), .DIN2 (______9__32435),
       .Q (______0__32445));
  nnd2s1 ___9___437772(.DIN1 (_________32432), .DIN2 (______0__32426),
       .Q (_________32439));
  nor2s1 ___9___437773(.DIN1 (_________32437), .DIN2 (_________32431),
       .Q (_________32438));
  nnd2s1 ___9___437774(.DIN1 (_________32430), .DIN2 (_________32440),
       .Q (______0__32436));
  nor2s1 ___9___437775(.DIN1 (_________32429), .DIN2 (______0__31211),
       .Q (______9__32435));
  xor2s1 ___9__437776(.DIN1 (________23905), .DIN2
       (_________________18734), .Q (_________32434));
  xor2s1 ___9___437777(.DIN1 (_________29563), .DIN2
       (_____________0___18740), .Q (_________32433));
  nnd2s1 ___9___437778(.DIN1 (_____9___31351), .DIN2 (_________32424),
       .Q (_________32432));
  or2s1 ___9___437779(.DIN1 (_____________0___18740), .DIN2
       (____9____32697), .Q (_________32431));
  xor2s1 ___9__437780(.DIN1 (______9__32425), .DIN2 (_____9___31352),
       .Q (_________32430));
  and2s1 ___9___437781(.DIN1 (_________32427), .DIN2
       (_____________0___18740), .Q (_________32429));
  nor2s1 ___9___437782(.DIN1 (_____________0___18740), .DIN2
       (_________32427), .Q (_________32428));
  nnd2s1 ___9__437783(.DIN1 (______9__32425), .DIN2
       (_________________18725), .Q (______0__32426));
  or2s1 ___9__437784(.DIN1 (_________________18725), .DIN2
       (______9__32425), .Q (_________32424));
  dffacs1 ___________________437785(.CLRB (reset), .CLK (clk), .DIN
       (_________32417), .Q (_________________18734));
  xor2s1 ___9___437786(.DIN1 (_________34457), .DIN2 (_________32420),
       .Q (_________32423));
  nnd2s1 ___9___437787(.DIN1 (______9__32415), .DIN2 (_________32440),
       .Q (_________32422));
  dffacs1 _________________0_437788(.CLRB (reset), .CLK (clk), .DIN
       (______0__32416), .QN (_____________0___18740));
  and2s1 ___9___437789(.DIN1 (_________32420), .DIN2 (_________34457),
       .Q (_________32421));
  nor2s1 ___9___437790(.DIN1 (_________34457), .DIN2 (_________32420),
       .Q (_________32419));
  nor2s1 ___9___437791(.DIN1 (_____0___29622), .DIN2 (_________32414),
       .Q (______9__32425));
  nnd2s1 ___9___437792(.DIN1 (_________32411), .DIN2 (_________32440),
       .Q (_________32418));
  nor2s1 ___9___437793(.DIN1 (_________32919), .DIN2 (_________32412),
       .Q (_________32417));
  nnd2s1 ___9___437794(.DIN1 (_________32409), .DIN2 (____99__23083),
       .Q (______0__32416));
  xor2s1 ___9___437795(.DIN1 (_________29640), .DIN2 (_________32413),
       .Q (______9__32415));
  xor2s1 ___9___437796(.DIN1 (______0__32406), .DIN2 (_____9___32383),
       .Q (______9__32505));
  nor2s1 ___9__437797(.DIN1 (_________29601), .DIN2 (_________32413),
       .Q (_________32414));
  dffacs1 _________________0_437798(.CLRB (reset), .CLK (clk), .DIN
       (_________32408), .QN (_________34457));
  xor2s1 ___9___437799(.DIN1 (_________32375), .DIN2 (_________32401),
       .Q (_________32412));
  xor2s1 ___9___437800(.DIN1 (_________32402), .DIN2 (_________32410),
       .Q (_________32411));
  nnd2s1 ___9___437801(.DIN1 (______9__32405), .DIN2 (_________32440),
       .Q (_________32409));
  nnd2s1 ___9__437802(.DIN1 (_________32404), .DIN2 (_________29458),
       .Q (_________32456));
  nnd2s1 ___9___437803(.DIN1 (_________32403), .DIN2 (_________32407),
       .Q (_________32408));
  nor2s1 ___9___437804(.DIN1 (_____0___31190), .DIN2 (_________32400),
       .Q (_________32413));
  xor2s1 ___9___437805(.DIN1 (_________18855), .DIN2 (_________29457),
       .Q (______0__32406));
  xor2s1 ___9___437806(.DIN1 (_________31212), .DIN2 (_________32399),
       .Q (______9__32405));
  nnd2s1 ___9___437807(.DIN1 (_________29510), .DIN2 (_________18855),
       .Q (_________32404));
  xor2s1 ___9___437808(.DIN1 (_________32398), .DIN2 (______0__32594),
       .Q (_________32403));
  xor2s1 ___9___437809(.DIN1 (______0__32396), .DIN2 (_________31373),
       .Q (_________32402));
  xor2s1 ___9__437810(.DIN1 (_________32397), .DIN2 (_________32554),
       .Q (_________32401));
  nor2s1 ___9___437811(.DIN1 (_________31209), .DIN2 (_________32399),
       .Q (_________32400));
  dffacs1 __________________437812(.CLRB (reset), .CLK (clk), .DIN
       (_____09__32395), .QN (_________18855));
  nor2s1 ___9___437813(.DIN1 (_________31372), .DIN2 (_____0___32394),
       .Q (_________32399));
  xor2s1 ___9___437814(.DIN1 (_____0___32391), .DIN2 (_____99__32385),
       .Q (_________32398));
  xor2s1 ___9___437815(.DIN1 (_____0___32390), .DIN2 (_________32374),
       .Q (_________32397));
  xor2s1 ___9___437816(.DIN1 (_________31423), .DIN2 (_____0___32393),
       .Q (______0__32396));
  nnd2s1 ___9___437817(.DIN1 (_____0___32392), .DIN2 (_________33279),
       .Q (_____09__32395));
  nor2s1 ___9___437818(.DIN1 (_________31374), .DIN2 (_____0___32393),
       .Q (_____0___32394));
  xor2s1 ___9___437819(.DIN1 (_____9___32384), .DIN2 (_____0___32387),
       .Q (_____0___32392));
  nnd2s1 ___9__437820(.DIN1 (_____0___32389), .DIN2 (____00___34533),
       .Q (_____0___32391));
  nnd2s1 ___9__437821(.DIN1 (_____00__32386), .DIN2 (_____0___32389),
       .Q (_____0___32390));
  nor2s1 ___9___437822(.DIN1 (_____9___32382), .DIN2 (_____0___32388),
       .Q (_____0___32393));
  nor2s1 ___9___437823(.DIN1 (_____0___32387), .DIN2 (_____9___32381),
       .Q (_____0___32388));
  dffacs1 __________________437824(.CLRB (reset), .CLK (clk), .DIN
       (_____9___32379), .QN (_________34485));
  nnd2s1 ___9___437825(.DIN1 (_____99__32385), .DIN2 (____00___34533),
       .Q (_____00__32386));
  xor2s1 ___9___437826(.DIN1 (_____9___32378), .DIN2 (_____90__31526),
       .Q (_____0___32389));
  xor2s1 ___9___437827(.DIN1 (_____9___32383), .DIN2 (_________34468),
       .Q (_____9___32384));
  nor2s1 ___9___437828(.DIN1 (_________34468), .DIN2 (_____9___32380),
       .Q (_____9___32382));
  and2s1 ___9___437829(.DIN1 (_____9___32380), .DIN2 (_________34468),
       .Q (_____9___32381));
  nnd2s1 ___9__437830(.DIN1 (_____90__32377), .DIN2 (_________32356),
       .Q (_____9___32379));
  nnd2s1 ___9___437831(.DIN1 (_________32376), .DIN2 (_________32306),
       .Q (_____9___32378));
  nor2s1 ___9___437832(.DIN1 (_________32372), .DIN2 (_________29387),
       .Q (_____90__32377));
  dffacs1 __________________437833(.CLRB (reset), .CLK (clk), .DIN
       (_________32373), .Q (_________34468));
  xor2s1 ___9___437834(.DIN1 (____00___34534), .DIN2
       (_________________18720), .Q (_________32375));
  xor2s1 ___9___437835(.DIN1 (_________32367), .DIN2 (_____0___31191),
       .Q (_________32376));
  nor2s1 ___9_9_437836(.DIN1 (_________32365), .DIN2 (_________32371),
       .Q (_________32374));
  dffacs1 __________________437837(.CLRB (reset), .CLK (clk), .DIN
       (______9__32369), .QN (________________18757));
  nnd2s1 ___9___437838(.DIN1 (____9____30840), .DIN2 (______0__32370),
       .Q (_________32373));
  nor2s1 ___9_437839(.DIN1 (_________32368), .DIN2 (_________32344), .Q
       (_________32372));
  nor2s1 ___9_9_437840(.DIN1 (_________32366), .DIN2 (_____0___31191),
       .Q (_________32371));
  nnd2s1 ___9___437841(.DIN1 (________19962), .DIN2 (_________32364),
       .Q (______0__32370));
  nnd2s1 ___9_9_437842(.DIN1 (______0__32360), .DIN2 (_________29504),
       .Q (______9__32369));
  xor2s1 ___9_9_437843(.DIN1 (_________32322), .DIN2 (_________18866),
       .Q (_________32368));
  xor2s1 ___9_9_437844(.DIN1 (_________18866), .DIN2
       (_____________9___18719), .Q (_________32367));
  nor2s1 ___9_0_437845(.DIN1 (_________18866), .DIN2
       (_____________9___18719), .Q (_________32366));
  and2s1 ___9_0_437846(.DIN1 (_____________9___18719), .DIN2
       (_________18866), .Q (_________32365));
  nnd2s1 ___9_9_437847(.DIN1 (_________32359), .DIN2 (inData[4]), .Q
       (_________32364));
  or2s1 ___9_9_437848(.DIN1 (_________32362), .DIN2 (_________32361),
       .Q (_________32363));
  nnd2s1 ___9_437849(.DIN1 (_________32358), .DIN2 (_________33186), .Q
       (______0__32360));
  dffacs1 _________________0_437850(.CLRB (reset), .CLK (clk), .DIN
       (_________32357), .QN (_________18866));
  nor2s1 ___9_437851(.DIN1 (_________32354), .DIN2 (_____0___32299), .Q
       (_________32359));
  nor2s1 ___9_0_437852(.DIN1 (_________32355), .DIN2 (_________32040),
       .Q (_________32361));
  xor2s1 ___9__437853(.DIN1 (______9__32350), .DIN2 (_________32352),
       .Q (_________32358));
  nnd2s1 ___9___437854(.DIN1 (_________32353), .DIN2 (_________32349),
       .Q (_________32530));
  nor2s1 ___9_0_437855(.DIN1 (_________34458), .DIN2 (_________32008),
       .Q (_________32362));
  nnd2s1 ___9___437856(.DIN1 (______0__32351), .DIN2 (_________32356),
       .Q (_________32357));
  hi1s1 ___9_0_437857(.DIN (_________34458), .Q (_________32355));
  xor2s1 ___9_437858(.DIN1 (_________________18733), .DIN2
       (______9__34460), .Q (_________32354));
  or2s1 ___9__437859(.DIN1 (_________32352), .DIN2 (_________32348), .Q
       (_________32353));
  dffacs1 _________________9_437860(.CLRB (reset), .CLK (clk), .DIN
       (_________32346), .QN (_________34458));
  dffacs1 _________________9_437861(.CLRB (reset), .CLK (clk), .DIN
       (_________32343), .QN (_____________9___18703));
  nor2s1 ___9___437862(.DIN1 (_________32345), .DIN2 (______9__32281),
       .Q (______0__32351));
  and2s1 ___9___437863(.DIN1 (_________32349), .DIN2 (_________32347),
       .Q (______9__32350));
  hi1s1 ___9___437864(.DIN (_________32347), .Q (_________32348));
  nnd2s1 ___9___437865(.DIN1 (_________32339), .DIN2 (_________32407),
       .Q (_________32346));
  dffacs1 __________________437866(.CLRB (reset), .CLK (clk), .DIN
       (______0__32341), .QN (________________18736));
  dffacs1 ___________________437867(.CLRB (reset), .CLK (clk), .DIN
       (______9__32340), .QN (______9__34460));
  nor2s1 ___9___437868(.DIN1 (_________32336), .DIN2 (_________32344),
       .Q (_________32345));
  nnd2s1 ___9___437869(.DIN1 (_________32303), .DIN2 (_________32335),
       .Q (_________32343));
  nnd2s1 ___9__437870(.DIN1 (_________32333), .DIN2 (_________31194),
       .Q (_________32347));
  xor2s1 ___9__437871(.DIN1 (_________18853), .DIN2 (_________32337),
       .Q (_________32342));
  nnd2s1 ___9__437872(.DIN1 (_________32332), .DIN2 (_________31195),
       .Q (_________32349));
  nnd2s1 ___9___437873(.DIN1 (_________30704), .DIN2 (______9__32330),
       .Q (______0__32341));
  nnd2s1 ___9___437874(.DIN1 (_________32250), .DIN2 (______0__32331),
       .Q (______9__32340));
  xor2s1 ___9___437875(.DIN1 (______0__32321), .DIN2 (_________32324),
       .Q (_________32339));
  nor2s1 ___9___437876(.DIN1 (_________18853), .DIN2 (_________32337),
       .Q (_________32338));
  nor2s1 ___9___437877(.DIN1 (_____0___31003), .DIN2 (_________32323),
       .Q (_________32336));
  nnd2s1 ___9__437878(.DIN1 (_________32329), .DIN2 (clk), .Q
       (_________32335));
  and2s1 ___9___437879(.DIN1 (_________32337), .DIN2 (_________18853),
       .Q (_________32334));
  hi1s1 ___9___437880(.DIN (_________32332), .Q (_________32333));
  nor2s1 ___9___437881(.DIN1 (_________32317), .DIN2 (_________32325),
       .Q (_____99__32385));
  dffacs1 ___________________437882(.CLRB (reset), .CLK (clk), .DIN
       (______9__32320), .QN (_________34486));
  xor2s1 ___9___437883(.DIN1 (______0__32311), .DIN2 (_________32304),
       .Q (_________32332));
  nnd2s1 ___9___437884(.DIN1 (________19962), .DIN2 (_________32318),
       .Q (______0__32331));
  nnd2s1 ___9___437885(.DIN1 (_________32319), .DIN2 (inData[24]), .Q
       (______9__32330));
  dffacs1 ___________________437886(.CLRB (reset), .CLK (clk), .DIN
       (_________32314), .Q (_________18853));
  nor2s1 ___9___437887(.DIN1 (_________32312), .DIN2 (_________32219),
       .Q (_________32329));
  nor2s1 ___9__437888(.DIN1 (_________32327), .DIN2 (_________32326),
       .Q (_________32328));
  nor2s1 ___9___437889(.DIN1 (_________32313), .DIN2 (_________32324),
       .Q (_________32325));
  xor2s1 ___9__437890(.DIN1 (_____________9___18703), .DIN2
       (_________32322), .Q (_________32323));
  xor2s1 ___9___437891(.DIN1 (_________32316), .DIN2 (_________32315),
       .Q (______0__32321));
  nnd2s1 ___9___437892(.DIN1 (_____0___32295), .DIN2 (_________32307),
       .Q (______9__32320));
  nnd2s1 ___9___437893(.DIN1 (_________32305), .DIN2 (______9__32310),
       .Q (_________32510));
  nor2s1 ___9___437894(.DIN1 (_____0___32296), .DIN2 (______0__32252),
       .Q (_________32319));
  nnd2s1 ___9___437895(.DIN1 (_____0___32300), .DIN2 (inData[28]), .Q
       (_________32318));
  nor2s1 ___9___437896(.DIN1 (_________32316), .DIN2 (_________32315),
       .Q (_________32317));
  nnd2s1 ___9___437897(.DIN1 (_____0___32297), .DIN2 (_________32407),
       .Q (_________32314));
  dffacs1 ___________________437898(.CLRB (reset), .CLK (clk), .DIN
       (_____0___32293), .Q (_________________18702));
  and2s1 ___9__437899(.DIN1 (_________32315), .DIN2 (_________32316),
       .Q (_________32313));
  xnr2s1 ___9___437900(.DIN1 (_________________18720), .DIN2
       (_________34485), .Q (_________32312));
  and2s1 ___9___437901(.DIN1 (______9__32310), .DIN2 (_____00__32292),
       .Q (______0__32311));
  and2s1 ___9___437902(.DIN1 (_________32309), .DIN2
       (_________________18733), .Q (_________32327));
  nor2s1 ___9___437903(.DIN1 (_________________18733), .DIN2
       (_________32309), .Q (_________32326));
  xor2s1 ___9___437904(.DIN1 (_____09__32301), .DIN2 (_________34459),
       .Q (_________32308));
  nnd2s1 ___9___437905(.DIN1 (_____9___32290), .DIN2 (____0___23981),
       .Q (_________32307));
  nor2s1 ___9__437906(.DIN1 (_________32258), .DIN2 (_____9___32289),
       .Q (_________32324));
  or2s1 ___9___437907(.DIN1 (_________32304), .DIN2 (_____99__32291),
       .Q (_________32305));
  nnd2s1 ___9_9_437908(.DIN1 (_____9___32287), .DIN2 (_____0___32294),
       .Q (_________32303));
  and2s1 ___9__437909(.DIN1 (_________34485), .DIN2
       (_________________18720), .Q (_________32322));
  and2s1 ___9___437910(.DIN1 (_____09__32301), .DIN2 (_________34459),
       .Q (______0__32302));
  nor2s1 ___9___437911(.DIN1 (_________34459), .DIN2 (_____0___32299),
       .Q (_____0___32300));
  nor2s1 ___9___437912(.DIN1 (_________34459), .DIN2 (_____09__32301),
       .Q (_____0___32298));
  xor2s1 ___9___437913(.DIN1 (_________32270), .DIN2 (_____9___32288),
       .Q (_____0___32297));
  dffacs1 ___________________437914(.CLRB (reset), .CLK (clk), .DIN
       (_____9___32285), .QN (_________________18733));
  xor2s1 ___9___437915(.DIN1 (________________18738), .DIN2
       (_________32228), .Q (_____0___32296));
  nnd2s1 ___990_(.DIN1 (_________32280), .DIN2 (_____0___32294), .Q
       (_____0___32295));
  nnd2s1 ___9_437916(.DIN1 (_____9___32283), .DIN2 (_________34850), .Q
       (_____0___32293));
  hi1s1 ___9___437917(.DIN (_____99__32291), .Q (_____00__32292));
  nnd2s1 ___9__437918(.DIN1 (_____9___32284), .DIN2 (_________32268),
       .Q (_________32306));
  xor2s1 ___9___437919(.DIN1 (_________32277), .DIN2 (____9____33599),
       .Q (_________32316));
  nnd2s1 ___9___437920(.DIN1 (________23906), .DIN2 (_________32279),
       .Q (_____9___32290));
  nor2s1 ___9___437921(.DIN1 (______9__32261), .DIN2 (_____9___32288),
       .Q (_____9___32289));
  nor2s1 ___9___437922(.DIN1 (________________18738), .DIN2
       (_____9___32286), .Q (_____99__32291));
  nnd2s1 ___99__(.DIN1 (_________32276), .DIN2 (___99___25264), .Q
       (_____9___32287));
  nnd2s1 ___9___437923(.DIN1 (_____9___32286), .DIN2
       (________________18738), .Q (______9__32310));
  dffacs1 ___________________437924(.CLRB (reset), .CLK (clk), .DIN
       (_________32278), .Q (_________________18720));
  nor2s1 ___9___437925(.DIN1 (_________32919), .DIN2 (_________32273),
       .Q (_____9___32285));
  or2s1 ___9___437926(.DIN1 (______0__32272), .DIN2 (____9____33599),
       .Q (_____9___32284));
  dffacs1 ___________________437927(.CLRB (reset), .CLK (clk), .DIN
       (_________32274), .Q (_________34459));
  nor2s1 ___99_9(.DIN1 (____9___24601), .DIN2 (_________32267), .Q
       (_____9___32283));
  xor2s1 ___9_9_437928(.DIN1 (______0__32262), .DIN2 (____9_9__31781),
       .Q (_____90__32282));
  nor2s1 ___9___437929(.DIN1 (_________29386), .DIN2 (_________32269),
       .Q (______9__32281));
  xnr2s1 ___99__437930(.DIN1 (_________32275), .DIN2 (___99___25265),
       .Q (_________32280));
  xor2s1 ___9___437931(.DIN1 (_____________9___18719), .DIN2
       (_________34473), .Q (_________32279));
  nor2s1 ___9___437932(.DIN1 (_________32231), .DIN2 (_________32266),
       .Q (_____9___32288));
  dffacs1 __________________437933(.CLRB (reset), .CLK (clk), .DIN
       (_________32264), .Q (________________18738));
  nnd2s1 ___9___437934(.DIN1 (_________32263), .DIN2 (_____9___34820),
       .Q (_________32278));
  xnr2s1 ___9___437935(.DIN1 (______9__32271), .DIN2
       (_____________9___18719), .Q (_________32277));
  nnd2s1 ___99__437936(.DIN1 (_________32275), .DIN2 (___99___25263),
       .Q (_________32276));
  xor2s1 ___9_9_437937(.DIN1 (_________32255), .DIN2 (______9__34369),
       .Q (______0__34055));
  nnd2s1 ___9___437938(.DIN1 (_________32257), .DIN2 (_________32407),
       .Q (_________32274));
  xor2s1 ___9___437939(.DIN1 (_________32244), .DIN2 (_________32265),
       .Q (_________32273));
  nor2s1 ___9___437940(.DIN1 (______9__32271), .DIN2
       (_____________9___18719), .Q (______0__32272));
  xor2s1 ___9_9_437941(.DIN1 (_________32259), .DIN2 (_________32260),
       .Q (_________32270));
  nor2s1 ___9_9_437942(.DIN1 (______9__32251), .DIN2 (_________32256),
       .Q (_________32269));
  nnd2s1 ___9__437943(.DIN1 (_____________9___18719), .DIN2
       (______9__32271), .Q (_________32268));
  nor2s1 ___99__437944(.DIN1 (_________32158), .DIN2 (_________32254),
       .Q (_________32267));
  and2s1 ___9___437945(.DIN1 (_________32265), .DIN2 (_________32237),
       .Q (_________32266));
  nnd2s1 ___9_437946(.DIN1 (_____0___31001), .DIN2 (_________32253), .Q
       (_________32264));
  nnd2s1 ___9900(.DIN1 (_________32245), .DIN2 (_____0___32294), .Q
       (_________32263));
  nor2s1 ___99__437947(.DIN1 (______0__31958), .DIN2 (_________32249),
       .Q (______0__32262));
  and2s1 ___990_437948(.DIN1 (_________32260), .DIN2 (_________32259),
       .Q (______9__32261));
  nor2s1 ___990_437949(.DIN1 (_________32259), .DIN2 (_________32260),
       .Q (_________32258));
  nor2s1 ___99__437950(.DIN1 (_________32166), .DIN2 (_________32247),
       .Q (_________32275));
  xor2s1 ___9_9_437951(.DIN1 (______0__32223), .DIN2 (_________32234),
       .Q (_________32257));
  dffacs1 ___________________437952(.CLRB (reset), .CLK (clk), .DIN
       (______0__32243), .QN (_________________18701));
  dffacs1 _________________9_437953(.CLRB (reset), .CLK (clk), .DIN
       (______9__32242), .QN (_____________9___18719));
  and2s1 ___990_437954(.DIN1 (_________32241), .DIN2 (____0____32777),
       .Q (_________32256));
  xor2s1 ___99__437955(.DIN1 (_________32248), .DIN2 (_________34069),
       .Q (_________32255));
  xor2s1 ___99_0(.DIN1 (_________32246), .DIN2 (_________32167), .Q
       (_________32254));
  or2s1 ___9909(.DIN1 (_________32229), .DIN2 (______0__32252), .Q
       (_________32253));
  nor2s1 ___99__437956(.DIN1 (____0____32777), .DIN2 (_________32224),
       .Q (______9__32251));
  nnd2s1 ___9_9_437957(.DIN1 (______0__32233), .DIN2 (___9____19692),
       .Q (_________32250));
  nor2s1 ___990_437958(.DIN1 (______9__32222), .DIN2 (_________32235),
       .Q (_________32265));
  and2s1 ___99__437959(.DIN1 (_________32248), .DIN2 (_________31961),
       .Q (_________32249));
  nor2s1 ___99__437960(.DIN1 (_________32165), .DIN2 (_________32246),
       .Q (_________32247));
  nnd2s1 ___99__437961(.DIN1 (_________32227), .DIN2 (___9____24281),
       .Q (_________32245));
  xor2s1 ___99__437962(.DIN1 (_________32217), .DIN2 (______0__32594),
       .Q (_________32259));
  xor2s1 ___99_437963(.DIN1 (____09___30994), .DIN2 (_________32236),
       .Q (_________32244));
  nnd2s1 ___99__437964(.DIN1 (_________32210), .DIN2 (_________32218),
       .Q (______0__32243));
  nnd2s1 ___99__437965(.DIN1 (_____0___32201), .DIN2 (_________32220),
       .Q (______9__32242));
  xor2s1 ___99__437966(.DIN1 (_________32225), .DIN2 (_________32226),
       .Q (_________32241));
  nnd2s1 ___99__437967(.DIN1 (_________32239), .DIN2 (_________32238),
       .Q (_________32240));
  xor2s1 ___99__437968(.DIN1 (______0__32213), .DIN2 (____9____30882),
       .Q (_________32315));
  or2s1 ___99__437969(.DIN1 (_________32230), .DIN2 (_________32236),
       .Q (_________32237));
  nor2s1 ___99__437970(.DIN1 (_________32221), .DIN2 (_________32234),
       .Q (_________32235));
  xor2s1 ___990_437971(.DIN1 (_________32211), .DIN2 (______9__32232),
       .Q (______0__32233));
  and2s1 ___99__437972(.DIN1 (_________32236), .DIN2 (_________32230),
       .Q (_________32231));
  xor2s1 ___99_437973(.DIN1 (______), .DIN2 (_________32228), .Q
       (_________32229));
  or2s1 ___99__437974(.DIN1 (_________32226), .DIN2 (_________32225),
       .Q (_________32227));
  nnd2s1 ___99_437975(.DIN1 (_________32225), .DIN2 (_________32226),
       .Q (_________32224));
  or2s1 ___99__437976(.DIN1 (______9__32222), .DIN2 (_________32221),
       .Q (______0__32223));
  nnd2s1 ___99__437977(.DIN1 (_________32214), .DIN2 (_________32204),
       .Q (_________32246));
  nor2s1 ___99__437978(.DIN1 (_________31913), .DIN2 (______9__32212),
       .Q (_________32248));
  or2s1 ___99__437979(.DIN1 (_________32207), .DIN2 (_________32219),
       .Q (_________32220));
  nnd2s1 ___99_437980(.DIN1 (_________32206), .DIN2 (inData[2]), .Q
       (_________32218));
  nnd2s1 ___99__437981(.DIN1 (_________32216), .DIN2 (______), .Q
       (_________32238));
  dffacs1 ___________________437982(.CLRB (reset), .CLK (clk), .DIN
       (_________32205), .QN (_________34487));
  nor2s1 ___99__437983(.DIN1 (_____90__32184), .DIN2 (_________32209),
       .Q (_________32217));
  or2s1 ___99__437984(.DIN1 (______), .DIN2 (_________32216), .Q
       (_________32239));
  xor2s1 ___99__437985(.DIN1 (_____0___32196), .DIN2 (_________32215),
       .Q (______9__34026));
  xor2s1 ___99__437986(.DIN1 (_____0___32199), .DIN2 (____9_0__33587),
       .Q (_________32260));
  or2s1 ___999_(.DIN1 (_____9___33026), .DIN2 (______0__32203), .Q
       (_________32214));
  xor2s1 ___99_437987(.DIN1 (_____9___32187), .DIN2 (_____0___32851),
       .Q (_________32221));
  xor2s1 ___99__437988(.DIN1 (_____9___32186), .DIN2 (_________32208),
       .Q (_________32236));
  nnd2s1 ___99__437989(.DIN1 (_____0___32200), .DIN2 (_____0___32197),
       .Q (______0__32213));
  xor2s1 ___99__437990(.DIN1 (_____99__32193), .DIN2 (_________32606),
       .Q (______9__32212));
  xor2s1 ___99__437991(.DIN1 (_________32182), .DIN2 (_________33144),
       .Q (_________32225));
  xnr2s1 ___99_437992(.DIN1 (_________32171), .DIN2 (_________32179),
       .Q (_________32211));
  nnd2s1 ___99_437993(.DIN1 (_____0___32195), .DIN2 (_____0___32294),
       .Q (_________32210));
  dffacs1 ___________________437994(.CLRB (reset), .CLK (clk), .DIN
       (_____9___32190), .QN (______));
  dffacs1 ___________________437995(.CLRB (reset), .CLK (clk), .DIN
       (_____9___32191), .QN (_________________18732));
  nor2s1 ___99__437996(.DIN1 (_____9___32189), .DIN2 (_________32208),
       .Q (_________32209));
  xor2s1 ___99_437997(.DIN1 (_________________18701), .DIN2
       (_________32170), .Q (_________32207));
  nor2s1 ___99__437998(.DIN1 (_____9___32188), .DIN2 (_________32219),
       .Q (_________32206));
  nnd2s1 ___99__437999(.DIN1 (_____00__32194), .DIN2 (_________32156),
       .Q (_________32205));
  nnd2s1 ___000_(.DIN1 (_________32175), .DIN2 (_____9___33026), .Q
       (_________32204));
  nor2s1 ___9999(.DIN1 (_________32111), .DIN2 (_________32177), .Q
       (______0__32203));
  dffacs1 ___________________438000(.CLRB (reset), .CLK (clk), .DIN
       (_________32169), .QN (_________________18718));
  nnd2s1 ___99__438001(.DIN1 (_________32168), .DIN2 (_____0___32294),
       .Q (_____0___32201));
  nnd2s1 ___99__438002(.DIN1 (____9_0__33587), .DIN2 (_____0___32198),
       .Q (_____0___32200));
  nnd2s1 ___99__438003(.DIN1 (_____0___32198), .DIN2 (_____0___32197),
       .Q (_____0___32199));
  xor2s1 ___99__438004(.DIN1 (_____9___32192), .DIN2 (______9__34369),
       .Q (_____0___32196));
  nor2s1 ___99_438005(.DIN1 (_________32178), .DIN2 (______9__32173),
       .Q (_________32234));
  xor2s1 ___000_438006(.DIN1 (_________32176), .DIN2 (______0__32174),
       .Q (_____0___32195));
  nor2s1 ___0000(.DIN1 (___9____24297), .DIN2 (______0__32164), .Q
       (_____00__32194));
  and2s1 ___999_438007(.DIN1 (_____9___32192), .DIN2 (____0____31877),
       .Q (_____99__32193));
  nnd2s1 ___99__438008(.DIN1 (______9__32163), .DIN2 (______0__32036),
       .Q (_____9___32191));
  nnd2s1 ___99__438009(.DIN1 (_________32162), .DIN2 (_____00__34728),
       .Q (_____9___32190));
  xor2s1 ___999_438010(.DIN1 (______0__32155), .DIN2 (_________34345),
       .Q (_____0___32202));
  and2s1 ___99__438011(.DIN1 (______9__32183), .DIN2 (_____9___32185),
       .Q (_____9___32189));
  xor2s1 ___99__438012(.DIN1 (_________34486), .DIN2 (_________34473),
       .Q (_____9___32188));
  nnd2s1 ___99__438013(.DIN1 (_________32180), .DIN2 (_________32181),
       .Q (_____9___32187));
  xnr2s1 ___99__438014(.DIN1 (_____9___32185), .DIN2 (_________34473),
       .Q (_____9___32186));
  nor2s1 ___99_438015(.DIN1 (_____9___32185), .DIN2 (______9__32183),
       .Q (_____90__32184));
  nnd2s1 ___99__438016(.DIN1 (_________32161), .DIN2 (_________31236),
       .Q (_________32182));
  nor2s1 ___99__438017(.DIN1 (_________32181), .DIN2 (_________32180),
       .Q (______9__32222));
  nor2s1 ___99__438018(.DIN1 (_________32172), .DIN2 (_________32178),
       .Q (_________32179));
  and2s1 ___00__(.DIN1 (_________32176), .DIN2 (_________32112), .Q
       (_________32177));
  nor2s1 ___00__438019(.DIN1 (______0__32174), .DIN2 (_________32176),
       .Q (_________32175));
  nor2s1 ___99_438020(.DIN1 (_________32172), .DIN2 (_________32171),
       .Q (______9__32173));
  dffacs1 ___________________438021(.CLRB (reset), .CLK (clk), .DIN
       (_________32157), .QN (_________34488));
  nor2s1 ___99__438022(.DIN1 (___9), .DIN2 (_________34473), .Q
       (_________32170));
  nnd2s1 ___99_438023(.DIN1 (_________32159), .DIN2 (___0____24396), .Q
       (_________32169));
  xor2s1 ___99_438024(.DIN1 (_________31258), .DIN2 (_________32160),
       .Q (_________32168));
  or2s1 ___99__438025(.DIN1 (______9__32271), .DIN2 (_________34473),
       .Q (_____0___32198));
  nnd2s1 ___99__438026(.DIN1 (______9__32271), .DIN2 (_________34473),
       .Q (_____0___32197));
  nor2s1 ___00_9(.DIN1 (_________32166), .DIN2 (_________32165), .Q
       (_________32167));
  nor2s1 ___00_0(.DIN1 (_________32122), .DIN2 (_________32147), .Q
       (______0__32164));
  nnd2s1 ___99__438027(.DIN1 (_________32148), .DIN2 (_________34966),
       .Q (______9__32163));
  nor2s1 ___000_438028(.DIN1 (______9__32154), .DIN2 (_________32152),
       .Q (_____9___32192));
  nnd2s1 ___99__438029(.DIN1 (_________32153), .DIN2 (_________34966),
       .Q (_________32162));
  nnd2s1 ___99__438030(.DIN1 (_________32160), .DIN2 (_________31235),
       .Q (_________32161));
  xor2s1 ___99__438031(.DIN1 (_________32137), .DIN2 (______9__32232),
       .Q (_________32181));
  or2s1 ___999_438032(.DIN1 (_________32158), .DIN2 (_________32142),
       .Q (_________32159));
  nnd2s1 ___9990(.DIN1 (_________32143), .DIN2 (_________32156), .Q
       (_________32157));
  nor2s1 ___999_438033(.DIN1 (_____00__32096), .DIN2 (_________32146),
       .Q (_________32171));
  dffacs2 ___________________438034(.CLRB (reset), .CLK (clk), .DIN
       (______9__32144), .Q (_________34473));
  or2s1 ___00__438035(.DIN1 (______9__32154), .DIN2 (_________32139),
       .Q (______0__32155));
  xor2s1 ___99__438036(.DIN1 (_________32132), .DIN2 (______0__30283),
       .Q (_________32178));
  nor2s1 ___00__438037(.DIN1 (_____0___32100), .DIN2 (_________32141),
       .Q (_________32176));
  dffacs1 ___________________438038(.CLRB (reset), .CLK (clk), .DIN
       (_________32136), .Q (_________________18700));
  xor2s1 ___999_438039(.DIN1 (______0__32145), .DIN2 (_____0___32097),
       .Q (_________32153));
  and2s1 ___00__438040(.DIN1 (_________32138), .DIN2 (_________34345),
       .Q (_________32152));
  nor2s1 ___000_438041(.DIN1 (_____0___31187), .DIN2 (______9__32134),
       .Q (_________32160));
  or2s1 ___00__438042(.DIN1 (_________32150), .DIN2 (_________32149),
       .Q (_________32151));
  xor2s1 ___99__438043(.DIN1 (_________32124), .DIN2 (_________32108),
       .Q (_________32148));
  xor2s1 ___00_438044(.DIN1 (_____0___32102), .DIN2 (_________32140),
       .Q (_________32147));
  xor2s1 ___00__438045(.DIN1 (______9__32115), .DIN2 (____9_9__33643),
       .Q (_________32165));
  nor2s1 ___000_438046(.DIN1 (______0__32145), .DIN2 (_____99__32095),
       .Q (_________32146));
  nnd2s1 ___000_438047(.DIN1 (_________32120), .DIN2 (____0___23982),
       .Q (______9__32144));
  nor2s1 ___000_438048(.DIN1 (_________32123), .DIN2 (_____0___32099),
       .Q (_________32143));
  xor2s1 ___0009(.DIN1 (_____0___31189), .DIN2 (_________32133), .Q
       (_________32142));
  nor2s1 ___00__438049(.DIN1 (_____0___32101), .DIN2 (_________32140),
       .Q (_________32141));
  hi1s1 ___00__438050(.DIN (_________32138), .Q (_________32139));
  nnd2s1 ___00_438051(.DIN1 (_________32121), .DIN2 (______0__32106),
       .Q (_________32137));
  or2s1 ___00__438052(.DIN1 (_________32072), .DIN2 (______0__32116),
       .Q (_________32136));
  xor2s1 ___00__438053(.DIN1 (_________32129), .DIN2 (_________32128),
       .Q (______0__32135));
  nor2s1 ___00__438054(.DIN1 (_____0___31188), .DIN2 (_________32133),
       .Q (______9__32134));
  nnd2s1 ___00__438055(.DIN1 (______0__34658), .DIN2 (_________32131),
       .Q (_________32132));
  nnd2s1 ___00__438056(.DIN1 (______9__32125), .DIN2 (_________32215),
       .Q (_________32138));
  nor2s1 ___000_438057(.DIN1 (_________32131), .DIN2 (______0__34658),
       .Q (_________32172));
  nor2s1 ___00__438058(.DIN1 (_________32129), .DIN2 (_________32128),
       .Q (_________32130));
  and2s1 ___00__438059(.DIN1 (_________32128), .DIN2 (_________32129),
       .Q (_________32127));
  nor2s1 ___00__438060(.DIN1 (_________________18797), .DIN2
       (______0__32126), .Q (_________32150));
  and2s1 ___00__438061(.DIN1 (______0__32126), .DIN2
       (_________________18797), .Q (_________32149));
  nor2s1 ___00_438062(.DIN1 (_________32215), .DIN2 (______9__32125),
       .Q (______9__32154));
  xor2s1 ___00__438063(.DIN1 (_____9___32091), .DIN2 (_________32070),
       .Q (_________32124));
  and2s1 ___00__438064(.DIN1 (_________32122), .DIN2 (_________32107),
       .Q (_________32123));
  nnd2s1 ___00_438065(.DIN1 (_____0___33226), .DIN2 (_____09__32105),
       .Q (_________32121));
  nnd2s1 ___00__438066(.DIN1 (_____0___32103), .DIN2 (_____0___32294),
       .Q (_________32120));
  nnd2s1 ___00__438067(.DIN1 (_________32109), .DIN2 (_________32071),
       .Q (______0__32145));
  xor2s1 ___00__438068(.DIN1 (_____9___32090), .DIN2 (_________34077),
       .Q (_________34006));
  nnd2s1 ___00__438069(.DIN1 (_________32118), .DIN2 (_________32117),
       .Q (_________32119));
  nor2s1 ___00_438070(.DIN1 (______0__32006), .DIN2 (_____0___32098),
       .Q (______0__32116));
  nnd2s1 ___00__438071(.DIN1 (_________32113), .DIN2 (_________32114),
       .Q (______9__32115));
  nor2s1 ___00__438072(.DIN1 (_________32114), .DIN2 (_________32113),
       .Q (_________32166));
  xnr2s1 ___00__438073(.DIN1 (_________32114), .DIN2 (_____9___34038),
       .Q (______0__32174));
  xor2s1 ___00__438074(.DIN1 (_____9___32089), .DIN2
       (_________________0___18633), .Q (_________32140));
  dffacs1 ___________________438075(.CLRB (reset), .CLK (clk), .DIN
       (_________32110), .QN (_________34474));
  or2s1 ___00__438076(.DIN1 (_________32114), .DIN2 (_____9___34038),
       .Q (_________32112));
  nor2s1 ___00__438077(.DIN1 (_________31165), .DIN2 (_____9___32094),
       .Q (_________32133));
  xor2s1 ___00__438078(.DIN1 (_____90__30810), .DIN2
       (_________________18717), .Q (_________32131));
  nor2s1 ___00__438079(.DIN1 (_________32044), .DIN2 (_____9___32087),
       .Q (______9__32125));
  and2s1 ___00__438080(.DIN1 (_____9___34038), .DIN2 (_________32114),
       .Q (_________32111));
  hi1s1 ___0_00(.DIN (_________32113), .Q (______0__32126));
  nnd2s1 ___00__438081(.DIN1 (_____9___32088), .DIN2 (_________32030),
       .Q (_________32128));
  dffacs1 ___________________438082(.CLRB (reset), .CLK (clk), .DIN
       (_____9___32092), .QN (_________________18699));
  nnd2s1 ___00__438083(.DIN1 (______9__32085), .DIN2 (_____0__23821),
       .Q (_________32110));
  nnd2s1 ___00__438084(.DIN1 (_________32108), .DIN2 (_________32084),
       .Q (_________32109));
  or2s1 ___00__438085(.DIN1 (_____09__31192), .DIN2
       (_________________18717), .Q (_________32107));
  or2s1 ___00__438086(.DIN1 (_________________18717), .DIN2
       (_____0___32104), .Q (______0__32106));
  nnd2s1 ___00__438087(.DIN1 (_____0___32104), .DIN2
       (_________________18717), .Q (_____09__32105));
  xor2s1 ___00_438088(.DIN1 (______9__31166), .DIN2 (_____9___32093),
       .Q (_____0___32103));
  or2s1 ___0_0_(.DIN1 (_____0___32101), .DIN2 (_____0___32100), .Q
       (_____0___32102));
  nor2s1 ___0090(.DIN1 (_________32122), .DIN2 (_________32080), .Q
       (_____0___32099));
  xor2s1 ___009_(.DIN1 (_________32064), .DIN2 (_________28828), .Q
       (_____0___32098));
  nor2s1 ___00__438089(.DIN1 (_____00__32096), .DIN2 (_____99__32095),
       .Q (_____0___32097));
  xor2s1 ___0099(.DIN1 (______0__32066), .DIN2 (_________31431), .Q
       (_________32118));
  nnd2s1 ___0_09(.DIN1 (_________32079), .DIN2 (_________31126), .Q
       (_________32113));
  dffacs1 ___________________438090(.CLRB (reset), .CLK (clk), .DIN
       (_________32082), .QN (_________34475));
  and2s1 ___00__438091(.DIN1 (_____9___32093), .DIN2 (_________31137),
       .Q (_____9___32094));
  nnd2s1 ___00__438092(.DIN1 (_________32007), .DIN2 (_________32073),
       .Q (_____9___32092));
  xor2s1 ___00__438093(.DIN1 (_________32083), .DIN2 (_________33925),
       .Q (_____9___32091));
  xor2s1 ___00__438094(.DIN1 (_________32057), .DIN2 (_________34345),
       .Q (_____9___32090));
  nor2s1 ___0_0_438095(.DIN1 (_____9___31991), .DIN2 (_________32068),
       .Q (_____9___32089));
  or2s1 ___0_0_438096(.DIN1 (_____________9___18751), .DIN2
       (______9__32065), .Q (_____9___32088));
  nor2s1 ___00__438097(.DIN1 (____0____31831), .DIN2 (_________32069),
       .Q (_____9___32087));
  xor2s1 ___0___(.DIN1 (________21853), .DIN2 (______0__32076), .Q
       (_____90__32086));
  xnr2s1 ___0___438098(.DIN1 (_____0___31902), .DIN2 (_________32078),
       .Q (_____9___34038));
  or2s1 ___00__438099(.DIN1 (_________32158), .DIN2 (______0__32056),
       .Q (______9__32085));
  nnd2s1 ___00__438100(.DIN1 (_________32083), .DIN2 (_________30682),
       .Q (_________32084));
  nnd2s1 ___00__438101(.DIN1 (_________32059), .DIN2 (_________32156),
       .Q (_________32082));
  xor2s1 ___00__438102(.DIN1 (_________32043), .DIN2 (_________32081),
       .Q (_____99__32095));
  dffacs1 ___________________438103(.CLRB (reset), .CLK (clk), .DIN
       (_________32060), .QN (_________________18717));
  xor2s1 ___0___438104(.DIN1 (_________32027), .DIN2 (_________32067),
       .Q (_________32080));
  nnd2s1 ___0__9(.DIN1 (_________32078), .DIN2 (_____9___31088), .Q
       (_________32079));
  nnd2s1 ___0___438105(.DIN1 (______0__32076), .DIN2 (_________32074),
       .Q (_________32077));
  nor2s1 ___0___438106(.DIN1 (_________32074), .DIN2 (______0__32076),
       .Q (______9__32075));
  nor2s1 ___0___438107(.DIN1
       (______________0______________________18824), .DIN2
       (______0__32076), .Q (_____0___32101));
  dffacs1 ___________________438108(.CLRB (reset), .CLK (clk), .DIN
       (_________32061), .QN (_________________18731));
  nnd2s1 ___00_438109(.DIN1 (_________32054), .DIN2 (inData[22]), .Q
       (_________32073));
  nor2s1 ___00_438110(.DIN1 (_________32050), .DIN2 (_________32053),
       .Q (_________32072));
  nnd2s1 ___00__438111(.DIN1 (_________32058), .DIN2 (_________32070),
       .Q (_________32071));
  nnd2s1 ___00_438112(.DIN1 (_________32047), .DIN2 (____9____31738),
       .Q (_________32069));
  nor2s1 ___00__438113(.DIN1 (____0____30944), .DIN2 (_________32052),
       .Q (_____9___32093));
  nor2s1 ___0___438114(.DIN1 (_________32010), .DIN2 (_________32067),
       .Q (_________32068));
  nor2s1 ___0___438115(.DIN1 (_________32062), .DIN2 (_________32063),
       .Q (______0__32066));
  xnr2s1 ___0__0(.DIN1 (_____9___33022), .DIN2 (_________32031), .Q
       (______9__32065));
  xor2s1 ___0___438116(.DIN1 (_________32024), .DIN2 (______9__32035),
       .Q (_________32064));
  nnd2s1 ___0___438117(.DIN1 (_________32063), .DIN2 (_________32062),
       .Q (_________32117));
  nor2s1 ___0___438118(.DIN1 (_________32114), .DIN2 (______9__32055),
       .Q (_____0___32100));
  nnd2s1 ___00__438119(.DIN1 (_________32038), .DIN2 (________23926),
       .Q (_________32061));
  nnd2s1 ___00_438120(.DIN1 (_________32039), .DIN2 (________25894), .Q
       (_________32060));
  nor2s1 ___00__438121(.DIN1 (_____9__24635), .DIN2 (_________32037),
       .Q (_________32059));
  hi1s1 ___00__438122(.DIN (_________32058), .Q (_________32083));
  xor2s1 ___009_438123(.DIN1 (______9__32045), .DIN2 (______0__32046),
       .Q (_________32057));
  xor2s1 ___00__438124(.DIN1 (____0____30967), .DIN2 (_________32051),
       .Q (______0__32056));
  nnd2s1 ___0___438125(.DIN1 (_________32033), .DIN2 (_________31925),
       .Q (_________32078));
  hi1s1 ___0__438126(.DIN (______9__32055), .Q (______0__32076));
  nor2s1 ___00__438127(.DIN1 (_________32028), .DIN2 (_________32053),
       .Q (_________32054));
  nor2s1 ___00_438128(.DIN1 (____0____30948), .DIN2 (_________32051),
       .Q (_________32052));
  xor2s1 ___00__438129(.DIN1 (____09__25760), .DIN2 (_________32017),
       .Q (_________32050));
  xor2s1 ___00__438130(.DIN1 (_________32018), .DIN2 (_________32049),
       .Q (_________32058));
  xor2s1 ___009_438131(.DIN1 (____9____31778), .DIN2 (_________32022),
       .Q (______9__33908));
  nor2s1 ___009_438132(.DIN1 (_________32041), .DIN2 (_________32042),
       .Q (_____00__32096));
  nnd2s1 ___0__438133(.DIN1 (_________32023), .DIN2 (_________28937),
       .Q (_________32048));
  nnd2s1 ___0_0_438134(.DIN1 (______0__32046), .DIN2 (______9__32045),
       .Q (_________32047));
  nor2s1 ___0_0_438135(.DIN1 (____0____31840), .DIN2 (______0__32046),
       .Q (_________32044));
  nnd2s1 ___009_438136(.DIN1 (_________32042), .DIN2 (_________32041),
       .Q (_________32043));
  nor2s1 ___0___438137(.DIN1 (_________32034), .DIN2 (______9__32025),
       .Q (_________32067));
  xor2s1 ___0___438138(.DIN1 (_________28962), .DIN2 (_________32040),
       .Q (_________32063));
  xor2s1 ___0___438139(.DIN1 (_________31944), .DIN2 (_________32032),
       .Q (______9__32055));
  nnd2s1 ___009_438140(.DIN1 (_________32020), .DIN2 (___9____24302),
       .Q (_________32039));
  nnd2s1 ___00_438141(.DIN1 (_________32019), .DIN2 (_________34966),
       .Q (_________32038));
  nnd2s1 ___00__438142(.DIN1 (_________32021), .DIN2 (________24874),
       .Q (_________32037));
  nnd2s1 ___009_438143(.DIN1 (______9__32015), .DIN2 (clk), .Q
       (______0__32036));
  nor2s1 ___0___438144(.DIN1 (_________32013), .DIN2 (_________32034),
       .Q (______9__32035));
  nnd2s1 ___0___438145(.DIN1 (_________32032), .DIN2 (______9__31957),
       .Q (_________32033));
  nor2s1 ___0___438146(.DIN1 (_________32029), .DIN2 (_________32040),
       .Q (_________32031));
  nnd2s1 ___0___438147(.DIN1 (_________32040), .DIN2 (_________32029),
       .Q (_________32030));
  xor2s1 ___0___438148(.DIN1 (_________28961), .DIN2 (_________32420),
       .Q (_________32129));
  xor2s1 ___0___438149(.DIN1 (______0__32016), .DIN2
       (_________________18685), .Q (_________32028));
  nor2s1 ___0___438150(.DIN1 (_________30476), .DIN2 (_____0___32003),
       .Q (_________32041));
  nor2s1 ___0_0_438151(.DIN1 (____90___30825), .DIN2 (_____09__32005),
       .Q (_________32051));
  nnd2s1 ___0___438152(.DIN1 (_____0___32002), .DIN2 (____9____31777),
       .Q (______0__32046));
  xor2s1 ___0___438153(.DIN1 (___00___20700), .DIN2 (______0__32026),
       .Q (_________32027));
  and2s1 ___0___438154(.DIN1 (_________32024), .DIN2 (_________32012),
       .Q (______9__32025));
  nnd2s1 ___0__438155(.DIN1 (_________32420), .DIN2 (_________28933),
       .Q (_________32023));
  dffacs1 ___________________438156(.CLRB (reset), .CLK (clk), .DIN
       (_____9___31994), .QN (_________________18730));
  xor2s1 ___0___438157(.DIN1 (_____9___33026), .DIN2 (_____0___32001),
       .Q (_________32022));
  nor2s1 ___0_0_438158(.DIN1 (________24637), .DIN2 (______9__31986),
       .Q (_________32021));
  xor2s1 ___0___438159(.DIN1 (_____0___32004), .DIN2 (____9____30843),
       .Q (_________32020));
  xor2s1 ___0___438160(.DIN1 (_________31981), .DIN2 (_________31971),
       .Q (_________32019));
  xor2s1 ___0___438161(.DIN1 (______9__30519), .DIN2 (_________34476),
       .Q (_________32018));
  nnd2s1 ___0___438162(.DIN1 (______0__32016), .DIN2
       (_________________18700), .Q (_________32017));
  nor2s1 ___0_0_438163(.DIN1 (_________31985), .DIN2 (______0__32252),
       .Q (______9__32015));
  xor2s1 ___0_9_(.DIN1 (_____9___31992), .DIN2 (_____0___34424), .Q
       (_________32014));
  hi1s1 ___0__438164(.DIN (_________32012), .Q (_________32013));
  nnd2s1 ___0___438165(.DIN1 (______0__32026), .DIN2 (_____9__19224),
       .Q (_________32011));
  nor2s1 ___0___438166(.DIN1 (______0__18865), .DIN2 (______0__32026),
       .Q (_________32010));
  xor2s1 ___0___438167(.DIN1 (_____00__31997), .DIN2 (_____99__31996),
       .Q (_________32009));
  nnd2s1 ___0___438168(.DIN1 (_________31984), .DIN2 (____0____31853),
       .Q (_________32032));
  hi1s1 ___0_90(.DIN (_________32008), .Q (_________32040));
  or2s1 ___0___438169(.DIN1 (______0__32006), .DIN2 (______9__31976),
       .Q (_________32007));
  nor2s1 ___0__438170(.DIN1 (____9_0__30828), .DIN2 (_____0___32004),
       .Q (_____09__32005));
  nor2s1 ___0__438171(.DIN1 (_________34476), .DIN2 (_____0___30546),
       .Q (_____0___32003));
  nnd2s1 ___0__438172(.DIN1 (_____0___32001), .DIN2 (____9_0__31782),
       .Q (_____0___32002));
  hi1s1 ___0___438173(.DIN (_____0___31999), .Q (_____0___32000));
  and2s1 ___0___438174(.DIN1 (_____00__31997), .DIN2 (_____99__31996),
       .Q (_____0___31998));
  nor2s1 ___0___438175(.DIN1 (_____99__31996), .DIN2 (_____00__31997),
       .Q (_____9___31995));
  nnd2s1 ___009_438176(.DIN1 (_________31982), .DIN2 (________23213),
       .Q (_____9___31994));
  and2s1 ___0_0_438177(.DIN1 (_____9___31992), .DIN2 (_____0___34424),
       .Q (_____9___31993));
  nor2s1 ___0___438178(.DIN1 (______18913), .DIN2 (_____9___31989), .Q
       (_____9___31991));
  nnd2s1 ___0___438179(.DIN1 (_____9___31989), .DIN2
       (_________________18795), .Q (_____9___31990));
  or2s1 ___0_0_438180(.DIN1 (_____0___34424), .DIN2 (_____9___31992),
       .Q (_____9___31988));
  xor2s1 ___0_9_438181(.DIN1 (_________31975), .DIN2 (________19986),
       .Q (_________32024));
  nor2s1 ___0___438182(.DIN1 (_________34496), .DIN2 (_____90__31987),
       .Q (_________32034));
  xor2s1 ___0_438183(.DIN1 (_________31969), .DIN2 (_____0___31906), .Q
       (_________32008));
  nnd2s1 ___0___438184(.DIN1 (_____90__31987), .DIN2 (_________34496),
       .Q (_________32012));
  xor2s1 ___0_0_438185(.DIN1 (_________31970), .DIN2
       (_______________18884), .Q (_________32420));
  nor2s1 ___0___438186(.DIN1 (_________32122), .DIN2 (_________31974),
       .Q (______9__31986));
  xor2s1 ___0___438187(.DIN1 (___9____19761), .DIN2
       (_____________0___18729), .Q (_________31985));
  hi1s1 ___0___438188(.DIN (_________34476), .Q (______0__32016));
  nor2s1 ___0_0_438189(.DIN1 (____0____31854), .DIN2 (______0__31968),
       .Q (_________31984));
  nor2s1 ___0___438190(.DIN1 (_________31980), .DIN2 (_________31973),
       .Q (_________32108));
  xor2s1 ___0___438191(.DIN1 (_________31962), .DIN2 (_________31983),
       .Q (_____0___31999));
  hi1s1 ___0___438192(.DIN (_____9___31989), .Q (______0__32026));
  nnd2s1 ___0__438193(.DIN1 (_________31963), .DIN2 (_________31920),
       .Q (_________31982));
  or2s1 ___0___438194(.DIN1 (_________31972), .DIN2 (_________31980),
       .Q (_________31981));
  or2s1 ___0___438195(.DIN1 (_____________0___18729), .DIN2
       (_________31978), .Q (_________31979));
  nnd2s1 ___0__438196(.DIN1 (_________31978), .DIN2
       (_____________0___18729), .Q (______0__31977));
  nor2s1 ___0___438197(.DIN1 (______0__30791), .DIN2 (_________31966),
       .Q (_____0___32004));
  dffacs1 ___________________438198(.CLRB (reset), .CLK (clk), .DIN
       (_________31964), .Q (_________34476));
  xor2s1 ___0_9_438199(.DIN1 (_________31954), .DIN2 (_________31959),
       .Q (______9__31976));
  xnr2s1 ___0___438200(.DIN1 (_________32049), .DIN2 (_________31955),
       .Q (_____0___32001));
  nor2s1 ___0___438201(.DIN1 (_________31953), .DIN2 (_________31960),
       .Q (_____90__31987));
  xor2s1 ___0__438202(.DIN1 (____0____31836), .DIN2 (______9__31967),
       .Q (_____9___31989));
  hi1s1 ___0___438203(.DIN (_________31975), .Q (_____9___31992));
  xor2s1 ___0_99(.DIN1 (_________31952), .DIN2 (_________18856), .Q
       (_____00__31997));
  xor2s1 ___0___438204(.DIN1 (_____9___30811), .DIN2 (_________31965),
       .Q (_________31974));
  nor2s1 ___0___438205(.DIN1 (_________31972), .DIN2 (_________31971),
       .Q (_________31973));
  xor2s1 ___0___438206(.DIN1 (_________31939), .DIN2 (_________31943),
       .Q (_________31970));
  xor2s1 ___0___438207(.DIN1 (_________31942), .DIN2 (_________31290),
       .Q (_________31969));
  nor2s1 ___0___438208(.DIN1 (____0_9__31823), .DIN2 (______9__31967),
       .Q (______0__31968));
  xor2s1 ___0___438209(.DIN1 (_________31941), .DIN2 (______0__30591),
       .Q (_________31975));
  nor2s1 ___0___438210(.DIN1 (_________30793), .DIN2 (_________31965),
       .Q (_________31966));
  or2s1 ___0___438211(.DIN1 (_________31949), .DIN2 (______9__31947),
       .Q (_________31964));
  xor2s1 ___0___438212(.DIN1 (_________31935), .DIN2 (_________31936),
       .Q (_________31963));
  xor2s1 ___0___438213(.DIN1 (____00___34536), .DIN2 (____0____32823),
       .Q (_________31980));
  dffacs1 _________________0_438214(.CLRB (reset), .CLK (clk), .DIN
       (______0__31948), .Q (_____________0___18729));
  xor2s1 ___0_9_438215(.DIN1 (_________31932), .DIN2 (_________31933),
       .Q (_________31962));
  nnd2s1 ___0___438216(.DIN1 (_________34069), .DIN2 (______9__34369),
       .Q (_________31961));
  and2s1 ___0___438217(.DIN1 (_________31946), .DIN2 (_________31959),
       .Q (_________31960));
  nor2s1 ___0__438218(.DIN1 (______9__34369), .DIN2 (_________34069),
       .Q (______0__31958));
  xnr2s1 ___0___438219(.DIN1 (_________31956), .DIN2 (_________31927),
       .Q (______9__31957));
  dffacs1 ___________________438220(.CLRB (reset), .CLK (clk), .DIN
       (_________31950), .QN (_________34477));
  nnd2s1 ___0_0_438221(.DIN1 (_________31934), .DIN2 (_________31930),
       .Q (_________31955));
  nnd2s1 ___0_9_438222(.DIN1 (_________31937), .DIN2 (____0____31884),
       .Q (_________31971));
  or2s1 ___0___438223(.DIN1 (_________31953), .DIN2 (_________31945),
       .Q (_________31954));
  xor2s1 ___0___438224(.DIN1 (_________31914), .DIN2 (____9____30860),
       .Q (_________31952));
  xor2s1 ___0___438225(.DIN1 (_________31915), .DIN2 (_________31951),
       .Q (______9__31967));
  or2s1 ___0__438226(.DIN1 (_________31949), .DIN2 (______0__31919), .Q
       (_________31950));
  nnd2s1 ___0__438227(.DIN1 (_________31921), .DIN2 (________22824), .Q
       (______0__31948));
  nnd2s1 ___0___438228(.DIN1 (_________31922), .DIN2 (________25885),
       .Q (______9__31947));
  hi1s1 ___0___438229(.DIN (_________31945), .Q (_________31946));
  xor2s1 ___0_9_438230(.DIN1 (_________31911), .DIN2 (_________30693),
       .Q (_________31965));
  nor2s1 ___0_0_438231(.DIN1 (____0____31859), .DIN2 (______9__31918),
       .Q (_____99__31996));
  xor2s1 ___0___438232(.DIN1 (_________31943), .DIN2 (_________31926),
       .Q (_________31944));
  nnd2s1 ___0___438233(.DIN1 (______0__31938), .DIN2 (____0____31838),
       .Q (_________31942));
  xor2s1 ___0___438234(.DIN1 (_____0___31904), .DIN2 (_________31940),
       .Q (_________31941));
  nnd2s1 ___0___438235(.DIN1 (______0__31938), .DIN2 (_____0___31907),
       .Q (_________31939));
  dffacs1 ___________________438236(.CLRB (reset), .CLK (clk), .DIN
       (_________31916), .QN (_________________18728));
  xor2s1 ___0___438237(.DIN1 (____0____30950), .DIN2 (_____0___31905),
       .Q (_________34069));
  nnd2s1 ___0_0_438238(.DIN1 (_________31936), .DIN2 (____0____31887),
       .Q (_________31937));
  xor2s1 ___0___438239(.DIN1 (____099__31899), .DIN2 (____0____31885),
       .Q (_________31935));
  nnd2s1 ___0___438240(.DIN1 (_________31931), .DIN2 (_________31933),
       .Q (_________31934));
  nnd2s1 ___0__438241(.DIN1 (_________31931), .DIN2 (_________31930),
       .Q (_________31932));
  nor2s1 ___0___438242(.DIN1 (______0__31910), .DIN2 (______9__31928),
       .Q (______0__31929));
  nnd2s1 ___0_438243(.DIN1 (_________31943), .DIN2 (_________31926), .Q
       (_________31927));
  or2s1 ___0_9_438244(.DIN1 (_________31926), .DIN2 (_________31943),
       .Q (_________31925));
  xor2s1 ___0__438245(.DIN1 (____0_9__31889), .DIN2 (_____0___31450),
       .Q (_________31945));
  nnd2s1 ___0___438246(.DIN1 (_____0___31908), .DIN2 (____9____29068),
       .Q (_________32062));
  hi1s1 ___0___438247(.DIN (_________31923), .Q (_________31924));
  or2s1 ___0___438248(.DIN1 (______0__32006), .DIN2 (_____0___31901),
       .Q (_________31922));
  nnd2s1 ___0___438249(.DIN1 (____09___31896), .DIN2 (_________31920),
       .Q (_________31921));
  nnd2s1 ___0_9_438250(.DIN1 (_____00__31900), .DIN2 (________24180),
       .Q (______0__31919));
  nor2s1 ___0___438251(.DIN1 (_________31917), .DIN2 (____09___31892),
       .Q (______9__31918));
  nnd2s1 ___0___438252(.DIN1 (____09___31895), .DIN2 (_____0__22826),
       .Q (_________31916));
  nor2s1 ___0___438253(.DIN1 (_________31912), .DIN2 (_________30575),
       .Q (_________31972));
  nnd2s1 ___0_438254(.DIN1 (____09___31894), .DIN2 (_____0___31903), .Q
       (_________31915));
  xor2s1 ___0___438255(.DIN1 (_________32337), .DIN2 (____9____29015),
       .Q (_________31914));
  xor2s1 ___0___438256(.DIN1 (____0____31878), .DIN2 (____0____31863),
       .Q (_________31913));
  nor2s1 ___0___438257(.DIN1 (____9____31784), .DIN2 (____090__31890),
       .Q (______0__31938));
  dffacs1 _________________9_438258(.CLRB (reset), .CLK (clk), .DIN
       (____09___31897), .QN (______0__34461));
  dffacs1 ___________________438259(.CLRB (reset), .CLK (clk), .DIN
       (____09___31891), .QN (_________________18698));
  dffacs1 _________________0_438260(.CLRB (reset), .CLK (clk), .DIN
       (____09___31898), .QN (_____________0___18697));
  nor2s1 ___0___438261(.DIN1 (_________30757), .DIN2 (____0____31881),
       .Q (_________31911));
  xor2s1 ___0___438262(.DIN1 (____0____31866), .DIN2 (____0____31858),
       .Q (_________31923));
  nnd2s1 ___0___438263(.DIN1 (____0_9__31880), .DIN2 (____9_0__31792),
       .Q (_________31931));
  nor2s1 ___0___438264(.DIN1 (____0____31847), .DIN2 (____0____31883),
       .Q (_________31936));
  hi1s1 ___0__438265(.DIN (_____09__31909), .Q (______0__31910));
  nnd2s1 ___0_9_438266(.DIN1 (_________32337), .DIN2 (____9____29070),
       .Q (_____0___31908));
  nnd2s1 ___0_0_438267(.DIN1 (____0____31875), .DIN2 (_____0___31906),
       .Q (_____0___31907));
  nor2s1 ___0___438268(.DIN1 (____0____30925), .DIN2 (____0____31876),
       .Q (_____0___31905));
  and2s1 ___0__438269(.DIN1 (____09___31893), .DIN2 (_____0___31903),
       .Q (_____0___31904));
  xor2s1 ___0___438270(.DIN1 (____0____31867), .DIN2 (_____0___31902),
       .Q (_________31943));
  xor2s1 ___0___438271(.DIN1 (_________30759), .DIN2 (____0____34614),
       .Q (_____0___31901));
  or2s1 ___0___438272(.DIN1 (______0__32006), .DIN2 (____0____31873),
       .Q (_____00__31900));
  xor2s1 ___0___438273(.DIN1 (____0____31886), .DIN2 (_________31431),
       .Q (____099__31899));
  nnd2s1 ___0___438274(.DIN1 (____9____31755), .DIN2 (____0_9__31870),
       .Q (____09___31898));
  nnd2s1 ___0_0_438275(.DIN1 (____0____31874), .DIN2 (____0____34616),
       .Q (____09___31897));
  xor2s1 ___0___438276(.DIN1 (____0____31848), .DIN2 (____0____31882),
       .Q (____09___31896));
  nnd2s1 ___0___438277(.DIN1 (____0____31864), .DIN2 (_________31920),
       .Q (____09___31895));
  nnd2s1 ___0___438278(.DIN1 (____0_0__31871), .DIN2 (____0____31845),
       .Q (_________31912));
  nnd2s1 ___0___438279(.DIN1 (____09___31893), .DIN2
       (_______________18881), .Q (____09___31894));
  xor2s1 ___0___438280(.DIN1 (____0____31857), .DIN2 (______0__33983),
       .Q (____09___31892));
  or2s1 ___0_9_438281(.DIN1 (________20246), .DIN2 (____0____31865), .Q
       (____09___31891));
  nor2s1 ___0___438282(.DIN1 (_________35111), .DIN2 (____0____31862),
       .Q (____090__31890));
  nnd2s1 ___0_0_438283(.DIN1 (____0____31888), .DIN2
       (_________________18685), .Q (____0_9__31889));
  nnd2s1 ___0___438284(.DIN1 (____0____31879), .DIN2 (____9____31793),
       .Q (_________31930));
  nnd2s1 ___0_438285(.DIN1 (____0____31888), .DIN2
       (_________________18794), .Q (_____09__31909));
  nor2s1 ___0_0_438286(.DIN1 (_________________18685), .DIN2
       (____0____31888), .Q (_________31953));
  nor2s1 ___0_9_438287(.DIN1 (_________________18794), .DIN2
       (____0____31888), .Q (______9__31928));
  nnd2s1 ___0___438288(.DIN1 (____0____31886), .DIN2 (____0____31885),
       .Q (____0____31887));
  or2s1 ___0___438289(.DIN1 (____0____31885), .DIN2 (____0____31886),
       .Q (____0____31884));
  nor2s1 ___0__438290(.DIN1 (____0____31846), .DIN2 (____0____31882),
       .Q (____0____31883));
  nor2s1 ___0___438291(.DIN1 (_________30758), .DIN2 (____0____34614),
       .Q (____0____31881));
  hi1s1 ___0___438292(.DIN (____0____31879), .Q (____0_9__31880));
  or2s1 ___0___438293(.DIN1 (_________32215), .DIN2 (______9__34369),
       .Q (____0____31878));
  nnd2s1 ___0___438294(.DIN1 (______9__34369), .DIN2 (_________32215),
       .Q (____0____31877));
  xor2s1 ___0___438295(.DIN1 (____0____31837), .DIN2 (_________32624),
       .Q (____0____31876));
  xor2s1 ___0___438296(.DIN1 (____0____31839), .DIN2 (_________31060),
       .Q (____0____31875));
  nnd2s1 ___0___438297(.DIN1 (____0____31856), .DIN2 (____00___31811),
       .Q (_____0___31903));
  xor2s1 ___0___438298(.DIN1 (____0____31822), .DIN2 (____0_0__31833),
       .Q (_________32337));
  dffacs1 __________________438299(.CLRB (reset), .CLK (clk), .DIN
       (____0_9__31860), .QN (________________18787));
  nnd2s1 ___0__438300(.DIN1 (____0____31843), .DIN2 (_________31920),
       .Q (____0____31874));
  xor2s1 ___0__438301(.DIN1 (____0____31828), .DIN2 (____0____31872),
       .Q (____0____31873));
  nnd2s1 ___0___438302(.DIN1 (_________30319), .DIN2 (____0_9__31850),
       .Q (____0_0__31871));
  nnd2s1 ___0__438303(.DIN1 (____0____31849), .DIN2 (clk), .Q
       (____0_9__31870));
  hi1s1 ___0___438304(.DIN (____0____31868), .Q (____0____31869));
  nnd2s1 ___0___438305(.DIN1 (____0_0__31842), .DIN2 (_________31589),
       .Q (____0____31879));
  nnd2s1 ___0__438306(.DIN1 (____0____31835), .DIN2 (____00___31813),
       .Q (____0____31867));
  xor2s1 ___0___438307(.DIN1 (_________31917), .DIN2 (_________32309),
       .Q (____0____31866));
  nor2s1 ___0___438308(.DIN1 (____9____31759), .DIN2 (____0____31834),
       .Q (____0____31865));
  xor2s1 ___0__438309(.DIN1 (____0_0__31824), .DIN2 (____0____31863),
       .Q (____0____31864));
  xor2s1 ___0__438310(.DIN1 (____0____31819), .DIN2 (____0_0__31861),
       .Q (____0____31862));
  nnd2s1 ___0___438311(.DIN1 (____0____31855), .DIN2 (____0_9__31832),
       .Q (____09___31893));
  xor2s1 ___0__438312(.DIN1 (____0____31821), .DIN2
       (______________________________________0_____________18885), .Q
       (____0____31888));
  or2s1 ___0__438313(.DIN1 (________23663), .DIN2 (____0____31830), .Q
       (____0_9__31860));
  and2s1 ___0_0_438314(.DIN1 (_________32309), .DIN2 (____0____31858),
       .Q (____0____31859));
  nor2s1 ___0__438315(.DIN1 (____000__31808), .DIN2 (____0____31826),
       .Q (____0____31882));
  xor2s1 ___0___438316(.DIN1 (_________31672), .DIN2 (____0_9__31841),
       .Q (____0____31868));
  xor2s1 ___0___438317(.DIN1 (_____0___30368), .DIN2
       (_________________18716), .Q (____0____31886));
  nor2s1 ___0___438318(.DIN1 (____0____31858), .DIN2 (_________32309),
       .Q (____0____31857));
  hi1s1 ___0___438319(.DIN (____0____31855), .Q (____0____31856));
  nor2s1 ___0___438320(.DIN1 (____0_0__31851), .DIN2 (____0____31852),
       .Q (____0____31854));
  nnd2s1 ___0___438321(.DIN1 (____0____31852), .DIN2 (____0_0__31851),
       .Q (____0____31853));
  dffacs1 ___________________438322(.CLRB (reset), .CLK (clk), .DIN
       (____0____31827), .QN (_________18864));
  xnr2s1 ___0___438323(.DIN1 (____09___34620), .DIN2 (____09___30990),
       .Q (______9__34369));
  or2s1 ___0__438324(.DIN1 (_________________18716), .DIN2
       (____0____31844), .Q (____0_9__31850));
  and2s1 ___0___438325(.DIN1 (________21313), .DIN2
       (_________________18716), .Q (____0____31849));
  or2s1 ___0__438326(.DIN1 (____0____31847), .DIN2 (____0____31846), .Q
       (____0____31848));
  nnd2s1 ___0___438327(.DIN1 (____0____31844), .DIN2
       (_________________18716), .Q (____0____31845));
  xor2s1 ___0___438328(.DIN1 (____0____31825), .DIN2 (____00___31809),
       .Q (____0____31843));
  nnd2s1 ___0_0_438329(.DIN1 (____0_9__31841), .DIN2 (_____9___31630),
       .Q (____0_0__31842));
  nor2s1 ___0___438330(.DIN1 (____9____31786), .DIN2 (____00___31814),
       .Q (____0____31840));
  and2s1 ___0_438331(.DIN1 (____0____31838), .DIN2 (_________35111), .Q
       (____0____31839));
  nnd2s1 ___0___438332(.DIN1 (____09___34620), .DIN2 (____00___30913),
       .Q (____0____31837));
  xor2s1 ___0_9_438333(.DIN1 (_____0___31906), .DIN2 (________21184),
       .Q (____0____31836));
  nnd2s1 ___0___438334(.DIN1 (____090__34618), .DIN2 (____00___31812),
       .Q (____0____31835));
  xor2s1 ___0___438335(.DIN1 (____9_9__31749), .DIN2 (____99___31802),
       .Q (____0____31834));
  xor2s1 ___0_0_438336(.DIN1 (_____0__24710), .DIN2 (____0_9__31832),
       .Q (____0_0__31833));
  xor2s1 ___0_9_438337(.DIN1 (____9____31800), .DIN2 (____0____31831),
       .Q (____0____31855));
  dffacs1 _________________9_438338(.CLRB (reset), .CLK (clk), .DIN
       (____0____31817), .QN (_________34489));
  nor2s1 ___0_9_438339(.DIN1 (____0____31829), .DIN2 (____99___31803),
       .Q (____0____31830));
  xor2s1 ___0___438340(.DIN1 (____9____31795), .DIN2 (____0____33715),
       .Q (____0____31828));
  nnd2s1 ___0_9_438341(.DIN1 (____09___34622), .DIN2 (____0____31816),
       .Q (____0____31827));
  nor2s1 ___0_0_438342(.DIN1 (____999__31807), .DIN2 (____0____31825),
       .Q (____0____31826));
  xor2s1 ___0___438343(.DIN1 (____9____31789), .DIN2 (_________30147),
       .Q (____0_0__31824));
  nor2s1 ___0___438344(.DIN1 (____0____31818), .DIN2 (_____0___31906),
       .Q (____0_9__31823));
  xor2s1 ___0_0_438345(.DIN1 (____9____31785), .DIN2
       (_________________0___18607), .Q (____0____31822));
  xor2s1 ___0_9_438346(.DIN1 (____9____31775), .DIN2 (____0____31820),
       .Q (____0____31821));
  nnd2s1 ___0___438347(.DIN1 (______0__31706), .DIN2 (____0_9__31832),
       .Q (____0____31819));
  nnd2s1 ___0___438348(.DIN1 (_____0___31906), .DIN2 (____0____31818),
       .Q (____0____31852));
  xor2s1 ___0___438349(.DIN1 (____9____31788), .DIN2 (____0____34551),
       .Q (_________32309));
  nnd2s1 ___0_9_438350(.DIN1 (____9____31796), .DIN2 (____0____31816),
       .Q (____0____31817));
  xor2s1 ___0___438351(.DIN1 (____9____31773), .DIN2 (______0__33983),
       .Q (____0____31846));
  xnr2s1 ___0__438352(.DIN1 (____009__31815), .DIN2 (____9____31772),
       .Q (____0_9__31841));
  dffacs1 ___________________438353(.CLRB (reset), .CLK (clk), .DIN
       (____9_9__31791), .Q (_________________18716));
  and2s1 ___0___438354(.DIN1 (____9____31776), .DIN2 (____0____31831),
       .Q (____00___31814));
  or2s1 ___0___438355(.DIN1 (____00___31812), .DIN2 (____9____31780),
       .Q (____00___31813));
  nnd2s1 ___0___438356(.DIN1 (____9____31783), .DIN2 (____00___31811),
       .Q (____0____31838));
  dffacs1 ___________________438357(.CLRB (reset), .CLK (clk), .DIN
       (____9____31790), .QN (_________________18727));
  nor2s1 ___0__438358(.DIN1 (____000__31808), .DIN2 (____999__31807),
       .Q (____00___31809));
  xor2s1 ___0___438359(.DIN1 (____9____31797), .DIN2 (____0____31863),
       .Q (____99___31804));
  xor2s1 ___0___438360(.DIN1 (____9____31756), .DIN2 (______0__31678),
       .Q (____99___31803));
  nnd2s1 ___0___438361(.DIN1 (____9____31764), .DIN2 (____9_9__31774),
       .Q (____99___31802));
  nnd2s1 ___0___438362(.DIN1 (____9____31770), .DIN2 (_________31655),
       .Q (____9____31800));
  nnd2s1 ___0___438363(.DIN1 (____9____31769), .DIN2 (_________30148),
       .Q (____0____31825));
  hi1s1 ___0___438364(.DIN (____00___31811), .Q (____0_9__31832));
  xor2s1 ___0___438365(.DIN1 (___9____25212), .DIN2 (____9____31779),
       .Q (_____0___31906));
  hi1s1 ___0___438366(.DIN (_________34350), .Q (_________32215));
  or2s1 ___0___438367(.DIN1 (____9____31798), .DIN2 (____9____31797),
       .Q (____9____31799));
  nor2s1 ___0___438368(.DIN1 (____9____31761), .DIN2 (_________31713),
       .Q (____9____31796));
  xor2s1 ___0___438369(.DIN1 (_________________18699), .DIN2
       (____9____31771), .Q (____9____31795));
  nor2s1 ___0___438370(.DIN1 (____9_9__31757), .DIN2 (_________35004),
       .Q (____9____31794));
  hi1s1 ___0___438371(.DIN (____9_0__31792), .Q (____9____31793));
  nnd2s1 ___0___438372(.DIN1 (____9____31760), .DIN2 (___0____20713),
       .Q (____9_9__31791));
  nnd2s1 ___0___438373(.DIN1 (____9____31754), .DIN2 (_____0__22375),
       .Q (____9____31790));
  xor2s1 ___0_9_438374(.DIN1 (_________30146), .DIN2 (____9____31768),
       .Q (____9____31789));
  xor2s1 ___0_0_438375(.DIN1 (____9____31787), .DIN2 (____9_9__31742),
       .Q (____9____31788));
  nor2s1 ___0_0_438376(.DIN1 (____0____31831), .DIN2 (______9__32045),
       .Q (____9____31786));
  nor2s1 ___0__438377(.DIN1 (____9____31758), .DIN2 (_________30297),
       .Q (____0____31847));
  or2s1 ___0___438378(.DIN1 (____9____31784), .DIN2 (____9____31783),
       .Q (____9____31785));
  xnr2s1 ___0__438379(.DIN1 (____9_9__31781), .DIN2 (____9____31747),
       .Q (____9_0__31782));
  nnd2s1 ___0_9_438380(.DIN1 (____9____31779), .DIN2 (___9_0__25211),
       .Q (____9____31780));
  nnd2s1 ___0___438381(.DIN1 (____9____31748), .DIN2 (____9____31777),
       .Q (____9____31778));
  and2s1 ___0___438382(.DIN1 (______9__32045), .DIN2 (_________34345),
       .Q (____9____31776));
  xor2s1 ___0___438383(.DIN1 (____0____34551), .DIN2 (____09___34626),
       .Q (____9____31775));
  nnd2s1 ___0___438384(.DIN1 (____9____31751), .DIN2 (____9_9__31774),
       .Q (_________31959));
  xor2s1 ___0___438385(.DIN1 (____9_0__31743), .DIN2 (_________30496),
       .Q (____00___31811));
  xor2s1 ___0__438386(.DIN1 (____9____31741), .DIN2
       (_____________18905), .Q (_________34350));
  nor2s1 ___0__438387(.DIN1 (____09___34624), .DIN2 (______9__30298),
       .Q (____9____31773));
  nnd2s1 ___0___438388(.DIN1 (____9____31745), .DIN2 (_________31507),
       .Q (____9____31772));
  xor2s1 ___0___438389(.DIN1 (____9_0__31733), .DIN2 (_________33174),
       .Q (____999__31807));
  nor2s1 ___0___438390(.DIN1 (_________30505), .DIN2 (____9____31771),
       .Q (____99___31806));
  xor2s1 ___0___438391(.DIN1 (____90___31731), .DIN2 (_________31461),
       .Q (_________33841));
  nnd2s1 ___0__438392(.DIN1 (____09___34626), .DIN2 (_________31654),
       .Q (____9____31770));
  nnd2s1 ___0___438393(.DIN1 (____9____31768), .DIN2 (_________30145),
       .Q (____9____31769));
  and2s1 ___0__438394(.DIN1 (____9____31763), .DIN2 (____9____31765),
       .Q (____9_0__31767));
  xor2s1 ___0_438395(.DIN1 (____9____31765), .DIN2 (_____09__32301), .Q
       (____9_9__31766));
  xor2s1 ___0___438396(.DIN1 (____9_0__31750), .DIN2 (______9__33828),
       .Q (____9____31764));
  or2s1 ___0___438397(.DIN1 (____9____31765), .DIN2 (____9____31763),
       .Q (____9_9__31801));
  xor2s1 ___0___438398(.DIN1 (____90___31725), .DIN2 (_________31478),
       .Q (____9_0__31792));
  nnd2s1 ___0___438399(.DIN1 (____9____31798), .DIN2 (____90___31730),
       .Q (____9____31762));
  nor2s1 ___0___438400(.DIN1 (_________31702), .DIN2 (____9____31734),
       .Q (____9____31761));
  or2s1 ___0__438401(.DIN1 (____9____31759), .DIN2 (____9____31735), .Q
       (____9____31760));
  hi1s1 ___0___438402(.DIN (____09___34624), .Q (____9____31758));
  xor2s1 ___0_438403(.DIN1 (_________________18727), .DIN2
       (_________34462), .Q (____9_9__31757));
  xor2s1 ___0__438404(.DIN1 (_____9___31722), .DIN2 (____00___33677),
       .Q (____9____31756));
  or2s1 ___0___438405(.DIN1 (____9____31759), .DIN2 (____900__31724),
       .Q (____9____31755));
  nnd2s1 ___0___438406(.DIN1 (____9____31737), .DIN2 (_________31920),
       .Q (____9____31754));
  xor2s1 ___0_0_438407(.DIN1 (_________34462), .DIN2 (______9__32514),
       .Q (____9____31797));
  nnd2s1 ___0_438408(.DIN1 (____9_0__31750), .DIN2 (____9_9__31749), .Q
       (____9____31751));
  hi1s1 ___0___438409(.DIN (____9____31747), .Q (____9____31748));
  xor2s1 ___0_438410(.DIN1 (_____9___31717), .DIN2 (____9____31746), .Q
       (____9____31784));
  nor2s1 ___0___438411(.DIN1 (________19081), .DIN2 (____90___31727),
       .Q (____9____31779));
  xor2s1 ___0__438412(.DIN1 (______9__31714), .DIN2
       (_________________0___18633), .Q (______9__32045));
  dffacs1 _________________0_438413(.CLRB (reset), .CLK (clk), .DIN
       (____9____31736), .QN (_____________0___18715));
  dffacs1 __________________438414(.CLRB (reset), .CLK (clk), .DIN
       (____909__31732), .Q (________________18771));
  nor2s1 ___0___438415(.DIN1 (_________31508), .DIN2 (_____9___31719),
       .Q (____9____31745));
  nor2s1 ___0___438416(.DIN1 (_____9___30451), .DIN2 (_____9___31721),
       .Q (____9____31771));
  hi1s1 ___0___438417(.DIN (_____09__32301), .Q (____9____31763));
  nor2s1 ___0___438418(.DIN1 (______9__31658), .DIN2 (_____9___31716),
       .Q (____9____31768));
  xor2s1 ___0___438419(.DIN1 (________19175), .DIN2 (____90___31726),
       .Q (____9_0__31743));
  xor2s1 ___0___438420(.DIN1 (_________31707), .DIN2 (____99___31805),
       .Q (____9_9__31742));
  xor2s1 ___0_9_438421(.DIN1 (_________30795), .DIN2 (_____99__31723),
       .Q (____9____31741));
  nor2s1 ___0___438422(.DIN1 (____9____31739), .DIN2 (____9____31740),
       .Q (____9____31747));
  nnd2s1 ___0___438423(.DIN1 (____9____31740), .DIN2 (____9____31739),
       .Q (____9____31777));
  hi1s1 ___0___438424(.DIN (____9____31738), .Q (_________34345));
  xor2s1 ___0__438425(.DIN1 (______0__31659), .DIN2 (_____90__31715),
       .Q (____9____31737));
  nnd2s1 ___0___438426(.DIN1 (_________31708), .DIN2 (________21314),
       .Q (____9____31736));
  xor2s1 ___0___438427(.DIN1 (_________30508), .DIN2 (_____9___31720),
       .Q (____9____31735));
  xor2s1 ___0__438428(.DIN1 (________19129), .DIN2 (_________31701), .Q
       (____9____31734));
  nnd2s1 ___0_9_438429(.DIN1 (____90___31728), .DIN2 (____90___31729),
       .Q (____9_0__31733));
  nnd2s1 ___0_9_438430(.DIN1 (_________31710), .DIN2 (________23606),
       .Q (____909__31732));
  xor2s1 ___0___438431(.DIN1 (_____9___31718), .DIN2 (_____0___31447),
       .Q (____90___31731));
  hi1s1 ___0___438432(.DIN (_________34462), .Q (____90___31730));
  nor2s1 ___0_9_438433(.DIN1 (____90___31729), .DIN2 (____90___31728),
       .Q (____000__31808));
  and2s1 ___0___438434(.DIN1 (____90___31726), .DIN2 (____90), .Q
       (____90___31727));
  xor2s1 ___0_9_438435(.DIN1 (_________31691), .DIN2 (outData[30]), .Q
       (____90___31725));
  xor2s1 ___0___438436(.DIN1 (_________31606), .DIN2 (_________31698),
       .Q (____900__31724));
  or2s1 ___0__438437(.DIN1 (_________30778), .DIN2 (_____99__31723), .Q
       (____9____31753));
  xor2s1 ___0___438438(.DIN1 (______9__31685), .DIN2 (_________31983),
       .Q (____9_0__31750));
  xnr2s1 ___0__438439(.DIN1 (_________35012), .DIN2 (_________31684),
       .Q (____9_9__31774));
  xor2s1 ___0_0_438440(.DIN1 (_________31689), .DIN2 (______0__31130),
       .Q (____9____31738));
  dffacs1 __________________438441(.CLRB (reset), .CLK (clk), .DIN
       (_________31709), .QN
       (_______________0____________________18829));
  xor2s1 ___0___438442(.DIN1 (_________31688), .DIN2 (_________31700),
       .Q (_____09__32301));
  nnd2s1 ___0___438443(.DIN1 (______9__31705), .DIN2 (______0__31650),
       .Q (_____9___31722));
  nor2s1 ___0_0_438444(.DIN1 (_________30483), .DIN2 (_____9___31720),
       .Q (_____9___31721));
  and2s1 ___0___438445(.DIN1 (_____9___31718), .DIN2 (_____0___31448),
       .Q (_____9___31719));
  nor2s1 ___0__438446(.DIN1 (_________31703), .DIN2 (_________31588),
       .Q (____9____31744));
  dffacs1 ___________________438447(.CLRB (reset), .CLK (clk), .DIN
       (______0__31696), .QN (_________34462));
  nnd2s1 ___0___438448(.DIN1 (_________31682), .DIN2 (______0__31612),
       .Q (_____9___31717));
  and2s1 ___0_9_438449(.DIN1 (_____90__31715), .DIN2 (_____0___31635),
       .Q (_____9___31716));
  nor2s1 ___0___438450(.DIN1 (_________28762), .DIN2 (_________31692),
       .Q (______9__31714));
  nor2s1 ___0__438451(.DIN1 (_________31587), .DIN2 (______9__31695),
       .Q (_________31713));
  nor2s1 ___0___438452(.DIN1 (_________31711), .DIN2 (_________31694),
       .Q (_________31712));
  nnd2s1 ___0___438453(.DIN1 (_________31687), .DIN2 (_________31690),
       .Q (____9____31740));
  nnd2s1 ___0___438454(.DIN1 (_________31680), .DIN2 (_________32639),
       .Q (_________31710));
  nnd2s1 ___0___438455(.DIN1 (______9__31677), .DIN2 (____90___32662),
       .Q (_________31709));
  or2s1 ___0___438456(.DIN1 (____9____31759), .DIN2 (_________31676),
       .Q (_________31708));
  xor2s1 ___0___438457(.DIN1 (_________30113), .DIN2
       (_____________9___18714), .Q (____90___31728));
  nor2s1 ___0___438458(.DIN1 (_________31679), .DIN2 (_________31704),
       .Q (_________32903));
  nnd2s1 ___0___438459(.DIN1 (_________31673), .DIN2 (_____9___31625),
       .Q (_________31707));
  hi1s1 ___0__438460(.DIN (______0__31706), .Q (____9____31783));
  nnd2s1 ___0___438461(.DIN1 (_________31675), .DIN2 (_________31607),
       .Q (____9_9__31749));
  xor2s1 ___0___438462(.DIN1 (_____00__34333), .DIN2 (____9____30893),
       .Q (____9____31739));
  nor2s1 ___0__438463(.DIN1 (______0__30774), .DIN2 (_________31671),
       .Q (_____99__31723));
  xor2s1 ___0_438464(.DIN1 (_________31657), .DIN2 (_________31983), .Q
       (____90___31726));
  hi1s1 ___0__438465(.DIN (_________31704), .Q (______9__31705));
  nor2s1 ___0___438466(.DIN1 (_____________9___18714), .DIN2
       (_________31702), .Q (_________31703));
  and2s1 ___0___438467(.DIN1 (_________34489), .DIN2
       (_____________9___18714), .Q (_________31701));
  xor2s1 ___0___438468(.DIN1 (_________31644), .DIN2 (_________32644),
       .Q (_________31700));
  and2s1 ___0___438469(.DIN1 (____0____30072), .DIN2
       (_____________9___18714), .Q (_________31699));
  xor2s1 ___0__438470(.DIN1 (_________31697), .DIN2 (_________31674),
       .Q (_________31698));
  nnd2s1 ___0___438471(.DIN1 (_________31661), .DIN2 (________23817),
       .Q (______0__31696));
  xor2s1 ___0___438472(.DIN1 (_________31645), .DIN2 (____0____32777),
       .Q (______9__31695));
  nnd2s1 ___0___438473(.DIN1 (_________31660), .DIN2 (_________31422),
       .Q (_____9___31718));
  nor2s1 ___0___438474(.DIN1 (______0__28686), .DIN2 (_________31666),
       .Q (_________32583));
  nor2s1 ___0___438475(.DIN1 (______9__30334), .DIN2 (_________31664),
       .Q (_____9___31720));
  xor2s1 ___0__438476(.DIN1 (_________31652), .DIN2 (_________31366),
       .Q (____09___33764));
  hi1s1 ___0__438477(.DIN (_________31693), .Q (_________31694));
  and2s1 ___0___438478(.DIN1 (_____00__34333), .DIN2 (_____0___28711),
       .Q (_________31692));
  and2s1 ___0___438479(.DIN1 (______0__31686), .DIN2 (_________31690),
       .Q (_________31691));
  xor2s1 ___0___438480(.DIN1 (_____________18905), .DIN2
       (_________31670), .Q (_________31689));
  xor2s1 ___0___438481(.DIN1 (_________31642), .DIN2 (_________31290),
       .Q (_________31688));
  nnd2s1 ___0___438482(.DIN1 (______0__31686), .DIN2 (outData[30]), .Q
       (_________31687));
  nnd2s1 ___0___438483(.DIN1 (_________31683), .DIN2
       (______________0____________________), .Q (______9__31685));
  nor2s1 ___0___438484(.DIN1 (______________0____________________),
       .DIN2 (_________31683), .Q (_________31684));
  nnd2s1 ___0_438485(.DIN1 (_________31656), .DIN2 (______0__31641), .Q
       (_________31682));
  nor2s1 ___0___438486(.DIN1 (______9__31490), .DIN2 (_________31662),
       .Q (______0__31706));
  nor2s1 ___0___438487(.DIN1 (_________31647), .DIN2 (______9__31668),
       .Q (_____90__31715));
  xor2s1 ___0___438488(.DIN1 (_________28743), .DIN2 (_________31665),
       .Q (_________31680));
  nor2s1 ___0___438489(.DIN1 (______0__31678), .DIN2 (_________31651),
       .Q (_________31679));
  nor2s1 ___0___438490(.DIN1 (________21527), .DIN2 (______9__31649),
       .Q (______9__31677));
  xor2s1 ___0__438491(.DIN1 (_____0___30366), .DIN2 (_________31663),
       .Q (_________31676));
  nnd2s1 ___0__438492(.DIN1 (_________31674), .DIN2 (_____99__31631),
       .Q (_________31675));
  xor2s1 ___0___438493(.DIN1 (_____0___31638), .DIN2 (________19986),
       .Q (_________31704));
  nnd2s1 ___0__438494(.DIN1 (_________31643), .DIN2 (_________31562),
       .Q (_________31673));
  xor2s1 ___0___438495(.DIN1 (_____9___31628), .DIN2 (_____9___32930),
       .Q (_________31672));
  nor2s1 ___0___438496(.DIN1 (_________30741), .DIN2 (_________31670),
       .Q (_________31671));
  nnd2s1 ___0___438497(.DIN1 (______0__31669), .DIN2 (_____0___34425),
       .Q (_________31693));
  nor2s1 ___0___438498(.DIN1 (_____0___34425), .DIN2 (______0__31669),
       .Q (_________31711));
  dffacs1 __________________438499(.CLRB (reset), .CLK (clk), .DIN
       (_________31646), .QN (_________34437));
  nor2s1 ___0___438500(.DIN1 (_________31667), .DIN2 (_____0___31639),
       .Q (______9__31668));
  nor2s1 ___0___438501(.DIN1 (______0__28714), .DIN2 (_________31665),
       .Q (_________31666));
  nor2s1 ___0__438502(.DIN1 (______9__30344), .DIN2 (_________31663),
       .Q (_________31664));
  and2s1 ___0___438503(.DIN1 (_____00__34628), .DIN2 (____0____34551),
       .Q (_________31662));
  nnd2s1 ___0_0_438504(.DIN1 (_____0___31637), .DIN2 (_________31920),
       .Q (_________31661));
  nor2s1 ___0_0_438505(.DIN1 (_________31412), .DIN2 (_____0___31634),
       .Q (_________31660));
  nor2s1 ___0_438506(.DIN1 (______9__31658), .DIN2 (_____0___31636), .Q
       (______0__31659));
  dffacs1 _________________9_438507(.CLRB (reset), .CLK (clk), .DIN
       (_____09__31640), .Q (_____________9___18714));
  xor2s1 ___0__438508(.DIN1 (_____9___31623), .DIN2
       (_________________0___18618), .Q (____0_9__32839));
  nnd2s1 ___0__438509(.DIN1 (_____9___31629), .DIN2 (_________31579),
       .Q (_________31657));
  nor2s1 ___0___438510(.DIN1 (_____0___31537), .DIN2 (____0____34551),
       .Q (_________31656));
  or2s1 ___0__438511(.DIN1
       (______________________________________0_____________18885),
       .DIN2 (____0____34551), .Q (_________31655));
  nnd2s1 ___0__438512(.DIN1 (____0____34551), .DIN2
       (______________________________________0_____________18885), .Q
       (_________31654));
  nor2s1 ___0___438513(.DIN1 (_________31580), .DIN2 (_____9___31624),
       .Q (_________31681));
  nnd2s1 ___0___438514(.DIN1 (_________34309), .DIN2 (_________31653),
       .Q (______0__31686));
  hi1s1 ___0__438515(.DIN (______0__31669), .Q (_________31683));
  or2s1 ___0___438516(.DIN1 (_________31653), .DIN2 (_________34309),
       .Q (_________31690));
  xor2s1 ___0__438517(.DIN1 (______9__30744), .DIN2 (______0__31602),
       .Q (_____00__34333));
  xor2s1 ___0___438518(.DIN1 (_________31367), .DIN2 (_____0___34630),
       .Q (_________31652));
  hi1s1 ___0___438519(.DIN (______0__31650), .Q (_________31651));
  nor2s1 ___0___438520(.DIN1 (_________31648), .DIN2 (_________31620),
       .Q (______9__31649));
  and2s1 ___0___438521(.DIN1 (_________31600), .DIN2 (_________31667),
       .Q (_________31647));
  nnd2s1 ___0___438522(.DIN1 (______9__31621), .DIN2 (_____90__31622),
       .Q (_________31646));
  nor2s1 ___0___438523(.DIN1 (_________31484), .DIN2 (_________31609),
       .Q (_________31933));
  nnd2s1 ___0___438524(.DIN1 (______9__31611), .DIN2 (_________31584),
       .Q (_________31674));
  xor2s1 ___0_0_438525(.DIN1 (_________31586), .DIN2 (_________31610),
       .Q (_________31645));
  nnd2s1 ___0_0_438526(.DIN1 (_____09__31543), .DIN2 (_________31613),
       .Q (_________31644));
  hi1s1 ___0_9_438527(.DIN (_____00__34628), .Q (_________31643));
  xor2s1 ___0___438528(.DIN1 (______0__31641), .DIN2 (____0_9__30961),
       .Q (_________31642));
  nor2s1 ___0___438529(.DIN1 (______9__31601), .DIN2 (_________31608),
       .Q (_________31670));
  xor2s1 ___0___438530(.DIN1 (_________31581), .DIN2 (______0__31641),
       .Q (______0__31669));
  dffacs1 ___________________438531(.CLRB (reset), .CLK (clk), .DIN
       (_________31615), .QN (_________________18713));
  nnd2s1 ___0_0_438532(.DIN1 (_________31594), .DIN2 (_________35044),
       .Q (_____09__31640));
  nor2s1 ___0___438533(.DIN1 (_____9___31527), .DIN2 (______0__31583),
       .Q (_____0___31639));
  nor2s1 ___0_9_438534(.DIN1 (_____00__31632), .DIN2 (_____0___31633),
       .Q (_____0___31638));
  nnd2s1 ___0__438535(.DIN1 (_________31599), .DIN2 (______9__31592),
       .Q (_____0___31637));
  hi1s1 ___0___438536(.DIN (_____0___31635), .Q (_____0___31636));
  nor2s1 ___0___438537(.DIN1 (_________31432), .DIN2 (_____0___34630),
       .Q (_____0___31634));
  nor2s1 ___0___438538(.DIN1 (______0__28406), .DIN2 (_________31598),
       .Q (_________31665));
  nnd2s1 ___0_9_438539(.DIN1 (_____0___31633), .DIN2 (_____00__31632),
       .Q (______0__31650));
  xor2s1 ___0___438540(.DIN1 (_________31572), .DIN2 (_________32554),
       .Q (_________31663));
  xor2s1 ___0_0_438541(.DIN1 (_________________0___18618), .DIN2
       (______9__31573), .Q (____0____32837));
  dffacs1 ___________________438542(.CLRB (reset), .CLK (clk), .DIN
       (_________31595), .QN (_________34478));
  nnd2s1 ___0___438543(.DIN1 (_________31697), .DIN2
       (_____________0___18684), .Q (_____99__31631));
  xor2s1 ___0_438544(.DIN1 (_____9___31627), .DIN2 (_________34362), .Q
       (_____9___31630));
  nnd2s1 ___0__438545(.DIN1 (_________31591), .DIN2 (_________31295),
       .Q (_____9___31629));
  nor2s1 ___0__438546(.DIN1 (_________31590), .DIN2 (_____9___31627),
       .Q (_____9___31628));
  or2s1 ___0___438547(.DIN1
       (______________________________________0_____________18886),
       .DIN2 (______0__31641), .Q (_____9___31626));
  nnd2s1 ___0_9_438548(.DIN1 (______0__31544), .DIN2 (______0__31641),
       .Q (_____9___31625));
  and2s1 ___0___438549(.DIN1 (______0__31641), .DIN2
       (______________________________________0_____________18886), .Q
       (_____9___31624));
  xor2s1 ___0___438550(.DIN1 (_________31566), .DIN2 (outData[31]), .Q
       (_________34309));
  dffacs1 ___________________438551(.CLRB (reset), .CLK (clk), .DIN
       (______0__31593), .QN (_________34465));
  xor2s1 ___0_9_438552(.DIN1 (_________31557), .DIN2 (_________31290),
       .Q (_____9___31623));
  nnd2s1 ___0_438553(.DIN1 (_________31575), .DIN2 (_________31618), .Q
       (_____90__31622));
  nor2s1 ___0___438554(.DIN1 (_________31570), .DIN2 (_________29463),
       .Q (______9__31621));
  xor2s1 ___0___438555(.DIN1 (_____9___28423), .DIN2 (_____0___34632),
       .Q (_________31620));
  nnd2s1 ___0_0_438556(.DIN1 (_________31576), .DIN2 (_________31618),
       .Q (_________31619));
  nor2s1 ___0_9_438557(.DIN1 (_________31616), .DIN2 (_________31596),
       .Q (_________31617));
  nnd2s1 ___0___438558(.DIN1 (_________31310), .DIN2 (_________31571),
       .Q (_________31615));
  nnd2s1 ___0___438559(.DIN1 (_________31577), .DIN2 (_________33103),
       .Q (_________31614));
  xnr2s1 ___0___438560(.DIN1 (_________31134), .DIN2 (_________31547),
       .Q (_____0___31635));
  or2s1 ___0_0_438561(.DIN1 (_________31559), .DIN2 (______0__31612),
       .Q (_________31613));
  nnd2s1 ___0___438562(.DIN1 (_________31610), .DIN2 (_________31585),
       .Q (______9__31611));
  nor2s1 ___0___438563(.DIN1 (________19961), .DIN2 (_________31568),
       .Q (_________31609));
  and2s1 ___0__438564(.DIN1 (______0__31564), .DIN2 (_________30743),
       .Q (_________31608));
  nnd2s1 ___0___438565(.DIN1 (_________31604), .DIN2 (_________31606),
       .Q (_________31607));
  nnd2s1 ___0___438566(.DIN1 (_________31604), .DIN2 (_____0___34426),
       .Q (_________31605));
  nor2s1 ___0___438567(.DIN1 (_____0___34426), .DIN2 (_________31604),
       .Q (_________31603));
  nor2s1 ___0___438568(.DIN1 (_________31565), .DIN2 (______9__31601),
       .Q (______0__31602));
  hi1s1 ___0__438569(.DIN (_________31599), .Q (_________31600));
  nor2s1 ___0___438570(.DIN1 (_________28400), .DIN2 (_____0___34632),
       .Q (_________31598));
  hi1s1 ___0__438571(.DIN (_________31596), .Q (_________31597));
  nnd2s1 ___0___438572(.DIN1 (______0__31554), .DIN2 (____0____31816),
       .Q (_________31595));
  nnd2s1 ___0___438573(.DIN1 (______9__31553), .DIN2 (_________31702),
       .Q (_________31594));
  nnd2s1 ___0___438574(.DIN1 (_________31558), .DIN2 (_____9___31443),
       .Q (______0__31593));
  nnd2s1 ___0_9_438575(.DIN1 (_____00__31536), .DIN2 (_________31552),
       .Q (______9__31592));
  nnd2s1 ___0_0_438576(.DIN1 (______9__31582), .DIN2 (_________31551),
       .Q (_________31599));
  xor2s1 ___0___438577(.DIN1 (_____9___31530), .DIN2 (_____9___31531),
       .Q (_____00__31632));
  nnd2s1 ___0___438578(.DIN1 (_____0___31538), .DIN2 (__9_____26879),
       .Q (_________31591));
  hi1s1 ___0___438579(.DIN (_________31589), .Q (_________31590));
  nor2s1 ___0__438580(.DIN1 (_________31587), .DIN2 (_____0___31540),
       .Q (_________31588));
  nnd2s1 ___0_438581(.DIN1 (_________31585), .DIN2 (_________31584), .Q
       (_________31586));
  nor2s1 ___0___438582(.DIN1 (_____9___31528), .DIN2 (______9__31582),
       .Q (______0__31583));
  xor2s1 ___0___438583(.DIN1 (_________31580), .DIN2
       (______________________________________0_____________18886), .Q
       (_________31581));
  nnd2s1 ___0___438584(.DIN1 (_____0___31542), .DIN2 (______0__35078),
       .Q (_________31579));
  hi1s1 ___0_0_438585(.DIN (_________31604), .Q (_________31697));
  xnr2s1 ___0___438586(.DIN1 (_________31578), .DIN2 (_________31524),
       .Q (______0__31641));
  xor2s1 ___0___438587(.DIN1 (_________31515), .DIN2 (______9__33247),
       .Q (_________31577));
  nnd2s1 ___0___438588(.DIN1 (______0__31574), .DIN2 (inData[14]), .Q
       (_________31576));
  nnd2s1 ___0___438589(.DIN1 (______0__31574), .DIN2 (_________31497),
       .Q (_________31575));
  nor2s1 ___0___438590(.DIN1 (_____9___31532), .DIN2 (_________31499),
       .Q (______9__31573));
  nor2s1 ___0___438591(.DIN1 (______0__30188), .DIN2 (_____9___31534),
       .Q (_________31572));
  nnd2s1 ___0_9_438592(.DIN1 (________20192), .DIN2 (______9__31525),
       .Q (_________31571));
  and2s1 ___0___438593(.DIN1 (_________31569), .DIN2 (_________34437),
       .Q (_________31570));
  xor2s1 ___0___438594(.DIN1 (_________31518), .DIN2 (_________31951),
       .Q (_________31596));
  nor2s1 ___0___438595(.DIN1 (_____0___31539), .DIN2 (_________31523),
       .Q (_________31610));
  nor2s1 ___0___438596(.DIN1 (____0___23530), .DIN2 (_________31521),
       .Q (_________31568));
  xor2s1 ___0__438597(.DIN1 (_____0___31541), .DIN2 (____009__31815),
       .Q (_________31567));
  nor2s1 ___0_0_438598(.DIN1 (______9__31563), .DIN2 (_________31565),
       .Q (_________31566));
  or2s1 ___0_9_438599(.DIN1 (_____________18905), .DIN2
       (_________31565), .Q (______0__31564));
  nor2s1 ___0_9_438600(.DIN1 (outData[31]), .DIN2 (______9__31563), .Q
       (______9__31601));
  nnd2s1 ___0___438601(.DIN1 (_________31560), .DIN2 (_________31561),
       .Q (_________31589));
  hi1s1 ___0___438602(.DIN (_________31562), .Q (______0__31612));
  nor2s1 ___0___438603(.DIN1 (_________31561), .DIN2 (_________31560),
       .Q (_____9___31627));
  dffacs1 __________________438604(.CLRB (reset), .CLK (clk), .DIN
       (_____99__31535), .QN (_________34469));
  xor2s1 ___0___438605(.DIN1 (______0__31501), .DIN2 (_________31559),
       .Q (_________31604));
  nor2s1 ___0___438606(.DIN1 (_________31516), .DIN2 (_________31105),
       .Q (_________31558));
  xor2s1 ___0___438607(.DIN1 (_________31492), .DIN2 (_________31559),
       .Q (_________31557));
  hi1s1 ___0_438608(.DIN (_________31555), .Q (_________31556));
  nor2s1 ___0_9_438609(.DIN1 (____9___20317), .DIN2 (_________31514),
       .Q (______0__31554));
  xor2s1 ___0_9_438610(.DIN1 (_________30192), .DIN2 (_____9___31533),
       .Q (______9__31553));
  hi1s1 ___0___438611(.DIN (_________31551), .Q (_________31552));
  or2s1 ___0__438612(.DIN1 (_________31549), .DIN2 (_________31548), .Q
       (_________31550));
  nor2s1 ___0___438613(.DIN1 (_________31545), .DIN2 (_________31546),
       .Q (______9__31658));
  nnd2s1 ___0___438614(.DIN1 (_________31546), .DIN2 (_________31545),
       .Q (_________31547));
  hi1s1 ___0__438615(.DIN (_____09__31543), .Q (______0__31544));
  nor2s1 ___0___438616(.DIN1 (__9_0___26991), .DIN2 (_____0___31541),
       .Q (_____0___31542));
  nor2s1 ___0__438617(.DIN1 (_____0___31539), .DIN2 (_________31522),
       .Q (_____0___31540));
  nnd2s1 ___0___438618(.DIN1 (_____0___31541), .DIN2 (__9_____26878),
       .Q (_____0___31538));
  nnd2s1 ___0___438619(.DIN1 (_________31504), .DIN2
       (______________0______________________18825), .Q
       (_________31585));
  nor2s1 ___0___438620(.DIN1 (_____0___35109), .DIN2 (_____0___31537),
       .Q (_________31562));
  hi1s1 ___0_0_438621(.DIN (_____00__31536), .Q (______9__31582));
  dffacs1 ___________________438622(.CLRB (reset), .CLK (clk), .DIN
       (_________31509), .QN (_________________18726));
  nnd2s1 ___0___438623(.DIN1 (_________31480), .DIN2 (_________31303),
       .Q (_____99__31535));
  and2s1 ___0___438624(.DIN1 (_____9___31533), .DIN2 (_____00__30178),
       .Q (_____9___31534));
  nor2s1 ___0_9_438625(.DIN1 (_____9___31531), .DIN2 (_________31496),
       .Q (_____9___31532));
  nnd2s1 ___0_9_438626(.DIN1 (_________31494), .DIN2 (_________31495),
       .Q (_____9___31530));
  and2s1 ___0_9_438627(.DIN1 (______9__32872), .DIN2 (_________33444),
       .Q (_____9___31529));
  nor2s1 ___0___438628(.DIN1 (_________31498), .DIN2 (_________33103),
       .Q (_________31569));
  nor2s1 ___0___438629(.DIN1 (_____9___31528), .DIN2 (_____9___31527),
       .Q (_________31551));
  xor2s1 ___0_0_438630(.DIN1 (_________31475), .DIN2 (_____90__31526),
       .Q (_________31555));
  nor2s1 ___0___438631(.DIN1 (_________31493), .DIN2 (________22915),
       .Q (______0__31574));
  xor2s1 ___0___438632(.DIN1 (____00___34537), .DIN2 (___0___18982), .Q
       (______9__31525));
  xor2s1 ___0_438633(.DIN1 (_________31469), .DIN2 (____0____31818), .Q
       (_________31524));
  nor2s1 ___0_9_438634(.DIN1 (_________________18683), .DIN2
       (_________31522), .Q (_________31523));
  nor2s1 ___0_0_438635(.DIN1 (____0____31820), .DIN2 (_________31485),
       .Q (_________31521));
  nor2s1 ___0___438636(.DIN1 (_________31433), .DIN2 (_________31483),
       .Q (_________31561));
  nor2s1 ___0___438637(.DIN1 (_________31519), .DIN2 (_________31520),
       .Q (______9__31563));
  nnd2s1 ___0___438638(.DIN1 (______0__31491), .DIN2 (______9__31500),
       .Q (_____09__31543));
  nor2s1 ___0___438639(.DIN1 (______9__31389), .DIN2 (______0__31482),
       .Q (_________31580));
  nnd2s1 ___0__438640(.DIN1 (_________31487), .DIN2 (_____9___31437),
       .Q (_____00__31536));
  and2s1 ___0___438641(.DIN1 (_________31520), .DIN2 (_________31519),
       .Q (_________31565));
  nnd2s1 ___0_0_438642(.DIN1 (_________31512), .DIN2 (_________31513),
       .Q (_________31518));
  and2s1 ___0___438643(.DIN1 (_________31464), .DIN2 (_________31476),
       .Q (_________31516));
  xor2s1 ___0_438644(.DIN1 (_________31457), .DIN2
       (________________18756), .Q (_________31515));
  nor2s1 ___0___438645(.DIN1 (_________31587), .DIN2 (_________31472),
       .Q (_________31514));
  nor2s1 ___0_0_438646(.DIN1 (_________31513), .DIN2 (_________31512),
       .Q (_________31616));
  and2s1 ___0__438647(.DIN1 (______9__31510), .DIN2 (______0__31511),
       .Q (_________31548));
  nor2s1 ___0___438648(.DIN1 (______0__31511), .DIN2 (______9__31510),
       .Q (_________31549));
  nnd2s1 ___0___438649(.DIN1 (______9__31465), .DIN2 (_________31403),
       .Q (_________31509));
  nor2s1 ___0___438650(.DIN1 (_________31505), .DIN2 (_________31506),
       .Q (_________31508));
  nnd2s1 ___0___438651(.DIN1 (_________31506), .DIN2 (_________31505),
       .Q (_________31507));
  xor2s1 ___0___438652(.DIN1 (_________31502), .DIN2 (_________35002),
       .Q (_________31504));
  xor2s1 ___0_9_438653(.DIN1 (_________31502), .DIN2 (_____0___34427),
       .Q (_________31503));
  xor2s1 ___0_9_438654(.DIN1 (______9__31481), .DIN2 (_________31388),
       .Q (______0__31501));
  hi1s1 ___0__438655(.DIN (______9__31500), .Q (_____0___31537));
  nor2s1 ___0___438656(.DIN1 (_________31398), .DIN2 (_________31471),
       .Q (_____0___31539));
  xor2s1 ___0___438657(.DIN1 (________20547), .DIN2 (_________34299),
       .Q (_________31560));
  nor2s1 ___0__438658(.DIN1 (_________29844), .DIN2 (_________31463),
       .Q (_________31545));
  nnd2s1 ___0___438659(.DIN1 (_________31467), .DIN2 (_________31468),
       .Q (_____0___31541));
  and2s1 ___0___438660(.DIN1 (_____9___28417), .DIN2
       (_______________0__________________0), .Q (_________31499));
  nnd2s1 ___0_0_438661(.DIN1 (_______________0__________________0),
       .DIN2 (_________________18766), .Q (_________31498));
  or2s1 ___0_0_438662(.DIN1 (_______________0__________________0),
       .DIN2 (_________34437), .Q (_________31497));
  nor2s1 ___0___438663(.DIN1 (_______________0__________________0),
       .DIN2 (______0__31456), .Q (_________31496));
  or2s1 ___0___438664(.DIN1 (_______________0__________________0),
       .DIN2 (____9_9__29949), .Q (_________31495));
  nnd2s1 ___0___438665(.DIN1 (______0__28475), .DIN2
       (_______________0__________________0), .Q (_________31494));
  nor2s1 ___0_0_438666(.DIN1 (_________________18766), .DIN2
       (_______________0__________________0), .Q (_________31493));
  nnd2s1 ___0__438667(.DIN1 (______0__31491), .DIN2 (_____9___31263),
       .Q (_________31492));
  nor2s1 ___0___438668(.DIN1 (_________35111), .DIN2 (______0__31491),
       .Q (______9__31490));
  nor2s1 ___0___438669(.DIN1 (_________34686), .DIN2 (_________31489),
       .Q (_____9___31528));
  and2s1 ___0__438670(.DIN1 (_________31489), .DIN2 (_________34686),
       .Q (_____9___31527));
  nor2s1 ___0___438671(.DIN1 (_________28754), .DIN2 (_________31458),
       .Q (______9__32872));
  nnd2s1 ___0_0_438672(.DIN1 (_________31502), .DIN2 (__9), .Q
       (_________31488));
  or2s1 ___0___438673(.DIN1 (_________31486), .DIN2 (_____00__31446),
       .Q (_________31487));
  or2s1 ___0___438674(.DIN1 (_________30807), .DIN2 (_________34299),
       .Q (_________31485));
  and2s1 ___0___438675(.DIN1 (_________34299), .DIN2 (________23870),
       .Q (_________31484));
  nor2s1 ___0___438676(.DIN1 (____0____32823), .DIN2 (_____99__31445),
       .Q (_________31483));
  nor2s1 ___0_0_438677(.DIN1 (_________31387), .DIN2 (______9__31481),
       .Q (______0__31482));
  nor2s1 ___0___438678(.DIN1 (_____0___31453), .DIN2 (_____99__30455),
       .Q (_________31480));
  nnd2s1 ___0___438679(.DIN1 (_____0___31449), .DIN2 (_________31417),
       .Q (_________31520));
  xor2s1 ___0_9_438680(.DIN1 (_________31429), .DIN2 (_________31479),
       .Q (______9__31500));
  nor2s1 ___0___438681(.DIN1 (_________31435), .DIN2 (_________31470),
       .Q (_________31522));
  nor2s1 ___0___438682(.DIN1 (_____0___30100), .DIN2 (_____0___31452),
       .Q (_____9___31533));
  dffacs1 ___________________438683(.CLRB (reset), .CLK (clk), .DIN
       (_____9___31444), .QN (_________34463));
  dffacs1 __________________438684(.CLRB (reset), .CLK (clk), .DIN
       (_____09__31455), .QN (_________34447));
  nnd2s1 ___0_9_438685(.DIN1 (_________31383), .DIN2 (_____9___31440),
       .Q (_________31476));
  xor2s1 ___0___438686(.DIN1 (_________31397), .DIN2 (_________31459),
       .Q (_________31475));
  xnr2s1 ___0__438687(.DIN1 (_________35110), .DIN2 (______9__31473),
       .Q (______0__31474));
  xor2s1 ___0___438688(.DIN1 (_________30116), .DIN2 (_____0___31451),
       .Q (_________31472));
  nor2s1 ___0___438689(.DIN1 (______9__31343), .DIN2 (_____9___31441),
       .Q (______0__31511));
  xor2s1 ___0___438690(.DIN1 (_________28755), .DIN2 (_________32216),
       .Q (_________31512));
  xor2s1 ___0___438691(.DIN1 (______9__31426), .DIN2 (______9__33856),
       .Q (_________31513));
  hi1s1 ___0__438692(.DIN (_________31470), .Q (_________31471));
  nnd2s1 ___0__438693(.DIN1 (______0__31466), .DIN2 (_________31468),
       .Q (_________31469));
  nnd2s1 ___0___438694(.DIN1 (______0__31466), .DIN2 (____0____31818),
       .Q (_________31467));
  or2s1 ___0___438695(.DIN1 (_________31464), .DIN2 (_________31430),
       .Q (______9__31465));
  nnd2s1 ___0_0_438696(.DIN1 (_____9___31439), .DIN2 (_________29852),
       .Q (_________31463));
  nnd2s1 ___0_0_438697(.DIN1 (_________31460), .DIN2 (_____0___34427),
       .Q (_________31462));
  nnd2s1 ___0___438698(.DIN1 (_____9___31442), .DIN2 (_________31461),
       .Q (_________31506));
  or2s1 ___0___438699(.DIN1
       (______________0______________________18825), .DIN2
       (_________31460), .Q (_________31584));
  nor2s1 ___0___438700(.DIN1 (_________31434), .DIN2 (_________31459),
       .Q (_________31517));
  dffacs1 ___________________438701(.CLRB (reset), .CLK (clk), .DIN
       (_____9___31438), .QN (_________________18696));
  nor2s1 ___0___438702(.DIN1 (_________28753), .DIN2 (_________32216),
       .Q (_________31458));
  xor2s1 ___0___438703(.DIN1 (_____0___34634), .DIN2 (______0__31456),
       .Q (_________31457));
  nnd2s1 ___0___438704(.DIN1 (_________31428), .DIN2 (_____0___31454),
       .Q (_____09__31455));
  nor2s1 ___0_0_438705(.DIN1 (_________31424), .DIN2 (_________31241),
       .Q (_____0___31453));
  and2s1 ___0_9_438706(.DIN1 (_____0___31451), .DIN2 (____09___30090),
       .Q (_____0___31452));
  xor2s1 ___0___438707(.DIN1 (_________31407), .DIN2 (______0__28597),
       .Q (______9__31510));
  xor2s1 ___0___438708(.DIN1 (_________18863), .DIN2 (____9____29918),
       .Q (_________31489));
  xor2s1 ___0___438709(.DIN1 (_________31402), .DIN2 (_____0___31450),
       .Q (______0__31491));
  dffacs1 __________________438710(.CLRB (reset), .CLK (clk), .DIN
       (______0__31427), .QN (_______________0__________________0));
  nor2s1 ___0_0_438711(.DIN1 (____0_9__30931), .DIN2 (______9__31418),
       .Q (_____0___31449));
  nnd2s1 ___0___438712(.DIN1 (_____0___31447), .DIN2 (_________31393),
       .Q (_____0___31448));
  nor2s1 ___0___438713(.DIN1 (_________29878), .DIN2 (_________31420),
       .Q (_____00__31446));
  nor2s1 ___0___438714(.DIN1 (_____9___31346), .DIN2 (_________31413),
       .Q (_____99__31445));
  nnd2s1 ___0___438715(.DIN1 (_________31425), .DIN2 (_____9___31443),
       .Q (_____9___31444));
  nor2s1 ___0__438716(.DIN1 (______9__31246), .DIN2 (_________31415),
       .Q (______9__31481));
  nnd2s1 ___0___438717(.DIN1 (_________31421), .DIN2 (_________31377),
       .Q (_________31470));
  hi1s1 ___0___438718(.DIN (_________31460), .Q (_________31502));
  xor2s1 ___0_9_438719(.DIN1 (_________31394), .DIN2 (____0____30930),
       .Q (_________34299));
  hi1s1 ___0___438720(.DIN (_____0___31447), .Q (_____9___31442));
  nnd2s1 ___0_9_438721(.DIN1 (_________31404), .DIN2 (_________31338),
       .Q (_____9___31441));
  or2s1 ___0___438722(.DIN1 (_________34469), .DIN2 (______0__31400),
       .Q (_____9___31440));
  nnd2s1 ___0___438723(.DIN1 (_________29888), .DIN2 (_________18863),
       .Q (_____9___31439));
  nnd2s1 ___0__438724(.DIN1 (_________31408), .DIN2 (________20959), .Q
       (_____9___31438));
  nnd2s1 ___0__438725(.DIN1 (_________31391), .DIN2 (_________31486),
       .Q (_____9___31437));
  and2s1 ___0__438726(.DIN1 (_________28367), .DIN2 (_____0___34634),
       .Q (_________31477));
  xor2s1 ___0___438727(.DIN1 (_________31435), .DIN2
       (_________________18793), .Q (______9__31436));
  xor2s1 ___0___438728(.DIN1 (_________31362), .DIN2
       (_________________0___18607), .Q (_________31434));
  and2s1 ___0__438729(.DIN1 (_________31396), .DIN2 (____0____32823),
       .Q (_________31433));
  xor2s1 ___0___438730(.DIN1 (_________31368), .DIN2 (_________31431),
       .Q (_________31432));
  xor2s1 ___0___438731(.DIN1 (______0__31419), .DIN2 (______0__31390),
       .Q (_________31430));
  nor2s1 ___0__438732(.DIN1 (_______________18884), .DIN2
       (_________31386), .Q (_________31429));
  nnd2s1 ___0___438733(.DIN1 (_________31385), .DIN2
       (______________________________________0_____________18885), .Q
       (______0__31466));
  xor2s1 ___0___438734(.DIN1 (_________31414), .DIN2 (_________31282),
       .Q (_________31460));
  nor2s1 ___0__438735(.DIN1 (___0____20744), .DIN2 (_________31381), .Q
       (_________31428));
  nnd2s1 ___0___438736(.DIN1 (_________31375), .DIN2 (________24033),
       .Q (______0__31427));
  nnd2s1 ___0_438737(.DIN1 (______0__31380), .DIN2 (_________28598), .Q
       (______9__31426));
  nor2s1 ___0___438738(.DIN1 (________22857), .DIN2 (______0__31370),
       .Q (_________31425));
  xor2s1 ___0___438739(.DIN1 (_________31423), .DIN2 (_________31382),
       .Q (_________31424));
  xor2s1 ___0___438740(.DIN1 (______0__34638), .DIN2 (_________32410),
       .Q (_____0___31451));
  xor2s1 ___0___438741(.DIN1 (_____0___31355), .DIN2 (______0__35008),
       .Q (______9__31473));
  xor2s1 ___0__438742(.DIN1 (_____0___31356), .DIN2 (____9___19200), .Q
       (_________31459));
  xor2s1 ___0__438743(.DIN1 (_________31284), .DIN2 (_________31401),
       .Q (_________32216));
  nnd2s1 ___0___438744(.DIN1 (_________31411), .DIN2 (_________32606),
       .Q (_________31422));
  nnd2s1 ___0_0_438745(.DIN1 (______9__31369), .DIN2 (_________31376),
       .Q (_________31421));
  nor2s1 ___0__438746(.DIN1 (_________29879), .DIN2 (______0__31419),
       .Q (_________31420));
  nor2s1 ___0___438747(.DIN1 (_________31431), .DIN2 (_________31416),
       .Q (______9__31418));
  nnd2s1 ___0___438748(.DIN1 (_________31416), .DIN2 (_________35110),
       .Q (_________31417));
  and2s1 ___0___438749(.DIN1 (_________31414), .DIN2 (______0__31247),
       .Q (_________31415));
  nor2s1 ___0___438750(.DIN1 (_________31395), .DIN2 (_________31361),
       .Q (_________31413));
  nor2s1 ___0___438751(.DIN1 (_________32606), .DIN2 (_________31411),
       .Q (_________31412));
  nnd2s1 ___0___438752(.DIN1 (_________31384), .DIN2 (_____00__30456),
       .Q (_________31468));
  xor2s1 ___0_9_438753(.DIN1 (_____9___31348), .DIN2 (_____9___31345),
       .Q (_____0___31447));
  dffacs1 ___________________438754(.CLRB (reset), .CLK (clk), .DIN
       (_________31371), .QN (_________34464));
  hi1s1 ___0__438755(.DIN (______9__31409), .Q (______0__31410));
  nnd2s1 ___0_438756(.DIN1 (_____9___31349), .DIN2 (__99____27118), .Q
       (_________31408));
  xor2s1 ___0___438757(.DIN1 (________18841), .DIN2 (_________31405),
       .Q (_________31407));
  xor2s1 ___0___438758(.DIN1 (_________________18732), .DIN2
       (_________31405), .Q (_________31406));
  or2s1 ___0___438759(.DIN1 (_________________18748), .DIN2
       (_____0___31357), .Q (_________31404));
  nnd2s1 ___0___438760(.DIN1 (___0____23477), .DIN2 (_____00__31354),
       .Q (_________31403));
  and2s1 ___0___438761(.DIN1 (_________31401), .DIN2 (_________31244),
       .Q (_________31402));
  nor2s1 ___0___438762(.DIN1 (_________34466), .DIN2 (_________31423),
       .Q (______0__31400));
  nor2s1 ___0___438763(.DIN1 (_____0___31358), .DIN2 (______0__31309),
       .Q (_________32352));
  dffacs1 ___________________438764(.CLRB (reset), .CLK (clk), .DIN
       (_____0___34636), .QN (_________18863));
  or2s1 ___0__438765(.DIN1 (_________________18793), .DIN2
       (_________31398), .Q (______9__31399));
  xor2s1 ___0___438766(.DIN1 (_________31364), .DIN2 (_________31363),
       .Q (_________31397));
  nor2s1 ___0___438767(.DIN1 (_________31395), .DIN2 (______0__31360),
       .Q (_________31396));
  xor2s1 ___0___438768(.DIN1 (____0____30949), .DIN2 (_________34640),
       .Q (_________31394));
  hi1s1 ___0___438769(.DIN (_________31461), .Q (_________31393));
  nnd2s1 ___0__438770(.DIN1 (_________31398), .DIN2
       (_________________18793), .Q (_________31392));
  nor2s1 ___0___438771(.DIN1 (______0__31390), .DIN2 (_____0___31359),
       .Q (_________31391));
  and2s1 ___0___438772(.DIN1 (_________31559), .DIN2 (_________31388),
       .Q (______9__31389));
  nor2s1 ___0___438773(.DIN1 (_________31388), .DIN2 (_________31559),
       .Q (_________31387));
  nor2s1 ___0_9_438774(.DIN1 (______9__31219), .DIN2 (_________31559),
       .Q (_________31386));
  hi1s1 ___09_0(.DIN (_________31384), .Q (_________31385));
  dffacs1 ___________________438775(.CLRB (reset), .CLK (clk), .DIN
       (_____9___31350), .Q (_________________18695));
  nnd2s1 ___0___438776(.DIN1 (_________31382), .DIN2 (_________34467),
       .Q (_________31383));
  and2s1 ___0___438777(.DIN1 (_________31341), .DIN2 (_________33186),
       .Q (_________31381));
  or2s1 ___0___438778(.DIN1 (_________28587), .DIN2 (_________31405),
       .Q (______0__31380));
  and2s1 ___0__438779(.DIN1 (_________31405), .DIN2
       (_________________18732), .Q (______9__31379));
  nor2s1 ___0__438780(.DIN1 (_________________18732), .DIN2
       (_________31405), .Q (_________31378));
  or2s1 ___0__438781(.DIN1 (_________31376), .DIN2 (_________31331), .Q
       (_________31377));
  nnd2s1 ___0___438782(.DIN1 (_________31342), .DIN2 (_________33103),
       .Q (_________31375));
  and2s1 ___0___438783(.DIN1 (_________31373), .DIN2 (_________34467),
       .Q (_________31374));
  nor2s1 ___0___438784(.DIN1 (_________34467), .DIN2 (_________31373),
       .Q (_________31372));
  nnd2s1 ___0_0_438785(.DIN1 (_________31340), .DIN2 (_____9___31443),
       .Q (_________31371));
  nor2s1 ___0___438786(.DIN1 (_________31464), .DIN2 (_________31329),
       .Q (______0__31370));
  xor2s1 ___0___438787(.DIN1 (_________31320), .DIN2
       (_________________18748), .Q (______9__31409));
  nor2s1 ___0__438788(.DIN1 (_________31297), .DIN2 (______9__31333),
       .Q (______9__31369));
  or2s1 ___090_(.DIN1 (_________31367), .DIN2 (_________31366), .Q
       (_________31368));
  nnd2s1 ___0___438789(.DIN1 (_________31364), .DIN2 (_________31363),
       .Q (_________31365));
  nor2s1 ___0__438790(.DIN1 (_________31363), .DIN2 (_________31364),
       .Q (_________31362));
  hi1s1 ___0_9_438791(.DIN (______0__31360), .Q (_________31361));
  nnd2s1 ___09__(.DIN1 (_________31327), .DIN2 (_________31162), .Q
       (_________31414));
  nor2s1 ___090_438792(.DIN1 (____0____30927), .DIN2 (_________34640),
       .Q (_________31416));
  nnd2s1 ___090_438793(.DIN1 (_________31366), .DIN2 (_________31367),
       .Q (_________31411));
  nnd2s1 ___09_9(.DIN1 (_________31335), .DIN2 (__9__9__26911), .Q
       (_________31384));
  hi1s1 ___0___438794(.DIN (_____0___31359), .Q (______0__31419));
  hi1s1 ___09__438795(.DIN (_________31398), .Q (_________31435));
  nor2s1 ___0__438796(.DIN1 (_________31225), .DIN2 (_________31328),
       .Q (_________31461));
  dffacs1 __________________438797(.CLRB (reset), .CLK (clk), .DIN
       (_________31339), .Q (________________18756));
  nor2s1 ___0__438798(.DIN1 (____00___34539), .DIN2 (_________31322),
       .Q (_____0___31358));
  xor2s1 ___0___438799(.DIN1 (_________31307), .DIN2 (_________32644),
       .Q (_____0___31357));
  nor2s1 ___0___438800(.DIN1 (_________31202), .DIN2 (______0__31317),
       .Q (_____0___31356));
  xor2s1 ___0___438801(.DIN1 (_________31301), .DIN2 (______9__31316),
       .Q (_____0___31355));
  xnr2s1 ___0___438802(.DIN1 (___0____19798), .DIN2
       (_________________18725), .Q (_____00__31354));
  xor2s1 ___0_9_438803(.DIN1 (_________31305), .DIN2 (_____99__31353),
       .Q (_________31401));
  hi1s1 ___0_438804(.DIN (_________34467), .Q (_________31423));
  xnr2s1 ___0___438805(.DIN1 (_________________18725), .DIN2
       (_____9___31351), .Q (_____9___31352));
  nnd2s1 ___0___438806(.DIN1 (_________31315), .DIN2 (_____0__20540),
       .Q (_____9___31350));
  xor2s1 ___0__438807(.DIN1 (_________31332), .DIN2 (_________31330),
       .Q (_____9___31349));
  xor2s1 ___0___438808(.DIN1 (_____9___31347), .DIN2 (_________31395),
       .Q (_____9___31348));
  nor2s1 ___0_9_438809(.DIN1 (_____9___31345), .DIN2 (_____90__31344),
       .Q (_____9___31346));
  nnd2s1 ___090_438810(.DIN1 (_____90__31344), .DIN2 (_____9___31345),
       .Q (______0__31360));
  nnd2s1 ___0___438811(.DIN1 (_________31314), .DIN2 (_________31079),
       .Q (_____0___31359));
  xor2s1 ___09__438812(.DIN1 (_________31135), .DIN2 (_________31300),
       .Q (_________31398));
  dffacs1 __________________438813(.CLRB (reset), .CLK (clk), .DIN
       (______9__31324), .QN (________________18754));
  xnr2s1 ___09__438814(.DIN1 (______0__31334), .DIN2 (__9__0__26912),
       .Q (_________31559));
  nor2s1 ___0_0_438815(.DIN1 (_________31336), .DIN2 (_________31337),
       .Q (______9__31343));
  xor2s1 ___0___438816(.DIN1 (_________31294), .DIN2 (_________34706),
       .Q (_________31342));
  xor2s1 ___0___438817(.DIN1 (______9__31308), .DIN2 (_________31321),
       .Q (_________31341));
  nor2s1 ___0___438818(.DIN1 (________22751), .DIN2 (_________31302),
       .Q (_________31340));
  nnd2s1 ___0__438819(.DIN1 (_________31312), .DIN2 (_____9__21316), .Q
       (_________31339));
  nnd2s1 ___0_438820(.DIN1 (_________31337), .DIN2 (_________31336), .Q
       (_________31338));
  dffacs1 ________________9_438821(.CLRB (reset), .CLK (clk), .DIN
       (_________31304), .Q (_________34467));
  xor2s1 ___0_9_438822(.DIN1 (_________31291), .DIN2 (_________31136),
       .Q (_________31405));
  or2s1 ___09__438823(.DIN1 (__9_____26761), .DIN2 (______0__31334), .Q
       (_________31335));
  and2s1 ___0___438824(.DIN1 (_________31332), .DIN2 (_________31216),
       .Q (______9__31333));
  nnd2s1 ___0___438825(.DIN1 (_________31332), .DIN2 (_________31330),
       .Q (_________31331));
  xor2s1 ___0__438826(.DIN1 (_____9___31091), .DIN2 (_________31313),
       .Q (_________31329));
  nor2s1 ___09__438827(.DIN1 (_____9__19881), .DIN2 (______9__31298),
       .Q (_________31328));
  xor2s1 ___09__438828(.DIN1 (______0__31286), .DIN2 (_________31486),
       .Q (_________31327));
  nor2s1 ___09__438829(.DIN1 (______9__31237), .DIN2 (______0__31299),
       .Q (_________31366));
  xor2s1 ___090_438830(.DIN1 (_________31283), .DIN2 (_________31326),
       .Q (_________31364));
  nnd2s1 ___0_9_438831(.DIN1 (______9__31024), .DIN2 (_________31296),
       .Q (______9__31324));
  nor2s1 ___0___438832(.DIN1 (_________31255), .DIN2 (_________31321),
       .Q (_________31322));
  xor2s1 ___0___438833(.DIN1 (_________31318), .DIN2 (_________31306),
       .Q (_________31320));
  xor2s1 ___0__438834(.DIN1 (____0___21450), .DIN2 (_________31318), .Q
       (_________31319));
  nor2s1 ___0___438835(.DIN1 (_____00__31269), .DIN2 (______9__31316),
       .Q (______0__31317));
  nnd2s1 ___0___438836(.DIN1 (_________31285), .DIN2 (__99____27118),
       .Q (_________31315));
  or2s1 ___0_438837(.DIN1 (_________31070), .DIN2 (_________31313), .Q
       (_________31314));
  xor2s1 ___0___438838(.DIN1 (_____0___31271), .DIN2 (_________31256),
       .Q (______0__33506));
  hi1s1 ___09__438839(.DIN (_____9___31347), .Q (_____90__31344));
  nnd2s1 ___0_438840(.DIN1 (_____09__31277), .DIN2 (_________33186), .Q
       (_________31312));
  nnd2s1 ___0___438841(.DIN1 (_________31318), .DIN2 (____0___21449),
       .Q (_________31311));
  nnd2s1 ___0___438842(.DIN1 (_____0___31273), .DIN2 (__99____27118),
       .Q (_________31310));
  and2s1 ___0___438843(.DIN1 (______9__31308), .DIN2 (______0__31254),
       .Q (______0__31309));
  nnd2s1 ___0___438844(.DIN1 (_________31318), .DIN2 (_________31306),
       .Q (_________31307));
  nor2s1 ___0___438845(.DIN1 (_________31116), .DIN2 (_____0___31276),
       .Q (_________31305));
  nnd2s1 ___0___438846(.DIN1 (_____0___31274), .DIN2 (_________31303),
       .Q (_________31304));
  nor2s1 ___0___438847(.DIN1 (_________31306), .DIN2 (_________31318),
       .Q (_________31337));
  dffacs1 ___________________438848(.CLRB (reset), .CLK (clk), .DIN
       (_________31279), .QN (_________________18725));
  nor2s1 ___0_9_438849(.DIN1 (_________31464), .DIN2 (_____99__31268),
       .Q (_________31302));
  xor2s1 ___090_438850(.DIN1 (____00___34538), .DIN2 (_________31203),
       .Q (_________31301));
  xnr2s1 ____00_(.DIN1 (_______________18879), .DIN2 (_________34642),
       .Q (_________31300));
  nor2s1 ___09__438851(.DIN1 (____0____30965), .DIN2 (_____9___31265),
       .Q (______0__31299));
  nor2s1 ___09__438852(.DIN1 (________22649), .DIN2 (_____9___31267),
       .Q (______9__31298));
  nor2s1 ___099_(.DIN1 (_________31218), .DIN2 (_____9___31264), .Q
       (______0__31334));
  nor2s1 ___099_438853(.DIN1 (_________31215), .DIN2 (_________31297),
       .Q (_________31330));
  xor2s1 ___09__438854(.DIN1 (_________31248), .DIN2 (____9____30848),
       .Q (_____9___31347));
  xor2s1 ___09__438855(.DIN1 (_________31249), .DIN2 (____9___19200),
       .Q (_________31332));
  nnd2s1 ___0___438856(.DIN1 (______9__31262), .DIN2 (inData[10]), .Q
       (_________31296));
  nnd2s1 ___0__438857(.DIN1 (______0__31278), .DIN2 (_________31288),
       .Q (_________31294));
  nnd2s1 ___0___438858(.DIN1 (_____0___31272), .DIN2
       (_________________18731), .Q (______0__31293));
  hi1s1 ___0___438859(.DIN (_________33440), .Q (______9__31292));
  xor2s1 ___0___438860(.DIN1 (_____0___31275), .DIN2 (_________31290),
       .Q (_________31291));
  nor2s1 ___0___438861(.DIN1 (_____0___31099), .DIN2 (_________31260),
       .Q (_________31321));
  nnd2s1 ___0___438862(.DIN1 (_________31288), .DIN2 (_________34706),
       .Q (_________31323));
  nnd2s1 ____0_0(.DIN1 (_________34642), .DIN2 (_________31112), .Q
       (______0__31286));
  xor2s1 ___09_438863(.DIN1 (____0____34556), .DIN2 (_________31151),
       .Q (_________31285));
  xor2s1 ____0_438864(.DIN1 (______9__31219), .DIN2 (________24537), .Q
       (_________31284));
  xor2s1 ___09__438865(.DIN1 (_________31224), .DIN2 (_________31220),
       .Q (_________31283));
  xnr2s1 ____00_438866(.DIN1 (_________31281), .DIN2 (______9__31219),
       .Q (_________31282));
  xor2s1 ____009(.DIN1 (_________31217), .DIN2 (____00___31810), .Q
       (_________31280));
  nor2s1 ___09_438867(.DIN1 (______0__31121), .DIN2 (_________31250),
       .Q (_________31313));
  nor2s1 ___090_438868(.DIN1 (_____0___31270), .DIN2 (_________31257),
       .Q (______9__31316));
  dffacs1 ___________________438869(.CLRB (reset), .CLK (clk), .DIN
       (_________31251), .QN (______9__34490));
  nnd2s1 ___09__438870(.DIN1 (_________31243), .DIN2 (___0____23478),
       .Q (_________31279));
  xor2s1 ___0___438871(.DIN1 (_____0___31100), .DIN2 (_________31259),
       .Q (_____09__31277));
  nor2s1 ___0900(.DIN1 (_________31115), .DIN2 (_____0___31275), .Q
       (_____0___31276));
  nor2s1 ___0___438872(.DIN1 (_________31242), .DIN2 (____0____30964),
       .Q (_____0___31274));
  xor2s1 ___0_9_438873(.DIN1 (____0____30015), .DIN2 (______9__31253),
       .Q (_____0___31273));
  nor2s1 ___0___438874(.DIN1 (____00___34539), .DIN2 (_________31234),
       .Q (______9__31308));
  xor2s1 ___0___438875(.DIN1 (______9__31210), .DIN2 (____0_0__30916),
       .Q (_________33440));
  hi1s1 ___0_9_438876(.DIN (_____0___31272), .Q (_________31318));
  nor2s1 ___09__438877(.DIN1 (_____0___31270), .DIN2 (_________31232),
       .Q (_____0___31271));
  xor2s1 ___09_438878(.DIN1 (_________31204), .DIN2 (____0_0__31851),
       .Q (_____00__31269));
  xor2s1 ___09__438879(.DIN1 (_________31124), .DIN2 (_________34644),
       .Q (_____99__31268));
  nor2s1 ___09__438880(.DIN1 (_________35002), .DIN2 (_________31227),
       .Q (_____9___31267));
  nor2s1 ___0999(.DIN1 (_________31223), .DIN2 (_________31221), .Q
       (_____9___31265));
  nor2s1 ____0__438881(.DIN1 (_________________0___18633), .DIN2
       (_________31222), .Q (_____9___31264));
  nnd2s1 ____0__438882(.DIN1 (______9__31219), .DIN2 (_____0___35109),
       .Q (_____9___31263));
  xor2s1 ____0__438883(.DIN1 (______9__31200), .DIN2 (______9__32232),
       .Q (_________31297));
  and2s1 ___0___438884(.DIN1 (_________31261), .DIN2
       (________________18755), .Q (______9__31262));
  nor2s1 ___0___438885(.DIN1 (_____0___31098), .DIN2 (_________31259),
       .Q (_________31260));
  xor2s1 ___09__438886(.DIN1 (___0____19818), .DIN2 (_____0___31191),
       .Q (_________31258));
  and2s1 ___09__438887(.DIN1 (_________31231), .DIN2 (_________31256),
       .Q (_________31257));
  nor2s1 ___0___438888(.DIN1 (______0__31254), .DIN2 (_________31233),
       .Q (_________31255));
  nor2s1 ___09_438889(.DIN1 (_______19027), .DIN2 (_________31213), .Q
       (_________31289));
  and2s1 ___09__438890(.DIN1 (______9__31253), .DIN2 (____9____29985),
       .Q (_________31287));
  xor2s1 ___0909(.DIN1 (_____0___31186), .DIN2 (_________30612), .Q
       (_____0___31272));
  nnd2s1 ___0_9_438891(.DIN1 (_________31252), .DIN2
       (________________18755), .Q (______0__31278));
  or2s1 ___0__438892(.DIN1 (________________18755), .DIN2
       (_________31252), .Q (_________31288));
  nnd2s1 ___09__438893(.DIN1 (_________31205), .DIN2 (________22067),
       .Q (_________31251));
  and2s1 ___09__438894(.DIN1 (_________34644), .DIN2 (_________31119),
       .Q (_________31250));
  nnd2s1 ___0990(.DIN1 (_________31206), .DIN2 (_________31150), .Q
       (_________31249));
  xor2s1 ____00_438895(.DIN1 (____9____30847), .DIN2 (_________31214),
       .Q (_________31248));
  nnd2s1 ____0__438896(.DIN1 (_________31245), .DIN2 (_________31281),
       .Q (______0__31247));
  nor2s1 ____0__438897(.DIN1 (_________31281), .DIN2 (_________31245),
       .Q (______9__31246));
  nnd2s1 ____0__438898(.DIN1 (_________31245), .DIN2
       (_______________18884), .Q (_________31244));
  or2s1 ___09_438899(.DIN1 (_________31464), .DIN2 (_____99__31182), .Q
       (_________31243));
  nor2s1 ___09__438900(.DIN1 (______0__31193), .DIN2 (_________31241),
       .Q (_________31242));
  nnd2s1 ___09__438901(.DIN1 (_________31239), .DIN2 (______0__31238),
       .Q (_________31240));
  nor2s1 ____0__438902(.DIN1 (_________30131), .DIN2 (_____00__31183),
       .Q (______9__31237));
  or2s1 ___09__438903(.DIN1 (_____________9___18703), .DIN2
       (_____0___31191), .Q (_________31236));
  nnd2s1 ___09__438904(.DIN1 (_____0___31191), .DIN2
       (_____________9___18703), .Q (_________31235));
  hi1s1 ___0___438905(.DIN (_________31233), .Q (_________31234));
  hi1s1 ___09_438906(.DIN (_________31231), .Q (_________31232));
  xnr2s1 ____0__438907(.DIN1 (_____0___34429), .DIN2 (_________31230),
       .Q (______0__31229));
  nnd2s1 ___09_438908(.DIN1 (_________31196), .DIN2 (_____0___31185),
       .Q (_____0___31275));
  xor2s1 ____0__438909(.DIN1 (________20581), .DIN2 (______9__31228),
       .Q (_________31367));
  nnd2s1 ____0__438910(.DIN1 (_________31226), .DIN2 (_________30710),
       .Q (_________31227));
  nor2s1 ____0__438911(.DIN1 (____99__22717), .DIN2 (_________31226),
       .Q (_________31225));
  nor2s1 ____0__438912(.DIN1 (_____9___31180), .DIN2 (_________31223),
       .Q (_________31224));
  nor2s1 ____0__438913(.DIN1 (____0__19007), .DIN2 (_____9___31176), .Q
       (_________31222));
  and2s1 ____0_438914(.DIN1 (_____9___31181), .DIN2 (_________31220),
       .Q (_________31221));
  hi1s1 ____0__438915(.DIN (_________31245), .Q (______9__31219));
  nor2s1 ____09_438916(.DIN1 (_________35106), .DIN2 (_____9___31179),
       .Q (_________31218));
  xor2s1 _____0_438917(.DIN1 (_____0___34428), .DIN2 (_________31199),
       .Q (_________31217));
  hi1s1 _______438918(.DIN (_________31215), .Q (_________31216));
  nor2s1 ____0_438919(.DIN1 (____9_9__30845), .DIN2 (_________31214),
       .Q (_____9___31266));
  nor2s1 ___09__438920(.DIN1 (_____________________18662), .DIN2
       (_________31170), .Q (_________31213));
  xor2s1 ___09__438921(.DIN1 (______0__31211), .DIN2 (_________34466),
       .Q (_________31212));
  xor2s1 ___09__438922(.DIN1 (____0____30928), .DIN2 (_________31155),
       .Q (______9__31210));
  nor2s1 ___09__438923(.DIN1 (_________31172), .DIN2 (______0__31211),
       .Q (_________31209));
  nnd2s1 ___09__438924(.DIN1 (_________31207), .DIN2 (_________31208),
       .Q (_________31231));
  nnd2s1 ___09__438925(.DIN1 (_________31171), .DIN2 (_________31168),
       .Q (______9__31253));
  xor2s1 ___0___438926(.DIN1 (______9__31158), .DIN2 (____0____32762),
       .Q (_________31233));
  nor2s1 ___09_438927(.DIN1 (_________31208), .DIN2 (_________31207),
       .Q (_____0___31270));
  xor2s1 ___0__438928(.DIN1 (_________31156), .DIN2 (____0_0__31851),
       .Q (_________31259));
  dffacs1 __________________438929(.CLRB (reset), .CLK (clk), .DIN
       (_____9___31175), .Q (________________18755));
  or2s1 ____0__438930(.DIN1 (____9____34519), .DIN2 (_________31152),
       .Q (_________31206));
  nor2s1 ___09__438931(.DIN1 (____9___20598), .DIN2 (_____90__31174),
       .Q (_________31205));
  nor2s1 ___09__438932(.DIN1 (_________31203), .DIN2 (______0__31201),
       .Q (_________31204));
  and2s1 ____000(.DIN1 (______0__31201), .DIN2 (_________31203), .Q
       (_________31202));
  nnd2s1 _______438933(.DIN1 (_________31199), .DIN2
       (_________________18682), .Q (______9__31200));
  nor2s1 _______438934(.DIN1 (_____9__23665), .DIN2 (_________31199),
       .Q (_________31197));
  nor2s1 _______438935(.DIN1 (_________________18682), .DIN2
       (_________31199), .Q (_________31215));
  xor2s1 ______438936(.DIN1 (_____9___31178), .DIN2 (___9____19720), .Q
       (_________31245));
  xor2s1 ___09__438937(.DIN1 (_________31147), .DIN2 (______0__32594),
       .Q (_________31196));
  hi1s1 ___09__438938(.DIN (_________31194), .Q (_________31195));
  nor2s1 ___09__438939(.DIN1 (_____09__31192), .DIN2 (_________34466),
       .Q (______0__31193));
  nor2s1 ___09__438940(.DIN1 (_________34466), .DIN2 (______0__29512),
       .Q (_____0___31190));
  or2s1 ___09__438941(.DIN1 (_____0___31188), .DIN2 (_____0___31187),
       .Q (_____0___31189));
  and2s1 ___09__438942(.DIN1 (_____0___31185), .DIN2 (_________31146),
       .Q (_____0___31186));
  hi1s1 ___099_438943(.DIN (____090__33759), .Q (_____0___31191));
  nor2s1 ___09__438944(.DIN1 (____0_0__30942), .DIN2 (_________34466),
       .Q (_________31382));
  xor2s1 ___09__438945(.DIN1 (_________31145), .DIN2 (_____0___31184),
       .Q (_________31239));
  dffacs1 ___________________438946(.CLRB (reset), .CLK (clk), .DIN
       (______0__31159), .QN (_________________18712));
  nnd2s1 ____09_438947(.DIN1 (_________34205), .DIN2 (____9___20416),
       .Q (_____00__31183));
  xor2s1 ____00_438948(.DIN1 (_________29673), .DIN2 (______0__31167),
       .Q (_____99__31182));
  hi1s1 ____0__438949(.DIN (_____9___31180), .Q (_____9___31181));
  nnd2s1 _______438950(.DIN1 (_____9___31178), .DIN2 (________25579),
       .Q (_____9___31179));
  nor2s1 _______438951(.DIN1 (_____0___34428), .DIN2 (_________31160),
       .Q (_____9___31177));
  nor2s1 _______438952(.DIN1 (______18947), .DIN2 (_____9___31178), .Q
       (_____9___31176));
  nor2s1 ____09_438953(.DIN1 (_________30592), .DIN2 (_________34205),
       .Q (_________31223));
  nor2s1 _____0_438954(.DIN1 (______9__30773), .DIN2 (______0__31149),
       .Q (_________31214));
  hi1s1 ____0__438955(.DIN (______9__31228), .Q (_________31226));
  nnd2s1 ___0___438956(.DIN1 (_________31141), .DIN2 (____00___29085),
       .Q (_____9___31175));
  nor2s1 ____0_438957(.DIN1 (____9___20597), .DIN2 (_________31133), .Q
       (_____90__31174));
  hi1s1 ___09__438958(.DIN (_________34466), .Q (_________31172));
  nnd2s1 ___09_438959(.DIN1 (_________31169), .DIN2
       (_________________18695), .Q (_________31171));
  and2s1 ____00_438960(.DIN1 (_________31169), .DIN2 (_________31168),
       .Q (_________31170));
  nor2s1 ___09_438961(.DIN1 (____0____30917), .DIN2 (_________31143),
       .Q (_________31207));
  xnr2s1 ___09__438962(.DIN1 (_________31486), .DIN2 (_________34646),
       .Q (_________31194));
  xor2s1 ____0__438963(.DIN1 (_________31127), .DIN2 (____0____31831),
       .Q (____090__33759));
  nor2s1 ____0__438964(.DIN1 (_________31165), .DIN2 (_________31138),
       .Q (______9__31166));
  xor2s1 ______438965(.DIN1 (_________31113), .DIN2 (____0____31863),
       .Q (_________31162));
  nor2s1 ____09_438966(.DIN1 (___0____19837), .DIN2 (_________31161),
       .Q (_____9___31180));
  xor2s1 ____0__438967(.DIN1 (_________31114), .DIN2 (_________33268),
       .Q (______0__31201));
  xor2s1 _____0_438968(.DIN1 (_________30796), .DIN2 (______9__31148),
       .Q (______9__31228));
  hi1s1 _______438969(.DIN (_________31160), .Q (_________31199));
  xor2s1 _____0_438970(.DIN1 (_________31117), .DIN2 (_________33835),
       .Q (_________31230));
  nnd2s1 ___09__438971(.DIN1 (______9__31129), .DIN2 (_________35102),
       .Q (______0__31159));
  nor2s1 ___09__438972(.DIN1 (_________31038), .DIN2 (_________31144),
       .Q (______9__31158));
  nnd2s1 ___09__438973(.DIN1 (_________31128), .DIN2 (_________32440),
       .Q (_________31157));
  nnd2s1 ___0___438974(.DIN1 (_________31123), .DIN2 (______0__31101),
       .Q (_________31156));
  xor2s1 ____00_438975(.DIN1 (_________31142), .DIN2 (_________31154),
       .Q (_________31155));
  xor2s1 ____0__438976(.DIN1 (_________31108), .DIN2 (_________31153),
       .Q (_____0___31185));
  dffacs1 _________________0_438977(.CLRB (reset), .CLK (clk), .DIN
       (_________31122), .Q (_________34466));
  and2s1 ____0__438978(.DIN1 (_________31151), .DIN2
       (_________________18681), .Q (_________31152));
  or2s1 ____0_9(.DIN1 (_________________18681), .DIN2 (_________31151),
       .Q (_________31150));
  nor2s1 _______438979(.DIN1 (_________30775), .DIN2 (______9__31148),
       .Q (______0__31149));
  nor2s1 ____0__438980(.DIN1 (_________34486), .DIN2 (____9____33599),
       .Q (_____0___31187));
  xor2s1 _______438981(.DIN1 (_________31059), .DIN2 (_________31132),
       .Q (_________31160));
  and2s1 ____0__438982(.DIN1 (____9____33599), .DIN2 (_________34486),
       .Q (_____0___31188));
  xor2s1 ______438983(.DIN1 (_________31103), .DIN2 (______9__34123),
       .Q (_____9___31178));
  hi1s1 ______438984(.DIN (_________31161), .Q (_________34205));
  and2s1 ____0_438985(.DIN1 (_________31146), .DIN2
       (___________0___18883), .Q (_________31147));
  nor2s1 ____0__438986(.DIN1 (_________________18783), .DIN2
       (______9__31139), .Q (_________31145));
  and2s1 ____0_438987(.DIN1 (_________31142), .DIN2 (____0____30982),
       .Q (_________31143));
  nnd2s1 ___090_438988(.DIN1 (______0__31111), .DIN2 (_________32604),
       .Q (_________31141));
  xor2s1 ____0__438989(.DIN1 (_____9___31086), .DIN2 (_________31067),
       .Q (_________33474));
  nnd2s1 ____0__438990(.DIN1 (______0__31140), .DIN2 (_________33330),
       .Q (_________31168));
  or2s1 ____0__438991(.DIN1 (_________33330), .DIN2 (______0__31140),
       .Q (_________31169));
  nnd2s1 ____0__438992(.DIN1 (______9__31139), .DIN2
       (_________________18783), .Q (______0__31238));
  hi1s1 ____0_438993(.DIN (_________31137), .Q (_________31138));
  xor2s1 _______438994(.DIN1 (_________31135), .DIN2 (_________31134),
       .Q (_________31136));
  xor2s1 ____09_438995(.DIN1 (_____90__31084), .DIN2 (______0__35008),
       .Q (_________31133));
  nnd2s1 ____0__438996(.DIN1 (____9____32668), .DIN2 (_________31131),
       .Q (_________31198));
  nnd2s1 _____9_438997(.DIN1 (_________31132), .DIN2 (______9__31043),
       .Q (_________31163));
  nor2s1 ____0__438998(.DIN1 (______0__31054), .DIN2 (_________31104),
       .Q (______0__31167));
  nor2s1 ____0_438999(.DIN1 (_________31131), .DIN2 (____9____32668),
       .Q (_________31173));
  xor2s1 _____0_439000(.DIN1 (_____9___31085), .DIN2 (_________33144),
       .Q (_________31363));
  xor2s1 _______439001(.DIN1 (______9__31083), .DIN2 (______0__31130),
       .Q (_________31161));
  dffacs1 ___________________439002(.CLRB (reset), .CLK (clk), .DIN
       (_________31109), .QN (_________34492));
  nnd2s1 ____0_439003(.DIN1 (_________31102), .DIN2 (_________31047),
       .Q (______9__31129));
  xor2s1 ___09__439004(.DIN1 (_________31075), .DIN2 (_________30491),
       .Q (_________31128));
  nnd2s1 ____0__439005(.DIN1 (_____9___31090), .DIN2 (_________31126),
       .Q (_________31127));
  nor2s1 ____0__439006(.DIN1 (___9____21556), .DIN2 (____9_0__33587),
       .Q (_________31125));
  xor2s1 ____0__439007(.DIN1 (_____99__31092), .DIN2 (______9__31120),
       .Q (_________31124));
  or2s1 ___09__439008(.DIN1 (_____00__29176), .DIN2 (_____0___31094),
       .Q (_________31123));
  nnd2s1 ____0__439009(.DIN1 (_____0___31095), .DIN2 (_____9___31443),
       .Q (_________31122));
  nor2s1 ____0__439010(.DIN1 (______9__31120), .DIN2 (_________31118),
       .Q (______0__31121));
  nnd2s1 ____0__439011(.DIN1 (_________31118), .DIN2 (______9__31120),
       .Q (_________31119));
  nor2s1 ___099_439012(.DIN1 (_________31050), .DIN2 (_____0___31097),
       .Q (_____0___32387));
  xor2s1 ___09__439013(.DIN1 (_________31076), .DIN2 (_________32606),
       .Q (_________31144));
  xor2s1 _______439014(.DIN1 (_________31057), .DIN2
       (_________________0___18633), .Q (_________31117));
  nor2s1 _____439015(.DIN1 (_____0___35109), .DIN2 (_________31135), .Q
       (_________31116));
  and2s1 _____9_439016(.DIN1 (_________31135), .DIN2 (_________31290),
       .Q (_________31115));
  xor2s1 _______439017(.DIN1 (_________31061), .DIN2 (_________31041),
       .Q (_________31114));
  and2s1 _____9_439018(.DIN1 (_________31135), .DIN2
       (_______________18879), .Q (_________31113));
  or2s1 _____9_439019(.DIN1 (_______________18879), .DIN2
       (_________31135), .Q (_________31112));
  nnd2s1 ____0__439020(.DIN1 (____9_0__33587), .DIN2
       (_________________18702), .Q (_________31137));
  nor2s1 _______439021(.DIN1 (_________31081), .DIN2 (_____9___31087),
       .Q (______9__31148));
  nor2s1 ____0__439022(.DIN1 (_________________18702), .DIN2
       (____9_0__33587), .Q (_________31165));
  dffacs1 ___________________439023(.CLRB (reset), .CLK (clk), .DIN
       (_____0___31096), .QN (_________________18711));
  xor2s1 _______439024(.DIN1 (_________31062), .DIN2 (_________31956),
       .Q (_________31151));
  hi1s1 ____0__439025(.DIN (______9__31139), .Q (____9____33599));
  xor2s1 ___09__439026(.DIN1 (____9____30841), .DIN2 (______0__34648),
       .Q (______0__31111));
  nor2s1 ____0__439027(.DIN1 (_________________18782), .DIN2
       (_________31080), .Q (______9__31110));
  or2s1 ____0__439028(.DIN1 (____9____30867), .DIN2 (_________31071),
       .Q (_________31109));
  nor2s1 ____099(.DIN1 (_________31106), .DIN2 (_________31107), .Q
       (_________31108));
  nnd2s1 _____00(.DIN1 (_________31107), .DIN2 (_________31106), .Q
       (_________31146));
  nnd2s1 ____0__439029(.DIN1 (______9__31073), .DIN2 (_________29837),
       .Q (______0__31140));
  nor2s1 _______439030(.DIN1 (_________31464), .DIN2 (______9__31063),
       .Q (_________31105));
  and2s1 ______439031(.DIN1 (______0__31064), .DIN2 (_____0___32851),
       .Q (_________31104));
  nor2s1 _______439032(.DIN1 (________25124), .DIN2 (_________31066),
       .Q (_________31103));
  nnd2s1 _____0_439033(.DIN1 (_________31069), .DIN2 (____009__34540),
       .Q (_________31142));
  nnd2s1 _______439034(.DIN1 (_________31056), .DIN2 (______0__31007),
       .Q (_________31132));
  xor2s1 _____439035(.DIN1 (___9_9__25210), .DIN2 (_____9___31089), .Q
       (______9__31139));
  xor2s1 _______439036(.DIN1 (_________31036), .DIN2 (_________31039),
       .Q (____9____32668));
  xor2s1 ____090(.DIN1 (______0__29813), .DIN2 (_________31072), .Q
       (_________31102));
  nnd2s1 ___09__439037(.DIN1 (______0__34648), .DIN2 (_____00__31093),
       .Q (______0__31101));
  or2s1 ___09__439038(.DIN1 (_____0___31099), .DIN2 (_____0___31098),
       .Q (_____0___31100));
  nor2s1 ____0__439039(.DIN1 (______0__31074), .DIN2 (_________31052),
       .Q (_____0___31097));
  nnd2s1 ____0__439040(.DIN1 (_________31048), .DIN2 (________23856),
       .Q (_____0___31096));
  nor2s1 ____0__439041(.DIN1 (________22836), .DIN2 (_________31049),
       .Q (_____0___31095));
  nor2s1 ___09__439042(.DIN1 (_____00__31093), .DIN2 (______0__34648),
       .Q (_____0___31094));
  hi1s1 ____0__439043(.DIN (_____99__31092), .Q (_________31118));
  xor2s1 ____09_439044(.DIN1 (_________31077), .DIN2 (_________31078),
       .Q (_____9___31091));
  nnd2s1 ______439045(.DIN1 (_____9___31089), .DIN2 (_____9___31088),
       .Q (_____9___31090));
  nor2s1 _____0_439046(.DIN1 (_________30740), .DIN2 (_________31082),
       .Q (_____9___31087));
  nnd2s1 _______439047(.DIN1 (_________31068), .DIN2 (____009__34540),
       .Q (_____9___31086));
  nor2s1 _______439048(.DIN1 (____0____30953), .DIN2 (_________31042),
       .Q (_____9___31085));
  xor2s1 _______439049(.DIN1 (______9__31034), .DIN2 (_________31031),
       .Q (_____90__31084));
  or2s1 _____9_439050(.DIN1 (_________31082), .DIN2 (_________31081),
       .Q (______9__31083));
  dffacs1 ___________________439051(.CLRB (reset), .CLK (clk), .DIN
       (_________31046), .QN (_________________18694));
  xor2s1 _______439052(.DIN1 (___0____25295), .DIN2 (_________31065),
       .Q (_________31135));
  hi1s1 _______439053(.DIN (_________31080), .Q (____9_0__33587));
  or2s1 _______439054(.DIN1 (_________31078), .DIN2 (_________31077),
       .Q (_________31079));
  xor2s1 ____0__439055(.DIN1 (________________18737), .DIN2
       (____0_9__29109), .Q (_________31076));
  xor2s1 ____0__439056(.DIN1 (______0__31074), .DIN2 (_________31051),
       .Q (_________31075));
  or2s1 ______439057(.DIN1 (_________29836), .DIN2 (_________31072), .Q
       (______9__31073));
  nnd2s1 _______439058(.DIN1 (_________30594), .DIN2 (______0__31035),
       .Q (_________31071));
  and2s1 _______439059(.DIN1 (_________31077), .DIN2 (_________31078),
       .Q (_________31070));
  nnd2s1 _______439060(.DIN1 (_________31068), .DIN2 (_________31067),
       .Q (_________31069));
  nor2s1 _______439061(.DIN1 (____09___30989), .DIN2 (_________31037),
       .Q (_________31107));
  xor2s1 _____0_439062(.DIN1 (_________31021), .DIN2 (______0__29502),
       .Q (_____99__31092));
  nor2s1 _______439063(.DIN1 (___9____25239), .DIN2 (_________31065),
       .Q (_________31066));
  nnd2s1 _______439064(.DIN1 (_________31026), .DIN2 (____9____30876),
       .Q (______0__31064));
  and2s1 _______439065(.DIN1 (_________31029), .DIN2 (______9__31053),
       .Q (______9__31063));
  nor2s1 _____9_439066(.DIN1 (_________31033), .DIN2 (_________31032),
       .Q (_________31062));
  xor2s1 _____0_439067(.DIN1 (_________31017), .DIN2 (_________31060),
       .Q (_________31061));
  xor2s1 _______439068(.DIN1 (_________31106), .DIN2 (_________31058),
       .Q (_________31059));
  xor2s1 _______439069(.DIN1 (______9__31015), .DIN2 (_________31027),
       .Q (_________31057));
  nor2s1 _______439070(.DIN1 (_________31008), .DIN2 (_________31028),
       .Q (_________31056));
  xor2s1 ______439071(.DIN1 (______0__31016), .DIN2
       (_________________0___18607), .Q (_________31080));
  or2s1 ____0_439072(.DIN1 (________________18737), .DIN2
       (____9____29058), .Q (_________31055));
  nor2s1 _______439073(.DIN1 (_____0___32851), .DIN2 (______9__31053),
       .Q (______0__31054));
  and2s1 ____0_439074(.DIN1 (_________31051), .DIN2
       (________________18724), .Q (_________31052));
  nor2s1 ____0_439075(.DIN1 (________________18724), .DIN2
       (_________31051), .Q (_________31050));
  nor2s1 _______439076(.DIN1 (_________31464), .DIN2 (_________31019),
       .Q (_________31049));
  nnd2s1 _______439077(.DIN1 (_________31018), .DIN2 (_________31047),
       .Q (_________31048));
  xor2s1 ____00_439078(.DIN1 (____099__30996), .DIN2 (_________33278),
       .Q (_____0___31098));
  nnd2s1 _______439079(.DIN1 (_________31009), .DIN2 (________19356),
       .Q (_________31046));
  nnd2s1 _______439080(.DIN1 (______0__31044), .DIN2 (____0____30969),
       .Q (_________31045));
  nnd2s1 _______439081(.DIN1 (_________31106), .DIN2 (_________31058),
       .Q (______9__31043));
  nor2s1 ______439082(.DIN1 (_________31041), .DIN2 (_________31014),
       .Q (_________31042));
  nor2s1 _______439083(.DIN1 (_________31058), .DIN2 (_________31106),
       .Q (_________31040));
  xor2s1 ______439084(.DIN1 (____0____30980), .DIN2 (_________31926),
       .Q (_________31039));
  nor2s1 ______439085(.DIN1 (_________30151), .DIN2 (_________31012),
       .Q (_________31082));
  xor2s1 _______439086(.DIN1 (_____0___31002), .DIN2 (_____0___30999),
       .Q (_____9___31089));
  and2s1 ______439087(.DIN1 (_________31036), .DIN2 (____0_0__30979),
       .Q (_________31037));
  nnd2s1 _______439088(.DIN1 (_____________________18662), .DIN2
       (_____0___31004), .Q (______0__31035));
  nor2s1 _______439089(.DIN1 (______0__29671), .DIN2 (_____0___30998),
       .Q (_________31072));
  nnd2s1 ______439090(.DIN1 (_________31010), .DIN2 (_________30615),
       .Q (_________31068));
  nnd2s1 ______439091(.DIN1 (____09___30995), .DIN2 (_________29503),
       .Q (_________31078));
  nor2s1 ______439092(.DIN1 (_________31030), .DIN2 (_________31033),
       .Q (______9__31034));
  nor2s1 _______439093(.DIN1 (_________31031), .DIN2 (_________31030),
       .Q (_________31032));
  nnd2s1 _______439094(.DIN1 (______0__31025), .DIN2 (____9____30895),
       .Q (_________31029));
  and2s1 _______439095(.DIN1 (____0_9__30987), .DIN2 (_________31027),
       .Q (_________31028));
  nnd2s1 _______439096(.DIN1 (______0__31025), .DIN2 (____9____30875),
       .Q (_________31026));
  nor2s1 _______439097(.DIN1 (_________30190), .DIN2 (_________31011),
       .Q (_________31081));
  nor2s1 _____9_439098(.DIN1 (________25506), .DIN2 (____0____30984),
       .Q (_________31065));
  nnd2s1 ___09__439099(.DIN1 (____0_9__30971), .DIN2 (_________32604),
       .Q (______9__31024));
  nnd2s1 ____0__439100(.DIN1 (____0____30975), .DIN2 (_________31022),
       .Q (_________31023));
  xor2s1 _______439101(.DIN1 (_________________18710), .DIN2
       (_________31020), .Q (_________31021));
  xor2s1 ______439102(.DIN1 (____0____30956), .DIN2 (____99___35108),
       .Q (_________31019));
  xor2s1 _______439103(.DIN1 (_____9___29704), .DIN2 (_____00__30997),
       .Q (_________31018));
  nnd2s1 _____9_439104(.DIN1 (____09___30993), .DIN2 (____9____30896),
       .Q (______9__31053));
  dffacs1 __________________439105(.CLRB (reset), .CLK (clk), .DIN
       (____0____30973), .QN (________________18737));
  xor2s1 _____0_439106(.DIN1 (____0____30958), .DIN2 (_________32442),
       .Q (_________31038));
  nor2s1 ______439107(.DIN1 (____0____30943), .DIN2 (____0_0__30972),
       .Q (_________31051));
  nnd2s1 _______439108(.DIN1 (_________31013), .DIN2 (____0____30963),
       .Q (_________31017));
  xor2s1 _____0_439109(.DIN1 (____0____30947), .DIN2 (________25102),
       .Q (______0__31016));
  xor2s1 _____0_439110(.DIN1 (____090__30988), .DIN2 (______0__33107),
       .Q (______9__31015));
  xor2s1 _______439111(.DIN1 (_________31013), .DIN2 (_________28828),
       .Q (_________31014));
  hi1s1 _______439112(.DIN (_________31011), .Q (_________31012));
  nnd2s1 _______439113(.DIN1 (____0____30966), .DIN2 (_________31047),
       .Q (_________31009));
  nor2s1 _______439114(.DIN1 (_____0___31005), .DIN2 (_____09__31006),
       .Q (_________31008));
  nnd2s1 _______439115(.DIN1 (_____09__31006), .DIN2 (_____0___31005),
       .Q (______0__31007));
  xor2s1 _____439116(.DIN1 (____0_9__30951), .DIN2 (_________33278), .Q
       (______0__31044));
  xor2s1 _______439117(.DIN1 (________25895), .DIN2 (____0____30983),
       .Q (_________31106));
  or2s1 _______439118(.DIN1 (_____0___31003), .DIN2
       (_________________18710), .Q (_____0___31004));
  nnd2s1 _______439119(.DIN1 (____0_0__30952), .DIN2 (____0____30946),
       .Q (_____0___31002));
  nnd2s1 _______439120(.DIN1 (____0____30957), .DIN2 (_________34966),
       .Q (_____0___31001));
  xor2s1 _______439121(.DIN1 (____0____30936), .DIN2 (_____0___30999),
       .Q (_____0___31000));
  nor2s1 _______439122(.DIN1 (______9__29670), .DIN2 (_____00__30997),
       .Q (_____0___30998));
  nnd2s1 ____09_439123(.DIN1 (____09___30991), .DIN2 (____09___30992),
       .Q (____099__30996));
  or2s1 _____0_439124(.DIN1 (_________________18710), .DIN2
       (_________29494), .Q (____09___30995));
  xnr2s1 _____0_439125(.DIN1 (_________35066), .DIN2 (_________32230),
       .Q (____09___30994));
  xnr2s1 _____0_439126(.DIN1 (_________34023), .DIN2 (_________34652),
       .Q (_________31010));
  hi1s1 ______439127(.DIN (____09___30993), .Q (______0__31025));
  nor2s1 ____09_439128(.DIN1 (____09___30992), .DIN2 (____09___30991),
       .Q (_____0___31099));
  xor2s1 _____0_439129(.DIN1 (____0____30926), .DIN2 (_________31431),
       .Q (____09___30990));
  nor2s1 _______439130(.DIN1
       (______________________________________0_____________18887),
       .DIN2 (____090__30988), .Q (____09___30989));
  nnd2s1 ______439131(.DIN1 (____090__30988), .DIN2
       (___________0___18877), .Q (____0_9__30987));
  xnr2s1 _______439132(.DIN1 (_________35110), .DIN2 (____0____30985),
       .Q (____0____30986));
  nor2s1 _______439133(.DIN1 (________25507), .DIN2 (____0____30983),
       .Q (____0____30984));
  xor2s1 _______439134(.DIN1 (____0____30929), .DIN2 (____0____30981),
       .Q (____0____30982));
  xor2s1 _____439135(.DIN1 (____0_0__30962), .DIN2 (________19986), .Q
       (____0____30980));
  nnd2s1 _______439136(.DIN1 (____090__30988), .DIN2
       (______________________________________0_____________18887), .Q
       (____0_0__30979));
  xor2s1 _______439137(.DIN1 (_________34654), .DIN2 (_________33174),
       .Q (_________31011));
  nor2s1 ______439138(.DIN1 (_________________18680), .DIN2
       (_________34650), .Q (_________31033));
  and2s1 _______439139(.DIN1 (_________34650), .DIN2
       (_________________18680), .Q (_________31030));
  xnr2s1 _______439140(.DIN1 (_________35086), .DIN2 (_________31978),
       .Q (____0____30978));
  hi1s1 _______439141(.DIN (____0____30974), .Q (____0____30975));
  nor2s1 _______439142(.DIN1 (_________33370), .DIN2 (____0____30937),
       .Q (____0____30973));
  nor2s1 _______439143(.DIN1 (____0____30940), .DIN2 (_____9___32286),
       .Q (____0_0__30972));
  xor2s1 ____0_439144(.DIN1 (____0_0__34550), .DIN2 (____0____30933),
       .Q (____0_9__30971));
  hi1s1 _______439145(.DIN (____0____30969), .Q (____0____30970));
  xnr2s1 _______439146(.DIN1 (_________34439), .DIN2 (_________32208),
       .Q (____0____30968));
  xor2s1 _______439147(.DIN1 (____9___22075), .DIN2 (_________32208),
       .Q (____0____30967));
  xor2s1 _______439148(.DIN1 (____0____30919), .DIN2 (____0____30965),
       .Q (____0____30966));
  nor2s1 _____439149(.DIN1 (_____9___30454), .DIN2 (____0____30934), .Q
       (____0____30964));
  nnd2s1 _____9_439150(.DIN1 (____0____30985), .DIN2 (______0__30418),
       .Q (____0____30963));
  nnd2s1 _______439151(.DIN1 (____0_0__30962), .DIN2 (_________33835),
       .Q (_____09__31006));
  xor2s1 _______439152(.DIN1 (____0_9__30923), .DIN2 (____0_9__30961),
       .Q (____09___30993));
  and2s1 _______439153(.DIN1 (_________32208), .DIN2 (_________34439),
       .Q (____0____30960));
  nor2s1 _______439154(.DIN1 (_________34439), .DIN2 (_________32208),
       .Q (____0____30959));
  nnd2s1 ______439155(.DIN1 (____0____30922), .DIN2 (____9_0__30889),
       .Q (____0____30958));
  xor2s1 ______439156(.DIN1 (______9__29338), .DIN2 (____0_9__30941),
       .Q (____0____30957));
  xor2s1 ______439157(.DIN1 (____99___30898), .DIN2 (_________34660),
       .Q (____0____30956));
  nnd2s1 _______439158(.DIN1 (____0____30954), .DIN2 (____0____30955),
       .Q (_________31022));
  nor2s1 _______439159(.DIN1 (____0____30955), .DIN2 (____0____30954),
       .Q (____0____30974));
  xor2s1 _______439160(.DIN1 (_________34656), .DIN2 (_________31479),
       .Q (_____00__30997));
  xor2s1 _______439161(.DIN1 (____000__30906), .DIN2 (_____9___33026),
       .Q (____09___30991));
  xor2s1 _______439162(.DIN1 (____99___30901), .DIN2 (_________30804),
       .Q (_____90__33391));
  dffacs1 ___________________439163(.CLRB (reset), .CLK (clk), .DIN
       (____0_0__30924), .QN (_________________18710));
  nor2s1 _______439164(.DIN1 (________21138), .DIN2 (____0____30945),
       .Q (____0____30953));
  nor2s1 _______439165(.DIN1 (___9____25244), .DIN2 (____0____30921),
       .Q (____0_0__30952));
  nor2s1 _______439166(.DIN1
       (_______________0_____________________18831), .DIN2
       (_________32208), .Q (____0_9__30951));
  xor2s1 _______439167(.DIN1 (____0____30949), .DIN2 (outData[31]), .Q
       (____0____30950));
  nor2s1 _______439168(.DIN1 (____9___22074), .DIN2 (_________32208),
       .Q (____0____30948));
  nnd2s1 _______439169(.DIN1 (____0____30946), .DIN2 (____0____30920),
       .Q (____0____30947));
  nnd2s1 ______439170(.DIN1 (____0____30945), .DIN2 (____0___20046), .Q
       (_________31013));
  nor2s1 _______439171(.DIN1 (________25921), .DIN2 (____009__30915),
       .Q (____0____30983));
  nnd2s1 _______439172(.DIN1 (_________32208), .DIN2
       (_______________0_____________________18831), .Q
       (____0____30969));
  xor2s1 _______439173(.DIN1 (____99___30899), .DIN2 (______0__30345),
       .Q (_________31208));
  hi1s1 ______439174(.DIN (____0_0__30962), .Q (____090__30988));
  nor2s1 _______439175(.DIN1 (_________________18701), .DIN2
       (____00___30911), .Q (____0____30944));
  nor2s1 _______439176(.DIN1 (____0_0__30942), .DIN2 (____0_9__30941),
       .Q (____0____30943));
  and2s1 _______439177(.DIN1 (____0_9__30941), .DIN2 (____0_0__30942),
       .Q (____0____30940));
  nnd2s1 _____439178(.DIN1 (____0____30935), .DIN2 (____0____30938), .Q
       (____0____30939));
  xor2s1 _____0_439179(.DIN1 (______9__34470), .DIN2 (____9____30887),
       .Q (____0____30937));
  nor2s1 _____0_439180(.DIN1 (____0____30938), .DIN2 (____0____30935),
       .Q (____0____30936));
  xor2s1 _______439181(.DIN1 (____9____30883), .DIN2 (_________30472),
       .Q (____0____30934));
  nor2s1 _______439182(.DIN1 (____00___30908), .DIN2 (____0____30933),
       .Q (____0____30976));
  xor2s1 _______439183(.DIN1 (____9____30885), .DIN2 (____0_0__30932),
       .Q (_________31036));
  and2s1 _______439184(.DIN1 (____0____30949), .DIN2 (____0____30930),
       .Q (____0_9__30931));
  nor2s1 _____0_439185(.DIN1 (____9____30851), .DIN2 (____0____30928),
       .Q (____0____30929));
  nor2s1 _______439186(.DIN1 (____0____30930), .DIN2 (____0____30949),
       .Q (____0____30927));
  nor2s1 _______439187(.DIN1 (____0____30925), .DIN2 (____00___30912),
       .Q (____0____30926));
  xor2s1 _______439188(.DIN1 (________26064), .DIN2 (____00___30914),
       .Q (____0_0__30962));
  or2s1 _______439189(.DIN1 (_________28823), .DIN2 (____999__30905),
       .Q (_________32230));
  hi1s1 _______439190(.DIN (____0____30945), .Q (____0____30985));
  nnd2s1 ______439191(.DIN1 (____9____30884), .DIN2 (___9____20639), .Q
       (____0_0__30924));
  nnd2s1 _____439192(.DIN1 (____9____30892), .DIN2 (_____9___30815), .Q
       (____0_9__30923));
  nnd2s1 _______439193(.DIN1 (_____9___30358), .DIN2 (____9____30890),
       .Q (____0____30922));
  nor2s1 _______439194(.DIN1
       (______________________________________0_____________18887),
       .DIN2 (____0____30920), .Q (____0____30921));
  nnd2s1 _____9_439195(.DIN1 (____9____30878), .DIN2 (_____0___35109),
       .Q (____0____30946));
  xor2s1 _______439196(.DIN1 (____9_9__30871), .DIN2 (_________28248),
       .Q (____0____30954));
  hi1s1 ______439197(.DIN (____0____30935), .Q (_________31978));
  xor2s1 _______439198(.DIN1 (____9____30862), .DIN2 (____0____30918),
       .Q (____0____30919));
  nor2s1 _____9_439199(.DIN1 (____0_0__30916), .DIN2 (____9____30894),
       .Q (____0____30917));
  and2s1 _____9_439200(.DIN1 (____00___30914), .DIN2 (________25922),
       .Q (____009__30915));
  hi1s1 _____0_439201(.DIN (____00___30912), .Q (____00___30913));
  nor2s1 ______439202(.DIN1 (________19923), .DIN2 (____9_9__30880), .Q
       (_________31203));
  xor2s1 _______439203(.DIN1 (____9____30833), .DIN2 (____9_9__30897),
       .Q (____0____30945));
  hi1s1 _____9_439204(.DIN (____00___30911), .Q (_________32208));
  nnd2s1 _______439205(.DIN1 (____00___30909), .DIN2 (____00___30907),
       .Q (____00___30910));
  nor2s1 _______439206(.DIN1 (____00___30907), .DIN2 (____00___30909),
       .Q (____00___30908));
  xor2s1 ______439207(.DIN1 (_________34455), .DIN2 (_____0___28902),
       .Q (____000__30906));
  nnd2s1 _______439208(.DIN1 (____9____30866), .DIN2 (____900__30820),
       .Q (____999__30905));
  or2s1 _______439209(.DIN1 (____99___30903), .DIN2 (____99___30902),
       .Q (____99___30904));
  xor2s1 _______439210(.DIN1 (____9____30861), .DIN2 (_________30805),
       .Q (____99___30901));
  hi1s1 _______439211(.DIN (____99___30900), .Q (____0____32791));
  nor2s1 _______439212(.DIN1 (____9____30886), .DIN2 (____9____30870),
       .Q (____0_9__30941));
  xor2s1 _______439213(.DIN1 (____9____30856), .DIN2 (____0____31818),
       .Q (____0____30935));
  xor2s1 _______439214(.DIN1 (_____0___34148), .DIN2 (________23324),
       .Q (____99___30899));
  xor2s1 _____0_439215(.DIN1 (_____9___30814), .DIN2 (____9____30891),
       .Q (____99___30898));
  hi1s1 _______439216(.DIN (____9____30895), .Q (____9____30896));
  nor2s1 _______439217(.DIN1 (________20551), .DIN2 (____9____30864),
       .Q (_________31256));
  hi1s1 _______439218(.DIN (____9____30894), .Q (____0____30928));
  xor2s1 _______439219(.DIN1 (____9_0__30846), .DIN2 (____0____32807),
       .Q (____00___30912));
  xor2s1 _______439220(.DIN1 (________24539), .DIN2 (____9____30877),
       .Q (____00___30911));
  xor2s1 _______439221(.DIN1 (____9____30850), .DIN2 (____9____30893),
       .Q (____0____30949));
  dffacs1 ___________________439222(.CLRB (reset), .CLK (clk), .DIN
       (____9____30868), .QN (______0__34491));
  nnd2s1 _______439223(.DIN1 (____9____30891), .DIN2 (_________30801),
       .Q (____9____30892));
  or2s1 _______439224(.DIN1 (_________34455), .DIN2 (____9_9__30888),
       .Q (____9____30890));
  nnd2s1 _______439225(.DIN1 (____9_9__30888), .DIN2 (_________34455),
       .Q (____9_0__30889));
  nor2s1 ______439226(.DIN1 (____9____30869), .DIN2 (____9____30886),
       .Q (____9____30887));
  nnd2s1 ______439227(.DIN1 (____9____30857), .DIN2 (____90___30822),
       .Q (____9____30885));
  nor2s1 _______439228(.DIN1 (________20366), .DIN2 (____9____30852),
       .Q (____9____30884));
  xor2s1 _____439229(.DIN1 (____9_9__30837), .DIN2 (______0__34668), .Q
       (____9____30883));
  xor2s1 _____0_439230(.DIN1 (____9____30865), .DIN2 (_____9___32185),
       .Q (_________32180));
  nnd2s1 _______439231(.DIN1 (____9____30859), .DIN2 (_________28249),
       .Q (____99___30900));
  nor2s1 ______439232(.DIN1 (________19897), .DIN2 (_____0___34148), .Q
       (____9_9__30880));
  xnr2s1 _______439233(.DIN1 (_________________18792), .DIN2
       (_________31031), .Q (____9____30879));
  nnd2s1 _______439234(.DIN1 (____9____30877), .DIN2 (____0____31818),
       .Q (____9____30878));
  or2s1 _______439235(.DIN1 (____0____31818), .DIN2 (____9____30877),
       .Q (____0____30920));
  nnd2s1 _______439236(.DIN1 (____9____30876), .DIN2 (____9____30875),
       .Q (____9____30895));
  xor2s1 ______439237(.DIN1 (________20552), .DIN2 (______9__34094), .Q
       (____9____30894));
  xor2s1 _______439238(.DIN1 (____9____30834), .DIN2 (_________28828),
       .Q (____00___30914));
  and2s1 ______439239(.DIN1 (_________31031), .DIN2
       (_________________18792), .Q (____9____30873));
  or2s1 _______439240(.DIN1 (_________________18792), .DIN2
       (_________31031), .Q (____9_0__30872));
  xor2s1 _______439241(.DIN1 (______0__34451), .DIN2 (____9____30858),
       .Q (____9_9__30871));
  nor2s1 ______439242(.DIN1 (______9__34470), .DIN2 (____9____30869),
       .Q (____9____30870));
  nor2s1 _______439243(.DIN1 (______0__34461), .DIN2 (____9____30842),
       .Q (____99___30903));
  xor2s1 _______439244(.DIN1 (____9____30830), .DIN2 (_____0___28617),
       .Q (____00___30909));
  or2s1 _____0_439245(.DIN1 (____9____30867), .DIN2 (____9____30835),
       .Q (____9____30868));
  or2s1 _______439246(.DIN1 (_________31956), .DIN2 (____9____30865),
       .Q (____9____30866));
  and2s1 _______439247(.DIN1 (______9__34094), .DIN2 (________20086),
       .Q (____9____30864));
  xor2s1 _____0_439248(.DIN1 (____9____30844), .DIN2
       (______________0___________________9__18827), .Q
       (____9____30862));
  nor2s1 _______439249(.DIN1 (______0__30465), .DIN2 (____9____30832),
       .Q (____9_9__30897));
  xor2s1 _______439250(.DIN1 (____9_0__30838), .DIN2 (____9____30860),
       .Q (____9____30861));
  nnd2s1 _______439251(.DIN1 (____9____30858), .DIN2 (_________28246),
       .Q (____9____30859));
  nnd2s1 ______439252(.DIN1 (____9____30855), .DIN2 (____0____31818),
       .Q (____9____30857));
  and2s1 _____0_439253(.DIN1 (____9____30855), .DIN2 (____90___30821),
       .Q (____9____30856));
  and2s1 _____0_439254(.DIN1 (____0_0__34541), .DIN2 (____9____30853),
       .Q (____9_0__30854));
  nor2s1 _______439255(.DIN1 (_____________________18662), .DIN2
       (____90___30824), .Q (____9____30852));
  nor2s1 _______439256(.DIN1 (___0__18915), .DIN2 (____9____30858), .Q
       (____99___30902));
  nor2s1 _____439257(.DIN1 (____0____29108), .DIN2 (____909__30827), .Q
       (____9____30886));
  dffacs1 ________________9_439258(.CLRB (reset), .CLK (clk), .DIN
       (____90___30823), .Q (____________9_));
  dffacs1 __________________439259(.CLRB (reset), .CLK (clk), .DIN
       (____9____30829), .QN (_________34455));
  hi1s1 _______439260(.DIN (____0_0__30916), .Q (____9____30851));
  nor2s1 _______439261(.DIN1 (________19094), .DIN2 (_________30808),
       .Q (____9____30850));
  nnd2s1 _____439262(.DIN1 (____9____30848), .DIN2 (____9____30847), .Q
       (____9____30849));
  nnd2s1 _______439263(.DIN1 (____9____30848), .DIN2 (outData[31]), .Q
       (____9_0__30846));
  nor2s1 _______439264(.DIN1 (____9____30847), .DIN2 (____9____30848),
       .Q (____9_9__30845));
  nor2s1 _______439265(.DIN1 (_________30686), .DIN2 (_____9___30817),
       .Q (____9____30891));
  nor2s1 _______439266(.DIN1 (outData[31]), .DIN2 (____9____30848), .Q
       (____0____30925));
  nnd2s1 _______439267(.DIN1 (_________29460), .DIN2 (_____9___30813),
       .Q (____9____30876));
  nor2s1 _______439268(.DIN1 (____9____30844), .DIN2 (______9__30809),
       .Q (____9_0__30881));
  xor2s1 _______439269(.DIN1 (_________30798), .DIN2 (_________31326),
       .Q (____9____30877));
  xor2s1 _______439270(.DIN1 (_________30572), .DIN2 (____9____30831),
       .Q (_____0___34148));
  xnr2s1 _______439271(.DIN1 (_________34487), .DIN2 (_________33852),
       .Q (____9____30843));
  hi1s1 _____9_439272(.DIN (____9____30858), .Q (____9____30842));
  xor2s1 _______439273(.DIN1 (_____0___29177), .DIN2 (_____00__31093),
       .Q (____9____30841));
  nnd2s1 _______439274(.DIN1 (_________30802), .DIN2 (___9____19692),
       .Q (____9____30840));
  nnd2s1 _______439275(.DIN1 (_________29461), .DIN2 (_____9___30812),
       .Q (____9____30875));
  nnd2s1 _______439276(.DIN1 (____9_0__30838), .DIN2 (_________30806),
       .Q (____9_9__30863));
  nor2s1 _____0_439277(.DIN1 (____9____29057), .DIN2 (____90___30826),
       .Q (____9____30869));
  xor2s1 _______439278(.DIN1 (_________30685), .DIN2 (_____9___30816),
       .Q (____9_9__30837));
  xnr2s1 ______439279(.DIN1 (______9__34440), .DIN2 (_________33852),
       .Q (____9____30836));
  nnd2s1 _______439280(.DIN1 (_________30797), .DIN2 (_____9__19561),
       .Q (____9____30835));
  nor2s1 _______439281(.DIN1 (_________30780), .DIN2 (_________30794),
       .Q (____9____30834));
  xor2s1 _______439282(.DIN1 (_________30782), .DIN2 (_____0___33866),
       .Q (____9____30833));
  nor2s1 _______439283(.DIN1 (_________30559), .DIN2 (____9____30831),
       .Q (____9____30832));
  xor2s1 _______439284(.DIN1 (_________33852), .DIN2 (_____0___32104),
       .Q (____9____30865));
  nnd2s1 _______439285(.DIN1 (_________30799), .DIN2 (________20251),
       .Q (____0_0__30916));
  xor2s1 _______439286(.DIN1 (_________30785), .DIN2 (________19986),
       .Q (______9__34094));
  xnr2s1 _____0_439287(.DIN1 (_________30738), .DIN2 (_________30777),
       .Q (_________31031));
  xor2s1 _______439288(.DIN1 (_________30766), .DIN2 (_________30587),
       .Q (____9____30830));
  nnd2s1 ______439289(.DIN1 (_________30792), .DIN2 (_________33279),
       .Q (____9____30829));
  nor2s1 _____439290(.DIN1 (_________34487), .DIN2 (_________33852), .Q
       (____9_0__30828));
  hi1s1 _______439291(.DIN (____90___30826), .Q (____909__30827));
  and2s1 ______439292(.DIN1 (_________33852), .DIN2 (_________34487),
       .Q (____90___30825));
  xor2s1 _______439293(.DIN1 (_________29682), .DIN2 (______9__30800),
       .Q (____90___30824));
  nnd2s1 _______439294(.DIN1 (_________30787), .DIN2 (__9_____26934),
       .Q (____90___30823));
  or2s1 ______439295(.DIN1 (____9_9__31781), .DIN2 (____90___30821), .Q
       (____90___30822));
  xor2s1 _______439296(.DIN1 (_________30756), .DIN2 (____9_9__31781),
       .Q (____9____30855));
  xor2s1 _______439297(.DIN1 (_________30761), .DIN2 (______9__30754),
       .Q (______0__33292));
  xor2s1 _______439298(.DIN1 (_________30762), .DIN2
       (_________________0___18607), .Q (____9____30858));
  nnd2s1 _____9_439299(.DIN1 (_________33852), .DIN2 (_________28880),
       .Q (____900__30820));
  nor2s1 _____9_439300(.DIN1 (______9__34440), .DIN2 (_________33852),
       .Q (_____99__30819));
  and2s1 _____9_439301(.DIN1 (_________33852), .DIN2 (______9__34440),
       .Q (_____9___30818));
  nor2s1 _____439302(.DIN1 (_________30663), .DIN2 (_____9___30816), .Q
       (_____9___30817));
  nnd2s1 _____439303(.DIN1 (_____9___30814), .DIN2 (_________30648), .Q
       (_____9___30815));
  hi1s1 _____0_439304(.DIN (_____9___30812), .Q (_____9___30813));
  xor2s1 ______439305(.DIN1 (_________34488), .DIN2 (_____0___33226),
       .Q (_____9___30811));
  xor2s1 _______439306(.DIN1 (_____0___33226), .DIN2 (_____0___32104),
       .Q (_____90__30810));
  xor2s1 _______439307(.DIN1 (_________30746), .DIN2 (_________28828),
       .Q (______9__30809));
  nor2s1 _______439308(.DIN1 (_________31653), .DIN2 (_________30771),
       .Q (_________30808));
  nnd2s1 _______439309(.DIN1 (_________30769), .DIN2 (_________30712),
       .Q (____9____30844));
  xor2s1 _______439310(.DIN1 (________20588), .DIN2 (_____9___34042),
       .Q (_________31067));
  xor2s1 _______439311(.DIN1 (_________30770), .DIN2 (_________30807),
       .Q (____9____30848));
  or2s1 _______439312(.DIN1 (_________30805), .DIN2 (_________30804),
       .Q (_________30806));
  and2s1 _____439313(.DIN1 (_________30804), .DIN2 (_________30805), .Q
       (_________30803));
  nnd2s1 _____9_439314(.DIN1 (_____9___30719), .DIN2 (_________30768),
       .Q (_________30802));
  nnd2s1 _______439315(.DIN1 (_________30786), .DIN2 (_________34660),
       .Q (_________30801));
  nnd2s1 _______439316(.DIN1 (______0__30764), .DIN2 (_________30405),
       .Q (____90___30826));
  or2s1 _____0_439317(.DIN1 (_________29664), .DIN2 (______9__30800),
       .Q (____9____30839));
  xor2s1 _______439318(.DIN1 (_____0___30734), .DIN2 (_____0___30728),
       .Q (_________32042));
  nnd2s1 _______439319(.DIN1 (_________30765), .DIN2 (_________30668),
       .Q (____0____30955));
  nnd2s1 ______439320(.DIN1 (_________30790), .DIN2 (_________30602),
       .Q (____9____30853));
  or2s1 _______439321(.DIN1 (________20587), .DIN2 (_____9___34042), .Q
       (_________30799));
  nnd2s1 _______439322(.DIN1 (_________30752), .DIN2 (__9_____26763),
       .Q (_________30798));
  nnd2s1 _______439323(.DIN1 (_________30753), .DIN2 (__99____27118),
       .Q (_________30797));
  xor2s1 _______439324(.DIN1 (_____0___30277), .DIN2 (_________30795),
       .Q (_________30796));
  nor2s1 _______439325(.DIN1 (_________30428), .DIN2 (_________30750),
       .Q (_________30794));
  nor2s1 _______439326(.DIN1 (_________30389), .DIN2 (_________30748),
       .Q (____9____30831));
  nnd2s1 _______439327(.DIN1 (_________30739), .DIN2 (_________30776),
       .Q (_________31027));
  nnd2s1 _______439328(.DIN1 (_________30755), .DIN2 (_________30760),
       .Q (____9_0__30838));
  xor2s1 ______439329(.DIN1 (_____0___30731), .DIN2 (_____90__31526),
       .Q (_____9___30812));
  dffacs1 ___________________439330(.CLRB (reset), .CLK (clk), .DIN
       (_________30767), .QN (_________________18709));
  nor2s1 _______439331(.DIN1 (_________34488), .DIN2 (____9____33600),
       .Q (_________30793));
  xor2s1 _______439332(.DIN1 (_________30406), .DIN2 (______9__30763),
       .Q (_________30792));
  and2s1 _______439333(.DIN1 (____9____33600), .DIN2 (_________34488),
       .Q (______0__30791));
  and2s1 _____9_439334(.DIN1 (_____0___30729), .DIN2 (_________34475),
       .Q (_________30788));
  nnd2s1 _____9_439335(.DIN1 (_____0___30732), .DIN2 (inData[12]), .Q
       (_________30787));
  hi1s1 ______439336(.DIN (_________30786), .Q (_____9___30814));
  nnd2s1 _______439337(.DIN1 (_____0___30727), .DIN2 (_____9___30722),
       .Q (_____9___30816));
  nnd2s1 _______439338(.DIN1 (______0__30736), .DIN2 (_________30711),
       .Q (____90___30821));
  nor2s1 ______439339(.DIN1 (_____9___28610), .DIN2 (_____0___30730),
       .Q (_____00__31093));
  xnr2s1 _______439340(.DIN1 (_________30751), .DIN2 (__9_____27029),
       .Q (_________33852));
  xor2s1 _____9_439341(.DIN1 (______0__30494), .DIN2 (_________30747),
       .Q (_________30785));
  nnd2s1 _____0_439342(.DIN1 (____0____30918), .DIN2 (______0__18849),
       .Q (______0__30784));
  nor2s1 _____0_439343(.DIN1 (______0__18849), .DIN2 (____0____30918),
       .Q (______9__30783));
  nor2s1 _______439344(.DIN1 (_________30781), .DIN2 (_________30742),
       .Q (_________30782));
  nor2s1 _______439345(.DIN1 (_________31578), .DIN2 (_____9___30725),
       .Q (_________30780));
  nor2s1 _______439346(.DIN1 (outData[31]), .DIN2 (_________30795), .Q
       (_________30779));
  and2s1 _______439347(.DIN1 (_________30795), .DIN2 (outData[31]), .Q
       (_________30778));
  and2s1 ______439348(.DIN1 (_________30737), .DIN2 (_________30776),
       .Q (_________30777));
  nor2s1 _______439349(.DIN1 (_________30772), .DIN2 (_________30795),
       .Q (_________30775));
  nor2s1 _______439350(.DIN1 (outData[31]), .DIN2 (______0__31130), .Q
       (______0__30774));
  and2s1 _______439351(.DIN1 (_________30795), .DIN2 (_________30772),
       .Q (______9__30773));
  hi1s1 _____9_439352(.DIN (_________30770), .Q (_________30771));
  nnd2s1 _______439353(.DIN1 (_____00__30726), .DIN2 (___0__18931), .Q
       (_________30769));
  nnd2s1 _______439354(.DIN1 (_________30669), .DIN2 (_____9___30723),
       .Q (_________30768));
  nnd2s1 _______439355(.DIN1 (_____90__30717), .DIN2 (________21868),
       .Q (_________30767));
  xor2s1 _______439356(.DIN1 (_________34456), .DIN2 (____0_0__31861),
       .Q (_________30766));
  or2s1 _______439357(.DIN1 (_________________18746), .DIN2
       (_____9___30720), .Q (_________30765));
  or2s1 _______439358(.DIN1 (_________30384), .DIN2 (______9__30763),
       .Q (______0__30764));
  xor2s1 ______439359(.DIN1 (______9__30707), .DIN2 (_________30654),
       .Q (_________30762));
  nnd2s1 _______439360(.DIN1 (____0____34542), .DIN2 (_________30760),
       .Q (_________30761));
  or2s1 _____0_439361(.DIN1 (_________30758), .DIN2 (_________30757),
       .Q (_________30759));
  nnd2s1 _______439362(.DIN1 (_____09__30735), .DIN2 (_____9___30724),
       .Q (_________30756));
  nnd2s1 _______439363(.DIN1 (____0____34542), .DIN2 (______9__30754),
       .Q (_________30755));
  xor2s1 _______439364(.DIN1 (_________30701), .DIN2 (_________33925),
       .Q (______9__30800));
  xor2s1 _______439365(.DIN1 (_________30695), .DIN2 (_____0___33031),
       .Q (_________30786));
  xor2s1 _______439366(.DIN1 (_________30706), .DIN2 (_________30667),
       .Q (_________30790));
  nnd2s1 ______439367(.DIN1 (____0____34543), .DIN2 (_________30696),
       .Q (_________30753));
  or2s1 ______439368(.DIN1 (__9_____26753), .DIN2 (_________30751), .Q
       (_________30752));
  nor2s1 ______439369(.DIN1 (_________30658), .DIN2 (______9__30716),
       .Q (_________30750));
  nor2s1 _____0_439370(.DIN1
       (______________0___________________9__18827), .DIN2
       (______0__30745), .Q (_________30749));
  nor2s1 ______439371(.DIN1 (_____0___30463), .DIN2 (_________30747),
       .Q (_________30748));
  nnd2s1 _______439372(.DIN1 (______0__30745), .DIN2
       (______________0___________________9__18827), .Q
       (_________30746));
  xor2s1 _______439373(.DIN1 (____0___21079), .DIN2 (_________30743),
       .Q (______9__30744));
  nor2s1 _______439374(.DIN1 (_____________18905), .DIN2
       (_________30740), .Q (_________30741));
  nnd2s1 _______439375(.DIN1 (_________30738), .DIN2 (_________30737),
       .Q (_________30739));
  nnd2s1 _______439376(.DIN1 (_________30714), .DIN2 (_______19047), .Q
       (_________30770));
  xor2s1 _______439377(.DIN1 (_________30699), .DIN2 (___90___23352),
       .Q (_________30804));
  xor2s1 _______439378(.DIN1 (______0__30698), .DIN2 (_________30678),
       .Q (_____9___34042));
  hi1s1 _______439379(.DIN (____9____33600), .Q (_____0___33226));
  hi1s1 _______439380(.DIN (_____09__30735), .Q (______0__30736));
  xor2s1 _______439381(.DIN1 (_________34475), .DIN2 (_____0___30733),
       .Q (_____0___30734));
  nor2s1 ______439382(.DIN1 (_________30703), .DIN2 (________20485), .Q
       (_____0___30732));
  nnd2s1 _____9_439383(.DIN1 (_________30700), .DIN2 (_________30694),
       .Q (_____0___30731));
  and2s1 _______439384(.DIN1 (_________28719), .DIN2 (_________34456),
       .Q (_____0___30730));
  or2s1 ______439385(.DIN1 (_____0___30728), .DIN2 (_____9___33396), .Q
       (_____0___30729));
  xor2s1 _____9_439386(.DIN1 (_____9___30718), .DIN2 (____9____30860),
       .Q (_____0___30727));
  nnd2s1 _______439387(.DIN1 (_____9___33396), .DIN2 (_____0___30728),
       .Q (_________30789));
  hi1s1 _______439388(.DIN (____0____34543), .Q (_____00__30726));
  nor2s1 ______439389(.DIN1 (______9__30651), .DIN2 (_________30702),
       .Q (_____9___30725));
  nor2s1 _______439390(.DIN1 (_____09__30102), .DIN2 (_________30743),
       .Q (_________30742));
  nnd2s1 _______439391(.DIN1 (_____9___30724), .DIN2
       (______________________________________0_____________18891), .Q
       (_________30776));
  hi1s1 _____9_439392(.DIN (_________30740), .Q (______0__31130));
  hi1s1 _______439393(.DIN (______0__30745), .Q (____0____30918));
  xor2s1 _____0_439394(.DIN1
       (______________________________________0_____________18885),
       .DIN2 (_________30681), .Q (____9____33600));
  xor2s1 _______439395(.DIN1 (_________30713), .DIN2 (____0___22082),
       .Q (_________30795));
  nnd2s1 ______439396(.DIN1 (_____9___30722), .DIN2 (_____9___30629),
       .Q (_____9___30723));
  or2s1 ______439397(.DIN1 (_________________18766), .DIN2
       (_____0___30733), .Q (_____9___30721));
  xor2s1 ______439398(.DIN1 (______9__30661), .DIN2 (______0__32594),
       .Q (_____9___30720));
  nnd2s1 ______439399(.DIN1 (_____9___30718), .DIN2 (_____9___30722),
       .Q (_____9___30719));
  nnd2s1 _______439400(.DIN1 (______0__30689), .DIN2 (__99____27118),
       .Q (_____90__30717));
  nor2s1 _____0_439401(.DIN1 (_________30645), .DIN2 (_________30690),
       .Q (______9__30763));
  nnd2s1 _______439402(.DIN1 (_________30692), .DIN2 (_____9___30625),
       .Q (_____09__30735));
  and2s1 _______439403(.DIN1 (_____0___30733), .DIN2
       (_________________18700), .Q (_________30757));
  nor2s1 _______439404(.DIN1 (_________________18700), .DIN2
       (_____0___30733), .Q (_________30758));
  dffacs1 __________________439405(.CLRB (reset), .CLK (clk), .DIN
       (_________30684), .QN (________________18724));
  nor2s1 _______439406(.DIN1 (_________33835), .DIN2 (_________30673),
       .Q (______9__30716));
  and2s1 ______439407(.DIN1 (_____0___30733), .DIN2
       (_________________18766), .Q (_________30715));
  or2s1 ______439408(.DIN1 (________19075), .DIN2 (_________30713), .Q
       (_________30714));
  nnd2s1 _______439409(.DIN1 (_________30677), .DIN2 (_________35110),
       .Q (_________30712));
  nor2s1 _______439410(.DIN1 (______0__30680), .DIN2 (_________30676),
       .Q (_________30751));
  nnd2s1 _______439411(.DIN1 (_________30711), .DIN2 (______9__30537),
       .Q (_________30737));
  nor2s1 _______439412(.DIN1 (_____99__30631), .DIN2 (______0__30671),
       .Q (_________30738));
  nor2s1 _______439413(.DIN1 (______9__30697), .DIN2 (______9__30679),
       .Q (_________30747));
  xor2s1 _______439414(.DIN1 (________25103), .DIN2 (_________30656),
       .Q (______0__30745));
  xor2s1 _______439415(.DIN1 (_________30650), .DIN2 (_________30710),
       .Q (_________30740));
  dffacs1 ___________________439416(.CLRB (reset), .CLK (clk), .DIN
       (_________30683), .QN (_________34479));
  xor2s1 _______439417(.DIN1 (_________________18728), .DIN2
       (_________30705), .Q (______0__30708));
  xor2s1 _______439418(.DIN1 (_________30691), .DIN2
       (_______________18881), .Q (______9__30707));
  xor2s1 ______439419(.DIN1 (_________________18746), .DIN2
       (_________30705), .Q (_________30706));
  nnd2s1 _____9_439420(.DIN1 (_________30666), .DIN2 (_________34966),
       .Q (_________30704));
  xor2s1 _____9_439421(.DIN1 (_________34497), .DIN2 (_____09__30641),
       .Q (_________30703));
  xor2s1 _____9_439422(.DIN1 (_________30621), .DIN2 (_________30643),
       .Q (______0__33258));
  dffacs1 __________________439423(.CLRB (reset), .CLK (clk), .DIN
       (______0__30662), .QN (_________34456));
  hi1s1 _______439424(.DIN (_____0___30733), .Q (_____9___33396));
  nor2s1 _______439425(.DIN1 (_________33835), .DIN2 (_________30672),
       .Q (_________30702));
  nnd2s1 _______439426(.DIN1 (_________30660), .DIN2 (_________29507),
       .Q (_________30701));
  nnd2s1 _______439427(.DIN1 (_____9___30360), .DIN2 (____0____34544),
       .Q (_________30700));
  xor2s1 _______439428(.DIN1 (_____0___30635), .DIN2 (_________32644),
       .Q (_________30699));
  nor2s1 _______439429(.DIN1 (______9__30697), .DIN2 (_________30653),
       .Q (______0__30698));
  nnd2s1 _______439430(.DIN1 (_________30674), .DIN2 (_____0___30633),
       .Q (_________30696));
  and2s1 _______439431(.DIN1 (_________30694), .DIN2 (____0____34544),
       .Q (_________30695));
  nnd2s1 _____439432(.DIN1 (_________30688), .DIN2 (_________30498), .Q
       (_________30760));
  hi1s1 _______439433(.DIN (_________30711), .Q (_____9___30724));
  xor2s1 _______439434(.DIN1 (______9__30670), .DIN2 (_________30693),
       .Q (_________30743));
  nnd2s1 _____9_439435(.DIN1 (_________30691), .DIN2 (_____9___30626),
       .Q (_________30692));
  nor2s1 _______439436(.DIN1 (_____90__28983), .DIN2 (_________30647),
       .Q (_________30690));
  xor2s1 _______439437(.DIN1 (_________29509), .DIN2 (_________30659),
       .Q (______0__30689));
  nnd2s1 _______439438(.DIN1 (_________30705), .DIN2 (____9___19109),
       .Q (_________30687));
  nor2s1 _______439439(.DIN1 (_________30556), .DIN2 (_________30685),
       .Q (_________30686));
  nnd2s1 _____0_439440(.DIN1 (_____0___30640), .DIN2 (_________30588),
       .Q (_________30684));
  nnd2s1 _____439441(.DIN1 (_____0___30639), .DIN2 (________21770), .Q
       (_________30683));
  xor2s1 ______439442(.DIN1 (_________30620), .DIN2 (_________32410),
       .Q (_________30709));
  xor2s1 ______439443(.DIN1 (_________30617), .DIN2 (_________28828),
       .Q (_____9___30722));
  dffacs1 ___________________439444(.CLRB (reset), .CLK (clk), .DIN
       (_________30644), .Q (_________________18693));
  xor2s1 _____0_439445(.DIN1 (_________30619), .DIN2 (___0____21656),
       .Q (_____0___30733));
  hi1s1 _______439446(.DIN (_________32070), .Q (_________30682));
  nor2s1 _______439447(.DIN1 (______0__30680), .DIN2 (_________30675),
       .Q (_________30681));
  and2s1 _______439448(.DIN1 (______0__30652), .DIN2 (_________30678),
       .Q (______9__30679));
  nnd2s1 _______439449(.DIN1 (_____0___30634), .DIN2 (_________30649),
       .Q (_________30677));
  nor2s1 _______439450(.DIN1
       (______________________________________0_____________18885),
       .DIN2 (_________30675), .Q (_________30676));
  hi1s1 _______439451(.DIN (_________30672), .Q (_________30673));
  and2s1 ______439452(.DIN1 (_________30655), .DIN2 (_____9___30628),
       .Q (______0__30671));
  nor2s1 ______439453(.DIN1 (________19104), .DIN2 (_____0___30637), .Q
       (_________30713));
  and2s1 _______439454(.DIN1 (______9__30670), .DIN2 (_________30156),
       .Q (_________30781));
  nor2s1 ______439455(.DIN1 (_____9___30630), .DIN2 (_________30669),
       .Q (_____9___30718));
  xor2s1 _______439456(.DIN1 (__9_____26368), .DIN2 (_________30657),
       .Q (_________30711));
  nnd2s1 ______439457(.DIN1 (_________30664), .DIN2 (_________30667),
       .Q (_________30668));
  xor2s1 _______439458(.DIN1 (_________30646), .DIN2 (_________28977),
       .Q (_________30666));
  nnd2s1 _______439459(.DIN1 (_________30664), .DIN2
       (_________________18728), .Q (_________30665));
  nor2s1 ______439460(.DIN1 (______0__34668), .DIN2 (_____0___30638),
       .Q (_________30663));
  nnd2s1 _______439461(.DIN1 (_________30618), .DIN2 (_________33279),
       .Q (______0__30662));
  or2s1 _____9_439462(.DIN1 (_________30667), .DIN2 (_________30664),
       .Q (______9__30661));
  nnd2s1 ______439463(.DIN1 (_________30659), .DIN2 (______9__29511),
       .Q (_________30660));
  nnd2s1 _______439464(.DIN1 (_____90__30623), .DIN2 (______0__30642),
       .Q (_________30688));
  nor2s1 _______439465(.DIN1 (________26070), .DIN2 (_________30657),
       .Q (_________30658));
  xor2s1 _______439466(.DIN1 (_________30655), .DIN2 (_________30654),
       .Q (_________30656));
  hi1s1 _______439467(.DIN (______0__30652), .Q (_________30653));
  and2s1 ______439468(.DIN1 (_________30657), .DIN2
       (_______________18879), .Q (______9__30651));
  xor2s1 _______439469(.DIN1 (_____0___30636), .DIN2 (______0__35098),
       .Q (_________30650));
  nnd2s1 _____0_439470(.DIN1 (_____00__30632), .DIN2 (_________30649),
       .Q (_________30674));
  nor2s1 _____439471(.DIN1 (_______________18879), .DIN2
       (_________30657), .Q (_________30672));
  nor2s1 _______439472(.DIN1 (_________30603), .DIN2 (_________30616),
       .Q (_________32070));
  hi1s1 _______439473(.DIN (_________34660), .Q (_________30648));
  and2s1 _______439474(.DIN1 (_________30646), .DIN2
       (________________18722), .Q (_________30647));
  nor2s1 _______439475(.DIN1 (________________18722), .DIN2
       (_________30646), .Q (_________30645));
  nnd2s1 _______439476(.DIN1 (_________30609), .DIN2 (________22376),
       .Q (_________30644));
  nnd2s1 _______439477(.DIN1 (______9__30622), .DIN2 (______0__30642),
       .Q (_________30643));
  nnd2s1 _______439478(.DIN1 (____________9___18692), .DIN2
       (_____________0___18708), .Q (_____09__30641));
  nnd2s1 _______439479(.DIN1 (_________30610), .DIN2 (___9____19692),
       .Q (_____0___30640));
  nnd2s1 ______439480(.DIN1 (_________30608), .DIN2 (__99____27118), .Q
       (_____0___30639));
  xor2s1 ______439481(.DIN1 (_________34664), .DIN2 (______0__30607),
       .Q (_________30691));
  nnd2s1 _______439482(.DIN1 (___0_____27729), .DIN2
       (_____________0___18708), .Q (_________30694));
  hi1s1 ______439483(.DIN (_____0___30638), .Q (_________30685));
  hi1s1 _______439484(.DIN (_________30664), .Q (_________30705));
  and2s1 _____439485(.DIN1 (_____0___30636), .DIN2 (_____0__19262), .Q
       (_____0___30637));
  xor2s1 _____0_439486(.DIN1 (_________30597), .DIN2 (___90___23353),
       .Q (_____0___30635));
  nnd2s1 _______439487(.DIN1 (_____0___30633), .DIN2 (_____00__30632),
       .Q (_____0___30634));
  nor2s1 _____9_439488(.DIN1 (_____9___30627), .DIN2 (_________30654),
       .Q (_____99__30631));
  hi1s1 _____9_439489(.DIN (_____9___30629), .Q (_____9___30630));
  nnd2s1 _______439490(.DIN1 (_________30654), .DIN2 (_____9___30627),
       .Q (_____9___30628));
  or2s1 _______439491(.DIN1 (_________31940), .DIN2 (_________30654),
       .Q (_____9___30626));
  nnd2s1 _______439492(.DIN1 (_________30654), .DIN2 (_________31940),
       .Q (_____9___30625));
  nnd2s1 ______439493(.DIN1 (_________34662), .DIN2 (____9____30847),
       .Q (______0__30652));
  xor2s1 _____9_439494(.DIN1 (_________30593), .DIN2 (_____9___30624),
       .Q (______9__30670));
  nor2s1 _____9_439495(.DIN1 (___________0___18883), .DIN2
       (______9__30606), .Q (_________30675));
  nor2s1 _______439496(.DIN1 (____9____30847), .DIN2 (_________34662),
       .Q (______9__30697));
  nnd2s1 ______439497(.DIN1 (______9__30622), .DIN2 (_________30621),
       .Q (_____90__30623));
  xor2s1 _______439498(.DIN1 (_________34452), .DIN2 (_________30585),
       .Q (_________30620));
  xor2s1 ______439499(.DIN1 (_________30580), .DIN2 (_____0___32570),
       .Q (_________30619));
  xor2s1 _______439500(.DIN1 (_________34666), .DIN2 (_________34740),
       .Q (_________30618));
  xor2s1 _______439501(.DIN1 (_________30583), .DIN2 (_________35076),
       .Q (_____0___30638));
  xor2s1 _______439502(.DIN1 (______0__30582), .DIN2 (______0__35098),
       .Q (_________30664));
  nor2s1 _____0_439503(.DIN1 (_________30613), .DIN2 (_________30614),
       .Q (_________30617));
  nor2s1 _______439504(.DIN1 (_________________0___18607), .DIN2
       (______9__30599), .Q (_________30616));
  nnd2s1 _____0_439505(.DIN1 (_________30614), .DIN2 (_________30613),
       .Q (_____9___30629));
  nor2s1 _____439506(.DIN1 (_________30612), .DIN2 (_________30605), .Q
       (______0__30680));
  nor2s1 _____9_439507(.DIN1 (_____09__29455), .DIN2 (_________30601),
       .Q (_________30659));
  nnd2s1 _______439508(.DIN1 (_________30611), .DIN2 (____0___22723),
       .Q (_________30649));
  xnr2s1 ______439509(.DIN1 (____9____31798), .DIN2 (_________30571),
       .Q (_________30657));
  xor2s1 _____9_439510(.DIN1 (_________30568), .DIN2 (_____90__31526),
       .Q (_________30610));
  nnd2s1 _______439511(.DIN1 (_________30577), .DIN2 (__99____27118),
       .Q (_________30609));
  xor2s1 _____0_439512(.DIN1 (______0__29456), .DIN2 (______0__30600),
       .Q (_________30608));
  nnd2s1 _____0_439513(.DIN1 (_____0___30549), .DIN2 (_________30579),
       .Q (______0__30642));
  xor2s1 _______439514(.DIN1 (_________30567), .DIN2 (______0__30607),
       .Q (_________30646));
  dffacs1 _________________0_439515(.CLRB (reset), .CLK (clk), .DIN
       (_________30589), .Q (_____________0___18708));
  hi1s1 _______439516(.DIN (_________30605), .Q (______9__30606));
  nnd2s1 _______439517(.DIN1 (_________30576), .DIN2 (___90___23354),
       .Q (_________30615));
  xor2s1 _______439518(.DIN1 (_________30557), .DIN2
       (_________________0___18633), .Q (_________30655));
  nnd2s1 _______439519(.DIN1 (_________30604), .DIN2
       (______________0______________________18826), .Q
       (_____00__30632));
  nnd2s1 _______439520(.DIN1 (______0__30574), .DIN2 (________19241),
       .Q (_____0___30636));
  xor2s1 _______439521(.DIN1 (_________30561), .DIN2
       (______________________________________0_____________18891), .Q
       (_________30654));
  nor2s1 _______439522(.DIN1 (_____0___33866), .DIN2 (_________30598),
       .Q (_________30603));
  nor2s1 _______439523(.DIN1 (_____0___29454), .DIN2 (______0__30600),
       .Q (_________30601));
  nor2s1 ______439524(.DIN1 (______0__30510), .DIN2 (_________30598),
       .Q (______9__30599));
  nnd2s1 _____0_439525(.DIN1 (_____0___30550), .DIN2 (_________30578),
       .Q (______9__30622));
  xor2s1 _______439526(.DIN1 (_________30596), .DIN2 (_________30595),
       .Q (_________30597));
  nnd2s1 _______439527(.DIN1 (______0__30555), .DIN2 (__99____27118),
       .Q (_________30594));
  xor2s1 ______439528(.DIN1 (_________30592), .DIN2 (______9__30573),
       .Q (_________30593));
  hi1s1 _____9_439529(.DIN (_________30604), .Q (_________30611));
  xor2s1 ______439530(.DIN1 (_____9___30540), .DIN2 (____99___32749),
       .Q (_________30614));
  xor2s1 _______439531(.DIN1 (_____99__30544), .DIN2 (______0__30591),
       .Q (_________30605));
  nnd2s1 ______439532(.DIN1 (_____0___30548), .DIN2 (inData[16]), .Q
       (______9__30590));
  nnd2s1 _______439533(.DIN1 (_____0___30547), .DIN2 (___0____20745),
       .Q (_________30589));
  or2s1 _______439534(.DIN1 (_____0___32299), .DIN2 (_____0___30552),
       .Q (_________30588));
  xor2s1 ______439535(.DIN1 (_________________18727), .DIN2
       (_________30584), .Q (_________30586));
  xor2s1 _____0_439536(.DIN1 (___09____28053), .DIN2 (_________30584),
       .Q (_________30585));
  xor2s1 _____0_439537(.DIN1 (____0____29140), .DIN2
       (____________9___18707), .Q (_________30583));
  xor2s1 _____439538(.DIN1 (_________30517), .DIN2 (_________30563), .Q
       (______0__30582));
  nnd2s1 ______439539(.DIN1 (_____0___30551), .DIN2 (___090___28046),
       .Q (_________30602));
  hi1s1 _______439540(.DIN (______9__30581), .Q (______0__33175));
  xor2s1 _______439541(.DIN1 (_________30534), .DIN2 (_________31926),
       .Q (_________30580));
  hi1s1 _______439542(.DIN (_________30578), .Q (_________30579));
  xor2s1 _______439543(.DIN1 (_________30523), .DIN2 (_________30431),
       .Q (_________30577));
  nnd2s1 _____9_439544(.DIN1 (_________30596), .DIN2 (________23242),
       .Q (_________30576));
  or2s1 _____9_439545(.DIN1 (________19614), .DIN2 (______9__30573), .Q
       (______0__30574));
  nor2s1 ______439546(.DIN1 (_________30558), .DIN2 (_________30536),
       .Q (_________30572));
  nnd2s1 _______439547(.DIN1 (_____9___30539), .DIN2 (_________30560),
       .Q (_________30571));
  xor2s1 _____0_439548(.DIN1 (_________30522), .DIN2 (_________30527),
       .Q (_________30604));
  nnd2s1 _____439549(.DIN1 (_____9___30543), .DIN2 (_________30440), .Q
       (_____0___30633));
  nnd2s1 _______439550(.DIN1 (_________30569), .DIN2 (_______19039), .Q
       (_________30570));
  xor2s1 _______439551(.DIN1 (_________30512), .DIN2 (_________30352),
       .Q (_________30568));
  nor2s1 _______439552(.DIN1 (_________30486), .DIN2 (_________30533),
       .Q (_________30567));
  nnd2s1 _______439553(.DIN1 (_________30584), .DIN2 (______0__30564),
       .Q (_________30566));
  nor2s1 _______439554(.DIN1 (______0__30564), .DIN2 (_________30584),
       .Q (_________30565));
  nnd2s1 _______439555(.DIN1 (____0____29107), .DIN2
       (____________9___18707), .Q (_________30562));
  xor2s1 _______439556(.DIN1 (_____09__30554), .DIN2 (_________30506),
       .Q (_________30575));
  xor2s1 _______439557(.DIN1 (_________30513), .DIN2 (_____0___30371),
       .Q (______9__30581));
  and2s1 _______439558(.DIN1 (_____90__30538), .DIN2 (_________30560),
       .Q (_________30561));
  nor2s1 _____9_439559(.DIN1 (_________30518), .DIN2 (_________30558),
       .Q (_________30559));
  nor2s1 ______439560(.DIN1 (______0__30520), .DIN2 (_________30528),
       .Q (_________30557));
  hi1s1 ______439561(.DIN (______0__34668), .Q (_________30556));
  xor2s1 _______439562(.DIN1 (_________30466), .DIN2 (_____9___30542),
       .Q (______0__30555));
  nor2s1 _______439563(.DIN1 (_________30477), .DIN2 (_________30532),
       .Q (______0__30600));
  xor2s1 ______439564(.DIN1 (_________30501), .DIN2 (_________30524),
       .Q (_________30578));
  nor2s1 ______439565(.DIN1 (______0__30500), .DIN2 (_________30525),
       .Q (______9__30754));
  and2s1 _______439566(.DIN1 (_________30569), .DIN2 (_____09__30554),
       .Q (_________30598));
  nnd2s1 _______439567(.DIN1 (______0__30530), .DIN2 (_________34436),
       .Q (_____0___30553));
  xor2s1 _____439568(.DIN1 (_________30387), .DIN2 (_________30492), .Q
       (_____0___30552));
  nnd2s1 _______439569(.DIN1 (______9__30529), .DIN2 (___09____28054),
       .Q (_____0___30551));
  hi1s1 _______439570(.DIN (_____0___30549), .Q (_____0___30550));
  nor2s1 _____439571(.DIN1 (______9__30509), .DIN2 (_____0___32299), .Q
       (_____0___30548));
  nnd2s1 ______439572(.DIN1 (_________30514), .DIN2 (__99____27118), .Q
       (_____0___30547));
  xor2s1 _______439573(.DIN1 (_________30471), .DIN2 (_____00__30545),
       .Q (_____0___30546));
  nor2s1 _____0_439574(.DIN1 (___9____25245), .DIN2 (_________30503),
       .Q (_____99__30544));
  nnd2s1 _______439575(.DIN1 (_____9___30542), .DIN2 (_________30438),
       .Q (_____9___30543));
  xor2s1 _______439576(.DIN1 (_________30467), .DIN2 (______9__28944),
       .Q (_____9___30540));
  nnd2s1 _______439577(.DIN1 (_____90__30538), .DIN2 (______9__30537),
       .Q (_____9___30539));
  and2s1 _______439578(.DIN1 (_________30495), .DIN2 (_____9___30624),
       .Q (_________30536));
  nor2s1 _______439579(.DIN1 (_________30433), .DIN2 (_________30497),
       .Q (______9__30573));
  hi1s1 _______439580(.DIN (_________30535), .Q (_________30596));
  xor2s1 ______439581(.DIN1 (_________30502), .DIN2
       (______________________________________0_____________18886), .Q
       (_________30534));
  and2s1 ______439582(.DIN1 (______0__30485), .DIN2 (_________30587),
       .Q (_________30533));
  and2s1 _____439583(.DIN1 (_________30479), .DIN2 (_________30531), .Q
       (_________30532));
  dffacs1 ________________9_439584(.CLRB (reset), .CLK (clk), .DIN
       (_________30480), .Q (____________9___18707));
  nnd2s1 ______439585(.DIN1 (_________30488), .DIN2 (______9__30353),
       .Q (_________30669));
  nnd2s1 _______439586(.DIN1 (_________30482), .DIN2 (_____09__30372),
       .Q (_____0___30549));
  xor2s1 _____9_439587(.DIN1 (_________30445), .DIN2 (______0__35098),
       .Q (_________30563));
  hi1s1 _______439588(.DIN (______0__30530), .Q (_________30569));
  hi1s1 _______439589(.DIN (______9__30529), .Q (_________30584));
  dffacs2 _____________________0_439590(.CLRB (reset), .CLK (clk), .DIN
       (______9__30484), .QN (_________________0___18660));
  nor2s1 _______439591(.DIN1 (_________30521), .DIN2 (_________30527),
       .Q (_________30528));
  xor2s1 _______439592(.DIN1 (______0__34441), .DIN2 (____0____33715),
       .Q (_________30526));
  and2s1 _______439593(.DIN1 (_________30469), .DIN2 (_________30524),
       .Q (_________30525));
  xor2s1 _______439594(.DIN1 (_________30443), .DIN2 (_________35076),
       .Q (_________30523));
  nor2s1 _______439595(.DIN1 (_________30521), .DIN2 (______0__30520),
       .Q (_________30522));
  xor2s1 _______439596(.DIN1 (______0__30475), .DIN2 (____0____33715),
       .Q (______9__30519));
  and2s1 _______439597(.DIN1 (_________30515), .DIN2 (_____9___30624),
       .Q (_________30518));
  nnd2s1 _______439598(.DIN1 (_________30499), .DIN2 (_________30516),
       .Q (_________30517));
  nnd2s1 _______439599(.DIN1 (_____0___30461), .DIN2
       (_______________18878), .Q (_________30560));
  nor2s1 _______439600(.DIN1 (_____9___30624), .DIN2 (_________30515),
       .Q (_________30558));
  xor2s1 _______439601(.DIN1 (______9__30326), .DIN2 (______9__30493),
       .Q (_________30535));
  xor2s1 _______439602(.DIN1 (_________29381), .DIN2 (_________30478),
       .Q (_________30514));
  xor2s1 _______439603(.DIN1 (______0__30399), .DIN2 (_________30481),
       .Q (_________30513));
  xor2s1 ______439604(.DIN1 (_________30377), .DIN2 (_________30487),
       .Q (_________30512));
  or2s1 _______439605(.DIN1 (_________________18699), .DIN2
       (____0____33715), .Q (_________30511));
  and2s1 _____0_439606(.DIN1 (_____9___30448), .DIN2 (_________34477),
       .Q (______0__30510));
  xor2s1 _______439607(.DIN1 (________________18723), .DIN2
       (________________18721), .Q (______9__30509));
  xor2s1 _______439608(.DIN1 (_____0__21085), .DIN2 (_________30507),
       .Q (_________30508));
  xnr2s1 _______439609(.DIN1 (_________34477), .DIN2 (_________30507),
       .Q (_________30506));
  and2s1 _______439610(.DIN1 (____0____33715), .DIN2
       (_________________18699), .Q (_________30505));
  xnr2s1 _______439611(.DIN1 (_____9___32930), .DIN2 (_________30507),
       .Q (______0__30530));
  xor2s1 _____9_439612(.DIN1 (_________30425), .DIN2 (_________30247),
       .Q (______9__30529));
  dffacs1 _______________439613(.CLRB (reset), .CLK (clk), .DIN
       (_____9___30452), .QN (__________));
  dffacs1 __________________439614(.CLRB (reset), .CLK (clk), .DIN
       (_____9___30453), .Q (______9__34470));
  nor2s1 _______439615(.DIN1 (________19221), .DIN2 (____0____33715),
       .Q (_________30504));
  nor2s1 _______439616(.DIN1 (________25125), .DIN2 (_________30502),
       .Q (_________30503));
  nor2s1 ______439617(.DIN1 (______0__30500), .DIN2 (_________30468),
       .Q (_________30501));
  and2s1 _______439618(.DIN1 (_________30434), .DIN2 (_________30496),
       .Q (_________30497));
  xor2s1 ______439619(.DIN1 (_________31519), .DIN2 (_____09__30464),
       .Q (_________30495));
  nnd2s1 _______439620(.DIN1 (_____0___30462), .DIN2 (_________30435),
       .Q (______0__30494));
  nnd2s1 ______439621(.DIN1 (_____0___30460), .DIN2 (_________31058),
       .Q (_____90__30538));
  nnd2s1 _____0_439622(.DIN1 (______9__30493), .DIN2 (_________30253),
       .Q (_____9___30541));
  nor2s1 _______439623(.DIN1 (_________30442), .DIN2 (_________30432),
       .Q (_____9___30542));
  nnd2s1 _______439624(.DIN1 (________________18721), .DIN2
       (_________30491), .Q (_________30492));
  nnd2s1 _______439625(.DIN1 (_________30507), .DIN2
       (_________________18765), .Q (_________30490));
  nor2s1 ______439626(.DIN1 (_________________18765), .DIN2
       (_________30507), .Q (_________30489));
  nnd2s1 _______439627(.DIN1 (_________30487), .DIN2 (_________30378),
       .Q (_________30488));
  nor2s1 _______439628(.DIN1 (________________18721), .DIN2
       (_________34740), .Q (_________30486));
  nnd2s1 _______439629(.DIN1 (_________34740), .DIN2
       (________________18721), .Q (______0__30485));
  nnd2s1 _______439630(.DIN1 (__9_____27031), .DIN2 (______0__30427),
       .Q (______9__30484));
  nor2s1 _______439631(.DIN1 (____09__21084), .DIN2 (_________30507),
       .Q (_________30483));
  nnd2s1 _______439632(.DIN1 (_________30481), .DIN2 (_________30400),
       .Q (_________30482));
  nor2s1 _____0_439633(.DIN1 (_________30374), .DIN2 (______9__30426),
       .Q (_________30480));
  nnd2s1 _______439634(.DIN1 (_________30478), .DIN2 (_________18862),
       .Q (_________30479));
  nor2s1 _______439635(.DIN1 (_________18862), .DIN2 (_________30478),
       .Q (_________30477));
  dffacs1 __________________439636(.CLRB (reset), .CLK (clk), .DIN
       (_________30423), .Q (________________18690));
  dffacs1 __________________439637(.CLRB (reset), .CLK (clk), .DIN
       (_________30422), .QN (_________34493));
  dffacs1 _________________0_439638(.CLRB (reset), .CLK (clk), .DIN
       (_________30424), .Q (_________18862));
  nor2s1 _______439639(.DIN1 (______0__30475), .DIN2 (_________30470),
       .Q (_________30476));
  xor2s1 ______439640(.DIN1 (_________30473), .DIN2 (_________30472),
       .Q (______9__30474));
  nnd2s1 _______439641(.DIN1 (_________30470), .DIN2 (______0__30475),
       .Q (_________30471));
  hi1s1 _______439642(.DIN (_________30468), .Q (_________30469));
  xor2s1 _____0_439643(.DIN1 (______9__34480), .DIN2 (_________31153),
       .Q (_________30467));
  xor2s1 _______439644(.DIN1 (______________0___________________9),
       .DIN2 (_________30439), .Q (_________30466));
  nor2s1 ______439645(.DIN1 (_____09__30464), .DIN2 (_________31519),
       .Q (______0__30465));
  and2s1 _______439646(.DIN1 (_____0___30462), .DIN2 (_________30421),
       .Q (_____0___30463));
  hi1s1 ____90_439647(.DIN (_____0___30460), .Q (_____0___30461));
  nor2s1 _______439648(.DIN1 (______0__34441), .DIN2 (_________30470),
       .Q (_____0___30459));
  nor2s1 ____9__439649(.DIN1 (_____0___30458), .DIN2 (_____0___30457),
       .Q (_________30521));
  xor2s1 _____0_439650(.DIN1 (_________________0___18618), .DIN2
       (_________34670), .Q (_________30621));
  nnd2s1 _______439651(.DIN1 (_________31519), .DIN2 (_____09__30464),
       .Q (_________30515));
  nnd2s1 _____9_439652(.DIN1 (_____0___30457), .DIN2 (_____00__30456),
       .Q (_________30499));
  xor2s1 _____0_439653(.DIN1 (______0__30409), .DIN2 (________22956),
       .Q (_________30498));
  nnd2s1 _______439654(.DIN1 (_________30420), .DIN2 (______0__30291),
       .Q (_________30527));
  nor2s1 _______439655(.DIN1 (_____9___30454), .DIN2 (_________30414),
       .Q (_____99__30455));
  nnd2s1 ______439656(.DIN1 (_________30415), .DIN2 (_________31303),
       .Q (_____9___30453));
  nor2s1 _____0_439657(.DIN1 (_____9___34419), .DIN2 (_____99__30363),
       .Q (_____9___30452));
  nor2s1 _______439658(.DIN1 (_________________18698), .DIN2
       (_____90__30447), .Q (_____9___30451));
  nnd2s1 _______439659(.DIN1 (______9__32514), .DIN2 (_____9___30449),
       .Q (_____9___30450));
  or2s1 _______439660(.DIN1 (_____09__30554), .DIN2 (_____90__30447),
       .Q (_____9___30448));
  nor2s1 _______439661(.DIN1 (___09____28076), .DIN2 (______9__32514),
       .Q (______9__30446));
  nnd2s1 _______439662(.DIN1 (______9__30417), .DIN2 (_________30229),
       .Q (_________30445));
  nor2s1 _______439663(.DIN1 (_____0__19096), .DIN2 (_________30413),
       .Q (_________30502));
  nor2s1 _______439664(.DIN1 (_________30444), .DIN2 (_________30473),
       .Q (_________30468));
  and2s1 _______439665(.DIN1 (_________30473), .DIN2 (_________30444),
       .Q (______0__30500));
  hi1s1 _____9_439666(.DIN (_________30470), .Q (____0____33715));
  or2s1 ______439667(.DIN1 (_________30442), .DIN2 (_________30430), .Q
       (_________30443));
  nnd2s1 _______439668(.DIN1 (______0__28955), .DIN2 (______9__34480),
       .Q (_________30441));
  nnd2s1 _______439669(.DIN1 (_________30439), .DIN2
       (______________0___________________9), .Q (_________30440));
  or2s1 _______439670(.DIN1 (______________0___________________9),
       .DIN2 (_________30439), .Q (_________30438));
  nnd2s1 _______439671(.DIN1 (_________30439), .DIN2 (_____09__34430),
       .Q (______0__30437));
  nor2s1 _______439672(.DIN1 (_____09__34430), .DIN2 (_________30439),
       .Q (______9__30436));
  nnd2s1 _______439673(.DIN1 (______9__30408), .DIN2 (________21041),
       .Q (_________30435));
  nnd2s1 ______439674(.DIN1 (_________30407), .DIN2 (_____0__19272), .Q
       (_________30434));
  nor2s1 _____9_439675(.DIN1 (_________30496), .DIN2 (_________30411),
       .Q (_________30433));
  nor2s1 _______439676(.DIN1 (_________30431), .DIN2 (_________30430),
       .Q (_________30432));
  nor2s1 ____9__439677(.DIN1 (_________34409), .DIN2 (_________30429),
       .Q (______0__30520));
  nnd2s1 _____9_439678(.DIN1 (_________30429), .DIN2
       (______________________________________0_____________18885), .Q
       (_________30516));
  xor2s1 ____9__439679(.DIN1 (_________30396), .DIN2 (_________30428),
       .Q (_____0___30460));
  xor2s1 _______439680(.DIN1 (_________30394), .DIN2 (_____0___33866),
       .Q (______9__30493));
  nor2s1 _____0_439681(.DIN1 (_________30402), .DIN2 (________25006),
       .Q (______0__30427));
  xor2s1 ______439682(.DIN1 (______0__30382), .DIN2 (_________34674),
       .Q (______9__30426));
  xor2s1 ______439683(.DIN1 (_________30416), .DIN2
       (______________________________________0_____________18886), .Q
       (_________30425));
  nnd2s1 _______439684(.DIN1 (_________30404), .DIN2 (____09___30085),
       .Q (_________30487));
  xor2s1 _______439685(.DIN1 (_________30385), .DIN2 (_________31431),
       .Q (_________30481));
  nor2s1 _____0_439686(.DIN1 (_____9___30359), .DIN2 (______9__30398),
       .Q (_________30478));
  xor2s1 ______439687(.DIN1 (_____0__23850), .DIN2 (_________30412), .Q
       (_________30470));
  dffacs1 __________________439688(.CLRB (reset), .CLK (clk), .DIN
       (_________30401), .Q (________________18721));
  hi1s1 _____9_439689(.DIN (_____90__30447), .Q (_________30507));
  nnd2s1 _______439690(.DIN1 (_________30397), .DIN2 (________21752),
       .Q (_________30424));
  nnd2s1 ______439691(.DIN1 (____9____29975), .DIN2 (_________30390),
       .Q (_________30423));
  nnd2s1 ______439692(.DIN1 (_________30395), .DIN2 (_____9___30173),
       .Q (_________30422));
  nnd2s1 ____9_439693(.DIN1 (_________30419), .DIN2 (________21041), .Q
       (_________30421));
  nor2s1 _______439694(.DIN1 (_____00__30274), .DIN2 (______0__30391),
       .Q (_________30420));
  hi1s1 ____9__439695(.DIN (_________30429), .Q (_____0___30457));
  or2s1 ____9__439696(.DIN1 (________21041), .DIN2 (_________30419), .Q
       (_____0___30462));
  nor2s1 _______439697(.DIN1 (________24164), .DIN2 (_________30393),
       .Q (_________30805));
  xor2s1 ____9__439698(.DIN1 (______0__30418), .DIN2 (_________30410),
       .Q (_________31519));
  dffacs1 ______________0____439699(.CLRB (reset), .CLK (clk), .DIN
       (_________30386), .Q (_____9___34419));
  or2s1 _____9_439700(.DIN1 (_________30228), .DIN2 (_________30416),
       .Q (______9__30417));
  nor2s1 _____0_439701(.DIN1 (________23721), .DIN2 (______9__30381),
       .Q (_________30415));
  xor2s1 ______439702(.DIN1 (_________30114), .DIN2 (_________30403),
       .Q (_________30414));
  and2s1 _______439703(.DIN1 (_________30412), .DIN2 (________19127),
       .Q (_________30413));
  xor2s1 _____439704(.DIN1 (_____0___30365), .DIN2
       (_______________18881), .Q (_____90__30447));
  xor2s1 ______439705(.DIN1 (____0____34545), .DIN2 (_____00__30545),
       .Q (_________30473));
  xor2s1 _____0_439706(.DIN1 (_____0___30370), .DIN2 (_________30338),
       .Q (______9__32514));
  nnd2s1 ____9__439707(.DIN1 (_________30410), .DIN2 (______0__30418),
       .Q (_________30411));
  xor2s1 _______439708(.DIN1 (________24165), .DIN2 (_________33937),
       .Q (______0__30409));
  xor2s1 ____90_439709(.DIN1 (____0____30930), .DIN2 (_________30388),
       .Q (______9__30408));
  or2s1 ____9_439710(.DIN1 (___9___19032), .DIN2 (_________30410), .Q
       (_________30407));
  and2s1 _______439711(.DIN1 (_________30376), .DIN2
       (______________0___________________), .Q (_________30430));
  dffacs1 __________________439712(.CLRB (reset), .CLK (clk), .DIN
       (_________30375), .QN (______9__34480));
  xor2s1 ____9__439713(.DIN1 (_____9___30356), .DIN2 (_________33835),
       .Q (_________30429));
  xor2s1 ____9__439714(.DIN1 (______9__30290), .DIN2 (_________34672),
       .Q (_________30439));
  nnd2s1 _______439715(.DIN1 (_________30383), .DIN2 (_________30405),
       .Q (_________30406));
  nnd2s1 ______439716(.DIN1 (_________30403), .DIN2 (____0_9__30083),
       .Q (_________30404));
  nor2s1 _______439717(.DIN1 (_____9___30362), .DIN2 (________24931),
       .Q (_________30402));
  nnd2s1 _______439718(.DIN1 (____9_0__29920), .DIN2 (_____0___30367),
       .Q (_________30401));
  nnd2s1 _______439719(.DIN1 (______0__30399), .DIN2 (____0____30020),
       .Q (_________30400));
  and2s1 _______439720(.DIN1 (_____9___30361), .DIN2 (_________34674),
       .Q (______9__30398));
  nnd2s1 _______439721(.DIN1 (_____90__30354), .DIN2 (__99____27118),
       .Q (_________30397));
  dffacs1 _______________439722(.CLRB (reset), .CLK (clk), .DIN
       (_____00__30364), .QN (outData[5]));
  nnd2s1 ____9__439723(.DIN1 (_________30348), .DIN2 (_____9___30355),
       .Q (_________30396));
  nor2s1 _______439724(.DIN1 (_________30351), .DIN2 (____90___29909),
       .Q (_________30395));
  nor2s1 _____9_439725(.DIN1 (______9__30254), .DIN2 (_________30350),
       .Q (_________30394));
  and2s1 ____90_439726(.DIN1 (_________33937), .DIN2 (________24166),
       .Q (_________30393));
  xor2s1 ____9__439727(.DIN1 (______0__34431), .DIN2 (_________30379),
       .Q (_________30392));
  nor2s1 ____9__439728(.DIN1 (______0__30237), .DIN2 (_________34672),
       .Q (______0__30391));
  nnd2s1 _______439729(.DIN1 (_________30349), .DIN2 (inData[4]), .Q
       (_________30390));
  nor2s1 ____9__439730(.DIN1 (_________30388), .DIN2 (____0____30930),
       .Q (_________30389));
  nnd2s1 ____9__439731(.DIN1 (____0____30930), .DIN2 (_________30388),
       .Q (_________30419));
  xor2s1 _______439732(.DIN1 (_____________18905), .DIN2
       (________________18723), .Q (_________30387));
  nnd2s1 _______439733(.DIN1 (_________30342), .DIN2 (_________34393),
       .Q (_________30386));
  nor2s1 ______439734(.DIN1 (_________30155), .DIN2 (_________30343),
       .Q (_________30385));
  hi1s1 _____439735(.DIN (_________30383), .Q (_________30384));
  xor2s1 _______439736(.DIN1 (____________9___18692), .DIN2
       (_____0___33031), .Q (______0__30382));
  nor2s1 _______439737(.DIN1 (_____9___30454), .DIN2 (_________30333),
       .Q (______9__30381));
  nnd2s1 ______439738(.DIN1 (_________30340), .DIN2 (_____0___30369),
       .Q (_________30416));
  nnd2s1 _______439739(.DIN1 (_________30331), .DIN2 (__9_____26746),
       .Q (_________30412));
  xor2s1 _______439740(.DIN1 (_________30322), .DIN2 (_________30115),
       .Q (_________33159));
  nor2s1 ____9__439741(.DIN1 (______0__34431), .DIN2 (_________30379),
       .Q (_________30380));
  nnd2s1 ____90_439742(.DIN1 (_________30377), .DIN2 (_________28789),
       .Q (_________30378));
  xor2s1 ____439743(.DIN1 (_________30323), .DIN2 (______0__30607), .Q
       (_________30376));
  or2s1 ______439744(.DIN1 (_________30374), .DIN2 (_________30325), .Q
       (_________30375));
  and2s1 ____9__439745(.DIN1 (_________30379), .DIN2 (______0__34431),
       .Q (______0__30373));
  nnd2s1 _______439746(.DIN1 (_________30346), .DIN2 (_____0___30371),
       .Q (_____09__30372));
  nor2s1 ____9_439747(.DIN1 (______________0___________________), .DIN2
       (_________30379), .Q (_________30442));
  nor2s1 ____9__439748(.DIN1 (________20559), .DIN2 (_________30329),
       .Q (_________30410));
  and2s1 _______439749(.DIN1 (_________30339), .DIN2 (_____0___30369),
       .Q (_____0___30370));
  xor2s1 _______439750(.DIN1 (____0____31844), .DIN2 (_________30319),
       .Q (_____0___30368));
  or2s1 _____9_439751(.DIN1 (________________18723), .DIN2
       (_____0___32299), .Q (_____0___30367));
  xor2s1 ______439752(.DIN1 (_____________0___18697), .DIN2
       (_________30319), .Q (_____0___30366));
  xnr2s1 _______439753(.DIN1 (_________31281), .DIN2 (_________30330),
       .Q (_____0___30365));
  or2s1 _______439754(.DIN1 (_________34503), .DIN2 (_____99__30363),
       .Q (_____00__30364));
  or2s1 _______439755(.DIN1 (________________18723), .DIN2
       (_____9__23142), .Q (_____9___30362));
  nnd2s1 _______439756(.DIN1 (_____9___30360), .DIN2
       (____________9___18692), .Q (_____9___30361));
  nor2s1 _______439757(.DIN1 (____________9___18692), .DIN2
       (_____9___30360), .Q (_____9___30359));
  or2s1 _____0_439758(.DIN1 (________________18723), .DIN2
       (_____9___30358), .Q (_________30405));
  nnd2s1 _____439759(.DIN1 (_____9___30358), .DIN2
       (________________18723), .Q (_________30383));
  nor2s1 _______439760(.DIN1 (_________30224), .DIN2 (_________30321),
       .Q (_________30403));
  xor2s1 _______439761(.DIN1 (________23323), .DIN2 (_________30319),
       .Q (_____9___30357));
  and2s1 ____0_439762(.DIN1 (_________30347), .DIN2 (_____9___30355),
       .Q (_____9___30356));
  xor2s1 ____90_439763(.DIN1 (_________30310), .DIN2 (_________31479),
       .Q (_____90__30354));
  nnd2s1 ____90_439764(.DIN1 (_________30324), .DIN2 (_________30352),
       .Q (______9__30353));
  and2s1 ____9_439765(.DIN1 (____0____30080), .DIN2 (_________30315),
       .Q (_________30351));
  nnd2s1 ____9__439766(.DIN1 (______0__30318), .DIN2 (_________30249),
       .Q (_________30350));
  nor2s1 ____9__439767(.DIN1 (_________30316), .DIN2 (_________29858),
       .Q (_________30349));
  nnd2s1 ____99_439768(.DIN1 (_________30347), .DIN2 (_________33835),
       .Q (_________30348));
  hi1s1 ____90_439769(.DIN (_________30346), .Q (______0__30399));
  xor2s1 ____9__439770(.DIN1 (______9__30317), .DIN2 (_________30307),
       .Q (_________33937));
  xor2s1 ____99_439771(.DIN1 (_________30328), .DIN2 (______0__30345),
       .Q (____0____30930));
  and2s1 _______439772(.DIN1 (_________30319), .DIN2
       (_____________0___18697), .Q (______9__30344));
  nnd2s1 _______439773(.DIN1 (_________30312), .DIN2 (_________30165),
       .Q (_________30343));
  xor2s1 ______439774(.DIN1 (_________30302), .DIN2 (_________30341),
       .Q (_________30342));
  nnd2s1 _______439775(.DIN1 (_________30339), .DIN2 (_________30338),
       .Q (_________30340));
  and2s1 ______439776(.DIN1 (_________30319), .DIN2 (_________34442),
       .Q (_________30337));
  nor2s1 _______439777(.DIN1 (_____________0___18779), .DIN2
       (_________30319), .Q (_________30336));
  and2s1 _______439778(.DIN1 (_________30319), .DIN2
       (_____________0___18779), .Q (______0__30335));
  nor2s1 _______439779(.DIN1 (_____________0___18697), .DIN2
       (_________30319), .Q (______9__30334));
  xor2s1 _____439780(.DIN1 (_________30320), .DIN2 (_________30225), .Q
       (_________30333));
  dffacs1 __________________439781(.CLRB (reset), .CLK (clk), .DIN
       (_________30313), .QN (________________18722));
  nor2s1 _______439782(.DIN1 (_________34442), .DIN2 (_________30319),
       .Q (_________30332));
  nnd2s1 _____439783(.DIN1 (_________30330), .DIN2 (__9_____26681), .Q
       (_________30331));
  nor2s1 ____99_439784(.DIN1 (____0___19406), .DIN2 (_________30328),
       .Q (_________30329));
  xor2s1 ____9__439785(.DIN1 (_________30292), .DIN2 (_____0___31184),
       .Q (______9__30326));
  xor2s1 ____9_439786(.DIN1 (________________18691), .DIN2
       (_________30294), .Q (_________30325));
  hi1s1 ____9__439787(.DIN (_________30324), .Q (_________30377));
  xor2s1 ____9__439788(.DIN1 (_________30304), .DIN2 (____0____32777),
       .Q (_________30346));
  hi1s1 ____9__439789(.DIN (_________30323), .Q (_________30379));
  dffacs1 ______________0____439790(.CLRB (reset), .CLK (clk), .DIN
       (_________30303), .Q (_________34503));
  xor2s1 _______439791(.DIN1 (_________30311), .DIN2 (_____0___30999),
       .Q (_________30322));
  and2s1 _______439792(.DIN1 (_________30320), .DIN2 (_____0___30179),
       .Q (_________30321));
  nnd2s1 _____9_439793(.DIN1 (_________30300), .DIN2 (_________31388),
       .Q (_____0___30369));
  dffacs1 ________________9_439794(.CLRB (reset), .CLK (clk), .DIN
       (_________30301), .QN (____________9___18692));
  dffacs1 __________________439795(.CLRB (reset), .CLK (clk), .DIN
       (_________30305), .QN (________________18723));
  nnd2s1 ____9__439796(.DIN1 (______9__30317), .DIN2 (_________30119),
       .Q (______0__30318));
  xnr2s1 ____9_439797(.DIN1 (_________34493), .DIN2 (_____0___30280),
       .Q (_________30316));
  nnd2s1 ____9__439798(.DIN1 (_________30295), .DIN2 (inData[24]), .Q
       (_________30315));
  nor2s1 ____9_439799(.DIN1 (_____9___30265), .DIN2 (_________30296),
       .Q (_________30613));
  xor2s1 ____99_439800(.DIN1 (_____0___30281), .DIN2 (_________30338),
       .Q (_________30323));
  or2s1 ____0_439801(.DIN1 (_____9___30627), .DIN2 (_________30314), .Q
       (_____9___30355));
  nnd2s1 ____0__439802(.DIN1 (_________30314), .DIN2 (_____9___30627),
       .Q (_________30347));
  xor2s1 ____9_439803(.DIN1 (_____0___30276), .DIN2 (_____9___30268),
       .Q (_________30324));
  nnd2s1 _______439804(.DIN1 (_________30287), .DIN2 (____0___23975),
       .Q (_________30313));
  nnd2s1 ______439805(.DIN1 (_________30311), .DIN2 (_________30110),
       .Q (_________30312));
  nor2s1 ____9_439806(.DIN1 (________25897), .DIN2 (_________30288), .Q
       (_________30330));
  nor2s1 ____9__439807(.DIN1 (_________30158), .DIN2 (_________30286),
       .Q (_____9___33482));
  nnd2s1 _____9_439808(.DIN1 (______0__30299), .DIN2
       (_______________18880), .Q (_________30339));
  xor2s1 ____9_439809(.DIN1 (_________30256), .DIN2 (_________30262),
       .Q (_________30310));
  xor2s1 ____9__439810(.DIN1 (_________30260), .DIN2 (______0__35008),
       .Q (______0__30309));
  xor2s1 ____9__439811(.DIN1 (_________30257), .DIN2
       (_________________0___18618), .Q (______9__30308));
  nor2s1 ____0__439812(.DIN1 (_____0___30275), .DIN2 (_________30233),
       .Q (_________30307));
  nor2s1 ____0_439813(.DIN1 (________19290), .DIN2 (_____99__30273), .Q
       (_________30328));
  nnd2s1 ____9_439814(.DIN1 (_________30284), .DIN2 (_________30231),
       .Q (______0__30327));
  hi1s1 ____9__439815(.DIN (_________30306), .Q (_________30319));
  or2s1 _______439816(.DIN1 (________19627), .DIN2 (_____9___30271), .Q
       (_________30305));
  xor2s1 ____9__439817(.DIN1 (_________30213), .DIN2 (_________30232),
       .Q (_________30304));
  nnd2s1 _____9_439818(.DIN1 (_____9___30267), .DIN2 (_________34365),
       .Q (_________30303));
  xor2s1 ____9__439819(.DIN1 (_________30160), .DIN2 (_________30285),
       .Q (_________30302));
  nor2s1 ____9__439820(.DIN1 (_________30374), .DIN2 (_____90__30264),
       .Q (_________30301));
  hi1s1 ____9__439821(.DIN (______0__30299), .Q (_________30300));
  hi1s1 ____9__439822(.DIN (_________30297), .Q (______9__30298));
  xor2s1 ____9__439823(.DIN1 (_________30244), .DIN2 (_________31326),
       .Q (_________30306));
  xor2s1 _______439824(.DIN1 (______9__30245), .DIN2 (_____9___32930),
       .Q (_________30320));
  nor2s1 ____00_439825(.DIN1 (_____9___30269), .DIN2 (_________32946),
       .Q (_________30296));
  xor2s1 ____00_439826(.DIN1 (_____0___30279), .DIN2 (_______19029), .Q
       (_________30295));
  nor2s1 ____439827(.DIN1 (_____0___30278), .DIN2 (_________30293), .Q
       (_________30294));
  nor2s1 ____0__439828(.DIN1 (_________30250), .DIN2 (_________30251),
       .Q (_________30292));
  nnd2s1 ____0__439829(.DIN1 (______9__30290), .DIN2 (_________33925),
       .Q (______0__30291));
  nor2s1 ____0__439830(.DIN1 (_________30211), .DIN2 (_________30258),
       .Q (_________30314));
  nnd2s1 ____0__439831(.DIN1 (_____9___30270), .DIN2 (_________30259),
       .Q (______9__30317));
  nnd2s1 ____00_439832(.DIN1 (_________30263), .DIN2 (_________30234),
       .Q (_________30431));
  xor2s1 ____0__439833(.DIN1 (_____9___30272), .DIN2 (________19960),
       .Q (____9____30847));
  xor2s1 ____9_439834(.DIN1 (_________30218), .DIN2 (____0____31863),
       .Q (_________30288));
  nnd2s1 ______439835(.DIN1 (_________30243), .DIN2 (_________31241),
       .Q (_________30287));
  nor2s1 ____9__439836(.DIN1 (_________30285), .DIN2 (_________30159),
       .Q (_________30286));
  xor2s1 ____00_439837(.DIN1 (_________30212), .DIN2 (______0__30283),
       .Q (_________30284));
  nnd2s1 _____439838(.DIN1 (_________30241), .DIN2 (____9____29955), .Q
       (_________30311));
  xor2s1 ____9__439839(.DIN1 (_________30219), .DIN2 (_____0___31005),
       .Q (______0__30299));
  xor2s1 ____9__439840(.DIN1 (______0__30227), .DIN2 (_________30220),
       .Q (_________30297));
  hi1s1 ____9__439841(.DIN (_____09__30282), .Q (_____9___32565));
  xor2s1 ____0__439842(.DIN1 (______0__34678), .DIN2
       (_______________18875), .Q (_____0___30281));
  nor2s1 ____0__439843(.DIN1 (______________0___________________0),
       .DIN2 (_____0___30279), .Q (_____0___30280));
  xor2s1 ____0__439844(.DIN1 (_________30772), .DIN2 (_________31154),
       .Q (_____0___30277));
  xor2s1 ____0__439845(.DIN1 (______0__34481), .DIN2 (_________32946),
       .Q (_____0___30276));
  nor2s1 ____0__439846(.DIN1 (____90___28993), .DIN2 (_________30230),
       .Q (_____0___30275));
  nor2s1 ____0_439847(.DIN1 (_______________18876), .DIN2
       (_________30238), .Q (_____00__30274));
  nor2s1 ____0__439848(.DIN1 (________19289), .DIN2 (_____9___30272),
       .Q (_____99__30273));
  nor2s1 ____9__439849(.DIN1 (________19962), .DIN2 (_________30223),
       .Q (_____9___30271));
  xor2s1 ____0__439850(.DIN1 (_________30194), .DIN2 (____0____31831),
       .Q (_____9___30270));
  and2s1 ____0__439851(.DIN1 (_____9___30268), .DIN2 (______0__34481),
       .Q (_____9___30269));
  xor2s1 ____9__439852(.DIN1 (_________30202), .DIN2 (_________30150),
       .Q (_____9___30267));
  xor2s1 ____9__439853(.DIN1 (_________________18726), .DIN2
       (_________32538), .Q (_____9___30266));
  nor2s1 ____0__439854(.DIN1 (______0__34481), .DIN2 (_____9___30268),
       .Q (_____9___30265));
  xor2s1 ____9__439855(.DIN1 (______9__30197), .DIN2 (___0__18931), .Q
       (_____90__30264));
  nnd2s1 ____0__439856(.DIN1 (_________30262), .DIN2 (______9__30216),
       .Q (_________30263));
  xor2s1 ____9_439857(.DIN1 (_________30209), .DIN2 (____0_0__31861),
       .Q (_____09__30282));
  xor2s1 ____9_439858(.DIN1 (____9____29988), .DIN2 (_________34680),
       .Q (_________33234));
  and2s1 ____0_439859(.DIN1 (______0__30246), .DIN2 (_____9___32650),
       .Q (_________30293));
  hi1s1 ____9__439860(.DIN (_________30261), .Q (_________32490));
  nnd2s1 ____00_439861(.DIN1 (_________30222), .DIN2 (______9__30226),
       .Q (____0____31885));
  nnd2s1 ____0_439862(.DIN1 (_________30259), .DIN2 (_________30193),
       .Q (_________30260));
  and2s1 _______439863(.DIN1 (_________34676), .DIN2 (_________31134),
       .Q (_________30258));
  xor2s1 ____0__439864(.DIN1 (____0___21451), .DIN2 (______0__30255),
       .Q (_________30257));
  xor2s1 ____0__439865(.DIN1 (_________30215), .DIN2 (______0__30255),
       .Q (_________30256));
  nor2s1 _______439866(.DIN1 (_________30472), .DIN2 (_________30248),
       .Q (______9__30254));
  nnd2s1 ____09_439867(.DIN1 (_________30772), .DIN2 (______9__29521),
       .Q (_________30253));
  or2s1 ____09_439868(.DIN1 (______9__29465), .DIN2 (_________30772),
       .Q (_________30252));
  nor2s1 ____09_439869(.DIN1 (_________29471), .DIN2 (_________30772),
       .Q (_________30251));
  and2s1 ____09_439870(.DIN1 (_________30772), .DIN2 (_________29477),
       .Q (_________30250));
  nnd2s1 _______439871(.DIN1 (_________30248), .DIN2 (_________30472),
       .Q (_________30249));
  xor2s1 _____0_439872(.DIN1 (_________30247), .DIN2
       (_______________18876), .Q (______9__30290));
  nnd2s1 ____0__439873(.DIN1 (______0__34678), .DIN2 (____09___30087),
       .Q (_________30289));
  nor2s1 ____0__439874(.DIN1 (_____9___32650), .DIN2 (______0__30246),
       .Q (_____0___30278));
  nnd2s1 ____9__439875(.DIN1 (_________30204), .DIN2 (____0____30061),
       .Q (______9__30245));
  xor2s1 ____0__439876(.DIN1 (______0__30217), .DIN2 (________25898),
       .Q (_________30244));
  xor2s1 ____9__439877(.DIN1 (_____09__30187), .DIN2 (____0____30050),
       .Q (_________30243));
  xor2s1 ____9_439878(.DIN1 (_________33093), .DIN2 (______0__30283),
       .Q (_________30242));
  nnd2s1 ____9__439879(.DIN1 (_________34680), .DIN2 (____9_9__29959),
       .Q (_________30241));
  and2s1 ____9__439880(.DIN1 (_________32538), .DIN2
       (_________________18726), .Q (_________30240));
  or2s1 ____9__439881(.DIN1 (_________________18726), .DIN2
       (_________32538), .Q (_________30239));
  nor2s1 ____9__439882(.DIN1 (_________30201), .DIN2 (_________30206),
       .Q (_________30285));
  xor2s1 ____9__439883(.DIN1 (_____0___30185), .DIN2 (___0_9___27843),
       .Q (_________30261));
  dffacs1 __________________439884(.CLRB (reset), .CLK (clk), .DIN
       (______0__30208), .QN (_________34434));
  dffacs1 _______________439885(.CLRB (reset), .CLK (clk), .DIN
       (_________30205), .QN (outData[4]));
  or2s1 _______439886(.DIN1 (_________33925), .DIN2 (_________30247),
       .Q (_________30238));
  and2s1 _______439887(.DIN1 (_________30247), .DIN2
       (_______________18876), .Q (______0__30237));
  nor2s1 ____0__439888(.DIN1 (_________18847), .DIN2 (______0__30255),
       .Q (______9__30236));
  and2s1 ____0_439889(.DIN1 (______0__30255), .DIN2 (_________18847),
       .Q (_________30235));
  nnd2s1 ____0__439890(.DIN1 (______0__30255), .DIN2
       (_____________0___18679), .Q (_________30234));
  nor2s1 _______439891(.DIN1 (_________30472), .DIN2 (_________30210),
       .Q (_________30233));
  xnr2s1 ____0_439892(.DIN1 (_________30231), .DIN2 (_____0___33872),
       .Q (_________30232));
  nor2s1 _______439893(.DIN1 (______0__30112), .DIN2 (_________30191),
       .Q (_________30230));
  nnd2s1 _______439894(.DIN1 (_________30247), .DIN2
       (______________________________________0_____________18886), .Q
       (_________30229));
  nor2s1 ______439895(.DIN1
       (______________________________________0_____________18886),
       .DIN2 (_________30247), .Q (_________30228));
  nor2s1 _______439896(.DIN1 (____9___19106), .DIN2 (_________30199),
       .Q (_____9___30272));
  hi1s1 ____0__439897(.DIN (______0__34481), .Q (_____0___30279));
  nnd2s1 ____0__439898(.DIN1 (_________30221), .DIN2 (______9__30226),
       .Q (______0__30227));
  nor2s1 ____439899(.DIN1 (_________30224), .DIN2 (_____0___30180), .Q
       (_________30225));
  xor2s1 ____9_439900(.DIN1 (_____0___30096), .DIN2 (_________30203),
       .Q (_________30223));
  nnd2s1 ____0__439901(.DIN1 (_________30221), .DIN2 (_________30220),
       .Q (_________30222));
  nor2s1 ____439902(.DIN1 (____0____30039), .DIN2 (_____0___30182), .Q
       (_________30219));
  or2s1 ____0__439903(.DIN1 (________25896), .DIN2 (______0__30217), .Q
       (_________30218));
  nnd2s1 ____0__439904(.DIN1 (_________30189), .DIN2 (_________30215),
       .Q (______9__30216));
  dffacs1 __________________439905(.CLRB (reset), .CLK (clk), .DIN
       (_____0___30183), .QN (________________18691));
  dffacs1 __________________439906(.CLRB (reset), .CLK (clk), .DIN
       (_____9___30174), .Q (______0__34481));
  or2s1 ____09_439907(.DIN1 (_________30213), .DIN2 (_____0___33872),
       .Q (_________30214));
  and2s1 _____439908(.DIN1 (_____0___33872), .DIN2 (_________30213), .Q
       (_________30212));
  nor2s1 _______439909(.DIN1 (_________31134), .DIN2 (_____9___30177),
       .Q (_________30211));
  xor2s1 ____09_439910(.DIN1 (_________30157), .DIN2 (____0____31872),
       .Q (_________30259));
  hi1s1 ______439911(.DIN (_________30210), .Q (_________30248));
  xnr2s1 _____0_439912(.DIN1 (______0__29851), .DIN2 (_________34682),
       .Q (______0__30246));
  xor2s1 _______439913(.DIN1 (______0__30198), .DIN2 (________19964),
       .Q (_________30772));
  nor2s1 ____00_439914(.DIN1 (___0_____27838), .DIN2 (_________30168),
       .Q (_________30209));
  or2s1 ____0_439915(.DIN1 (______9__30207), .DIN2 (_____9___30172), .Q
       (______0__30208));
  nor2s1 ____99_439916(.DIN1 (_________30149), .DIN2 (_________30200),
       .Q (_________30206));
  or2s1 ____99_439917(.DIN1 (_________34502), .DIN2 (_____99__30363),
       .Q (_________30205));
  nnd2s1 ____9__439918(.DIN1 (_________30203), .DIN2 (____0____30069),
       .Q (_________30204));
  or2s1 ____0__439919(.DIN1 (_________30201), .DIN2 (_________30200),
       .Q (_________30202));
  xor2s1 ____0__439920(.DIN1 (____0____30041), .DIN2 (_____0___30181),
       .Q (_________32538));
  and2s1 _______439921(.DIN1 (______0__30198), .DIN2 (________19432),
       .Q (_________30199));
  xor2s1 ____0__439922(.DIN1 (_________30138), .DIN2 (_____0___33222),
       .Q (______9__30197));
  nnd2s1 ____0__439923(.DIN1 (_________30164), .DIN2 (_________30195),
       .Q (_________30196));
  nnd2s1 _______439924(.DIN1 (_________30141), .DIN2 (_________30193),
       .Q (_________30194));
  xor2s1 ____0__439925(.DIN1 (____99__21445), .DIN2 (_________33206),
       .Q (_________30192));
  nor2s1 _______439926(.DIN1 (______9__30111), .DIN2 (_________30190),
       .Q (_________30191));
  nnd2s1 _____9_439927(.DIN1 (_________30190), .DIN2 (_________30118),
       .Q (_________30210));
  hi1s1 _______439928(.DIN (_________30189), .Q (______0__30255));
  xor2s1 _____439929(.DIN1 (_____9___30176), .DIN2 (_____9___30175), .Q
       (_________30247));
  nor2s1 ____0__439930(.DIN1 (_________34489), .DIN2 (_________33206),
       .Q (______0__30188));
  xor2s1 ____9__439931(.DIN1 (_________30130), .DIN2 (______0__35098),
       .Q (_____09__30187));
  xor2s1 ____0__439932(.DIN1 (_________34463), .DIN2 (_____0___30184),
       .Q (_____0___30186));
  xor2s1 ____0__439933(.DIN1 (_________________18744), .DIN2
       (_____0___30184), .Q (_____0___30185));
  nor2s1 ____0__439934(.DIN1 (_________30374), .DIN2 (______0__30143),
       .Q (_____0___30183));
  nor2s1 ____0__439935(.DIN1 (____0____30040), .DIN2 (_____0___30181),
       .Q (_____0___30182));
  hi1s1 ____0__439936(.DIN (_____0___30179), .Q (_____0___30180));
  nnd2s1 ____0__439937(.DIN1 (_________33206), .DIN2 (_________34489),
       .Q (_____00__30178));
  xor2s1 ____439938(.DIN1 (____0____34546), .DIN2 (____0_9__30073), .Q
       (_________33093));
  nnd2s1 ______439939(.DIN1 (_____9___30176), .DIN2 (_____9___30175),
       .Q (_____9___30177));
  nnd2s1 ______439940(.DIN1 (_________30140), .DIN2 (_____9___30173),
       .Q (_____9___30174));
  nnd2s1 ____0_439941(.DIN1 (_________33206), .DIN2
       (_____________0___18715), .Q (_________30221));
  or2s1 ____0__439942(.DIN1 (_____________0___18715), .DIN2
       (_________33206), .Q (______9__30226));
  xor2s1 ______439943(.DIN1 (_________30105), .DIN2 (____99___29996),
       .Q (_________30189));
  nnd2s1 ____0__439944(.DIN1 (_________30144), .DIN2 (______0__30136),
       .Q (_________30262));
  nnd2s1 _____0_439945(.DIN1 (______9__30142), .DIN2 (________25932),
       .Q (______0__30217));
  xor2s1 _______439946(.DIN1 (_________30108), .DIN2 (____9____29971),
       .Q (_____0___33872));
  dffacs1 ______________0____439947(.CLRB (reset), .CLK (clk), .DIN
       (_________30128), .Q (_________34502));
  nnd2s1 ____0__439948(.DIN1 (_________30124), .DIN2 (_____0__23009),
       .Q (_____9___30172));
  nor2s1 ____0__439949(.DIN1 (______9__30169), .DIN2 (_____0___30184),
       .Q (_____9___30171));
  nnd2s1 ____0__439950(.DIN1 (_____0___30184), .DIN2 (______9__30169),
       .Q (_____90__30170));
  nor2s1 ____0_439951(.DIN1 (___0_9___27844), .DIN2 (_____0___30184),
       .Q (_________30168));
  nnd2s1 ____0__439952(.DIN1 (______9__30161), .DIN2 (______0__35078),
       .Q (_________30167));
  xor2s1 ____0__439953(.DIN1 (_____0___30095), .DIN2
       (_________________0___18607), .Q (_____0___30179));
  xor2s1 ____0__439954(.DIN1 (_____0___30101), .DIN2
       (_________________0___18618), .Q (_________30200));
  xor2s1 ____0__439955(.DIN1 (_____0___30099), .DIN2 (_________30166),
       .Q (_________30201));
  nor2s1 ____0__439956(.DIN1 (_________30129), .DIN2 (_________30132),
       .Q (_________30203));
  nnd2s1 _______439957(.DIN1 (_________30154), .DIN2 (_________33895),
       .Q (_________30165));
  hi1s1 ____0__439958(.DIN (_________30163), .Q (_________30164));
  nor2s1 ____09_439959(.DIN1 (______0__35078), .DIN2 (______9__30161),
       .Q (______0__30162));
  or2s1 ____09_439960(.DIN1 (_________30159), .DIN2 (_________30158),
       .Q (_________30160));
  and2s1 _____9_439961(.DIN1 (_________30156), .DIN2 (_____9___29263),
       .Q (_________30157));
  nor2s1 _______439962(.DIN1 (_________33895), .DIN2 (_________30154),
       .Q (_________30155));
  nor2s1 ____0_439963(.DIN1 (_________30133), .DIN2 (______0__30152),
       .Q (_________30153));
  xor2s1 ______439964(.DIN1 (____09___30089), .DIN2 (____90___33582),
       .Q (______0__30198));
  xor2s1 _____0_439965(.DIN1 (____09___30088), .DIN2 (_________30595),
       .Q (____90___31729));
  xor2s1 _____439966(.DIN1 (____0____30078), .DIN2 (_________31486), .Q
       (_________30193));
  hi1s1 _______439967(.DIN (_________30151), .Q (_________30190));
  xor2s1 _____0_439968(.DIN1 (_________30149), .DIN2 (________19986),
       .Q (_________30150));
  or2s1 ____0_439969(.DIN1 (_________30147), .DIN2 (_________30146), .Q
       (_________30148));
  nnd2s1 ____439970(.DIN1 (_________30146), .DIN2 (_________30147), .Q
       (_________30145));
  nnd2s1 _______439971(.DIN1 (_________30137), .DIN2 (_____0___33222),
       .Q (_________30144));
  xor2s1 ____0__439972(.DIN1 (____0____30059), .DIN2 (____0____32762),
       .Q (______0__30143));
  nor2s1 ______439973(.DIN1 (________25935), .DIN2 (_____0___30097), .Q
       (______9__30142));
  nnd2s1 _____0_439974(.DIN1 (_____00__30094), .DIN2 (____99___29993),
       .Q (_____0___30181));
  xor2s1 ____439975(.DIN1 (____0____30065), .DIN2 (_____0___31005), .Q
       (_________30163));
  nor2s1 _______439976(.DIN1 (_____00__35028), .DIN2 (____0____30081),
       .Q (_________30140));
  and2s1 ______439977(.DIN1 (_________30137), .DIN2 (______0__30136),
       .Q (_________30138));
  xor2s1 _______439978(.DIN1 (_________30117), .DIN2
       (_________________0___18618), .Q (_________30151));
  xor2s1 _______439979(.DIN1 (____0____30060), .DIN2 (_________33007),
       .Q (_____9___30176));
  hi1s1 _______439980(.DIN (______9__30135), .Q (_________33206));
  hi1s1 _____439981(.DIN (_________30133), .Q (_________30134));
  xor2s1 ____0__439982(.DIN1 (____0____30052), .DIN2 (_________30131),
       .Q (_________30132));
  or2s1 ____0__439983(.DIN1 (____0____30051), .DIN2 (_________30129),
       .Q (_________30130));
  nnd2s1 ____0__439984(.DIN1 (____0____30066), .DIN2 (_________34365),
       .Q (_________30128));
  nor2s1 ____0__439985(.DIN1 (_________30126), .DIN2 (____0_0__30074),
       .Q (______9__30127));
  nnd2s1 ______439986(.DIN1 (____0____30062), .DIN2 (_________32925),
       .Q (_________30124));
  nor2s1 ______439987(.DIN1 (_________30122), .DIN2 (______0__30121),
       .Q (_________30123));
  nnd2s1 _______439988(.DIN1 (______0__30121), .DIN2 (_________30122),
       .Q (______9__30161));
  nor2s1 _______439989(.DIN1 (___9___18979), .DIN2 (______0__30121), .Q
       (______0__30152));
  xor2s1 _____0_439990(.DIN1 (____0_9__30046), .DIN2
       (_______________18879), .Q (_____0___30184));
  or2s1 _______439991(.DIN1 (_________30118), .DIN2 (_________30117),
       .Q (_________30119));
  xor2s1 _______439992(.DIN1 (________24041), .DIN2 (_____90__33117),
       .Q (_________30116));
  xor2s1 _______439993(.DIN1 (____0____30057), .DIN2 (_________30109),
       .Q (_________30115));
  xor2s1 ______439994(.DIN1 (_________28883), .DIN2 (____090__30084),
       .Q (_________30114));
  xor2s1 _______439995(.DIN1 (_____90__33117), .DIN2 (____0____30071),
       .Q (_________30113));
  and2s1 ______439996(.DIN1 (_________30117), .DIN2 (______9__30111),
       .Q (______0__30112));
  nnd2s1 ______439997(.DIN1 (______0__30103), .DIN2 (_________30109),
       .Q (_________30110));
  xor2s1 _______439998(.DIN1 (____0_9__30036), .DIN2 (____000__32751),
       .Q (_________30108));
  nnd2s1 _____0_439999(.DIN1 (_________30106), .DIN2 (____90__19196),
       .Q (_________30107));
  xor2s1 _______440000(.DIN1 (____0____30076), .DIN2 (_________30104),
       .Q (_________30105));
  nor2s1 _____9_440001(.DIN1 (_________30109), .DIN2 (______0__30103),
       .Q (_________30154));
  xnr2s1 ______440002(.DIN1 (____9____30882), .DIN2 (____0____30035),
       .Q (_________30141));
  xor2s1 _______440003(.DIN1 (_____09__30102), .DIN2 (_________33007),
       .Q (_________30156));
  xor2s1 _______440004(.DIN1 (____0____30049), .DIN2 (_________30496),
       .Q (_________30158));
  xor2s1 ______440005(.DIN1 (__9__9), .DIN2 (_________34684), .Q
       (______9__30135));
  nnd2s1 _______440006(.DIN1 (_____0___29182), .DIN2 (_____0___30098),
       .Q (_____0___30101));
  and2s1 _______440007(.DIN1 (_____90__33117), .DIN2 (_________18864),
       .Q (_____0___30100));
  nor2s1 _______440008(.DIN1 (_____0___30098), .DIN2 (_____0___29181),
       .Q (_____0___30099));
  and2s1 _______440009(.DIN1 (_________34684), .DIN2 (_____9__25938),
       .Q (_____0___30097));
  xor2s1 ______440010(.DIN1 (____0____30067), .DIN2 (____0____30068),
       .Q (_____0___30096));
  nnd2s1 _______440011(.DIN1 (____09___30091), .DIN2 (____09___30092),
       .Q (_____0___30095));
  xor2s1 _______440012(.DIN1 (____0_0__30028), .DIN2 (____099__30093),
       .Q (_____00__30094));
  nor2s1 _______440013(.DIN1 (____09___30092), .DIN2 (____09___30091),
       .Q (_________30224));
  nor2s1 _______440014(.DIN1 (_________34464), .DIN2 (____0_9__30063),
       .Q (_________30133));
  xor2s1 _______440015(.DIN1 (_________34478), .DIN2 (____0____30032),
       .Q (_________30146));
  dffacs1 __________________440016(.CLRB (reset), .CLK (clk), .DIN
       (____0____30033), .QN (________________18706));
  dffacs1 _______________440017(.CLRB (reset), .CLK (clk), .DIN
       (____0____30048), .QN (outData[3]));
  or2s1 ______440018(.DIN1 (_________18864), .DIN2 (_____90__33117), .Q
       (____09___30090));
  nnd2s1 _____0_440019(.DIN1 (____0____30038), .DIN2 (________19268),
       .Q (____09___30089));
  nor2s1 _______440020(.DIN1 (____0____30031), .DIN2 (____0_0__30047),
       .Q (____09___30088));
  nnd2s1 _____9_440021(.DIN1 (_________30338), .DIN2 (____09___30086),
       .Q (____09___30087));
  nnd2s1 _______440022(.DIN1 (____0____30082), .DIN2 (____090__30084),
       .Q (____09___30085));
  or2s1 _______440023(.DIN1 (____090__30084), .DIN2 (____0____30082),
       .Q (____0_9__30083));
  nor2s1 _____0_440024(.DIN1 (____0____30080), .DIN2 (____0____30042),
       .Q (____0____30081));
  nor2s1 _____9_440025(.DIN1 (____09___30086), .DIN2 (_________30338),
       .Q (____0____30079));
  or2s1 ______440026(.DIN1 (_________29307), .DIN2 (_____09__30102), .Q
       (____0____30078));
  or2s1 _______440027(.DIN1 (____________9_), .DIN2 (____0____30077),
       .Q (______0__30136));
  nnd2s1 _______440028(.DIN1 (____0____30077), .DIN2 (____________9_),
       .Q (_________30137));
  nnd2s1 ______440029(.DIN1 (____0____30076), .DIN2 (____99___29995),
       .Q (_________30139));
  xor2s1 _______440030(.DIN1 (____0____30022), .DIN2 (____0____30075),
       .Q (_____0___33222));
  nor2s1 ____0__440031(.DIN1 (____0_9__30073), .DIN2 (____0_0__30064),
       .Q (____0_0__30074));
  or2s1 _______440032(.DIN1 (____0____30071), .DIN2 (____0____30070),
       .Q (____0____30072));
  or2s1 _______440033(.DIN1 (____0____30068), .DIN2 (____0____30067),
       .Q (____0____30069));
  xor2s1 _______440034(.DIN1 (____0____30016), .DIN2 (____0____30029),
       .Q (____0____30066));
  nor2s1 ______440035(.DIN1 (_________________18777), .DIN2
       (____0____30070), .Q (____0____30065));
  nnd2s1 _______440036(.DIN1 (____0____30070), .DIN2
       (_________________18777), .Q (_________30195));
  nnd2s1 ____0__440037(.DIN1 (____0_0__30064), .DIN2 (____0_9__30073),
       .Q (_________30120));
  nnd2s1 _______440038(.DIN1 (____0____30030), .DIN2 (____9____29984),
       .Q (_________30149));
  xor2s1 _____0_440039(.DIN1 (____0____30014), .DIN2 (_________35002),
       .Q (_________30129));
  hi1s1 _______440040(.DIN (____0_9__30063), .Q (______0__30121));
  xor2s1 _______440041(.DIN1 (____009__30008), .DIN2 (____9____29981),
       .Q (____0____30062));
  nnd2s1 _______440042(.DIN1 (____0____30067), .DIN2 (____0____30068),
       .Q (____0____30061));
  nor2s1 _______440043(.DIN1 (__99____27112), .DIN2 (____0____30024),
       .Q (____0____30060));
  xor2s1 _____9_440044(.DIN1 (____00___30007), .DIN2 (____0_0__30009),
       .Q (____0____30059));
  hi1s1 _______440045(.DIN (____0____30057), .Q (______0__30103));
  nnd2s1 _____9_440046(.DIN1 (____0____30070), .DIN2 (____0____30071),
       .Q (_________30125));
  nor2s1 _______440047(.DIN1 (____0_0__30056), .DIN2 (____0____30026),
       .Q (_________30106));
  xor2s1 _______440048(.DIN1 (________22793), .DIN2 (____0_0__30037),
       .Q (_________30117));
  nor2s1 _______440049(.DIN1 (____0____30054), .DIN2 (____0____30053),
       .Q (____0_9__30055));
  or2s1 _______440050(.DIN1 (____0____30051), .DIN2 (____0____30050),
       .Q (____0____30052));
  nnd2s1 _______440051(.DIN1 (_________29415), .DIN2 (____0____30043),
       .Q (____0____30049));
  or2s1 _______440052(.DIN1 (_________34504), .DIN2 (_____99__30363),
       .Q (____0____30048));
  and2s1 _____0_440053(.DIN1 (____0____30012), .DIN2 (_________34478),
       .Q (____0_0__30047));
  xor2s1 _____9_440054(.DIN1 (____0____30021), .DIN2 (____0_9__30027),
       .Q (____0_9__30046));
  hi1s1 _______440055(.DIN (____0____30045), .Q (_________33070));
  xor2s1 _____440056(.DIN1 (_______________18878), .DIN2
       (____99___29992), .Q (____0_9__30063));
  xor2s1 _____9_440057(.DIN1 (____9_9__29979), .DIN2 (____0____30044),
       .Q (_____0___30098));
  xor2s1 _____9_440058(.DIN1 (____9____29978), .DIN2 (____9____29964),
       .Q (____09___30092));
  nor2s1 _______440059(.DIN1 (____0____30043), .DIN2 (_________29416),
       .Q (_________30159));
  xor2s1 _______440060(.DIN1 (____99___29991), .DIN2
       (_________________0___18633), .Q (_________30126));
  nnd2s1 ______440061(.DIN1 (____0_9__30017), .DIN2 (_____9___29895),
       .Q (_________30147));
  xor2s1 _______440062(.DIN1 (____9____29006), .DIN2 (____0____30019),
       .Q (____0____30042));
  or2s1 _______440063(.DIN1 (____0____30040), .DIN2 (____0____30039),
       .Q (____0____30041));
  or2s1 _______440064(.DIN1 (_______19043), .DIN2 (____0_0__30037), .Q
       (____0____30038));
  nor2s1 _______440065(.DIN1 (____9_9__29939), .DIN2 (____999__29999),
       .Q (____0_9__30036));
  nnd2s1 _____440066(.DIN1 (____9____29972), .DIN2 (____99___29998), .Q
       (____0____30035));
  nor2s1 _______440067(.DIN1 (____90__19196), .DIN2 (____0____30025),
       .Q (____0____30034));
  nnd2s1 _______440068(.DIN1 (____00___30002), .DIN2 (_________29857),
       .Q (____0____30033));
  nor2s1 _______440069(.DIN1 (____00___30006), .DIN2 (____0____30010),
       .Q (____0____30077));
  nnd2s1 ______440070(.DIN1 (____00___30001), .DIN2 (____9____29922),
       .Q (____0____30076));
  xor2s1 _______440071(.DIN1 (____9____29974), .DIN2 (____9____29953),
       .Q (____0____30057));
  nor2s1 ______440072(.DIN1 (____9____29948), .DIN2 (____0_0__30018),
       .Q (____090__30084));
  xor2s1 _______440073(.DIN1 (____9____29987), .DIN2 (_____9__23791),
       .Q (_____09__30102));
  xor2s1 _______440074(.DIN1 (___0_99__27363), .DIN2 (____0____30023),
       .Q (_________30338));
  hi1s1 _______440075(.DIN (____0____30070), .Q (_____90__33117));
  nor2s1 _______440076(.DIN1 (____0____30011), .DIN2 (____0____30031),
       .Q (____0____30032));
  nnd2s1 _____440077(.DIN1 (____990__29990), .DIN2 (____0____30029), .Q
       (____0____30030));
  nnd2s1 _______440078(.DIN1 (____0_9__30027), .DIN2 (____90___29906),
       .Q (____0_0__30028));
  nor2s1 _______440079(.DIN1 (____0____34547), .DIN2 (____9____29982),
       .Q (______0__31678));
  xor2s1 _______440080(.DIN1 (____9_0__29960), .DIN2 (_________29692),
       .Q (____0____30045));
  xor2s1 _______440081(.DIN1 (____9_0__29950), .DIN2 (_________28476),
       .Q (____0____30067));
  xor2s1 _______440082(.DIN1 (____9____29968), .DIN2 (____0____31872),
       .Q (____0_0__30064));
  hi1s1 _______440083(.DIN (____0____30025), .Q (____0____30026));
  nor2s1 _____0_440084(.DIN1 (___00____27193), .DIN2 (____0____30023),
       .Q (____0____30024));
  xnr2s1 _______440085(.DIN1 (____0____30021), .DIN2 (____000__30000),
       .Q (____0____30022));
  hi1s1 _______440086(.DIN (____0____30020), .Q (_____0___30371));
  and2s1 _____0_440087(.DIN1 (____9____29004), .DIN2 (____0____30019),
       .Q (____0____30058));
  nor2s1 _______440088(.DIN1 (_____9__23991), .DIN2 (____9____29977),
       .Q (_________33415));
  xor2s1 _______440089(.DIN1 (____9____29952), .DIN2 (____0____32762),
       .Q (_________30109));
  xor2s1 _______440090(.DIN1 (___9_0__24306), .DIN2 (____0____30013),
       .Q (____0____30070));
  nor2s1 _______440091(.DIN1 (____9____29965), .DIN2 (____0____32816),
       .Q (____0_0__30018));
  or2s1 _____0_440092(.DIN1 (_________________18713), .DIN2
       (____9____29961), .Q (____0_9__30017));
  dffacs1 ______________0____440093(.CLRB (reset), .CLK (clk), .DIN
       (____9____29956), .Q (_________34504));
  xor2s1 _______440094(.DIN1 (____9_9__29989), .DIN2 (____0_9__29137),
       .Q (____0____30016));
  xor2s1 _______440095(.DIN1 (_________________18696), .DIN2
       (_________33388), .Q (____0____30015));
  nnd2s1 _______440096(.DIN1 (____00___30003), .DIN2 (____00___30004),
       .Q (____0____30014));
  hi1s1 _______440097(.DIN (____0____30011), .Q (____0____30012));
  nor2s1 _______440098(.DIN1 (____0_0__30009), .DIN2 (____00___30005),
       .Q (____0____30010));
  nor2s1 _______440099(.DIN1 (____0____34547), .DIN2 (____9_0__29980),
       .Q (____009__30008));
  nor2s1 ______440100(.DIN1 (____00___30006), .DIN2 (____00___30005),
       .Q (____00___30007));
  xor2s1 _______440101(.DIN1 (_____0__23992), .DIN2 (____9____29976),
       .Q (____0____30043));
  nor2s1 _______440102(.DIN1 (____00___30004), .DIN2 (____00___30003),
       .Q (____0____30051));
  or2s1 ______440103(.DIN1 (____0____30080), .DIN2 (____9____29951), .Q
       (____00___30002));
  nnd2s1 _______440104(.DIN1 (____000__30000), .DIN2 (____9____29923),
       .Q (____00___30001));
  nor2s1 _______440105(.DIN1 (____9____29942), .DIN2 (_____09__30464),
       .Q (____999__29999));
  nnd2s1 ______440106(.DIN1 (_____09__30464), .DIN2 (____9____29938),
       .Q (____99___29998));
  and2s1 _______440107(.DIN1 (____99___29996), .DIN2
       (______________________________________0_____________18890), .Q
       (____99___29997));
  or2s1 _______440108(.DIN1
       (______________________________________0_____________18890),
       .DIN2 (____99___29996), .Q (____99___29995));
  nor2s1 _______440109(.DIN1 (_________29675), .DIN2 (____9____29947),
       .Q (____0____30054));
  nnd2s1 _____9_440110(.DIN1 (____0_0__30009), .DIN2 (_________34432),
       .Q (____0____30025));
  nor2s1 _____0_440111(.DIN1 (_________34432), .DIN2 (____0_0__30009),
       .Q (____0_0__30056));
  nnd2s1 _______440112(.DIN1 (____9____29954), .DIN2 (____9____29973),
       .Q (____0____30020));
  and2s1 _______440113(.DIN1 (____99___29996), .DIN2 (_________31281),
       .Q (____0____30040));
  nor2s1 _______440114(.DIN1 (_________31281), .DIN2 (____99___29996),
       .Q (____0____30039));
  nor2s1 _____9_440115(.DIN1 (_______19020), .DIN2 (____9____29967), .Q
       (____0_0__30037));
  or2s1 _______440116(.DIN1 (_________________18696), .DIN2
       (_________33388), .Q (____99___29994));
  xor2s1 _______440117(.DIN1 (____9____29921), .DIN2 (_________33007),
       .Q (____99___29993));
  nnd2s1 _______440118(.DIN1 (____9_9__29969), .DIN2 (____9____29913),
       .Q (____99___29992));
  nor2s1 ______440119(.DIN1 (_________29887), .DIN2 (____9____29937),
       .Q (____99___29991));
  nnd2s1 _______440120(.DIN1 (____9____29983), .DIN2 (____9_9__29989),
       .Q (____990__29990));
  xor2s1 _______440121(.DIN1 (____9____29957), .DIN2 (____9____29958),
       .Q (____9____29988));
  xor2s1 _______440122(.DIN1 (____9____29986), .DIN2 (____9____29966),
       .Q (____9____29987));
  nnd2s1 _______440123(.DIN1 (_________33388), .DIN2
       (_________________18696), .Q (____9____29985));
  or2s1 _______440124(.DIN1 (____9_9__29989), .DIN2 (____9____29983),
       .Q (____9____29984));
  nor2s1 _______440125(.DIN1 (____9____29981), .DIN2 (____9_0__29980),
       .Q (____9____29982));
  xor2s1 _______440126(.DIN1 (____9____29917), .DIN2
       (_________________18713), .Q (_________31546));
  nor2s1 _______440127(.DIN1 (__99____27138), .DIN2 (____9____29941),
       .Q (____0____30023));
  xor2s1 _______440128(.DIN1 (____9____29916), .DIN2 (_________29585),
       .Q (____9_9__29979));
  xor2s1 _______440129(.DIN1 (________________18705), .DIN2
       (____0____32816), .Q (____9____29978));
  and2s1 _____440130(.DIN1 (____9____29976), .DIN2 (________19101), .Q
       (____9____29977));
  or2s1 _____9_440131(.DIN1 (____0____30080), .DIN2 (____9____29928),
       .Q (____9____29975));
  and2s1 _______440132(.DIN1 (____9____29973), .DIN2 (____9____29927),
       .Q (____9____29974));
  nnd2s1 _______440133(.DIN1 (____9____29971), .DIN2 (____9____29944),
       .Q (____9____29972));
  nnd2s1 _______440134(.DIN1 (____9____29935), .DIN2 (____9____29934),
       .Q (____0____30029));
  nor2s1 _______440135(.DIN1 (____9_0__29970), .DIN2 (_________33388),
       .Q (____0____30011));
  and2s1 _______440136(.DIN1 (_________33388), .DIN2 (____9_0__29970),
       .Q (____0____30031));
  nor2s1 _____0_440137(.DIN1 (_________28477), .DIN2 (____9_9__29929),
       .Q (____09___30091));
  nnd2s1 _______440138(.DIN1 (____9_9__29969), .DIN2 (____9____29914),
       .Q (____0_9__30027));
  nor2s1 _______440139(.DIN1 (_________29676), .DIN2 (____9____29946),
       .Q (____0____30053));
  nnd2s1 _______440140(.DIN1 (____9____29931), .DIN2 (_____99__28799),
       .Q (____0____30019));
  xor2s1 _______440141(.DIN1 (____90___29902), .DIN2 (___9____22478),
       .Q (____9____29968));
  nor2s1 _______440142(.DIN1 (_______18960), .DIN2 (____9____29966), .Q
       (____9____29967));
  nor2s1 _____9_440143(.DIN1 (________________18705), .DIN2
       (____9____29964), .Q (____9____29965));
  hi1s1 _______440144(.DIN (____9____29962), .Q (____9____29963));
  xor2s1 _______440145(.DIN1 (_____99__29900), .DIN2 (____0_0__31861),
       .Q (____9____29961));
  xor2s1 _______440146(.DIN1 (____9____29936), .DIN2 (_________29889),
       .Q (____9_0__29960));
  or2s1 _______440147(.DIN1 (____9____29958), .DIN2 (____9____29957),
       .Q (____9_9__29959));
  nnd2s1 _______440148(.DIN1 (____9_9__29919), .DIN2 (_________34393),
       .Q (____9____29956));
  nnd2s1 ______440149(.DIN1 (____9____29957), .DIN2 (____9____29958),
       .Q (____9____29955));
  xor2s1 ______440150(.DIN1 (____90___29903), .DIN2 (_________32410),
       .Q (____00___30003));
  xor2s1 _______440151(.DIN1 (____9____29943), .DIN2 (____99___31805),
       .Q (_____09__30464));
  xor2s1 _______440152(.DIN1 (__99____27140), .DIN2 (____9_0__29940),
       .Q (____99___29996));
  or2s1 _______440153(.DIN1 (____9____29953), .DIN2 (____9____29926),
       .Q (____9____29954));
  nor2s1 _____440154(.DIN1 (______9__29822), .DIN2 (____9____29915), .Q
       (____9____29952));
  xor2s1 _______440155(.DIN1 (____9_0__29930), .DIN2 (_________28825),
       .Q (____9____29951));
  xor2s1 ______440156(.DIN1 (_________34482), .DIN2 (____9_9__29949),
       .Q (____9_0__29950));
  and2s1 _____9_440157(.DIN1 (____9____29964), .DIN2
       (________________18705), .Q (____9____29948));
  hi1s1 _______440158(.DIN (____9____29946), .Q (____9____29947));
  nor2s1 _____440159(.DIN1 (___9___18952), .DIN2 (____9____29912), .Q
       (____0____30013));
  and2s1 _______440160(.DIN1 (____9____29945), .DIN2 (_________34497),
       .Q (____00___30005));
  nor2s1 _____0_440161(.DIN1 (_________34497), .DIN2 (____9____29945),
       .Q (____00___30006));
  nnd2s1 _____9_440162(.DIN1 (____9____29925), .DIN2 (_____90__29793),
       .Q (____000__30000));
  xor2s1 _______440163(.DIN1 (____90___29907), .DIN2 (______9__28578),
       .Q (____0_0__30009));
  nnd2s1 _______440164(.DIN1 (____9____29943), .DIN2 (____9____29942),
       .Q (____9____29944));
  nor2s1 _______440165(.DIN1 (__99____27139), .DIN2 (____9_0__29940),
       .Q (____9____29941));
  nor2s1 _______440166(.DIN1 (____9____29938), .DIN2 (____9____29943),
       .Q (____9_9__29939));
  nor2s1 _______440167(.DIN1 (______9__29890), .DIN2 (____9____29936),
       .Q (____9____29937));
  nnd2s1 _____9_440168(.DIN1 (_____9___29898), .DIN2 (____9____31752),
       .Q (____9____29935));
  nnd2s1 _____9_440169(.DIN1 (_____9___29896), .DIN2 (_________33333),
       .Q (____9____29934));
  xor2s1 _______440170(.DIN1 (______0__29881), .DIN2 (_________29733),
       .Q (____9____29962));
  nor2s1 _____0_440171(.DIN1 (____909__29910), .DIN2 (____0_9__34549),
       .Q (____9_0__29980));
  dffacs1 __________________440172(.CLRB (reset), .CLK (clk), .DIN
       (____900__29901), .Q (________________18677));
  xor2s1 _______440173(.DIN1 (____9____29932), .DIN2 (_________30131),
       .Q (____9____29933));
  nnd2s1 _______440174(.DIN1 (_____9___28798), .DIN2 (____9_0__29930),
       .Q (____9____29931));
  nor2s1 _______440175(.DIN1 (_________34482), .DIN2 (_________28449),
       .Q (____9_9__29929));
  xor2s1 _______440176(.DIN1 (_________29884), .DIN2 (_________29868),
       .Q (____9____29928));
  hi1s1 _______440177(.DIN (____9____29926), .Q (____9____29927));
  xnr2s1 _______440178(.DIN1 (______0__31325), .DIN2 (_________29872),
       .Q (____9_9__29969));
  nor2s1 _______440179(.DIN1 (_______19011), .DIN2 (_____9___29894), .Q
       (____9____29976));
  xor2s1 _______440180(.DIN1 (_____90__29891), .DIN2 (___0__0__27685),
       .Q (____9____29946));
  xor2s1 ______440181(.DIN1 (______0__29871), .DIN2 (____0____30981),
       .Q (____9_9__29989));
  xnr2s1 _______440182(.DIN1 (____9____29911), .DIN2 (____9___22259),
       .Q (_________33388));
  nnd2s1 _______440183(.DIN1 (_________29885), .DIN2 (_________29817),
       .Q (____9____29925));
  xor2s1 _______440184(.DIN1 (_________________18763), .DIN2
       (_________33330), .Q (____9____29924));
  or2s1 ______440185(.DIN1 (_______________18874), .DIN2
       (____0____30021), .Q (____9____29923));
  nnd2s1 ______440186(.DIN1 (____0____30021), .DIN2
       (_______________18874), .Q (____9____29922));
  nnd2s1 ______440187(.DIN1 (____0____30021), .DIN2 (_____9__26006), .Q
       (____9____29921));
  nnd2s1 ______440188(.DIN1 (______9__29880), .DIN2 (___9____19692), .Q
       (____9_0__29920));
  xor2s1 _______440189(.DIN1 (_____9___29897), .DIN2 (______0__29757),
       .Q (____9_9__29919));
  xor2s1 _______440190(.DIN1 (_________29855), .DIN2 (___0__18931), .Q
       (____9____29918));
  xor2s1 _______440191(.DIN1 (_____9___29899), .DIN2 (_________33330),
       .Q (____9____29917));
  nor2s1 _______440192(.DIN1 (________19422), .DIN2 (_________29883),
       .Q (____9____29966));
  xor2s1 ______440193(.DIN1 (_____9___29893), .DIN2
       (_________9______18801), .Q (____9____29916));
  nor2s1 _______440194(.DIN1 (________21942), .DIN2 (_________29874),
       .Q (____9____29915));
  nnd2s1 ______440195(.DIN1 (____9____29913), .DIN2 (_________31058),
       .Q (____9____29914));
  nor2s1 ______440196(.DIN1 (________19138), .DIN2 (____9____29911), .Q
       (____9____29912));
  nor2s1 _______440197(.DIN1 (____0____30080), .DIN2 (_________29867),
       .Q (____90___29909));
  nor2s1 _______440198(.DIN1 (____90___29908), .DIN2 (____9____29932),
       .Q (____9____29926));
  nnd2s1 _______440199(.DIN1 (____9____29932), .DIN2 (____90___29908),
       .Q (____9____29973));
  nnd2s1 _______440200(.DIN1 (______9__29870), .DIN2 (_________29819),
       .Q (____9____29945));
  xor2s1 ______440201(.DIN1 (_________29839), .DIN2 (_________29873),
       .Q (____9____29957));
  dffacs1 __________________440202(.CLRB (reset), .CLK (clk), .DIN
       (_________29875), .Q (________________18705));
  xor2s1 _______440203(.DIN1 (_________29818), .DIN2 (_________31951),
       .Q (____90___29907));
  nnd2s1 _______440204(.DIN1 (_________29877), .DIN2
       (_______________18879), .Q (____90___29906));
  and2s1 _______440205(.DIN1 (_________33330), .DIN2 (____90___29904),
       .Q (____90___29905));
  xor2s1 _______440206(.DIN1 (_________29814), .DIN2 (_________31252),
       .Q (____90___29903));
  xor2s1 _______440207(.DIN1 (_________29815), .DIN2 (_________29330),
       .Q (____90___29902));
  xor2s1 _______440208(.DIN1 (_________29816), .DIN2 (_________33564),
       .Q (____9_0__29940));
  nor2s1 _____0_440209(.DIN1 (_________29731), .DIN2 (_________29849),
       .Q (____9____29936));
  nnd2s1 _______440210(.DIN1 (_________29842), .DIN2 (_____9___29794),
       .Q (____9_0__29930));
  dffacs1 _____________9____440211(.CLRB (reset), .CLK (clk), .DIN
       (______0__29841), .Q (_________9______18802));
  xor2s1 _____0_440212(.DIN1 (_________29882), .DIN2 (_________30524),
       .Q (____9____29943));
  dffacs1 _______________440213(.CLRB (reset), .CLK (clk), .DIN
       (______9__29860), .QN (outData[2]));
  or2s1 ______440214(.DIN1 (_________29859), .DIN2 (___9____21582), .Q
       (____900__29901));
  nnd2s1 _______440215(.DIN1 (_________33330), .DIN2 (_____9___29899),
       .Q (_____99__29900));
  nor2s1 _______440216(.DIN1 (_________29846), .DIN2 (_____9___29897),
       .Q (_____9___29898));
  nnd2s1 _______440217(.DIN1 (_________29847), .DIN2 (_________29853),
       .Q (_____9___29896));
  or2s1 _______440218(.DIN1 (_____9___29899), .DIN2 (_________33330),
       .Q (_____9___29895));
  and2s1 _______440219(.DIN1 (_____9___29893), .DIN2 (_______19025), .Q
       (_____9___29894));
  nor2s1 _______440220(.DIN1 (____90___29904), .DIN2 (_________33330),
       .Q (_____9___29892));
  xor2s1 _______440221(.DIN1 (_________29829), .DIN2 (_________31252),
       .Q (____909__29910));
  xor2s1 ______440222(.DIN1 (_________29826), .DIN2 (___0__18931), .Q
       (____0____30050));
  nnd2s1 _____9_440223(.DIN1 (_________29862), .DIN2 (_________29753),
       .Q (____9____29971));
  dffacs1 __________________440224(.CLRB (reset), .CLK (clk), .DIN
       (_________29856), .Q (_________34482));
  xor2s1 _______440225(.DIN1 (_________________18742), .DIN2
       (_____9___31351), .Q (_____90__29891));
  and2s1 ______440226(.DIN1 (_________29889), .DIN2 (_________29886),
       .Q (______9__29890));
  xor2s1 _______440227(.DIN1 (_____0___29810), .DIN2 (_____0___31184),
       .Q (_________29888));
  nor2s1 _______440228(.DIN1 (_________29886), .DIN2 (_________29889),
       .Q (_________29887));
  xnr2s1 _____9_440229(.DIN1 (____90___33582), .DIN2 (______9__29792),
       .Q (_________29885));
  nor2s1 _____440230(.DIN1 (_________29820), .DIN2 (_________29869), .Q
       (_________29884));
  nor2s1 _______440231(.DIN1 (________19421), .DIN2 (_________29882),
       .Q (_________29883));
  xor2s1 ______440232(.DIN1 (_________29734), .DIN2 (_________29848),
       .Q (______0__29881));
  xor2s1 _______440233(.DIN1 (_________29791), .DIN2 (_________29784),
       .Q (______9__29880));
  or2s1 _______440234(.DIN1 (_________29879), .DIN2 (_________29878),
       .Q (______0__31390));
  nor2s1 _______440235(.DIN1 (___9____22479), .DIN2 (_________29824),
       .Q (____9____29958));
  xor2s1 _______440236(.DIN1 (______0__29861), .DIN2 (_____9___29801),
       .Q (____9____29932));
  hi1s1 _______440237(.DIN (_________29877), .Q (____0____30021));
  nor2s1 _______440238(.DIN1 (_________29825), .DIN2 (_________32639),
       .Q (_________29876));
  nor2s1 _______440239(.DIN1 (_________________0___18660), .DIN2
       (_________29821), .Q (_________29875));
  and2s1 _______440240(.DIN1 (_________29838), .DIN2 (_________29873),
       .Q (_________29874));
  nor2s1 _______440241(.DIN1 (_________29863), .DIN2 (_________29864),
       .Q (_________29872));
  xor2s1 _____0_440242(.DIN1 (_____0___29804), .DIN2
       (___________0___18872), .Q (______0__29871));
  or2s1 _____0_440243(.DIN1 (_________29869), .DIN2 (_________29868),
       .Q (______9__29870));
  xor2s1 _____440244(.DIN1 (_________29787), .DIN2 (_____0___29806), .Q
       (_________29867));
  hi1s1 _____9_440245(.DIN (_________29865), .Q (_________29866));
  nor2s1 _____9_440246(.DIN1 (_________29827), .DIN2 (_________29834),
       .Q (_____9___31531));
  nor2s1 _____9_440247(.DIN1 (________25503), .DIN2 (______0__29833),
       .Q (____9____29911));
  nor2s1 ______440248(.DIN1 (___0_____27686), .DIN2 (_________29835),
       .Q (______0__32496));
  nnd2s1 _______440249(.DIN1 (_________29864), .DIN2 (_________29863),
       .Q (____9____29913));
  nnd2s1 _______440250(.DIN1 (______0__29861), .DIN2 (_________29761),
       .Q (_________29862));
  or2s1 ______440251(.DIN1 (_________34501), .DIN2 (_____99__30363), .Q
       (______9__29860));
  nor2s1 _______440252(.DIN1 (_____9___29798), .DIN2 (_________29858),
       .Q (_________29859));
  or2s1 _______440253(.DIN1 (_________29858), .DIN2 (_____9___29799),
       .Q (_________29857));
  nnd2s1 ______440254(.DIN1 (_____9___29800), .DIN2 (_________34393),
       .Q (_________29856));
  xor2s1 _______440255(.DIN1 (_____0___29809), .DIN2 (_________29854),
       .Q (_________29855));
  nnd2s1 _______440256(.DIN1 (_____09__29812), .DIN2 (_____99__29802),
       .Q (_____9___29893));
  nnd2s1 _______440257(.DIN1 (_________29845), .DIN2 (_________29853),
       .Q (_____9___29897));
  xor2s1 _______440258(.DIN1 (______9__29775), .DIN2 (____099__30093),
       .Q (_________33114));
  nor2s1 ______440259(.DIN1 (___09____28063), .DIN2 (_____0___29811),
       .Q (____0____30068));
  xnr2s1 _______440260(.DIN1 (______9__29832), .DIN2 (________25505),
       .Q (_________33330));
  nnd2s1 ______440261(.DIN1 (_________29843), .DIN2 (______0__29851),
       .Q (_________29852));
  xor2s1 _____0_440262(.DIN1 (_________29854), .DIN2 (____0___22720),
       .Q (______9__29850));
  nor2s1 _______440263(.DIN1 (_________29735), .DIN2 (_________29848),
       .Q (_________29849));
  nnd2s1 _______440264(.DIN1 (_________29846), .DIN2 (_________29845),
       .Q (_________29847));
  nor2s1 _______440265(.DIN1 (______0__29851), .DIN2 (_________29843),
       .Q (_________29844));
  nnd2s1 ______440266(.DIN1 (_____9___29796), .DIN2 (_________28645),
       .Q (_________29842));
  nnd2s1 _______440267(.DIN1 (_____0___29808), .DIN2 (________19987),
       .Q (______0__29841));
  xor2s1 _____0_440268(.DIN1 (____0___21721), .DIN2 (_________29840),
       .Q (_________29839));
  xor2s1 _____0_440269(.DIN1 (______0__29823), .DIN2 (______0__35098),
       .Q (_________29865));
  xor2s1 _______440270(.DIN1 (_________29780), .DIN2 (_________30104),
       .Q (_________29877));
  nnd2s1 _______440271(.DIN1 (_________29840), .DIN2 (___0_____27735),
       .Q (_________29838));
  nnd2s1 _______440272(.DIN1 (_________29854), .DIN2 (______9__34490),
       .Q (_________29837));
  nor2s1 _______440273(.DIN1 (______9__34490), .DIN2 (_________29854),
       .Q (_________29836));
  nor2s1 ______440274(.DIN1 (___0__9__27684), .DIN2 (_________29790),
       .Q (_________29835));
  nor2s1 _______440275(.DIN1 (_________31252), .DIN2 (_________29828),
       .Q (_________29834));
  nor2s1 _______440276(.DIN1 (________25504), .DIN2 (______9__29832),
       .Q (______0__29833));
  nor2s1 _______440277(.DIN1 (_________________18774), .DIN2
       (_________29854), .Q (_________29831));
  and2s1 _______440278(.DIN1 (_________29854), .DIN2
       (_________________18774), .Q (_________29830));
  or2s1 _______440279(.DIN1 (_________29828), .DIN2 (_________29827),
       .Q (_________29829));
  nor2s1 _______440280(.DIN1 (_________29744), .DIN2 (_________29785),
       .Q (_________29826));
  nor2s1 _______440281(.DIN1 (______9__29728), .DIN2 (______0__29776),
       .Q (_________29864));
  xor2s1 _______440282(.DIN1 (______9__29765), .DIN2 (_____9___33022),
       .Q (_________29889));
  nor2s1 _______440283(.DIN1 (_________32437), .DIN2 (_________29789),
       .Q (_________29825));
  nor2s1 ______440284(.DIN1 (___9____22476), .DIN2 (______0__29823), .Q
       (_________29824));
  nor2s1 ______440285(.DIN1 (___0____22551), .DIN2 (_________29840), .Q
       (______9__29822));
  xor2s1 _______440286(.DIN1 (_____9___29795), .DIN2 (_________29758),
       .Q (_________29821));
  hi1s1 _______440287(.DIN (_________29819), .Q (_________29820));
  xnr2s1 _______440288(.DIN1 (_________29817), .DIN2 (_________29863),
       .Q (_________29818));
  nnd2s1 _____9_440289(.DIN1 (_________29778), .DIN2 (_________29779),
       .Q (_________29816));
  xor2s1 _____0_440290(.DIN1 (_________29774), .DIN2 (_________35050),
       .Q (_________29815));
  xor2s1 _____0_440291(.DIN1 (___09____28062), .DIN2 (_________34483),
       .Q (_________29814));
  xor2s1 _____440292(.DIN1 (______9__34490), .DIN2 (______0__32899), .Q
       (______0__29813));
  nor2s1 _______440293(.DIN1 (_________29722), .DIN2 (_________29782),
       .Q (_________29878));
  xor2s1 _______440294(.DIN1 (______9__29756), .DIN2 (______9__32232),
       .Q (_________29882));
  nor2s1 _______440295(.DIN1 (_____0___29805), .DIN2 (_________29788),
       .Q (_________29868));
  nnd2s1 _______440296(.DIN1 (_____00__29803), .DIN2
       (___________0___18872), .Q (_____09__29812));
  nor2s1 _______440297(.DIN1 (_________34483), .DIN2 (____0____28161),
       .Q (_____0___29811));
  nor2s1 _______440298(.DIN1 (_____0___29809), .DIN2 (______0__32899),
       .Q (_____0___29810));
  dffacs1 ______________0____440299(.CLRB (reset), .CLK (clk), .DIN
       (_________29771), .Q (_________34501));
  or2s1 ______440300(.DIN1 (______0__33373), .DIN2 (_________29768), .Q
       (_____0___29808));
  nor2s1 _______440301(.DIN1 (_________29760), .DIN2 (_____00__33220),
       .Q (_____0___29807));
  nor2s1 ______440302(.DIN1 (_____0___29805), .DIN2 (_________29767),
       .Q (_____0___29806));
  and2s1 ______440303(.DIN1 (_____00__29803), .DIN2 (_____99__29802),
       .Q (_____0___29804));
  nnd2s1 ______440304(.DIN1 (_________28921), .DIN2 (_________29770),
       .Q (_________29845));
  and2s1 ______440305(.DIN1 (______0__32899), .DIN2 (_____0___29809),
       .Q (_________29843));
  nor2s1 _______440306(.DIN1 (______0__29624), .DIN2 (_________29773),
       .Q (_________29848));
  nor2s1 _______440307(.DIN1 (_________29723), .DIN2 (_________29781),
       .Q (_________29879));
  nor2s1 _______440308(.DIN1 (_________29754), .DIN2 (_________29755),
       .Q (_____9___29801));
  xor2s1 _____9_440309(.DIN1 (_________29740), .DIN2 (_________34494),
       .Q (_____9___29800));
  xor2s1 _____9_440310(.DIN1 (________________18677), .DIN2
       (_____9___29797), .Q (_____9___29799));
  xor2s1 _____9_440311(.DIN1 (________________18676), .DIN2
       (_____9___29797), .Q (_____9___29798));
  or2s1 _______440312(.DIN1 (________________18689), .DIN2
       (_____9___29795), .Q (_____9___29796));
  nnd2s1 _______440313(.DIN1 (_____9___29795), .DIN2
       (________________18689), .Q (_____9___29794));
  or2s1 _______440314(.DIN1 (_______________18873), .DIN2
       (_________29863), .Q (_____90__29793));
  and2s1 _______440315(.DIN1 (_________29863), .DIN2
       (_______________18873), .Q (______9__29792));
  xor2s1 _______440316(.DIN1 (_________29746), .DIN2 (_________29745),
       .Q (_________29791));
  nnd2s1 _______440317(.DIN1 (_________29764), .DIN2 (_________29572),
       .Q (______0__29861));
  xor2s1 ______440318(.DIN1 (_________29737), .DIN2 (_________31505),
       .Q (_________29869));
  xor2s1 _______440319(.DIN1 (_________29741), .DIN2 (____0____31863),
       .Q (_________29819));
  hi1s1 ______440320(.DIN (_________29790), .Q (_____9___31351));
  nor2s1 ______440321(.DIN1 (_________18860), .DIN2 (________21366), .Q
       (_________29789));
  and2s1 _______440322(.DIN1 (______0__29766), .DIN2 (_________29787),
       .Q (_________29788));
  nnd2s1 _______440323(.DIN1 (_________29668), .DIN2 (_________18860),
       .Q (_________29786));
  nor2s1 _______440324(.DIN1 (______9__29747), .DIN2 (_________29784),
       .Q (_________29785));
  nnd2s1 _______440325(.DIN1 (_____0___28899), .DIN2 (_________29769),
       .Q (_________29853));
  and2s1 _______440326(.DIN1 (_________34752), .DIN2 (_________18860),
       .Q (_________29827));
  nor2s1 _______440327(.DIN1 (_________18860), .DIN2 (_________34752),
       .Q (_________29828));
  nor2s1 _______440328(.DIN1 (__9__9__26458), .DIN2 (_________29748),
       .Q (______9__29832));
  hi1s1 _______440329(.DIN (_________29781), .Q (_________29782));
  and2s1 _______440330(.DIN1 (_________29777), .DIN2 (_________29779),
       .Q (_________29780));
  nnd2s1 _______440331(.DIN1 (_________29777), .DIN2 (_________30104),
       .Q (_________29778));
  xnr2s1 _____9_440332(.DIN1 (_____00__30545), .DIN2 (_________29727),
       .Q (______0__29776));
  nnd2s1 _______440333(.DIN1 (______0__29739), .DIN2 (______9__29689),
       .Q (______9__29775));
  xor2s1 ______440334(.DIN1 (_________29693), .DIN2 (_________29772),
       .Q (_________33003));
  hi1s1 _______440335(.DIN (_________29774), .Q (______0__29823));
  xor2s1 _____0_440336(.DIN1 (___________0___18877), .DIN2
       (______0__29729), .Q (_________29790));
  xnr2s1 _____0_440337(.DIN1 (_________29674), .DIN2 (_________29763),
       .Q (_________29840));
  hi1s1 _____440338(.DIN (______0__32899), .Q (_________29854));
  and2s1 _______440339(.DIN1 (_________29772), .DIN2 (______9__29579),
       .Q (_________29773));
  nnd2s1 _______440340(.DIN1 (_________29721), .DIN2 (_________34393),
       .Q (_________29771));
  hi1s1 _______440341(.DIN (_________29769), .Q (_________29770));
  xor2s1 _____9_440342(.DIN1 (_____9___29706), .DIN2 (______9__29738),
       .Q (_________29768));
  hi1s1 ______440343(.DIN (______0__29766), .Q (_________29767));
  xor2s1 _____440344(.DIN1 (_____0___29714), .DIN2 (_____0___29715), .Q
       (______9__29765));
  nnd2s1 _______440345(.DIN1 (_________29763), .DIN2 (______9__29661),
       .Q (_________29764));
  xor2s1 _____0_440346(.DIN1 (_____9___29702), .DIN2 (_________29762),
       .Q (_________29774));
  xor2s1 _____9_440347(.DIN1 (_________________18712), .DIN2
       (_____99__29709), .Q (_________29781));
  dffacs1 __________________440348(.CLRB (reset), .CLK (clk), .DIN
       (_________29732), .Q (_________34483));
  xor2s1 ______440349(.DIN1 (_____0___29711), .DIN2 (_________34702),
       .Q (_________32965));
  xor2s1 _____0_440350(.DIN1 (_________29697), .DIN2 (___0__18931), .Q
       (_________32446));
  xor2s1 _____440351(.DIN1 (______0__34688), .DIN2 (__9__0__26825), .Q
       (______0__32899));
  or2s1 _____0_440352(.DIN1 (____9____29071), .DIN2 (_________30388),
       .Q (_________29761));
  hi1s1 _______440353(.DIN (_________29759), .Q (_________29760));
  xnr2s1 _______440354(.DIN1 (________________18689), .DIN2
       (_________28645), .Q (_________29758));
  xnr2s1 _______440355(.DIN1 (______0__32594), .DIN2 (_________29846),
       .Q (______0__29757));
  nnd2s1 _______440356(.DIN1 (_____09__29718), .DIN2 (_________29655),
       .Q (______9__29756));
  and2s1 _____0_440357(.DIN1 (_________30388), .DIN2 (____90___28994),
       .Q (_________29755));
  nor2s1 _____0_440358(.DIN1 (____999__29082), .DIN2 (_________30388),
       .Q (_________29754));
  nnd2s1 _____0_440359(.DIN1 (_________30388), .DIN2 (_____0___28905),
       .Q (_________29753));
  nnd2s1 _______440360(.DIN1 (_________29751), .DIN2 (_________29750),
       .Q (_________29752));
  or2s1 ______440361(.DIN1 (_________9______18800), .DIN2
       (_________29749), .Q (_____99__29802));
  nnd2s1 ______440362(.DIN1 (_________29749), .DIN2
       (_________9______18800), .Q (_____00__29803));
  nnd2s1 _______440363(.DIN1 (_________29720), .DIN2 (______0__29652),
       .Q (_____9___29795));
  xnr2s1 ______440364(.DIN1 (_________28593), .DIN2 (_____90__29700),
       .Q (_________29863));
  nor2s1 _______440365(.DIN1 (__9_____26731), .DIN2 (______0__34688),
       .Q (_________29748));
  nor2s1 _______440366(.DIN1 (_________29743), .DIN2 (_________29746),
       .Q (______9__29747));
  xor2s1 _____0_440367(.DIN1 (_____9___29703), .DIN2 (_________35012),
       .Q (_________29745));
  and2s1 _______440368(.DIN1 (_________29746), .DIN2 (_________29743),
       .Q (_________29744));
  nnd2s1 _______440369(.DIN1 (_____0___29717), .DIN2
       (______________0___________________0), .Q (______0__29766));
  nor2s1 _______440370(.DIN1 (_____9___29708), .DIN2 (_________29742),
       .Q (_________29783));
  xor2s1 _____9_440371(.DIN1 (_________29694), .DIN2 (_________35094),
       .Q (_________29769));
  nor2s1 _______440372(.DIN1 (_____0___29712), .DIN2 (_____0___29716),
       .Q (____0_9__30073));
  nor2s1 _______440373(.DIN1 (_________18845), .DIN2 (_________29742),
       .Q (_____00__33220));
  dffacs1 __________________440374(.CLRB (reset), .CLK (clk), .DIN
       (_____00__29710), .QN (_________18860));
  nor2s1 _______440375(.DIN1 (________________18678), .DIN2
       (_________33098), .Q (_________29741));
  xor2s1 ______440376(.DIN1 (______0__29719), .DIN2 (____0____32816),
       .Q (_________29740));
  or2s1 _______440377(.DIN1 (______9__29738), .DIN2 (_________29695),
       .Q (______0__29739));
  and2s1 _______440378(.DIN1 (_________33098), .DIN2
       (________________18678), .Q (_________29737));
  nnd2s1 ______440379(.DIN1 (________________18689), .DIN2
       (______18920), .Q (_____9___29797));
  xor2s1 _______440380(.DIN1 (_________29681), .DIN2 (_________29736),
       .Q (____00___30004));
  nnd2s1 _____9_440381(.DIN1 (______9__29699), .DIN2 (____9_0__29047),
       .Q (_________29777));
  xnr2s1 _______440382(.DIN1 (_____00__30545), .DIN2 (_________29691),
       .Q (_________29759));
  xor2s1 _______440383(.DIN1 (______0__29680), .DIN2 (____0_9__28157),
       .Q (_________31077));
  dffacs1 _____________9____440384(.CLRB (reset), .CLK (clk), .DIN
       (_____9___29701), .Q (_________9______18801));
  nor2s1 ______440385(.DIN1 (_________29734), .DIN2 (_________29733),
       .Q (_________29735));
  nnd2s1 _______440386(.DIN1 (______0__29690), .DIN2 (_________34365),
       .Q (_________29732));
  and2s1 _______440387(.DIN1 (_________29734), .DIN2 (_________29733),
       .Q (_________29731));
  or2s1 _______440388(.DIN1 (_________________18712), .DIN2
       (_________29677), .Q (_________29730));
  nor2s1 _______440389(.DIN1 (______9__29728), .DIN2 (_________29726),
       .Q (______0__29729));
  nor2s1 _______440390(.DIN1 (_________33835), .DIN2 (_________29726),
       .Q (_________29727));
  nor2s1 _______440391(.DIN1 (_________29642), .DIN2 (_________29687),
       .Q (_________29749));
  xor2s1 _____0_440392(.DIN1 (_________29672), .DIN2 (____00___31810),
       .Q (_________29772));
  nor2s1 _____9_440393(.DIN1 (_________29724), .DIN2 (_________29684),
       .Q (_________29725));
  hi1s1 _______440394(.DIN (_________29722), .Q (_________29723));
  xor2s1 _______440395(.DIN1 (_________29648), .DIN2 (_________29649),
       .Q (_________29721));
  or2s1 _____0_440396(.DIN1 (_________29653), .DIN2 (______0__29719),
       .Q (_________29720));
  nnd2s1 _______440397(.DIN1 (_________29678), .DIN2 (outData[20]), .Q
       (_____09__29718));
  nnd2s1 _____9_440398(.DIN1 (_________29698), .DIN2
       (_______________18876), .Q (_________29779));
  nnd2s1 ______440399(.DIN1 (_________29686), .DIN2 (_________29520),
       .Q (_________29763));
  xor2s1 _______440400(.DIN1 (_________29659), .DIN2 (_________32049),
       .Q (_________29751));
  xor2s1 _______440401(.DIN1 (_________29658), .DIN2 (___0____21689),
       .Q (_________30388));
  xor2s1 _______440402(.DIN1 (_____9___29705), .DIN2 (_____0___33866),
       .Q (_____0___29717));
  nor2s1 ______440403(.DIN1 (_____0___29715), .DIN2 (_____0___29713),
       .Q (_____0___29716));
  nor2s1 _______440404(.DIN1 (_____0___29713), .DIN2 (_____0___29712),
       .Q (_____0___29714));
  xor2s1 _____0_440405(.DIN1 (_________29641), .DIN2 (_________29583),
       .Q (_____0___29711));
  nnd2s1 _______440406(.DIN1 (_________29669), .DIN2 (____90___32662),
       .Q (_____00__29710));
  xor2s1 ______440407(.DIN1 (_____9___29708), .DIN2 (_____9___29707),
       .Q (_____99__29709));
  xor2s1 _______440408(.DIN1 (________21852), .DIN2 (_____9___29705),
       .Q (_____9___29706));
  xor2s1 _______440409(.DIN1 (_________________18694), .DIN2
       (_____9___29707), .Q (_____9___29704));
  hi1s1 _______440410(.DIN (_____9___29703), .Q (_________29743));
  xor2s1 _______440411(.DIN1 (_____9___29707), .DIN2 (____099__30093),
       .Q (_________29742));
  xor2s1 ______440412(.DIN1 (_________29685), .DIN2 (_________29552),
       .Q (_____9___29702));
  nnd2s1 _____9_440413(.DIN1 (_________29667), .DIN2 (________20550),
       .Q (_____9___29701));
  xor2s1 _____0_440414(.DIN1 (_________29636), .DIN2 (____09___30086),
       .Q (_____90__29700));
  hi1s1 _______440415(.DIN (_________29698), .Q (______9__29699));
  xor2s1 _______440416(.DIN1 (_________29644), .DIN2 (_________29696),
       .Q (_________29697));
  nnd2s1 ______440417(.DIN1 (_________29657), .DIN2 (_________29629),
       .Q (_________29817));
  nor2s1 _____9_440418(.DIN1 (______________0___________________0),
       .DIN2 (_________29654), .Q (_____0___29805));
  xor2s1 _______440419(.DIN1 (______9__29633), .DIN2 (____9____32728),
       .Q (______9__29738));
  nnd2s1 _____9_440420(.DIN1 (_________29663), .DIN2 (____0_0__28158),
       .Q (_________29722));
  nor2s1 _____440421(.DIN1 (_________29647), .DIN2 (_________29650), .Q
       (_________29846));
  dffacs1 __________________440422(.CLRB (reset), .CLK (clk), .DIN
       (_________29666), .Q (________________18689));
  xor2s1 _______440423(.DIN1 (_________29630), .DIN2 (_________29656),
       .Q (_________33098));
  nor2s1 _______440424(.DIN1 (_________29688), .DIN2 (_____9___29705),
       .Q (_________29695));
  xor2s1 _______440425(.DIN1 (_____0___29621), .DIN2 (_________29592),
       .Q (_________29694));
  xor2s1 _______440426(.DIN1 (_________29625), .DIN2
       (_________________0___18607), .Q (_________29693));
  xnr2s1 _______440427(.DIN1 (____9____31798), .DIN2 (_________29886),
       .Q (_________29692));
  nnd2s1 _____9_440428(.DIN1 (_____9___29707), .DIN2 (_________18845),
       .Q (_________29691));
  xor2s1 _______440429(.DIN1 (_____0___29620), .DIN2 (_________34700),
       .Q (______0__29690));
  nnd2s1 ______440430(.DIN1 (_____9___29705), .DIN2 (_________29688),
       .Q (______9__29689));
  and2s1 _____440431(.DIN1 (_________34690), .DIN2 (_________32410), .Q
       (_________29687));
  nnd2s1 _____9_440432(.DIN1 (_________29685), .DIN2 (_________29467),
       .Q (_________29686));
  xor2s1 _______440433(.DIN1 (_____0___29619), .DIN2 (_________29637),
       .Q (_____9___29703));
  nor2s1 _____440434(.DIN1 (_________29540), .DIN2 (______9__29643), .Q
       (_________29733));
  hi1s1 ______440435(.DIN (_________29683), .Q (_________29684));
  xor2s1 _____440436(.DIN1 (______0__34491), .DIN2 (______9__29679), .Q
       (_________29682));
  nor2s1 _______440437(.DIN1 (_________29603), .DIN2 (_________29638),
       .Q (_________29681));
  xor2s1 _______440438(.DIN1 (_________________18711), .DIN2
       (______9__29679), .Q (______0__29680));
  nnd2s1 _____440439(.DIN1 (_________29627), .DIN2 (outData[18]), .Q
       (_________29678));
  and2s1 _____0_440440(.DIN1 (_____9___29707), .DIN2 (_____9___29708),
       .Q (_________29677));
  hi1s1 _______440441(.DIN (_________29675), .Q (_________29676));
  nor2s1 _____9_440442(.DIN1 (_________29660), .DIN2 (_________29628),
       .Q (_________29674));
  nor2s1 ______440443(.DIN1 (_________29591), .DIN2 (______0__29634),
       .Q (______0__29719));
  nnd2s1 _______440444(.DIN1 (_________29632), .DIN2 (_________29635),
       .Q (_________29698));
  xnr2s1 _______440445(.DIN1 (____000__32751), .DIN2 (_____9___29613),
       .Q (_________29726));
  xor2s1 _______440446(.DIN1 (______9__29605), .DIN2 (_________31578),
       .Q (_________29673));
  nnd2s1 _______440447(.DIN1 (_____0___29618), .DIN2 (_________29584),
       .Q (_________29672));
  nor2s1 _______440448(.DIN1 (_________________18694), .DIN2
       (_________32956), .Q (______0__29671));
  and2s1 _______440449(.DIN1 (_________32956), .DIN2
       (_________________18694), .Q (______9__29670));
  nor2s1 _______440450(.DIN1 (_________29668), .DIN2 (_____09__29623),
       .Q (_________29669));
  or2s1 _______440451(.DIN1 (______0__33373), .DIN2 (_____99__29614),
       .Q (_________29667));
  nor2s1 ______440452(.DIN1 (_________________0___18660), .DIN2
       (_____00__29615), .Q (_________29666));
  and2s1 _______440453(.DIN1 (______9__29679), .DIN2 (______0__34491),
       .Q (_________29665));
  nor2s1 _______440454(.DIN1 (______0__34491), .DIN2 (______9__29679),
       .Q (_________29664));
  or2s1 _______440455(.DIN1 (____0____28156), .DIN2 (______9__29679),
       .Q (_________29663));
  nor2s1 _______440456(.DIN1 (______0__29662), .DIN2 (____9____33624),
       .Q (_____0___29713));
  and2s1 ______440457(.DIN1 (____9____33624), .DIN2 (______0__29662),
       .Q (_____0___29712));
  or2s1 ______440458(.DIN1 (_____0___29616), .DIN2 (_________29660), .Q
       (______9__29661));
  nor2s1 _______440459(.DIN1 (_________29646), .DIN2 (______9__29679),
       .Q (_________29659));
  nnd2s1 _______440460(.DIN1 (_____9___29609), .DIN2 (_____9___29607),
       .Q (_________29658));
  or2s1 _______440461(.DIN1 (_________29656), .DIN2 (_____9___29611),
       .Q (_________29657));
  nnd2s1 _____0_440462(.DIN1 (_________29626), .DIN2
       (_____________18897), .Q (_________29655));
  hi1s1 _______440463(.DIN (_____9___29705), .Q (_________29654));
  and2s1 _______440464(.DIN1 (______9__29651), .DIN2 (_________34494),
       .Q (_________29653));
  or2s1 _______440465(.DIN1 (_________34494), .DIN2 (______9__29651),
       .Q (______0__29652));
  nor2s1 ______440466(.DIN1 (_________29649), .DIN2 (_________34692),
       .Q (_________29650));
  or2s1 _______440467(.DIN1 (_________29647), .DIN2 (_________34692),
       .Q (_________29648));
  nnd2s1 _______440468(.DIN1 (______9__29679), .DIN2 (_________29646),
       .Q (_________29750));
  nor2s1 _______440469(.DIN1 (______0__18842), .DIN2 (_________29645),
       .Q (_________29724));
  nnd2s1 _______440470(.DIN1 (_____0___29617), .DIN2 (___0_____27408),
       .Q (_________29675));
  nnd2s1 _______440471(.DIN1 (_________29645), .DIN2 (______0__18842),
       .Q (_________29683));
  xor2s1 _______440472(.DIN1 (___0_____27419), .DIN2 (_________29639),
       .Q (_________29644));
  nor2s1 _______440473(.DIN1 (_____9__19991), .DIN2 (______9__29596),
       .Q (______9__29643));
  nor2s1 ______440474(.DIN1 (_________32410), .DIN2 (_________29593),
       .Q (_________29642));
  xor2s1 ______440475(.DIN1 (_________34694), .DIN2 (______0__30591),
       .Q (_________29641));
  xor2s1 _______440476(.DIN1 (_________34465), .DIN2 (_________29639),
       .Q (_________29640));
  nor2s1 _______440477(.DIN1 (_________29595), .DIN2 (_________29637),
       .Q (_________29638));
  nnd2s1 ______440478(.DIN1 (_________29600), .DIN2 (_________29397),
       .Q (_________29685));
  hi1s1 _______440479(.DIN (_________32956), .Q (_____9___29707));
  and2s1 ______440480(.DIN1 (_________29631), .DIN2 (_________29635),
       .Q (_________29636));
  nor2s1 _______440481(.DIN1 (______0__31456), .DIN2 (_________29590),
       .Q (______0__29634));
  nor2s1 _______440482(.DIN1 (_________29421), .DIN2 (_________29589),
       .Q (______9__29633));
  nnd2s1 ______440483(.DIN1 (_________29631), .DIN2
       (_______________18875), .Q (_________29632));
  nnd2s1 _______440484(.DIN1 (_____9___29610), .DIN2 (_________29629),
       .Q (_________29630));
  and2s1 _______440485(.DIN1 (_________29586), .DIN2 (______0__30283),
       .Q (_________29628));
  hi1s1 _______440486(.DIN (_________29626), .Q (_________29627));
  nnd2s1 _______440487(.DIN1 (______9__29588), .DIN2 (_________29478),
       .Q (_________29787));
  xor2s1 _______440488(.DIN1 (_________29573), .DIN2 (_________35066),
       .Q (_____9___29705));
  nor2s1 ______440489(.DIN1 (______0__29624), .DIN2 (______0__29580),
       .Q (_________29625));
  nnd2s1 _______440490(.DIN1 (_________29578), .DIN2 (___0_9__21648),
       .Q (_____09__29623));
  nor2s1 _______440491(.DIN1 (______18918), .DIN2 (_________29639), .Q
       (_____0___29622));
  xor2s1 _______440492(.DIN1 (_________29602), .DIN2 (_________35066),
       .Q (_____0___29621));
  xor2s1 _______440493(.DIN1 (_________28303), .DIN2 (______0__29562),
       .Q (_____0___29620));
  xor2s1 _______440494(.DIN1 (_________34484), .DIN2 (_____99__29445),
       .Q (_____0___29619));
  nnd2s1 _____9_440495(.DIN1 (_________34694), .DIN2 (_________29582),
       .Q (_____0___29618));
  nnd2s1 _______440496(.DIN1 (_________29639), .DIN2 (___0_____27420),
       .Q (_____0___29617));
  nor2s1 _______440497(.DIN1 (_________29656), .DIN2 (_____9___29612),
       .Q (______9__29728));
  nnd2s1 _______440498(.DIN1 (_________29581), .DIN2 (________19976),
       .Q (_________29886));
  xor2s1 _______440499(.DIN1 (___0_____27417), .DIN2 (______0__29597),
       .Q (_________32956));
  xor2s1 _______440500(.DIN1 (_________29388), .DIN2 (_________29599),
       .Q (____9____33624));
  and2s1 _______440501(.DIN1 (_____9___29608), .DIN2 (______0__30283),
       .Q (_____0___29616));
  xor2s1 _______440502(.DIN1 (_________29480), .DIN2 (_________29587),
       .Q (_____00__29615));
  xor2s1 _____440503(.DIN1 (_________29433), .DIN2 (______0__34698), .Q
       (_____99__29614));
  nnd2s1 _______440504(.DIN1 (_____9___29612), .DIN2 (_________29656),
       .Q (_____9___29613));
  hi1s1 _______440505(.DIN (_____9___29610), .Q (_____9___29611));
  nnd2s1 _______440506(.DIN1 (_________34696), .DIN2 (_________35110),
       .Q (_____9___29609));
  nor2s1 ______440507(.DIN1 (______0__30283), .DIN2 (_____9___29608),
       .Q (_________29660));
  hi1s1 _______440508(.DIN (_____90__29606), .Q (_________29645));
  nnd2s1 _______440509(.DIN1 (_________34696), .DIN2 (_____9___29607),
       .Q (_________29626));
  dffacs1 __________________440510(.CLRB (reset), .CLK (clk), .DIN
       (_________29577), .Q (_________34494));
  nb1s1 _______440511(.DIN (_____90__29606), .Q (______9__29679));
  nnd2s1 _______440512(.DIN1 (_________29604), .DIN2 (_________29555),
       .Q (______9__29605));
  nor2s1 _____9_440513(.DIN1 (_________34484), .DIN2 (_________29594),
       .Q (_________29603));
  nor2s1 _______440514(.DIN1 (_________34465), .DIN2 (______9__29570),
       .Q (_________29601));
  nnd2s1 _______440515(.DIN1 (_________29599), .DIN2 (_________29401),
       .Q (_________29600));
  nor2s1 ______440516(.DIN1 (___0_____27416), .DIN2 (______0__29597),
       .Q (_________29598));
  nor2s1 ______440517(.DIN1 (________22650), .DIN2 (_________29569), .Q
       (______9__29596));
  and2s1 _____9_440518(.DIN1 (_________29594), .DIN2 (_________34484),
       .Q (_________29595));
  nnd2s1 _____9_440519(.DIN1 (_________29602), .DIN2 (_________29592),
       .Q (_________29593));
  xor2s1 _______440520(.DIN1 (________19977), .DIN2 (_____9___33572),
       .Q (_________29734));
  nor2s1 _______440521(.DIN1 (_________34495), .DIN2 (_________34700),
       .Q (_________29591));
  and2s1 _______440522(.DIN1 (_________34700), .DIN2 (_________34495),
       .Q (_________29590));
  nor2s1 _____0_440523(.DIN1 (_________29398), .DIN2 (______0__34698),
       .Q (_________29589));
  nnd2s1 _______440524(.DIN1 (_________29587), .DIN2 (_________29479),
       .Q (______9__29588));
  xor2s1 _______440525(.DIN1 (______0__29571), .DIN2 (_________30678),
       .Q (_________29586));
  xor2s1 _____0_440526(.DIN1 (_________29550), .DIN2
       (______________________________________0_____________18891), .Q
       (_____90__29606));
  nnd2s1 _______440527(.DIN1 (______9__29561), .DIN2 (_________29585),
       .Q (_____9___29610));
  nor2s1 _____440528(.DIN1 (_________29574), .DIN2 (______0__28925), .Q
       (_________29647));
  nnd2s1 _______440529(.DIN1 (_________29565), .DIN2
       (_______________18874), .Q (_________29631));
  dffacs1 _____________9____440530(.CLRB (reset), .CLK (clk), .DIN
       (_________29568), .Q (_________9______18799));
  nnd2s1 _______440531(.DIN1 (_________34702), .DIN2 (_________29583),
       .Q (_________29584));
  or2s1 ______440532(.DIN1 (_________29583), .DIN2 (_________34702), .Q
       (_________29582));
  nnd2s1 _______440533(.DIN1 (_____9___33572), .DIN2 (_____0__19975),
       .Q (_________29581));
  hi1s1 _______440534(.DIN (______9__29579), .Q (______0__29580));
  nnd2s1 _______440535(.DIN1 (_________29554), .DIN2 (_________32639),
       .Q (_________29578));
  nnd2s1 _____0_440536(.DIN1 (_________29551), .DIN2 (_________34393),
       .Q (_________29577));
  hi1s1 _______440537(.DIN (_________29575), .Q (_________29576));
  nor2s1 _______440538(.DIN1 (_________29377), .DIN2 (_________29557),
       .Q (_____9___29612));
  xor2s1 _______440539(.DIN1 (_____09__29536), .DIN2
       (___________0___18872), .Q (_________29573));
  or2s1 _____0_440540(.DIN1 (______0__29571), .DIN2 (_________30678),
       .Q (_________29572));
  nnd2s1 ______440541(.DIN1 (_________30678), .DIN2 (______0__29571),
       .Q (_____9___29608));
  nnd2s1 _______440542(.DIN1 (_________29564), .DIN2 (____0____30075),
       .Q (_________29635));
  nnd2s1 ______440543(.DIN1 (_________29560), .DIN2
       (______________________________________0__________0__18892), .Q
       (_________29629));
  hi1s1 _______440544(.DIN (______9__29570), .Q (_________29639));
  dffacs1 _____________9____440545(.CLRB (reset), .CLK (clk), .DIN
       (______9__29553), .Q (_________9______18800));
  nor2s1 ______440546(.DIN1 (_________35002), .DIN2 (_____0___29535),
       .Q (_________29569));
  nnd2s1 _____0_440547(.DIN1 (_________29547), .DIN2 (_____0__20059),
       .Q (_________29568));
  xor2s1 ______440548(.DIN1 (____0____34548), .DIN2 (_________29495),
       .Q (_________29575));
  nnd2s1 _____9_440549(.DIN1 (_________29566), .DIN2 (_________29567),
       .Q (______9__29579));
  nnd2s1 ______440550(.DIN1 (_________29546), .DIN2 (_________29549),
       .Q (______0__29597));
  nnd2s1 ______440551(.DIN1 (______9__29544), .DIN2 (______9__29292),
       .Q (_________29599));
  nor2s1 _____9_440552(.DIN1 (_________29567), .DIN2 (_________29566),
       .Q (______0__29624));
  xor2s1 _______440553(.DIN1 (_____0___29533), .DIN2 (___0__18931), .Q
       (_________29604));
  dffacs1 __________________440554(.CLRB (reset), .CLK (clk), .DIN
       (_________29542), .QN (_________34484));
  hi1s1 _______440555(.DIN (_________29564), .Q (_________29565));
  xor2s1 ______440556(.DIN1 (______0__31211), .DIN2 (_________32427),
       .Q (_________29563));
  xor2s1 _______440557(.DIN1 (_________34495), .DIN2 (____0____30044),
       .Q (______0__29562));
  hi1s1 _____0_440558(.DIN (_________29560), .Q (______9__29561));
  xor2s1 _______440559(.DIN1 (_________29390), .DIN2 (_________29556),
       .Q (______9__29570));
  xor2s1 _______440560(.DIN1 (_____00__29532), .DIN2 (_________29468),
       .Q (_________29574));
  nnd2s1 _______440561(.DIN1 (_________29538), .DIN2 (_____0___29449),
       .Q (_________29587));
  xor2s1 _______440562(.DIN1 (_____9___29526), .DIN2 (____0____32807),
       .Q (_________29602));
  and2s1 _______440563(.DIN1 (_________29558), .DIN2 (_____99__29531),
       .Q (_________29559));
  nor2s1 _______440564(.DIN1 (_________29376), .DIN2 (_________29556),
       .Q (_________29557));
  xor2s1 _______440565(.DIN1 (________________18754), .DIN2
       (_________29498), .Q (_________29554));
  nnd2s1 _______440566(.DIN1 (_____9___29529), .DIN2 (________20542),
       .Q (______9__29553));
  xor2s1 _______440567(.DIN1 (_________29543), .DIN2 (_________29378),
       .Q (_____9___33572));
  nor2s1 _______440568(.DIN1 (_________29473), .DIN2 (_____90__29522),
       .Q (_________29552));
  xor2s1 ______440569(.DIN1 (______0__29537), .DIN2 (_____0___29450),
       .Q (_________29551));
  and2s1 ______440570(.DIN1 (______0__29545), .DIN2 (_________29549),
       .Q (_________29550));
  nnd2s1 _______440571(.DIN1 (_________29519), .DIN2 (______9__29374),
       .Q (_________29560));
  nnd2s1 _______440572(.DIN1 (_________29515), .DIN2 (_______19009), .Q
       (_________29564));
  nnd2s1 _______440573(.DIN1 (_________29548), .DIN2 (___0__18931), .Q
       (_____9___29607));
  nor2s1 _______440574(.DIN1 (_____9___29523), .DIN2 (_________29548),
       .Q (_________30678));
  dffacs1 ____0__________________(.CLRB (reset), .CLK (clk), .DIN
       (_____9___29524), .QN (____0________________18649));
  nnd2s1 _______440575(.DIN1 (______9__29501), .DIN2 (_________34071),
       .Q (_________29547));
  nnd2s1 _______440576(.DIN1 (______0__29545), .DIN2 (______9__30537),
       .Q (_________29546));
  nnd2s1 _______440577(.DIN1 (_________29543), .DIN2 (_____9___29351),
       .Q (______9__29544));
  nnd2s1 _______440578(.DIN1 (_________29499), .DIN2 (_________34365),
       .Q (_________29542));
  xor2s1 _______440579(.DIN1 (_____9__20584), .DIN2 (_________29541),
       .Q (_________29566));
  nnd2s1 ______440580(.DIN1 (_________29506), .DIN2 (_________29412),
       .Q (_________29555));
  nor2s1 _______440581(.DIN1 (____9___22716), .DIN2 (_________29539),
       .Q (_________29540));
  or2s1 _____0_440582(.DIN1 (_________29418), .DIN2 (______0__29537),
       .Q (_________29538));
  xor2s1 ______440583(.DIN1 (_________29389), .DIN2 (_________29518),
       .Q (_____09__29536));
  nnd2s1 _______440584(.DIN1 (_________29539), .DIN2 (______9__28887),
       .Q (_____0___29535));
  xor2s1 _______440585(.DIN1 (_________29514), .DIN2 (___0____22550),
       .Q (_________29656));
  nnd2s1 _______440586(.DIN1 (_________29505), .DIN2 (_________29413),
       .Q (_____0___29533));
  nor2s1 _____9_440587(.DIN1 (_________29469), .DIN2 (_____9___29525),
       .Q (_____00__29532));
  or2s1 _______440588(.DIN1 (_____9___29527), .DIN2 (_________31373),
       .Q (_____99__29531));
  or2s1 ______440589(.DIN1 (___0__0__27384), .DIN2 (_________31373), .Q
       (_____9___29530));
  nnd2s1 _____9_440590(.DIN1 (_________29482), .DIN2 (_________34071),
       .Q (_____9___29529));
  xor2s1 _______440591(.DIN1 (_________________18761), .DIN2
       (_________31020), .Q (_____9___29528));
  nnd2s1 _______440592(.DIN1 (_________31373), .DIN2 (_____9___29527),
       .Q (_________29558));
  nor2s1 _____9_440593(.DIN1 (_____9___29525), .DIN2 (_________29470),
       .Q (_____9___29526));
  or2s1 ____90_440594(.DIN1 (__90____26287), .DIN2 (_________29481), .Q
       (_____9___29524));
  nor2s1 ______440595(.DIN1 (_________29513), .DIN2 (_________29516),
       .Q (_____9___29523));
  nor2s1 _______440596(.DIN1 (______0__29466), .DIN2 (______9__29521),
       .Q (_____90__29522));
  nnd2s1 _______440597(.DIN1 (______9__29521), .DIN2 (_________29472),
       .Q (_________29520));
  nnd2s1 ______440598(.DIN1 (_________29518), .DIN2 (_________29373),
       .Q (_________29519));
  and2s1 ______440599(.DIN1 (_________29516), .DIN2 (________19288), .Q
       (_________29517));
  or2s1 _______440600(.DIN1 (________19452), .DIN2 (_________29514), .Q
       (_________29515));
  and2s1 _____9_440601(.DIN1 (_________29516), .DIN2 (_________29513),
       .Q (_________29548));
  nnd2s1 _____440602(.DIN1 (_________29488), .DIN2 (____09___30086), .Q
       (_________29549));
  nor2s1 _____440603(.DIN1 (_____9___29261), .DIN2 (_________29485), .Q
       (_________29556));
  dffacs1 __________________440604(.CLRB (reset), .CLK (clk), .DIN
       (_________29486), .Q (_________34495));
  hi1s1 _____0_440605(.DIN (______0__29512), .Q (______0__31211));
  nnd2s1 _______440606(.DIN1 (_________31020), .DIN2 (_________34492),
       .Q (______9__29511));
  xnr2s1 _______440607(.DIN1 (_________34023), .DIN2 (_____0___29453),
       .Q (_________29510));
  xor2s1 _______440608(.DIN1 (_________34492), .DIN2 (_________29508),
       .Q (_________29509));
  or2s1 _______440609(.DIN1 (_________34492), .DIN2 (_________31020),
       .Q (_________29507));
  hi1s1 _______440610(.DIN (_________29505), .Q (_________29506));
  nnd2s1 _____0_440611(.DIN1 (______0__29476), .DIN2 (inData[0]), .Q
       (_________29504));
  nnd2s1 _____0_440612(.DIN1 (______9__29475), .DIN2 (____09___29170),
       .Q (_________29543));
  nnd2s1 _____9_440613(.DIN1 (_________29487), .DIN2
       (_______________18875), .Q (______0__29545));
  hi1s1 _____0_440614(.DIN (_________29541), .Q (_________29539));
  or2s1 _____440615(.DIN1 (______0__29502), .DIN2 (_________31020), .Q
       (_________29503));
  xor2s1 _______440616(.DIN1 (_____0___29452), .DIN2 (_________29500),
       .Q (______9__29501));
  xor2s1 _______440617(.DIN1 (_____0___29447), .DIN2 (_________31252),
       .Q (_________29499));
  nor2s1 _______440618(.DIN1 (_________29483), .DIN2 (______9__29491),
       .Q (_________29498));
  xor2s1 _______440619(.DIN1 (_____00__29446), .DIN2 (_________30166),
       .Q (______0__29537));
  xor2s1 _______440620(.DIN1 (_____0___29268), .DIN2 (______0__29484),
       .Q (______0__29512));
  nor2s1 ______440621(.DIN1 (_________28257), .DIN2 (_________29508),
       .Q (_________29494));
  xor2s1 _______440622(.DIN1 (_____9___29444), .DIN2 (_________34444),
       .Q (_________29493));
  or2s1 ______440623(.DIN1 (_________________18761), .DIN2
       (_________29508), .Q (_________29492));
  and2s1 _______440624(.DIN1 (_________29508), .DIN2
       (_________________18761), .Q (_________29490));
  nnd2s1 _______440625(.DIN1 (_________29459), .DIN2 (___9____20635),
       .Q (_________29567));
  nnd2s1 _______440626(.DIN1 (_________29489), .DIN2 (_________29495),
       .Q (_____0___29534));
  xor2s1 _______440627(.DIN1 (_________________18709), .DIN2
       (_____9___29442), .Q (_________29505));
  xor2s1 _______440628(.DIN1 (____09___29171), .DIN2 (_________29474),
       .Q (_________29541));
  xor2s1 _______440629(.DIN1 (_________29434), .DIN2 (______0__30607),
       .Q (_________31373));
  hi1s1 _______440630(.DIN (_________29487), .Q (_________29488));
  nnd2s1 _______440631(.DIN1 (_____0___29448), .DIN2 (_________34365),
       .Q (_________29486));
  nor2s1 _______440632(.DIN1 (_________29252), .DIN2 (______0__29484),
       .Q (_________29485));
  xor2s1 _______440633(.DIN1 (_________29336), .DIN2 (_________29464),
       .Q (_________29482));
  nnd2s1 ____9__440634(.DIN1 (_____0___29451), .DIN2 (__9_____26942),
       .Q (_________29481));
  nnd2s1 _______440635(.DIN1 (_________29479), .DIN2 (_________29478),
       .Q (_________29480));
  xor2s1 ____9__440636(.DIN1 (_________29431), .DIN2 (______0__29851),
       .Q (_________29514));
  xnr2s1 _____9_440637(.DIN1 (____0____30044), .DIN2 (_________34714),
       .Q (_________29518));
  xnr2s1 _______440638(.DIN1 (____90___33582), .DIN2 (_________29435),
       .Q (_____9___29525));
  xor2s1 ____9__440639(.DIN1 (_________29432), .DIN2 (____009__31815),
       .Q (_________29516));
  hi1s1 ____9__440640(.DIN (_________29477), .Q (______9__29521));
  nor2s1 _______440641(.DIN1 (_____9___29439), .DIN2 (_________33186),
       .Q (______0__29476));
  nnd2s1 _______440642(.DIN1 (_________29474), .DIN2 (____09___29169),
       .Q (______9__29475));
  nor2s1 ______440643(.DIN1 (____9___24978), .DIN2 (_____9___29438), .Q
       (_________29487));
  xor2s1 _______440644(.DIN1 (___9____20636), .DIN2 (_________33459),
       .Q (_________29583));
  hi1s1 _______440645(.DIN (_________29508), .Q (_________31020));
  nor2s1 ____9__440646(.DIN1 (_________29472), .DIN2 (_________29471),
       .Q (_________29473));
  nor2s1 _______440647(.DIN1 (_________29469), .DIN2 (_________29468),
       .Q (_________29470));
  nnd2s1 ____9__440648(.DIN1 (_________29471), .DIN2 (______0__29466),
       .Q (_________29467));
  nor2s1 _______440649(.DIN1 (_____9___29441), .DIN2 (_________29594),
       .Q (_________29483));
  xor2s1 ____9__440650(.DIN1 (______9__29465), .DIN2 (_________32644),
       .Q (_________29477));
  nnd2s1 _______440651(.DIN1 (_________29464), .DIN2 (______0__29320),
       .Q (_________29497));
  nor2s1 _____9_440652(.DIN1 (_________31618), .DIN2 (______0__29429),
       .Q (_________29463));
  xor2s1 _______440653(.DIN1 (_________29405), .DIN2 (____9____30874),
       .Q (_________29462));
  hi1s1 _______440654(.DIN (_________29460), .Q (_________29461));
  nnd2s1 _______440655(.DIN1 (_________33459), .DIN2 (___9_0__20634),
       .Q (_________29459));
  nnd2s1 _______440656(.DIN1 (_____9___32380), .DIN2 (_________29457),
       .Q (_________29458));
  nor2s1 ______440657(.DIN1 (_____09__29455), .DIN2 (_____0___29454),
       .Q (______0__29456));
  nor2s1 _______440658(.DIN1 (_________29457), .DIN2 (_____9___32380),
       .Q (_____0___29453));
  xor2s1 _______440659(.DIN1 (_________29414), .DIN2 (_________28601),
       .Q (_________29489));
  nnd2s1 _______440660(.DIN1 (______9__29428), .DIN2 (___0_____28009),
       .Q (______9__31120));
  xor2s1 _____9_440661(.DIN1 (_________29409), .DIN2 (_____90__34718),
       .Q (_____0___29452));
  nnd2s1 ____9__440662(.DIN1 (_________29425), .DIN2 (__9__0__26854),
       .Q (_____0___29451));
  nnd2s1 ____9__440663(.DIN1 (______9__29419), .DIN2 (_____0___29449),
       .Q (_____0___29450));
  xor2s1 _______440664(.DIN1 (_________29400), .DIN2
       (________________18675), .Q (_____0___29448));
  xor2s1 _____9_440665(.DIN1 (_____09__29365), .DIN2
       (________________18688), .Q (_____0___29447));
  nor2s1 ____9__440666(.DIN1 (_________29399), .DIN2 (_________29422),
       .Q (_____00__29446));
  nor2s1 ______440667(.DIN1 (_________29193), .DIN2 (_________29424),
       .Q (______0__29484));
  nor2s1 ______440668(.DIN1 (_____9___29440), .DIN2 (_____99__29445),
       .Q (______9__29491));
  xor2s1 ____9__440669(.DIN1 (_________29395), .DIN2 (_____0___33866),
       .Q (_________29479));
  dffacs1 ____0__________________440670(.CLRB (reset), .CLK (clk), .DIN
       (_________29426), .Q (____0________________18646));
  xor2s1 _______440671(.DIN1 (_____9__24915), .DIN2 (_____90__29437),
       .Q (_________29508));
  xor2s1 _______440672(.DIN1 (____0____32835), .DIN2 (_________31060),
       .Q (_____9___29444));
  xor2s1 _____440673(.DIN1 (______0__31074), .DIN2 (_________29406), .Q
       (_____9___29443));
  xor2s1 ______440674(.DIN1 (___0_____28008), .DIN2 (____0____32835),
       .Q (_____9___29442));
  hi1s1 _______440675(.DIN (_____9___29440), .Q (_____9___29441));
  nnd2s1 _____9_440676(.DIN1 (___0____21680), .DIN2 (_________29417),
       .Q (_____9___29439));
  nor2s1 ______440677(.DIN1 (____0___24795), .DIN2 (_____90__29437), .Q
       (_____9___29438));
  hi1s1 _______440678(.DIN (_____9___32380), .Q (_____9___32383));
  nnd2s1 ______440679(.DIN1 (_________29411), .DIN2 (____990__29073),
       .Q (_________29474));
  xor2s1 _______440680(.DIN1 (_________29380), .DIN2 (___0_____27828),
       .Q (_________29460));
  xor2s1 _______440681(.DIN1 (_________29379), .DIN2 (_________29222),
       .Q (_________32882));
  nnd2s1 ____90_440682(.DIN1 (_________31252), .DIN2
       (________________18688), .Q (_________29436));
  nnd2s1 ____9__440683(.DIN1
       (______________________________________0__________0), .DIN2
       (_________9____), .Q (_________29435));
  xor2s1 _____9_440684(.DIN1 (_________29210), .DIN2 (_________29423),
       .Q (_________29434));
  xor2s1 ____9_440685(.DIN1 (______0__29420), .DIN2
       (________________18788), .Q (_________29433));
  nnd2s1 ____9__440686(.DIN1 (_________29393), .DIN2 (_____9__19418),
       .Q (_________29432));
  nnd2s1 ____99_440687(.DIN1 (_________29391), .DIN2 (_____0___29357),
       .Q (_________29431));
  nor2s1 ____9__440688(.DIN1 (_________9____), .DIN2
       (______________________________________0__________0), .Q
       (_________29469));
  nnd2s1 ____9__440689(.DIN1 (______0__29403), .DIN2 (_________29408),
       .Q (_________29464));
  hi1s1 ____9__440690(.DIN (______9__29465), .Q (_________29471));
  or2s1 _______440691(.DIN1 (_________34444), .DIN2 (____0____32835),
       .Q (_________29430));
  xor2s1 _______440692(.DIN1 (_________29382), .DIN2 (_________29367),
       .Q (______0__29429));
  or2s1 _______440693(.DIN1 (___0_____28007), .DIN2 (____0____32835),
       .Q (______9__29428));
  nnd2s1 _______440694(.DIN1 (____0____32835), .DIN2 (_________34444),
       .Q (_________29427));
  and2s1 _______440695(.DIN1 (____0____32835), .DIN2
       (_________________18693), .Q (_____09__29455));
  nnd2s1 _____9_440696(.DIN1 (_________29383), .DIN2 (_________29366),
       .Q (_____9___29440));
  nor2s1 _______440697(.DIN1 (_________________18693), .DIN2
       (____0____32835), .Q (_____0___29454));
  nnd2s1 ____0__440698(.DIN1 (______0__29375), .DIN2 (____90___28999),
       .Q (_________29426));
  nor2s1 ____00_440699(.DIN1 (___0_____27430), .DIN2 (_________29372),
       .Q (_________29425));
  nor2s1 ____90_440700(.DIN1 (_________29192), .DIN2 (_________29423),
       .Q (_________29424));
  and2s1 ____9__440701(.DIN1 (______0__29385), .DIN2
       (________________18675), .Q (_________29422));
  nor2s1 ____9__440702(.DIN1 (_____18906), .DIN2 (______0__29420), .Q
       (_________29421));
  hi1s1 ____9__440703(.DIN (_________29418), .Q (______9__29419));
  xor2s1 ____440704(.DIN1 (_________29392), .DIN2 (_________29873), .Q
       (______9__29465));
  xor2s1 _____440705(.DIN1 (_________34716), .DIN2 (____0_0__29156), .Q
       (_________33459));
  xor2s1 ____900(.DIN1 (_____0___29359), .DIN2 (_______________18876),
       .Q (_____9___32380));
  xor2s1 _______440706(.DIN1 (______0__29339), .DIN2 (____0__18997), .Q
       (_________29417));
  xor2s1 _______440707(.DIN1 (_________29415), .DIN2 (______9__33828),
       .Q (_________29416));
  xor2s1 _____9_440708(.DIN1 (_________29415), .DIN2 (_________29370),
       .Q (_________29414));
  hi1s1 ____90_440709(.DIN (_________29412), .Q (_________29413));
  nnd2s1 ____440710(.DIN1 (_________34716), .DIN2 (____090__29166), .Q
       (_________29411));
  nnd2s1 ____9__440711(.DIN1 (_________29408), .DIN2 (______9__29402),
       .Q (_________29409));
  or2s1 ____9_440712(.DIN1 (_________29406), .DIN2 (_________29404), .Q
       (_________29407));
  and2s1 ____9__440713(.DIN1 (_________29404), .DIN2 (_________29406),
       .Q (_________29405));
  nnd2s1 ____9__440714(.DIN1 (______9__29402), .DIN2 (_____90__34718),
       .Q (______0__29403));
  dffacs1 _____________9____440715(.CLRB (reset), .CLK (clk), .DIN
       (_____99__29355), .Q (_________9____));
  nor2s1 ____9__440716(.DIN1 (__9_____26546), .DIN2 (_____0___29361),
       .Q (_____90__29437));
  nnd2s1 ____0__440717(.DIN1 (_________30118), .DIN2 (_________29396),
       .Q (_________29401));
  nor2s1 ____9_440718(.DIN1 (_________29399), .DIN2 (______9__29384),
       .Q (_________29400));
  nor2s1 ____9_440719(.DIN1 (________________18788), .DIN2
       (______0__29394), .Q (_________29398));
  or2s1 ____0__440720(.DIN1 (_________29396), .DIN2 (_________30118),
       .Q (_________29397));
  nor2s1 ____9__440721(.DIN1 (________________18677), .DIN2
       (______0__29394), .Q (_________29395));
  or2s1 ____00_440722(.DIN1 (________19131), .DIN2 (_________29392), .Q
       (_________29393));
  nnd2s1 ____00_440723(.DIN1 (_____9___29354), .DIN2 (_____9___30624),
       .Q (_________29391));
  xor2s1 ____99_440724(.DIN1
       (______________________________________0_____________18891),
       .DIN2 (_________29389), .Q (_________29390));
  xor2s1 ____99_440725(.DIN1 (_________29396), .DIN2 (______9__30111),
       .Q (_________29388));
  nor2s1 ____99_440726(.DIN1 (________________18676), .DIN2
       (_____9___29353), .Q (_________29418));
  xor2s1 ____99_440727(.DIN1 (_________29334), .DIN2 (____00___31810),
       .Q (_____0___29449));
  nnd2s1 ____9_440728(.DIN1 (______0__29394), .DIN2
       (________________18677), .Q (_________29478));
  dffacs1 __________________440729(.CLRB (reset), .CLK (clk), .DIN
       (_____00__29356), .Q (________________18688));
  nor2s1 ____90_440730(.DIN1 (_________29386), .DIN2 (_________29340),
       .Q (_________29387));
  hi1s1 ____9__440731(.DIN (______9__29384), .Q (______0__29385));
  or2s1 ____9_440732(.DIN1 (_________29382), .DIN2 (_________29343), .Q
       (_________29383));
  xor2s1 ____9__440733(.DIN1 (_________18862), .DIN2 (_________30531),
       .Q (_________29381));
  xor2s1 ____9__440734(.DIN1 (_________34479), .DIN2 (_________30531),
       .Q (_________29380));
  xor2s1 ____9_440735(.DIN1 (_____0___29358), .DIN2 (_____9___29259),
       .Q (_________29379));
  nor2s1 ____9__440736(.DIN1 (____9____29048), .DIN2 (_________29347),
       .Q (_________29423));
  nnd2s1 ____9__440737(.DIN1 (_________29344), .DIN2 (___0__9__27829),
       .Q (_________29412));
  hi1s1 ____9_440738(.DIN (_________29404), .Q (______0__31074));
  xnr2s1 ____9__440739(.DIN1 (_____0___29360), .DIN2 (__9_____26826),
       .Q (____0____32835));
  nor2s1 ____440740(.DIN1 (_____9___29350), .DIN2 (_________29337), .Q
       (_________29378));
  and2s1 ____00_440741(.DIN1 (_________29389), .DIN2 (______9__30537),
       .Q (_________29377));
  nor2s1 ____440742(.DIN1 (______9__30537), .DIN2 (_________29389), .Q
       (_________29376));
  nor2s1 ____0__440743(.DIN1 (__9_9___26986), .DIN2 (_________29335),
       .Q (______0__29375));
  nnd2s1 ____0__440744(.DIN1 (_________29389), .DIN2
       (___________0___18872), .Q (______9__29374));
  or2s1 ____0__440745(.DIN1 (___________0___18872), .DIN2
       (_________29389), .Q (_________29373));
  nnd2s1 ____0__440746(.DIN1 (_________29331), .DIN2 (__9_____26406),
       .Q (_________29372));
  hi1s1 ____0_440747(.DIN (______0__29394), .Q (______0__29420));
  dffacs1 __________________440748(.CLRB (reset), .CLK (clk), .DIN
       (_________29341), .QN (_________18846));
  dffacs1 ____0__________________440749(.CLRB (reset), .CLK (clk), .DIN
       (_________29332), .QN (____0________________18592));
  and2s1 ____90_440750(.DIN1 (_________29368), .DIN2 (_________29370),
       .Q (_________29371));
  nor2s1 ____9__440751(.DIN1 (_________29370), .DIN2 (_________29368),
       .Q (_________29369));
  nnd2s1 ____9__440752(.DIN1 (_________29366), .DIN2 (_________29342),
       .Q (_________29367));
  xor2s1 ____9_440753(.DIN1 (________19479), .DIN2 (____9____32693), .Q
       (_____0___29364));
  nor2s1 ____9_440754(.DIN1 (_____0___29362), .DIN2 (_________30531),
       .Q (_____0___29363));
  nor2s1 ____9__440755(.DIN1 (__9_____26545), .DIN2 (_____0___29360),
       .Q (_____0___29361));
  xor2s1 ____9__440756(.DIN1 (____99___29078), .DIN2 (_________29346),
       .Q (_____0___29359));
  xor2s1 ____9__440757(.DIN1 (_________29313), .DIN2 (_____0___29272),
       .Q (_____0___31633));
  nnd2s1 ____9__440758(.DIN1 (_____0___29358), .DIN2 (_________29302),
       .Q (_________29410));
  or2s1 ____9__440759(.DIN1 (________________18787), .DIN2
       (_____90__29349), .Q (_________29408));
  xor2s1 ____9__440760(.DIN1 (_________29312), .DIN2 (____09___30086),
       .Q (_________29404));
  or2s1 ____0__440761(.DIN1 (_____9___30624), .DIN2 (_________29324),
       .Q (_____0___29357));
  nor2s1 ____9__440762(.DIN1 (_________________0___18660), .DIN2
       (_________29325), .Q (_____00__29356));
  nor2s1 ____9__440763(.DIN1 (_________________0___18660), .DIN2
       (______0__29329), .Q (_____99__29355));
  nnd2s1 ____0__440764(.DIN1 (_________29316), .DIN2 (________25612),
       .Q (_____9___29354));
  xor2s1 ____0__440765(.DIN1 (_________29333), .DIN2 (_________35050),
       .Q (_____9___29353));
  or2s1 ____0__440766(.DIN1 (______9__29319), .DIN2 (_____9___29350),
       .Q (_____9___29351));
  nnd2s1 ____9__440767(.DIN1 (_____90__29349), .DIN2
       (________________18787), .Q (______9__29402));
  nor2s1 ____0__440768(.DIN1 (___9_9), .DIN2 (_________29318), .Q
       (_________29392));
  and2s1 ____99_440769(.DIN1 (_____90__29349), .DIN2 (______9__29348),
       .Q (_________29399));
  nor2s1 ____99_440770(.DIN1 (______9__29348), .DIN2 (_____90__29349),
       .Q (______9__29384));
  xor2s1 ____0__440771(.DIN1 (_________29306), .DIN2 (_________29253),
       .Q (______0__29394));
  hi1s1 ____0__440772(.DIN (______9__30111), .Q (_________30118));
  nor2s1 ____9__440773(.DIN1 (____9_9__29046), .DIN2 (_________29346),
       .Q (_________29347));
  nor2s1 ____9__440774(.DIN1
       (_______________0_____________________18833), .DIN2
       (____9____32693), .Q (_________29345));
  nnd2s1 ____9__440775(.DIN1 (____9____32693), .DIN2 (___0_____27827),
       .Q (_________29344));
  hi1s1 ____9__440776(.DIN (_________29342), .Q (_________29343));
  or2s1 ____90_440777(.DIN1 (______9__30207), .DIN2 (_________29314),
       .Q (_________29341));
  xor2s1 ____9__440778(.DIN1 (______0__29293), .DIN2 (_________29287),
       .Q (_________29340));
  xor2s1 ____9__440779(.DIN1 (_________34447), .DIN2 (______0__18857),
       .Q (______0__29339));
  nnd2s1 ____9__440780(.DIN1 (_________29311), .DIN2 (_________29288),
       .Q (_____09__29365));
  hi1s1 ____9_440781(.DIN (_________29368), .Q (_________29415));
  xor2s1 ____99_440782(.DIN1 (_________34469), .DIN2 (_____9___32286),
       .Q (______9__29338));
  and2s1 ____0__440783(.DIN1 (_________29308), .DIN2 (_________34362),
       .Q (_________29337));
  xor2s1 ____0__440784(.DIN1 (_________34433), .DIN2 (_________29321),
       .Q (_________29336));
  nnd2s1 ____0__440785(.DIN1 (______9__29309), .DIN2 (__909___26330),
       .Q (_________29335));
  nnd2s1 ____0_440786(.DIN1 (_________29333), .DIN2
       (________________18676), .Q (_________29334));
  nnd2s1 ____0__440787(.DIN1 (_________29304), .DIN2 (___0_____27998),
       .Q (_________29332));
  nor2s1 ____0__440788(.DIN1 (__9_____27023), .DIN2 (_________29303),
       .Q (_________29331));
  xor2s1 ____0__440789(.DIN1 (_________29317), .DIN2 (_________29330),
       .Q (______9__30111));
  xor2s1 ____0__440790(.DIN1 (_________29323), .DIN2 (________26063),
       .Q (_________29389));
  xor2s1 ____0__440791(.DIN1 (_________29290), .DIN2 (______9__29255),
       .Q (______0__29329));
  nor2s1 ____9__440792(.DIN1 (_________29327), .DIN2 (______0__29301),
       .Q (_________29328));
  nnd2s1 ____9__440793(.DIN1 (_________29297), .DIN2 (_________29285),
       .Q (_____0___29358));
  nor2s1 ____9__440794(.DIN1 (___0_____27309), .DIN2 (_________29299),
       .Q (_____0___29360));
  or2s1 ____9__440795(.DIN1 (______0__18857), .DIN2 (_________29326),
       .Q (_________29366));
  nnd2s1 ____9__440796(.DIN1 (_________29326), .DIN2 (______0__18857),
       .Q (_________29342));
  xor2s1 ____9__440797(.DIN1 (_________29286), .DIN2 (_____0___28807),
       .Q (_________29368));
  hi1s1 ____9__440798(.DIN (____9____32693), .Q (_________30531));
  xor2s1 ____0__440799(.DIN1 (_________29278), .DIN2 (_________29234),
       .Q (_________29325));
  or2s1 ____0__440800(.DIN1 (________26062), .DIN2 (_________29323), .Q
       (_________29324));
  and2s1 ____0__440801(.DIN1 (_________29321), .DIN2 (_________34433),
       .Q (_________29322));
  or2s1 ____0_440802(.DIN1 (_________34433), .DIN2 (_________29321), .Q
       (______0__29320));
  and2s1 ____0__440803(.DIN1 (_________29315), .DIN2 (_________34362),
       .Q (______9__29319));
  and2s1 ____0__440804(.DIN1 (_________29317), .DIN2 (_____9__19233),
       .Q (_________29318));
  nnd2s1 ____0_440805(.DIN1 (_________29323), .DIN2 (________25613), .Q
       (_________29316));
  nor2s1 ____0__440806(.DIN1 (_________29305), .DIN2 (_________29294),
       .Q (_____9___29352));
  nor2s1 ____0_440807(.DIN1 (_________34362), .DIN2 (_________29315),
       .Q (_____9___29350));
  xor2s1 ____0__440808(.DIN1 (_________29281), .DIN2 (____99___29077),
       .Q (_____90__29349));
  nnd2s1 ____9_440809(.DIN1 (_________29289), .DIN2 (____9___23077), .Q
       (_________29314));
  xnr2s1 ____9_440810(.DIN1 (_________29284), .DIN2 (_________29296),
       .Q (_________29313));
  nor2s1 ____0__440811(.DIN1 (_____0___29269), .DIN2 (______0__29310),
       .Q (_________29312));
  nnd2s1 ____00_440812(.DIN1 (_____99__29445), .DIN2 (______0__29283),
       .Q (_________29311));
  nor2s1 ____0__440813(.DIN1 (_____0___29270), .DIN2 (______0__29310),
       .Q (_________29346));
  xnr2s1 ____440814(.DIN1 (_________29298), .DIN2 (___0_____27311), .Q
       (____9____32693));
  nnd2s1 _____0_440815(.DIN1 (_________29276), .DIN2 (__9_____27021),
       .Q (______9__29309));
  xor2s1 ____0__440816(.DIN1 (_________29291), .DIN2 (_________29307),
       .Q (_________29308));
  xor2s1 ____09_440817(.DIN1 (_____0___29267), .DIN2 (_________29305),
       .Q (_________29306));
  nor2s1 _____0_440818(.DIN1 (___0_0___27561), .DIN2 (_________29277),
       .Q (_________29304));
  nnd2s1 _____0_440819(.DIN1 (______9__29282), .DIN2 (_________34982),
       .Q (_________29303));
  hi1s1 ____0__440820(.DIN (_________29321), .Q (_________29333));
  xor2s1 ____0_440821(.DIN1 (_____9___29260), .DIN2 (_____0___30999),
       .Q (_________29302));
  hi1s1 ____00_440822(.DIN (______9__29300), .Q (______0__29301));
  nor2s1 ____00_440823(.DIN1 (___0_____27310), .DIN2 (_________29298),
       .Q (_________29299));
  nnd2s1 ____0__440824(.DIN1 (_____0___29273), .DIN2 (_________29296),
       .Q (_________29297));
  dffacs1 __________________440825(.CLRB (reset), .CLK (clk), .DIN
       (_____09__29274), .Q (______0__18857));
  xor2s1 ____440826(.DIN1 (_________29254), .DIN2 (______0__35098), .Q
       (_________29294));
  xor2s1 ____0__440827(.DIN1 (________________18687), .DIN2
       (_____99__29445), .Q (______0__29293));
  or2s1 ____0_440828(.DIN1 (_________29291), .DIN2 (_________29307), .Q
       (______9__29292));
  nnd2s1 ______440829(.DIN1 (_____0___29266), .DIN2 (_________29236),
       .Q (_________29317));
  nnd2s1 ____0__440830(.DIN1 (_________29307), .DIN2 (_________29291),
       .Q (_________29315));
  xor2s1 ______440831(.DIN1 (_________29245), .DIN2 (____9____29986),
       .Q (_________29323));
  xor2s1 _____440832(.DIN1 (_________29209), .DIN2 (_________29250), .Q
       (_________29321));
  xor2s1 ____0__440833(.DIN1
       (______________________________________0_____________18890),
       .DIN2 (_____9___34511), .Q (_____9___32286));
  xor2s1 ____09_440834(.DIN1 (_________29232), .DIN2 (_________34434),
       .Q (_________29290));
  nnd2s1 ____9__440835(.DIN1 (_____9___29262), .DIN2 (_________32925),
       .Q (_________29289));
  or2s1 ____0__440836(.DIN1 (________________18687), .DIN2
       (_________29287), .Q (_________29288));
  xor2s1 ____0__440837(.DIN1 (_____00__29265), .DIN2 (______0__29571),
       .Q (_________29286));
  nnd2s1 ____0__440838(.DIN1 (_____9___29258), .DIN2 (_________29284),
       .Q (_________29285));
  nnd2s1 ____0_440839(.DIN1 (_________29287), .DIN2
       (________________18687), .Q (______0__29283));
  xnr2s1 ____0__440840(.DIN1 (_________31983), .DIN2 (_________29237),
       .Q (______0__29310));
  nor2s1 ____0__440841(.DIN1 (_____________0___18759), .DIN2
       (_____9___30360), .Q (_________29327));
  nnd2s1 ____0__440842(.DIN1 (_____9___30360), .DIN2
       (_____________0___18759), .Q (______9__29300));
  nor2s1 _______440843(.DIN1 (___0_9___27848), .DIN2 (______9__29246),
       .Q (______9__29282));
  xor2s1 ____09_440844(.DIN1 (_________29231), .DIN2 (_________33144),
       .Q (_________29281));
  nnd2s1 ____09_440845(.DIN1 (______0__29275), .DIN2 (_________29233),
       .Q (_________29278));
  nnd2s1 _______440846(.DIN1 (______0__29247), .DIN2 (_____0___28337),
       .Q (_________29277));
  nor2s1 _______440847(.DIN1 (__9_____26597), .DIN2 (_________29249),
       .Q (_________29276));
  nnd2s1 ____09_440848(.DIN1 (______0__29275), .DIN2 (_________29235),
       .Q (______9__29348));
  dffacs1 ____0___________________(.CLRB (reset), .CLK (clk), .DIN
       (_________29248), .QN (____0_________________18659));
  nnd2s1 ____0_440849(.DIN1 (_________29243), .DIN2 (_____0___31454),
       .Q (_____09__29274));
  nnd2s1 ____0__440850(.DIN1 (_____0___29272), .DIN2 (____0____29095),
       .Q (_____0___29273));
  nnd2s1 ____0__440851(.DIN1 (_________29242), .DIN2 (_________34071),
       .Q (_____0___29271));
  nnd2s1 ____0_440852(.DIN1 (_________29244), .DIN2 (____0____29164),
       .Q (_________29296));
  nor2s1 ____0_440853(.DIN1 (__9_____26918), .DIN2 (_________29241), .Q
       (_________29298));
  hi1s1 ____0__440854(.DIN (_____9___30360), .Q (_____0___33031));
  nor2s1 ____0__440855(.DIN1 (_______________18875), .DIN2
       (_____0___29269), .Q (_____0___29270));
  xor2s1 _______440856(.DIN1 (_____0___29267), .DIN2 (_____9___30627),
       .Q (_____0___29268));
  or2s1 _______440857(.DIN1 (_________31667), .DIN2 (_____9___34720),
       .Q (_____0___29266));
  nor2s1 _______440858(.DIN1 (_________29189), .DIN2 (______0__29239),
       .Q (_________29305));
  or2s1 ____0__440859(.DIN1 (_________28779), .DIN2 (_____00__29265),
       .Q (_________29295));
  xnr2s1 _______440860(.DIN1 (_____99__29264), .DIN2 (_____9___29263),
       .Q (_________29307));
  xor2s1 ____0_440861(.DIN1 (_________29214), .DIN2 (_____9___34722),
       .Q (_____9___29262));
  nor2s1 _______440862(.DIN1 (_____9___30627), .DIN2 (_____0___29267),
       .Q (_____9___29261));
  nor2s1 ____0__440863(.DIN1 (_____9___29259), .DIN2 (_____90__29256),
       .Q (_____9___29260));
  hi1s1 ____0__440864(.DIN (_____0___29272), .Q (_____9___29258));
  and2s1 ____0__440865(.DIN1 (_____90__29256), .DIN2 (_____9___29259),
       .Q (_____9___29257));
  or2s1 ______440866(.DIN1 (_________29224), .DIN2 (______9__29255), .Q
       (_________29279));
  nnd2s1 _______440867(.DIN1 (_________29228), .DIN2
       (________________18674), .Q (______0__29275));
  dffacs1 __________________440868(.CLRB (reset), .CLK (clk), .DIN
       (_________29227), .QN (________________18687));
  xor2s1 ____0_440869(.DIN1 (___0_____27278), .DIN2 (_________29240),
       .Q (_____9___30360));
  and2s1 _______440870(.DIN1 (_____0___29267), .DIN2 (_________29253),
       .Q (_________29254));
  and2s1 _______440871(.DIN1 (_____0___29267), .DIN2 (_____9___30627),
       .Q (_________29252));
  or2s1 _______440872(.DIN1 (_________29253), .DIN2 (_____0___29267),
       .Q (_________29251));
  xnr2s1 _______440873(.DIN1
       (______________________________________0__________0), .DIN2
       (______9__29238), .Q (_________29250));
  nnd2s1 _______440874(.DIN1 (_________29217), .DIN2 (___00____27196),
       .Q (_________29249));
  nnd2s1 _______440875(.DIN1 (_________29218), .DIN2 (__99_9__27162),
       .Q (_________29248));
  and2s1 _______440876(.DIN1 (______0__29221), .DIN2 (________23130),
       .Q (______0__29247));
  nnd2s1 _______440877(.DIN1 (_________29219), .DIN2 (_____9__25634),
       .Q (______9__29246));
  nor2s1 _______440878(.DIN1 (_________29194), .DIN2 (______9__29220),
       .Q (_________29245));
  dffacs1 ______________________0_(.CLRB (reset), .CLK (clk), .DIN
       (_________29223), .QN (__________________0___18628));
  nnd2s1 ____0__440879(.DIN1 (______9__29211), .DIN2 (_____0___29184),
       .Q (_________29244));
  nor2s1 ____0__440880(.DIN1 (___0____20714), .DIN2 (_________29215),
       .Q (_________29243));
  xor2s1 ____0_440881(.DIN1 (_________29204), .DIN2 (____9____29007),
       .Q (_________29242));
  and2s1 ____0_440882(.DIN1 (_________29240), .DIN2 (___0_____27300),
       .Q (_________29241));
  xor2s1 ____09_440883(.DIN1 (______9__29202), .DIN2 (_____0___32570),
       .Q (_____00__29265));
  nor2s1 ____0__440884(.DIN1 (_________29213), .DIN2 (_________29216),
       .Q (____9____29981));
  xor2s1 ____09_440885(.DIN1 (_________29200), .DIN2 (_____0___29178),
       .Q (_____0___29272));
  nor2s1 ______440886(.DIN1 (______9__29238), .DIN2 (_________29198),
       .Q (______0__29239));
  nnd2s1 _____0_440887(.DIN1 (______9__29229), .DIN2 (______0__29230),
       .Q (_________29237));
  nnd2s1 _______440888(.DIN1 (_________29208), .DIN2 (_________31667),
       .Q (_________29236));
  nnd2s1 _______440889(.DIN1 (_________29234), .DIN2 (_________29233),
       .Q (_________29235));
  xor2s1 _______440890(.DIN1 (_________29225), .DIN2 (______0__31254),
       .Q (_________29232));
  xor2s1 _______440891(.DIN1 (_________29191), .DIN2 (____9____29052),
       .Q (_________29231));
  nor2s1 _____0_440892(.DIN1 (______0__29230), .DIN2 (______9__29229),
       .Q (_____0___29269));
  xor2s1 ____440893(.DIN1 (______0__29203), .DIN2 (____0____30981), .Q
       (_________29495));
  xor2s1 ______440894(.DIN1 (_________29206), .DIN2 (_________31505),
       .Q (_________29228));
  nor2s1 _____0_440895(.DIN1 (_________34187), .DIN2 (_________29201),
       .Q (_________29227));
  and2s1 _______440896(.DIN1 (_________29225), .DIN2 (_________34434),
       .Q (_________29226));
  nor2s1 _______440897(.DIN1 (_________34434), .DIN2 (_________29225),
       .Q (_________29224));
  nnd2s1 ______440898(.DIN1 (______0__29196), .DIN2 (__9_90__26504), .Q
       (_________29223));
  hi1s1 _______440899(.DIN (_________29222), .Q (_____90__29256));
  nor2s1 _____440900(.DIN1 (___0____24377), .DIN2 (_________29187), .Q
       (______0__29221));
  and2s1 _______440901(.DIN1 (______0__29186), .DIN2 (_________31951),
       .Q (______9__29220));
  nor2s1 _______440902(.DIN1 (__9_9___26511), .DIN2 (______9__29195),
       .Q (_________29219));
  and2s1 ______440903(.DIN1 (_________29190), .DIN2 (___090__25357), .Q
       (_________29218));
  nor2s1 _____9_440904(.DIN1 (______0__28751), .DIN2 (_________29188),
       .Q (_________29217));
  xnr2s1 _______440905(.DIN1 (______0__29662), .DIN2 (_________29207),
       .Q (_____9___29263));
  xor2s1 _______440906(.DIN1 (____09___29168), .DIN2 (____0____29150),
       .Q (_____0___29267));
  dffacs1 _____________________9_(.CLRB (reset), .CLK (clk), .DIN
       (_________29197), .QN (_________________9___18606));
  nor2s1 ____0__440907(.DIN1 (_____9___34722), .DIN2 (______0__29212),
       .Q (_________29216));
  and2s1 ____0__440908(.DIN1 (_____0___29183), .DIN2 (_________33186),
       .Q (_________29215));
  nor2s1 ____09_440909(.DIN1 (_________29213), .DIN2 (______0__29212),
       .Q (_________29214));
  xor2s1 _______440910(.DIN1 (____0____29162), .DIN2 (____0____31820),
       .Q (______9__29211));
  nnd2s1 ______440911(.DIN1 (_____0___29180), .DIN2 (_________29199),
       .Q (_________29222));
  xor2s1 _______440912(.DIN1 (____0____29159), .DIN2 (____0____30044),
       .Q (_________29240));
  xor2s1 ______440913(.DIN1 (_________29209), .DIN2 (_________34409),
       .Q (_________29210));
  nor2s1 _______440914(.DIN1 (___9____19713), .DIN2 (_________29207),
       .Q (_________29208));
  nnd2s1 _______440915(.DIN1 (____09___29173), .DIN2 (____0____29135),
       .Q (_________29234));
  or2s1 _______440916(.DIN1 (________________18674), .DIN2
       (_________29206), .Q (_________29233));
  nor2s1 _____0_440917(.DIN1 (____9____29051), .DIN2 (____099__29175),
       .Q (______9__29238));
  nnd2s1 _______440918(.DIN1 (____09___29167), .DIN2 (_________29205),
       .Q (______9__29229));
  xor2s1 _______440919(.DIN1 (____0____29143), .DIN2 (_________31153),
       .Q (_________29204));
  nnd2s1 _______440920(.DIN1 (____0____29157), .DIN2 (________20173),
       .Q (______0__29203));
  nnd2s1 ______440921(.DIN1 (____0____29160), .DIN2 (_________28778),
       .Q (______9__29202));
  xor2s1 _______440922(.DIN1 (____0____29139), .DIN2 (____09___29172),
       .Q (_________29201));
  and2s1 _______440923(.DIN1 (_____0___29179), .DIN2 (_________29199),
       .Q (_________29200));
  and2s1 _____9_440924(.DIN1 (_________29209), .DIN2
       (______________________________________0__________0), .Q
       (_________29198));
  nnd2s1 _____9_440925(.DIN1 (____0_9__29145), .DIN2 (__99____27136),
       .Q (_________29197));
  nor2s1 _____9_440926(.DIN1 (___0_____27381), .DIN2 (____0____29152),
       .Q (______0__29196));
  dffacs1 _______________________(.CLRB (reset), .CLK (clk), .DIN
       (____0____29158), .QN (_____________________18624));
  nnd2s1 ______440927(.DIN1 (____0____29147), .DIN2 (__9_____26875), .Q
       (______9__29195));
  nor2s1 ______440928(.DIN1 (_________31951), .DIN2 (____0____29151),
       .Q (_________29194));
  nor2s1 ______440929(.DIN1 (_____0___30458), .DIN2 (_________29209),
       .Q (_________29193));
  and2s1 _______440930(.DIN1 (_________29209), .DIN2 (_____0___30458),
       .Q (_________29192));
  xnr2s1 _______440931(.DIN1 (_____99__29264), .DIN2 (____09___29174),
       .Q (_________29191));
  nnd2s1 _______440932(.DIN1 (____0____29148), .DIN2 (_____9___28891),
       .Q (_________29190));
  nor2s1 _____9_440933(.DIN1
       (______________________________________0__________0), .DIN2
       (_________29209), .Q (_________29189));
  nnd2s1 _______440934(.DIN1 (____0_0__29146), .DIN2 (____9___25170),
       .Q (_________29188));
  nnd2s1 _______440935(.DIN1 (____0____29153), .DIN2 (___990__22526),
       .Q (_________29187));
  nnd2s1 _______440936(.DIN1 (____0____29144), .DIN2 (________25610),
       .Q (______0__29186));
  hi1s1 _____0_440937(.DIN (_________29206), .Q (_________29225));
  dffacs1 ________________0_440938(.CLRB (reset), .CLK (clk), .DIN
       (____0_9__29165), .QN (____________0___18686));
  xor2s1 _______440939(.DIN1 (_____0___29184), .DIN2 (____0____29163),
       .Q (_____09__29185));
  xor2s1 _______440940(.DIN1 (____0____29122), .DIN2 (_________35050),
       .Q (_____0___29183));
  xnr2s1 ______440941(.DIN1 (______0__30283), .DIN2 (_____0___29181),
       .Q (_____0___29182));
  nnd2s1 _______440942(.DIN1 (_____0___29179), .DIN2 (_____0___29178),
       .Q (_____0___29180));
  xor2s1 _______440943(.DIN1 (_____00__29176), .DIN2 (____9____32728),
       .Q (_____0___29177));
  xor2s1 _______440944(.DIN1 (____0_0__29128), .DIN2 (____099__30093),
       .Q (______0__29212));
  xor2s1 ______440945(.DIN1 (____09__20894), .DIN2 (_____0___29181), .Q
       (_____9___29259));
  nor2s1 _______440946(.DIN1 (____9____29053), .DIN2 (____09___29174),
       .Q (____099__29175));
  nnd2s1 _______440947(.DIN1 (____0____29134), .DIN2 (____09___29172),
       .Q (____09___29173));
  nnd2s1 _______440948(.DIN1 (____09___29170), .DIN2 (____09___29169),
       .Q (____09___29171));
  xor2s1 _______440949(.DIN1 (____0____29149), .DIN2 (______0__29851),
       .Q (____09___29168));
  nnd2s1 _______440950(.DIN1 (____0____29154), .DIN2 (_________30104),
       .Q (____09___29167));
  or2s1 _______440951(.DIN1 (____0____29132), .DIN2 (____0_9__29155),
       .Q (____090__29166));
  nnd2s1 _______440952(.DIN1 (____0____29136), .DIN2 (____0_0__29119),
       .Q (_________29207));
  xor2s1 _______440953(.DIN1 (____0____29114), .DIN2 (______0__29230),
       .Q (_________29206));
  nnd2s1 _____9_440954(.DIN1 (____0_9__29127), .DIN2 (___09____28126),
       .Q (____0_9__29165));
  nnd2s1 _______440955(.DIN1 (____0____29161), .DIN2 (____0____29163),
       .Q (____0____29164));
  nor2s1 _______440956(.DIN1 (____0____29163), .DIN2 (____0____29161),
       .Q (____0____29162));
  xor2s1 ______440957(.DIN1 (____0____29104), .DIN2 (_________33894),
       .Q (____0____29160));
  nnd2s1 _______440958(.DIN1 (____0____29126), .DIN2 (____00___29087),
       .Q (____0____29159));
  nnd2s1 _______440959(.DIN1 (____0____29120), .DIN2 (__9_99__27082),
       .Q (____0____29158));
  or2s1 _______440960(.DIN1 (____0___20893), .DIN2 (_____0___29181), .Q
       (____0____29157));
  nor2s1 _____440961(.DIN1 (____0_9__29155), .DIN2 (____0____29123), .Q
       (____0_0__29156));
  nor2s1 _____440962(.DIN1 (____9____29008), .DIN2 (____0____29131), .Q
       (______9__29255));
  nnd2s1 _______440963(.DIN1 (____0____29125), .DIN2 (_________28865),
       .Q (_________29205));
  nnd2s1 _______440964(.DIN1 (____9____29983), .DIN2 (___0_____28026),
       .Q (_________29199));
  nor2s1 _______440965(.DIN1 (________23331), .DIN2 (____0____29111),
       .Q (____0____29153));
  nor2s1 _______440966(.DIN1 (___0__9__27771), .DIN2 (____0____29115),
       .Q (____0____29152));
  or2s1 _____9_440967(.DIN1 (____0____29150), .DIN2 (____0____29149),
       .Q (____0____29151));
  nor2s1 _______440968(.DIN1 (___0_____27291), .DIN2 (____0____29110),
       .Q (____0____29148));
  nor2s1 _______440969(.DIN1 (________25963), .DIN2 (____0____29112),
       .Q (____0____29147));
  nor2s1 _______440970(.DIN1 (___0____25336), .DIN2 (____0____29113),
       .Q (____0_0__29146));
  nnd2s1 _______440971(.DIN1 (____0____29117), .DIN2 (__9_____26962),
       .Q (____0_9__29145));
  nnd2s1 ______440972(.DIN1 (____0____29149), .DIN2 (________25611), .Q
       (____0____29144));
  dffacs1 _____________9__0_(.CLRB (reset), .CLK (clk), .DIN
       (____0_9__29118), .QN (___________________________________));
  xor2s1 _______440973(.DIN1 (____0____29097), .DIN2 (_________29585),
       .Q (_________29209));
  dffacs1 _______________________440974(.CLRB (reset), .CLK (clk), .DIN
       (____0____29121), .QN (_____________________18623));
  dffacs1 _______________________440975(.CLRB (reset), .CLK (clk), .DIN
       (____0____29116), .QN (_____________________18604));
  xor2s1 ______440976(.DIN1 (_________18846), .DIN2 (____0_0__29138),
       .Q (____0____29143));
  xor2s1 _______440977(.DIN1 (________21399), .DIN2 (_____9___32650),
       .Q (____0____29141));
  xor2s1 ______440978(.DIN1 (____0____29106), .DIN2 (_____9___32650),
       .Q (____0____29140));
  xor2s1 ______440979(.DIN1 (________________18673), .DIN2
       (____0_0__29138), .Q (____0____29139));
  nnd2s1 _______440980(.DIN1 (____0_9__29137), .DIN2 (________19216),
       .Q (_____0___29179));
  nnd2s1 _______440981(.DIN1 (____0____29096), .DIN2 (_________33204),
       .Q (____0____29136));
  or2s1 _______440982(.DIN1 (________________18673), .DIN2
       (____0____29133), .Q (____0____29135));
  nnd2s1 _______440983(.DIN1 (____0____29133), .DIN2
       (________________18673), .Q (____0____29134));
  nor2s1 _______440984(.DIN1 (_________________0___18633), .DIN2
       (____0____29094), .Q (____0____29132));
  nnd2s1 _______440985(.DIN1 (____0____29124), .DIN2 (_________28911),
       .Q (____0____29154));
  xor2s1 ______440986(.DIN1 (____9____29069), .DIN2 (____0_9__30961),
       .Q (____09___29170));
  nor2s1 _______440987(.DIN1 (_________28940), .DIN2 (____0_0__29101),
       .Q (____09___29174));
  nor2s1 _______440988(.DIN1 (____9____29034), .DIN2 (____0_0__29138),
       .Q (____0____29131));
  nnd2s1 _____9_440989(.DIN1 (_____9___32650), .DIN2 (_________18861),
       .Q (____0____29130));
  nor2s1 _____9_440990(.DIN1 (_________18861), .DIN2 (_____9___32650),
       .Q (____0____29129));
  nor2s1 _______440991(.DIN1 (___0_____28015), .DIN2 (____00___29090),
       .Q (____0_0__29128));
  or2s1 ______440992(.DIN1 (_________32158), .DIN2 (____99___29081), .Q
       (____0_9__29127));
  nnd2s1 _____0_440993(.DIN1 (____009__29091), .DIN2 (_________35086),
       .Q (____0____29126));
  hi1s1 _______440994(.DIN (____0____29124), .Q (____0____29125));
  nor2s1 _______440995(.DIN1 (_________________0___18633), .DIN2
       (____000__29083), .Q (____0____29123));
  xor2s1 _______440996(.DIN1 (____9____29060), .DIN2 (_____9___28989),
       .Q (____0____29122));
  xor2s1 _______440997(.DIN1 (____9____29061), .DIN2 (_________30496),
       .Q (_____00__29176));
  xor2s1 _______440998(.DIN1 (____9_9__29054), .DIN2 (_________33204),
       .Q (____09___29169));
  hi1s1 _____0_440999(.DIN (____0_9__29137), .Q (____9____29983));
  nor2s1 _____0_441000(.DIN1 (_________28764), .DIN2 (____00___29086),
       .Q (____0____29163));
  xnr2s1 _______441001(.DIN1 (____0____29103), .DIN2 (_________28835),
       .Q (_____0___29181));
  nnd2s1 _______441002(.DIN1 (____99___29075), .DIN2 (__9__9__26882),
       .Q (____0____29121));
  and2s1 _______441003(.DIN1 (____99___29074), .DIN2 (__9__9__27063),
       .Q (____0____29120));
  nnd2s1 _______441004(.DIN1 (____00___29084), .DIN2 (__9_00__26989),
       .Q (____0_0__29119));
  nnd2s1 ______441005(.DIN1 (____99___29080), .DIN2 (_________35042),
       .Q (____0_9__29118));
  nnd2s1 _______441006(.DIN1 (____0_0__29092), .DIN2 (___9____25208),
       .Q (____0____29117));
  nnd2s1 _______441007(.DIN1 (____99___29076), .DIN2 (___0_____27485),
       .Q (____0____29116));
  nnd2s1 _______441008(.DIN1 (____99___29079), .DIN2 (__99____27091),
       .Q (____0____29115));
  xor2s1 _____0_441009(.DIN1 (____0_9__29100), .DIN2 (_________28939),
       .Q (____0____29114));
  nnd2s1 _______441010(.DIN1 (____9____29062), .DIN2 (________25798),
       .Q (____0____29113));
  nnd2s1 _______441011(.DIN1 (____9____29066), .DIN2 (________22969),
       .Q (____0____29112));
  nnd2s1 _______441012(.DIN1 (____9_9__29063), .DIN2 (___0__0__27802),
       .Q (____0____29111));
  nnd2s1 _______441013(.DIN1 (_____9___34724), .DIN2 (__9_9___26507),
       .Q (____0____29110));
  nor2s1 _______441014(.DIN1 (_________35106), .DIN2 (____0____29093),
       .Q (____0_9__29155));
  nnd2s1 _______441015(.DIN1 (____9____29065), .DIN2 (__900___26253),
       .Q (____0____29149));
  xor2s1 _______441016(.DIN1 (____0____29108), .DIN2 (____9____29056),
       .Q (____0_9__29109));
  nnd2s1 _____441017(.DIN1 (____0____29102), .DIN2 (____0____29106), .Q
       (____0____29107));
  nor2s1 _______441018(.DIN1 (_________28693), .DIN2 (____0____29103),
       .Q (____0____29104));
  nor2s1 _______441019(.DIN1 (___0_____28016), .DIN2 (____00___29089),
       .Q (_________29213));
  nor2s1 _______441020(.DIN1 (____0____29106), .DIN2 (____0____29102),
       .Q (____0____29142));
  xor2s1 _______441021(.DIN1 (____9____29033), .DIN2 (____0____31831),
       .Q (_____0___29184));
  xor2s1 ______441022(.DIN1 (_____9___34726), .DIN2 (_____0___31450),
       .Q (____0____29124));
  xor2s1 _______441023(.DIN1 (____9____29035), .DIN2 (_________28549),
       .Q (____0_9__29137));
  nor2s1 _______441024(.DIN1 (_________28938), .DIN2 (____0_9__29100),
       .Q (____0_0__29101));
  nnd2s1 ______441025(.DIN1 (____0____29098), .DIN2 (____9____29059),
       .Q (____0____29099));
  xor2s1 _______441026(.DIN1 (____9_0__29064), .DIN2 (_________29253),
       .Q (____0____29097));
  nnd2s1 ______441027(.DIN1 (____9____29050), .DIN2 (_________28963),
       .Q (____0____29096));
  hi1s1 _______441028(.DIN (_________29284), .Q (____0____29095));
  hi1s1 _______441029(.DIN (____0____29093), .Q (____0____29094));
  hi1s1 _______441030(.DIN (____0_0__29138), .Q (____0____29133));
  dffacs1 ____0________________0_(.CLRB (reset), .CLK (clk), .DIN
       (____9____29043), .Q (____0____________0___18645));
  dffacs1 ____0___________________441031(.CLRB (reset), .CLK (clk),
       .DIN (____9____29045), .QN (____0_________________18656));
  dffacs1 ____0__________________441032(.CLRB (reset), .CLK (clk), .DIN
       (____9____29044), .QN (____0________________18653));
  nor2s1 ______441033(.DIN1 (________23729), .DIN2 (____9_9__29018), .Q
       (____0_0__29092));
  nnd2s1 _______441034(.DIN1 (____9____29040), .DIN2 (________25408),
       .Q (____009__29091));
  hi1s1 _____0_441035(.DIN (____00___29089), .Q (____00___29090));
  nnd2s1 _______441036(.DIN1 (____9____29036), .DIN2 (_________33442),
       .Q (____00___29088));
  or2s1 _______441037(.DIN1 (_________35086), .DIN2 (____9____29039),
       .Q (____00___29087));
  nor2s1 _______441038(.DIN1 (_________29280), .DIN2 (____9_9__29037),
       .Q (____00___29086));
  nnd2s1 ______441039(.DIN1 (____9____29030), .DIN2 (inData[16]), .Q
       (____00___29085));
  nnd2s1 _____441040(.DIN1 (____9_9__29028), .DIN2 (_________28971), .Q
       (____00___29084));
  xor2s1 _____9_441041(.DIN1 (____999__29082), .DIN2 (____9_9__29072),
       .Q (____000__29083));
  xor2s1 _____9_441042(.DIN1 (____9____29014), .DIN2 (____9_0__29019),
       .Q (____99___29081));
  nnd2s1 _____0_441043(.DIN1 (____9____29026), .DIN2 (_________34071),
       .Q (____99___29080));
  nor2s1 _____0_441044(.DIN1 (__9__9__26757), .DIN2 (____9_0__29029),
       .Q (____99___29079));
  nor2s1 _______441045(.DIN1 (____9____29041), .DIN2 (____9____29032),
       .Q (_________29284));
  xor2s1 _____0_441046(.DIN1 (____9_0__29002), .DIN2 (_________28866),
       .Q (____0_0__29138));
  hi1s1 _______441047(.DIN (____0____29102), .Q (_____9___32650));
  xor2s1 _______441048(.DIN1 (____99___29077), .DIN2 (_________31431),
       .Q (____99___29078));
  nor2s1 _______441049(.DIN1 (__90____26316), .DIN2 (____9____29023),
       .Q (____99___29076));
  nor2s1 _______441050(.DIN1 (__9_9___27078), .DIN2 (____9____29024),
       .Q (____99___29075));
  nnd2s1 ______441051(.DIN1 (____9____29027), .DIN2 (_________35010),
       .Q (____99___29074));
  or2s1 _______441052(.DIN1 (____9_9__29072), .DIN2 (____9____29071),
       .Q (____990__29073));
  or2s1 _______441053(.DIN1 (_________18856), .DIN2 (____9____29067),
       .Q (____9____29070));
  nnd2s1 _______441054(.DIN1 (____9____29942), .DIN2 (_________28641),
       .Q (____9____29069));
  nnd2s1 _______441055(.DIN1 (____9____29067), .DIN2 (_________18856),
       .Q (____9____29068));
  nor2s1 _______441056(.DIN1 (________25027), .DIN2 (____9____29021),
       .Q (____9____29066));
  or2s1 _______441057(.DIN1 (__900___26252), .DIN2 (____9_0__29064), .Q
       (____9____29065));
  nor2s1 _______441058(.DIN1 (___09____28117), .DIN2 (____9____29022),
       .Q (____9_9__29063));
  nor2s1 _______441059(.DIN1 (_________28775), .DIN2 (____9____29016),
       .Q (____9____29062));
  nnd2s1 ______441060(.DIN1 (____9____29020), .DIN2 (____9____29013),
       .Q (____09___29172));
  nnd2s1 _______441061(.DIN1 (____9____29071), .DIN2 (____9_9__29072),
       .Q (____0____29093));
  dffacs1 _______________________441062(.CLRB (reset), .CLK (clk), .DIN
       (____9____29017), .QN (_____________________18611));
  xor2s1 _____441063(.DIN1 (________________18736), .DIN2
       (_____9___28984), .Q (____9____29061));
  nor2s1 ______441064(.DIN1 (_____9___28988), .DIN2 (____9_0__29055),
       .Q (____9____29060));
  and2s1 _______441065(.DIN1 (____9____29009), .DIN2 (inData[14]), .Q
       (____9____29059));
  and2s1 _____9_441066(.DIN1 (____9____29057), .DIN2 (____9____29056),
       .Q (____9____29058));
  nor2s1 _____441067(.DIN1 (____9____29056), .DIN2 (____9____29057), .Q
       (____0____29105));
  nor2s1 _____0_441068(.DIN1 (_________28550), .DIN2 (____9_9__29011),
       .Q (____0____29103));
  nor2s1 ______441069(.DIN1 (_____9___28990), .DIN2 (____9_0__29055),
       .Q (____0____30933));
  xor2s1 _______441070(.DIN1 (_____99__28991), .DIN2 (_________28930),
       .Q (____00___29089));
  xor2s1 _______441071(.DIN1 (____9_0__29038), .DIN2 (_____0___34730),
       .Q (____0____29102));
  xor2s1 _____0_441072(.DIN1 (____9____29031), .DIN2 (_________28979),
       .Q (____0____29161));
  nnd2s1 _______441073(.DIN1 (____9____29938), .DIN2 (____0____28175),
       .Q (____9_9__29054));
  nor2s1 ______441074(.DIN1 (____9____29052), .DIN2 (____99___29077),
       .Q (____9____29053));
  and2s1 ______441075(.DIN1 (____99___29077), .DIN2 (____9____29052),
       .Q (____9____29051));
  nnd2s1 ______441076(.DIN1 (____90___28998), .DIN2 (outData[15]), .Q
       (____9____29050));
  and2s1 ______441077(.DIN1 (____99___29077), .DIN2 (____9_0__29047),
       .Q (____9____29048));
  nor2s1 _____441078(.DIN1 (____9_0__29047), .DIN2 (____99___29077), .Q
       (____9_9__29046));
  nnd2s1 _______441079(.DIN1 (____909__29001), .DIN2 (_________28942),
       .Q (____9____29045));
  nnd2s1 ______441080(.DIN1 (____90___29000), .DIN2 (____9____29042),
       .Q (____9____29044));
  nnd2s1 ______441081(.DIN1 (____90___28995), .DIN2 (____9____29042),
       .Q (____9____29043));
  nor2s1 _______441082(.DIN1 (_________28855), .DIN2 (____90___28996),
       .Q (____0_9__29100));
  nnd2s1 _______441083(.DIN1 (_________28947), .DIN2 (_________28980),
       .Q (____9____29041));
  or2s1 _______441084(.DIN1 (________25409), .DIN2 (_____0___34730), .Q
       (____9____29040));
  nnd2s1 _____441085(.DIN1 (_____0___34730), .DIN2 (____9_0__29038), .Q
       (____9____29039));
  nnd2s1 _____9_441086(.DIN1 (_____9___28987), .DIN2 (______0__28850),
       .Q (____9_9__29037));
  xor2s1 _____9_441087(.DIN1 (______9__28954), .DIN2 (____9____29003),
       .Q (____9____29036));
  xor2s1 _____0_441088(.DIN1 (____9____29010), .DIN2 (_________29396),
       .Q (____9____29035));
  nor2s1 _______441089(.DIN1 (_________18846), .DIN2 (____9____29025),
       .Q (____9____29034));
  nnd2s1 _______441090(.DIN1 (____900__28992), .DIN2 (_________28932),
       .Q (____9____29033));
  and2s1 _______441091(.DIN1 (____9____29031), .DIN2 (_____9__21392),
       .Q (____9____29032));
  and2s1 _______441092(.DIN1 (_________31261), .DIN2 (_________28981),
       .Q (____9____29030));
  nnd2s1 _______441093(.DIN1 (_________28970), .DIN2 (______0__28974),
       .Q (____9_0__29029));
  nnd2s1 _______441094(.DIN1 (____90___28997), .DIN2 (outData[15]), .Q
       (____9_9__29028));
  nor2s1 _______441095(.DIN1 (__9_0___26897), .DIN2 (______9__28973),
       .Q (____9____29027));
  hi1s1 ______441096(.DIN (____9____29057), .Q (____0____29108));
  or2s1 _____9_441097(.DIN1 (_________28950), .DIN2 (____9____29025),
       .Q (____9____29026));
  nor2s1 _______441098(.DIN1 (__9_____26743), .DIN2 (_________28975),
       .Q (____9____29024));
  nnd2s1 _______441099(.DIN1 (______9__28964), .DIN2 (__9_____26577),
       .Q (____9____29023));
  nnd2s1 _______441100(.DIN1 (_________28957), .DIN2 (___0_____27800),
       .Q (____9____29022));
  nnd2s1 ______441101(.DIN1 (_________28959), .DIN2 (________22698), .Q
       (____9____29021));
  or2s1 _______441102(.DIN1 (____9_0__29019), .DIN2 (_________28966),
       .Q (____9____29020));
  nnd2s1 _______441103(.DIN1 (_____9___28985), .DIN2 (________23219),
       .Q (____9_9__29018));
  nnd2s1 _______441104(.DIN1 (_________28972), .DIN2 (_________28832),
       .Q (____9____29017));
  nnd2s1 _______441105(.DIN1 (_________28960), .DIN2 (___0_09__27665),
       .Q (____9____29016));
  nor2s1 _______441106(.DIN1 (_____9__25615), .DIN2 (_________28968),
       .Q (____9_0__29064));
  xor2s1 _____0_441107(.DIN1 (____9____29015), .DIN2 (_________35094),
       .Q (____9____29067));
  hi1s1 ______441108(.DIN (____999__29082), .Q (____9____29071));
  hi1s1 _______441109(.DIN (____9____29938), .Q (____9____29942));
  dffacs1 ________________________(.CLRB (reset), .CLK (clk), .DIN
       (_________28969), .QN (______________________18630));
  and2s1 _____441110(.DIN1 (____9____29013), .DIN2 (______0__28965), .Q
       (____9____29014));
  nor2s1 _______441111(.DIN1 (_________28577), .DIN2 (____9____29010),
       .Q (____9_9__29011));
  nnd2s1 _______441112(.DIN1 (_________28952), .DIN2 (_____0___28904),
       .Q (____9____29009));
  nor2s1 _______441113(.DIN1 (________19191), .DIN2 (____9____29007),
       .Q (____9____29008));
  and2s1 _______441114(.DIN1 (____9____29005), .DIN2 (____9____29004),
       .Q (____9____29006));
  nor2s1 _____0_441115(.DIN1 (____9____29003), .DIN2 (_________28949),
       .Q (____9____29049));
  xnr2s1 _____9_441116(.DIN1 (____0____31831), .DIN2 (_________28928),
       .Q (____9_0__29055));
  xor2s1 _______441117(.DIN1 (_________28978), .DIN2 (_____9___28701),
       .Q (____9____29057));
  xor2s1 _____0_441118(.DIN1 (_________28912), .DIN2 (_________29500),
       .Q (____9_0__29002));
  nor2s1 _______441119(.DIN1 (________26104), .DIN2 (_________28936),
       .Q (____909__29001));
  and2s1 _______441120(.DIN1 (______9__28934), .DIN2 (____90___28999),
       .Q (____90___29000));
  hi1s1 ______441121(.DIN (____90___28997), .Q (____90___28998));
  nor2s1 _______441122(.DIN1 (_________28910), .DIN2 (_________28941),
       .Q (____90___28996));
  nor2s1 _______441123(.DIN1 (____00__26047), .DIN2 (______0__28935),
       .Q (____90___28995));
  xor2s1 _____0_441124(.DIN1 (____90___28994), .DIN2 (____90___28993),
       .Q (____999__29082));
  xor2s1 _____441125(.DIN1 (________19443), .DIN2 (_____0___34732), .Q
       (____9____29938));
  dffacs1 ____0___________________441126(.CLRB (reset), .CLK (clk),
       .DIN (_________28943), .QN (____0_________________18658));
  xor2s1 _______441127(.DIN1 (_________28967), .DIN2 (__9_00__26514),
       .Q (____99___29077));
  nnd2s1 _____9_441128(.DIN1 (_________28929), .DIN2 (_____0___34734),
       .Q (____900__28992));
  xor2s1 _____0_441129(.DIN1 (_____0___28901), .DIN2 (_________28931),
       .Q (_____99__28991));
  nor2s1 _______441130(.DIN1 (_____9___28989), .DIN2 (_____9___28988),
       .Q (_____9___28990));
  nor2s1 _______441131(.DIN1 (_____0__21130), .DIN2 (_________28926),
       .Q (_____9___28987));
  xor2s1 _______441132(.DIN1 (____0___22719), .DIN2 (____99___32749),
       .Q (_____9___28986));
  nor2s1 _______441133(.DIN1 (__9_0___26427), .DIN2 (_________28922),
       .Q (_____9___28985));
  xor2s1 _____441134(.DIN1 (________25959), .DIN2 (_____90__28983), .Q
       (_____9___28984));
  nnd2s1 _______441135(.DIN1 (_________28923), .DIN2 (_________33279),
       .Q (______9__28982));
  xor2s1 _______441136(.DIN1 (_________________18749), .DIN2
       (_________28951), .Q (_________28981));
  or2s1 _____9_441137(.DIN1 (_________28979), .DIN2 (_________28976),
       .Q (_________28980));
  xnr2s1 _____9_441138(.DIN1 (________________18722), .DIN2
       (_____90__28983), .Q (_________28977));
  nor2s1 _______441139(.DIN1 (________25960), .DIN2 (_________28924),
       .Q (____09___30992));
  hi1s1 _______441140(.DIN (____9____29007), .Q (____9____29025));
  nor2s1 _____0_441141(.DIN1 (_________28976), .DIN2 (_________28946),
       .Q (____9____29031));
  nnd2s1 _______441142(.DIN1 (_________28918), .DIN2 (______0__28974),
       .Q (_________28975));
  nnd2s1 _______441143(.DIN1 (______0__28917), .DIN2 (________25734),
       .Q (______9__28973));
  nor2s1 _______441144(.DIN1 (_________28461), .DIN2 (______9__28916),
       .Q (_________28972));
  or2s1 _______441145(.DIN1 (outData[13]), .DIN2 (_____0___34732), .Q
       (_________28971));
  nor2s1 _______441146(.DIN1 (______0__28551), .DIN2 (_________28927),
       .Q (_________28970));
  nnd2s1 ______441147(.DIN1 (_________28915), .DIN2 (___00_9__27217),
       .Q (_________28969));
  nor2s1 ______441148(.DIN1 (________25614), .DIN2 (_________28967), .Q
       (_________28968));
  hi1s1 _______441149(.DIN (______0__28965), .Q (_________28966));
  nnd2s1 _______441150(.DIN1 (_________28913), .DIN2 (________21886),
       .Q (______9__28964));
  nnd2s1 _______441151(.DIN1 (_____0___34732), .DIN2 (_____0___29715),
       .Q (_________28963));
  xnr2s1 ______441152(.DIN1 (_____________9___18751), .DIN2
       (_________32029), .Q (_________28962));
  xnr2s1 ______441153(.DIN1 (_________34448), .DIN2 (_________32029),
       .Q (_________28961));
  nor2s1 ______441154(.DIN1 (___0_9___27748), .DIN2 (_________28908),
       .Q (_________28960));
  nor2s1 _______441155(.DIN1 (________24642), .DIN2 (_________28909),
       .Q (_________28959));
  nor2s1 _______441156(.DIN1 (__9_9___26698), .DIN2 (_____09__28906),
       .Q (_________28958));
  and2s1 ______441157(.DIN1 (_________28914), .DIN2 (___0__0__27792),
       .Q (_________28957));
  nnd2s1 _______441158(.DIN1 (_____0___34732), .DIN2 (outData[13]), .Q
       (____90___28997));
  nnd2s1 ______441159(.DIN1 (_________28948), .DIN2 (_________28953),
       .Q (_________28956));
  nnd2s1 _______441160(.DIN1 (____99___32749), .DIN2 (___0_____27790),
       .Q (______0__28955));
  xor2s1 _____9_441161(.DIN1 (_____0___28900), .DIN2 (_________28953),
       .Q (______9__28954));
  or2s1 _______441162(.DIN1 (_________________18749), .DIN2
       (_________28951), .Q (_________28952));
  nor2s1 _______441163(.DIN1 (____________0___18786), .DIN2
       (______0__28945), .Q (_________28950));
  nor2s1 _______441164(.DIN1 (_________28953), .DIN2 (_________28948),
       .Q (_________28949));
  nnd2s1 _______441165(.DIN1 (_________28946), .DIN2 (________21041),
       .Q (_________28947));
  or2s1 _______441166(.DIN1 (________________18690), .DIN2
       (____99___32749), .Q (____9____29004));
  nnd2s1 ______441167(.DIN1 (____99___32749), .DIN2
       (________________18690), .Q (____9____29005));
  or2s1 _______441168(.DIN1 (____________0_), .DIN2 (______0__28945),
       .Q (____9____29013));
  nor2s1 _____0_441169(.DIN1 (______9__28944), .DIN2 (____99___32749),
       .Q (____9_0__29012));
  xor2s1 _____0_441170(.DIN1 (_________28881), .DIN2 (_________33325),
       .Q (____9____29010));
  nnd2s1 _______441171(.DIN1 (______0__28945), .DIN2
       (____________0___18786), .Q (____9____29007));
  nnd2s1 _______441172(.DIN1 (_____9___28895), .DIN2 (_________28942),
       .Q (_________28943));
  xor2s1 _______441173(.DIN1 (_________28867), .DIN2 (____9_9__31781),
       .Q (_________28941));
  and2s1 _______441174(.DIN1 (______0__29230), .DIN2 (_________28939),
       .Q (_________28940));
  nor2s1 _______441175(.DIN1 (_________28939), .DIN2 (______0__29230),
       .Q (_________28938));
  nnd2s1 _______441176(.DIN1 (_________32029), .DIN2 (_________34448),
       .Q (_________28937));
  nnd2s1 _____0_441177(.DIN1 (_____9___28892), .DIN2 (__9_____27040),
       .Q (_________28936));
  nnd2s1 _______441178(.DIN1 (_____9___28889), .DIN2 (___0_____27587),
       .Q (______0__28935));
  and2s1 _______441179(.DIN1 (_____90__28888), .DIN2 (__9_9___26885),
       .Q (______9__28934));
  or2s1 ______441180(.DIN1 (_________34448), .DIN2 (_________32029), .Q
       (_________28933));
  nnd2s1 _____9_441181(.DIN1 (_____9___28893), .DIN2 (______9__28732),
       .Q (____9_0__29019));
  nnd2s1 _____9_441182(.DIN1 (_________28885), .DIN2 (_____9___28894),
       .Q (____9____29015));
  nnd2s1 _______441183(.DIN1 (______0__28945), .DIN2 (____________0_),
       .Q (______0__28965));
  dffacs1 _______________441184(.CLRB (reset), .CLK (clk), .DIN
       (_____0___28903), .QN (outData[1]));
  dffacs1 ____0_________________0_(.CLRB (reset), .CLK (clk), .DIN
       (_____9___28890), .QN (____0_____________0___18655));
  nnd2s1 ______441185(.DIN1 (_________28931), .DIN2 (_________28930),
       .Q (_________28932));
  or2s1 ______441186(.DIN1 (_________28930), .DIN2 (_________28931), .Q
       (_________28929));
  nnd2s1 _______441187(.DIN1 (_________28919), .DIN2 (_________28920),
       .Q (_________28928));
  nnd2s1 _______441188(.DIN1 (_________28872), .DIN2 (___00____27220),
       .Q (_________28927));
  and2s1 _______441189(.DIN1 (_________28882), .DIN2 (______0__28925),
       .Q (_________28926));
  nor2s1 ______441190(.DIN1 (________25958), .DIN2 (_____99__28897), .Q
       (_________28924));
  xor2s1 _______441191(.DIN1 (____________0___18753), .DIN2
       (_____00__28898), .Q (_________28923));
  or2s1 _______441192(.DIN1 (________22302), .DIN2 (_________28875), .Q
       (_________28922));
  xnr2s1 _______441193(.DIN1 (______0__31325), .DIN2 (_________28861),
       .Q (_________28978));
  nor2s1 _______441194(.DIN1 (________23567), .DIN2 (_________28921),
       .Q (_________28976));
  nor2s1 _______441195(.DIN1 (_________28920), .DIN2 (_________28919),
       .Q (_____9___28988));
  nor2s1 ______441196(.DIN1 (__9_____26713), .DIN2 (______0__28878), .Q
       (_________28918));
  nor2s1 _______441197(.DIN1 (__9_____26905), .DIN2 (______9__28877),
       .Q (______0__28917));
  nnd2s1 _______441198(.DIN1 (_________28874), .DIN2 (____0____28153),
       .Q (______9__28916));
  nor2s1 _______441199(.DIN1 (__9__9__26636), .DIN2 (_________28884),
       .Q (_________28915));
  nor2s1 ______441200(.DIN1 (______9__28320), .DIN2 (_________28870),
       .Q (_________28914));
  nor2s1 _______441201(.DIN1 (________26032), .DIN2 (_________28876),
       .Q (_________28913));
  xor2s1 _____9_441202(.DIN1 (_________28911), .DIN2 (_________28910),
       .Q (_________28912));
  nnd2s1 _______441203(.DIN1 (______0__28907), .DIN2 (__90____26286),
       .Q (_________28909));
  nnd2s1 _____0_441204(.DIN1 (______0__28907), .DIN2 (__9_9___26985),
       .Q (_________28908));
  nnd2s1 _____0_441205(.DIN1 (_________28871), .DIN2 (___0_____27410),
       .Q (_____09__28906));
  nor2s1 _______441206(.DIN1 (__9_____26432), .DIN2 (______0__28869),
       .Q (_________28967));
  hi1s1 _______441207(.DIN (_____0___28905), .Q (____90___28994));
  or2s1 _______441208(.DIN1 (____________0___18753), .DIN2 (____9), .Q
       (_____0___28904));
  or2s1 _____9_441209(.DIN1 (_________34500), .DIN2 (_____99__30363),
       .Q (_____0___28903));
  xnr2s1 _______441210(.DIN1 (____9_9__30888), .DIN2 (_____9___30358),
       .Q (_____0___28902));
  xnr2s1 _______441211(.DIN1 (____0____31820), .DIN2 (_____0___34734),
       .Q (_____0___28901));
  nnd2s1 _______441212(.DIN1 (____________0___18753), .DIN2
       (_____0__20049), .Q (_________28951));
  hi1s1 ______441213(.DIN (_____0___28900), .Q (_________28948));
  nor2s1 _______441214(.DIN1 (________23566), .DIN2 (_____0___28899),
       .Q (_________28946));
  or2s1 _____9_441215(.DIN1 (____________0___18753), .DIN2
       (_____00__28898), .Q (_________29382));
  hi1s1 _______441216(.DIN (_____99__28897), .Q (_____90__28983));
  xor2s1 _____441217(.DIN1 (_________28834), .DIN2 (_________28637), .Q
       (______0__28945));
  hi1s1 _______441218(.DIN (_____9___28896), .Q (____99___32749));
  and2s1 _______441219(.DIN1 (_________28857), .DIN2 (__9__9__26738),
       .Q (_____9___28895));
  nnd2s1 _______441220(.DIN1 (_________28886), .DIN2 (outData[31]), .Q
       (_____9___28894));
  nor2s1 _______441221(.DIN1 (_________28864), .DIN2 (______0__28860),
       .Q (_____9___28893));
  nnd2s1 _______441222(.DIN1 (_________28854), .DIN2 (_____9___28891),
       .Q (_____9___28892));
  nnd2s1 _______441223(.DIN1 (_________28858), .DIN2 (____9____29042),
       .Q (_____9___28890));
  nnd2s1 _______441224(.DIN1 (_________28856), .DIN2 (_____9___28891),
       .Q (_____9___28889));
  nor2s1 _______441225(.DIN1 (__9__9__26484), .DIN2 (______9__28859),
       .Q (_____90__28888));
  xor2s1 _____0_441226(.DIN1 (_________28873), .DIN2 (______9__28887),
       .Q (_____0___28905));
  nor2s1 _______441227(.DIN1 (______0__28840), .DIN2 (_________28886),
       .Q (____0____31858));
  xor2s1 _______441228(.DIN1 (__9_____26727), .DIN2 (______9__28868),
       .Q (______0__29230));
  hi1s1 ______441229(.DIN (_________28885), .Q (_________32029));
  nor2s1 ______441230(.DIN1 (________22146), .DIN2 (_________28852), .Q
       (_________28884));
  xor2s1 _____9_441231(.DIN1 (____0____30082), .DIN2 (____9____29986),
       .Q (_________28883));
  nnd2s1 _______441232(.DIN1 (_________28851), .DIN2 (_____9__21129),
       .Q (_________28882));
  nor2s1 _____9_441233(.DIN1 (_____09__28531), .DIN2 (_________28845),
       .Q (_________28881));
  nnd2s1 _______441234(.DIN1 (_________28846), .DIN2 (_____9___32185),
       .Q (_________28880));
  and2s1 _______441235(.DIN1 (_________28847), .DIN2 (_________32228),
       .Q (_________28879));
  xor2s1 _____9_441236(.DIN1 (_____90__28791), .DIN2 (_________28824),
       .Q (_____0___28900));
  xor2s1 _______441237(.DIN1 (______0__28820), .DIN2 (_________30166),
       .Q (_________28919));
  hi1s1 ______441238(.DIN (_____0___28899), .Q (_________28921));
  xor2s1 _______441239(.DIN1 (_________28827), .DIN2 (____0____32823),
       .Q (____9____29003));
  xor2s1 _______441240(.DIN1 (__9_____26733), .DIN2 (_________28862),
       .Q (_____9___28896));
  xor2s1 _____0_441241(.DIN1 (_________28816), .DIN2
       (______________________________________0__________0__18892), .Q
       (_____99__28897));
  xor2s1 _____0_441242(.DIN1 (_________28826), .DIN2 (_________35094),
       .Q (_________28931));
  xor2s1 _______441243(.DIN1 (______9__28819), .DIN2 (_________34023),
       .Q (_____0___30728));
  nnd2s1 ______441244(.DIN1 (_________28841), .DIN2 (___90___23350), .Q
       (______0__28878));
  nnd2s1 _______441245(.DIN1 (_________28842), .DIN2 (__9_00__26798),
       .Q (______9__28877));
  nnd2s1 _______441246(.DIN1 (______9__28839), .DIN2 (_________28837),
       .Q (_________28876));
  nnd2s1 _______441247(.DIN1 (_________28838), .DIN2 (___9____21622),
       .Q (_________28875));
  nor2s1 _______441248(.DIN1 (________23907), .DIN2 (_________28836),
       .Q (_________28874));
  nor2s1 _______441249(.DIN1 (________23589), .DIN2 (_________28843),
       .Q (_________28872));
  nor2s1 _______441250(.DIN1 (____90__23965), .DIN2 (_________28831),
       .Q (_________28871));
  nnd2s1 _______441251(.DIN1 (______9__28829), .DIN2 (________22694),
       .Q (_________28870));
  nor2s1 ______441252(.DIN1 (__9_____26431), .DIN2 (______9__28868), .Q
       (______0__28869));
  nor2s1 _______441253(.DIN1 (_________28866), .DIN2 (_________28865),
       .Q (_________28867));
  nor2s1 _______441254(.DIN1 (_____0___28805), .DIN2 (______0__28830),
       .Q (______0__28907));
  nnd2s1 _______441255(.DIN1 (_________28853), .DIN2
       (_____________18905), .Q (_________28885));
  xor2s1 ______441256(.DIN1 (_____09__28809), .DIN2 (_____0___32570),
       .Q (____9____31765));
  dffacs1 _______________________441257(.CLRB (reset), .CLK (clk), .DIN
       (_________28833), .QN (_____________________18612));
  nnd2s1 _______441258(.DIN1 (_________28813), .DIN2 (__9_____26810),
       .Q (_________28864));
  nor2s1 _______441259(.DIN1 (__9_____26732), .DIN2 (_________28862),
       .Q (_________28863));
  nnd2s1 _______441260(.DIN1 (_________28818), .DIN2 (_____9___28614),
       .Q (_________28861));
  dffacs1 ______________0____441261(.CLRB (reset), .CLK (clk), .DIN
       (_________28821), .Q (_________34500));
  nnd2s1 _______441262(.DIN1 (_________28812), .DIN2 (__9_____26808),
       .Q (______0__28860));
  xor2s1 _____0_441263(.DIN1 (_________28765), .DIN2 (_________28844),
       .Q (_____0___28899));
  dffacs1 ________________0_441264(.CLRB (reset), .CLK (clk), .DIN
       (_________28822), .QN (____________0___18753));
  nor2s1 ______441265(.DIN1 (__990___27084), .DIN2 (_____0___28803), .Q
       (______9__28859));
  nor2s1 _______441266(.DIN1 (__9_____26861), .DIN2 (_____0___28802),
       .Q (_________28858));
  nor2s1 _______441267(.DIN1 (__9__0__26864), .DIN2 (_____0___28806),
       .Q (_________28857));
  nor2s1 _______441268(.DIN1 (_____9__22699), .DIN2 (_____0___28804),
       .Q (_________28856));
  nor2s1 _______441269(.DIN1 (______________18869), .DIN2
       (_________28911), .Q (_________28855));
  nor2s1 ______441270(.DIN1 (____9___22349), .DIN2 (_____0___28801), .Q
       (_________28854));
  hi1s1 _______441271(.DIN (_________28853), .Q (_________28886));
  nor2s1 _______441272(.DIN1 (_________28638), .DIN2 (_________28815),
       .Q (_________28910));
  nnd2s1 _______441273(.DIN1 (______9__28780), .DIN2 (__9_____26877),
       .Q (_________28852));
  nnd2s1 _______441274(.DIN1 (_____9___28797), .DIN2 (_________28734),
       .Q (_________28851));
  nnd2s1 _____441275(.DIN1 (_____9___28795), .DIN2 (________19986), .Q
       (______0__28850));
  nnd2s1 _______441276(.DIN1 (_________28848), .DIN2 (_____9___28703),
       .Q (______9__28849));
  nor2s1 _______441277(.DIN1 (_____00__28800), .DIN2 (___9____23393),
       .Q (_________28847));
  nnd2s1 _______441278(.DIN1 (______9__28790), .DIN2 (_________31956),
       .Q (_________28846));
  nor2s1 ______441279(.DIN1 (_________28664), .DIN2 (_________28844),
       .Q (_________28845));
  nnd2s1 ______441280(.DIN1 (_________28786), .DIN2 (___9____26200), .Q
       (_________28843));
  nor2s1 ______441281(.DIN1 (____9___25943), .DIN2 (_____9___28794), .Q
       (_________28842));
  nor2s1 _______441282(.DIN1 (___9____23407), .DIN2 (_____9___28793),
       .Q (_________28841));
  xor2s1 _____0_441283(.DIN1 (_________28767), .DIN2 (____0_0__30932),
       .Q (_____09__30554));
  nnd2s1 ______441284(.DIN1 (_____9___28792), .DIN2 (_________28490),
       .Q (____00___30907));
  xor2s1 _______441285(.DIN1 (_____00__28616), .DIN2 (_________28817),
       .Q (_____9___30358));
  xor2s1 _______441286(.DIN1 (_________28756), .DIN2 (_________31326),
       .Q (______0__28840));
  nor2s1 _______441287(.DIN1 (__9_____26632), .DIN2 (_________28784),
       .Q (______9__28839));
  nnd2s1 _______441288(.DIN1 (_________28782), .DIN2 (_________28837),
       .Q (_________28838));
  nnd2s1 _____9_441289(.DIN1 (_________28785), .DIN2 (_________28298),
       .Q (_________28836));
  nnd2s1 _____9_441290(.DIN1 (_________28749), .DIN2 (_________28787),
       .Q (_________28835));
  xor2s1 _____441291(.DIN1 (_________28814), .DIN2 (_________28661), .Q
       (_________28834));
  nnd2s1 _______441292(.DIN1 (_________28783), .DIN2 (_________28832),
       .Q (_________28833));
  nnd2s1 _______441293(.DIN1 (_________28776), .DIN2 (________26089),
       .Q (_________28831));
  nnd2s1 _______441294(.DIN1 (_________28772), .DIN2 (_________35064),
       .Q (______0__28830));
  nor2s1 ______441295(.DIN1 (________23105), .DIN2 (_________28777), .Q
       (______9__28829));
  xor2s1 _____0_441296(.DIN1 (_________28758), .DIN2 (_________28828),
       .Q (_________28853));
  nor2s1 _______441297(.DIN1 (________19091), .DIN2 (_________28774),
       .Q (______9__28868));
  hi1s1 _______441298(.DIN (_________28911), .Q (_________28865));
  xor2s1 _____0_441299(.DIN1 (_________28759), .DIN2 (____0____30044),
       .Q (_________28873));
  dffacs1 _______________________441300(.CLRB (reset), .CLK (clk), .DIN
       (______0__28781), .QN (_____________________18610));
  nnd2s1 _______441301(.DIN1 (_________28763), .DIN2 (___0_____27342),
       .Q (_________28827));
  xor2s1 _____9_441302(.DIN1 (___090___28044), .DIN2 (_____9___28796),
       .Q (_________28826));
  xnr2s1 _____9_441303(.DIN1 (_________34493), .DIN2 (_________32946),
       .Q (_________28825));
  xor2s1 _____9_441304(.DIN1 (_________28727), .DIN2 (_________32049),
       .Q (_________28824));
  nor2s1 _____441305(.DIN1 (_____9___32185), .DIN2 (_____0___32104), .Q
       (_________28823));
  nnd2s1 _____441306(.DIN1 (______9__28770), .DIN2 (________20537), .Q
       (_________28822));
  nnd2s1 _______441307(.DIN1 (______0__28771), .DIN2 (_________34365),
       .Q (_________28821));
  xor2s1 _______441308(.DIN1 (_________28491), .DIN2
       (________________18735), .Q (______0__28820));
  nnd2s1 _______441309(.DIN1 (_____0___32104), .DIN2 (_____0___28712),
       .Q (______9__28819));
  nnd2s1 _______441310(.DIN1 (_________28817), .DIN2 (_________28580),
       .Q (_________28818));
  nnd2s1 _______441311(.DIN1 (_________28768), .DIN2 (________23744),
       .Q (_________28862));
  xor2s1 _____441312(.DIN1 (_________28742), .DIN2 (___0__0__27589), .Q
       (____0____30082));
  xor2s1 _____9_441313(.DIN1 (_________28729), .DIN2 (____099__30093),
       .Q (_________28816));
  nor2s1 _______441314(.DIN1 (_________28662), .DIN2 (_________28814),
       .Q (_________28815));
  or2s1 _______441315(.DIN1 (______0__28810), .DIN2 (_________28811),
       .Q (_________28813));
  nnd2s1 _______441316(.DIN1 (_________28811), .DIN2 (______0__28810),
       .Q (_________28812));
  and2s1 ______441317(.DIN1 (______9__28760), .DIN2 (_________28766),
       .Q (_____09__28809));
  nor2s1 _______441318(.DIN1 (_____0___28807), .DIN2 (______9__28750),
       .Q (_____0___28808));
  nor2s1 _______441319(.DIN1 (_____0___28805), .DIN2 (_________28752),
       .Q (_____0___28806));
  nnd2s1 ______441320(.DIN1 (_________28747), .DIN2 (__9_____26525), .Q
       (_____0___28804));
  nnd2s1 _______441321(.DIN1 (______0__28761), .DIN2 (________22953),
       .Q (_____0___28803));
  nnd2s1 _______441322(.DIN1 (_________28746), .DIN2 (___0_9___27356),
       .Q (_____0___28802));
  nnd2s1 ______441323(.DIN1 (_________28745), .DIN2 (_________28602),
       .Q (_____0___28801));
  xor2s1 _______441324(.DIN1 (_________28773), .DIN2 (________20433),
       .Q (_________28911));
  dffacs1 __________________441325(.CLRB (reset), .CLK (clk), .DIN
       (_________28769), .QN (______0__34471));
  nor2s1 _______441326(.DIN1 (________________18735), .DIN2
       (_________28788), .Q (_____00__28800));
  nnd2s1 _______441327(.DIN1 (_________32946), .DIN2 (_________34493),
       .Q (_____99__28799));
  or2s1 _______441328(.DIN1 (_________34493), .DIN2 (_________32946),
       .Q (_____9___28798));
  or2s1 _______441329(.DIN1 (_____0__19985), .DIN2 (_____9___28796), .Q
       (_____9___28797));
  and2s1 _______441330(.DIN1 (_____9___28796), .DIN2 (_____9__20381),
       .Q (_____9___28795));
  nnd2s1 _______441331(.DIN1 (_________28740), .DIN2 (___9____24253),
       .Q (_____9___28794));
  nnd2s1 _______441332(.DIN1 (______9__28741), .DIN2 (________24970),
       .Q (_____9___28793));
  nnd2s1 _____9_441333(.DIN1 (_________28489), .DIN2
       (________________18735), .Q (_____9___28792));
  hi1s1 _______441334(.DIN (_____0___32104), .Q (______9__28790));
  hi1s1 _______441335(.DIN (_________28789), .Q (_________30352));
  xor2s1 _______441336(.DIN1 (_____09__28713), .DIN2 (____009__31815),
       .Q (_________28848));
  xor2s1 _____0_441337(.DIN1 (_____0___34736), .DIN2 (_________33384),
       .Q (_________28844));
  nnd2s1 ______441338(.DIN1 (_________28788), .DIN2
       (________________18735), .Q (_________32228));
  dffacs1 ____0__________________441339(.CLRB (reset), .CLK (clk), .DIN
       (_________28724), .QN (____0________________18589));
  nnd2s1 _______441340(.DIN1 (_________28730), .DIN2 (_________31956),
       .Q (_________28787));
  nor2s1 _______441341(.DIN1 (__9__9__27073), .DIN2 (_________28735),
       .Q (_________28786));
  nor2s1 _______441342(.DIN1 (_________28671), .DIN2 (______0__28733),
       .Q (_________28785));
  nnd2s1 _______441343(.DIN1 (_________28738), .DIN2 (___09___23522),
       .Q (_________28784));
  nor2s1 _______441344(.DIN1 (_________28667), .DIN2 (_________28736),
       .Q (_________28783));
  nor2s1 _______441345(.DIN1 (___90___26154), .DIN2 (_________28725),
       .Q (_________28782));
  nnd2s1 _______441346(.DIN1 (_________28731), .DIN2 (______9__28444),
       .Q (______0__28781));
  nor2s1 _______441347(.DIN1 (__9_____26350), .DIN2 (_________28739),
       .Q (______9__28780));
  nor2s1 ______441348(.DIN1 (___09____28064), .DIN2 (______0__29571),
       .Q (_________28779));
  xor2s1 _______441349(.DIN1 (_________28748), .DIN2 (_________31956),
       .Q (_________28778));
  nnd2s1 _______441350(.DIN1 (_________28721), .DIN2 (___0_9__24418),
       .Q (_________28777));
  nor2s1 _______441351(.DIN1 (_________28775), .DIN2 (______9__28722),
       .Q (_________28776));
  nor2s1 ______441352(.DIN1 (_______19005), .DIN2 (_________28773), .Q
       (_________28774));
  nor2s1 _____441353(.DIN1 (__9_____26838), .DIN2 (______0__28723), .Q
       (_________28772));
  dffacs1 ________________________441354(.CLRB (reset), .CLK (clk),
       .DIN (_________28720), .Q (______________________18644));
  xor2s1 ______441355(.DIN1 (_________28683), .DIN2 (_________28684),
       .Q (______0__28771));
  or2s1 _______441356(.DIN1 (____9____32723), .DIN2 (_________28690),
       .Q (______9__28770));
  nnd2s1 _______441357(.DIN1 (_________28718), .DIN2 (_________31303),
       .Q (_________28769));
  nor2s1 ______441358(.DIN1 (___09___24427), .DIN2 (_____0___28707), .Q
       (_________28768));
  nnd2s1 _______441359(.DIN1 (_________28716), .DIN2 (_________28766),
       .Q (_________28767));
  xor2s1 _____9_441360(.DIN1 (______0__28677), .DIN2 (_____0___31450),
       .Q (_________28765));
  nor2s1 _______441361(.DIN1 (_________31153), .DIN2 (_____0___28708),
       .Q (_________28764));
  xnr2s1 ______441362(.DIN1 (_________31505), .DIN2 (_________28678),
       .Q (_________28763));
  nnd2s1 _______441363(.DIN1 (_________28717), .DIN2 (___0_____27590),
       .Q (_________28789));
  nnd2s1 _______441364(.DIN1 (_____00__28705), .DIN2 (_________28728),
       .Q (_________28817));
  nor2s1 _____0_441365(.DIN1 (______9__28596), .DIN2 (_____0___28709),
       .Q (_________30220));
  xor2s1 _______441366(.DIN1 (_________28680), .DIN2 (_________31154),
       .Q (____0____31844));
  nor2s1 _____0_441367(.DIN1 (_________28762), .DIN2 (_____0___28710),
       .Q (_____0___32104));
  nor2s1 _______441368(.DIN1 (__9_____26935), .DIN2 (_____90__28696),
       .Q (______0__28761));
  and2s1 _______441369(.DIN1 (_________28757), .DIN2 (_____9___28612),
       .Q (______9__28760));
  nnd2s1 _______441370(.DIN1 (_____9___28698), .DIN2 (_____9__19428),
       .Q (_________28759));
  nor2s1 _______441371(.DIN1 (outData[30]), .DIN2 (_________28757), .Q
       (_________28758));
  nnd2s1 _______441372(.DIN1 (_________28757), .DIN2 (outData[30]), .Q
       (_________28756));
  nor2s1 _______441373(.DIN1 (_________28754), .DIN2 (_________28753),
       .Q (_________28755));
  or2s1 ______441374(.DIN1 (______0__28751), .DIN2 (_________28688), .Q
       (_________28752));
  hi1s1 _______441375(.DIN (______0__29571), .Q (______9__28750));
  nnd2s1 _____9_441376(.DIN1 (_________28748), .DIN2 (___0____22546),
       .Q (_________28749));
  nor2s1 _______441377(.DIN1 (_____0__22242), .DIN2 (_________28689),
       .Q (_________28747));
  or2s1 ______441378(.DIN1 (_____0___28805), .DIN2 (_________28691), .Q
       (_________28746));
  nor2s1 ______441379(.DIN1 (__9_____27037), .DIN2 (______9__28695), .Q
       (_________28745));
  nor2s1 ______441380(.DIN1 (_________28654), .DIN2 (_________28744),
       .Q (_________28814));
  nor2s1 _______441381(.DIN1 (_________28653), .DIN2 (_________28744),
       .Q (_________28811));
  xor2s1 _____9_441382(.DIN1 (________________18757), .DIN2
       (_________28645), .Q (_________28743));
  xor2s1 _____441383(.DIN1 (________________18706), .DIN2
       (_________28645), .Q (_________28742));
  nor2s1 _______441384(.DIN1 (___00___24340), .DIN2 (______0__34738),
       .Q (______9__28741));
  nor2s1 _______441385(.DIN1 (________24806), .DIN2 (______9__28676),
       .Q (_________28740));
  nnd2s1 _______441386(.DIN1 (_________28666), .DIN2 (___9____26218),
       .Q (_________28739));
  nor2s1 _______441387(.DIN1 (__9_____26650), .DIN2 (_________34742),
       .Q (_________28738));
  nnd2s1 _______441388(.DIN1 (_________28672), .DIN2 (________24146),
       .Q (_________28736));
  nnd2s1 ______441389(.DIN1 (_________28675), .DIN2 (__9_____26591), .Q
       (_________28735));
  xor2s1 _______441390(.DIN1 (_________28628), .DIN2 (_________28648),
       .Q (_____90__28791));
  nor2s1 _____0_441391(.DIN1 (_________28681), .DIN2 (______9__28685),
       .Q (_________29649));
  xnr2s1 _____0_441392(.DIN1 (outData[30]), .DIN2 (_________28715), .Q
       (______0__30475));
  xnr2s1 _____0_441393(.DIN1 (_________28734), .DIN2 (______0__28925),
       .Q (_____9___28796));
  dffacs1 __________________441394(.CLRB (reset), .CLK (clk), .DIN
       (_________28679), .Q (________________18735));
  xnr2s1 _____441395(.DIN1 (_____0___28706), .DIN2 (____0___24794), .Q
       (_________32946));
  nnd2s1 _____9_441396(.DIN1 (_________28674), .DIN2 (_________28278),
       .Q (______0__28733));
  xor2s1 _____9_441397(.DIN1 (_________28640), .DIN2 (____90___28993),
       .Q (______9__28732));
  nor2s1 _____9_441398(.DIN1 (______9__28588), .DIN2 (______9__28668),
       .Q (_________28731));
  xor2s1 _____441399(.DIN1 (_________28692), .DIN2 (______0__29466), .Q
       (_________28730));
  nnd2s1 _____0_441400(.DIN1 (_____99__28704), .DIN2 (_________28728),
       .Q (_________28729));
  nor2s1 _____0_441401(.DIN1 (_________28726), .DIN2 (_____9___28699),
       .Q (_________28727));
  nnd2s1 _____9_441402(.DIN1 (_________28669), .DIN2 (__9_____26871),
       .Q (_________28725));
  nnd2s1 _______441403(.DIN1 (______0__28659), .DIN2 (_________28626),
       .Q (_________28724));
  nnd2s1 _______441404(.DIN1 (______9__28658), .DIN2 (___0_____27897),
       .Q (______0__28723));
  nnd2s1 _______441405(.DIN1 (_________28657), .DIN2 (________23760),
       .Q (______9__28722));
  nor2s1 _______441406(.DIN1 (________25544), .DIN2 (_________28655),
       .Q (_________28721));
  nnd2s1 _______441407(.DIN1 (_________28660), .DIN2 (_____9___28517),
       .Q (_________28720));
  xor2s1 ______441408(.DIN1 (_________28639), .DIN2 (_________33541),
       .Q (_________28773));
  dffacs1 _____________________9_441409(.CLRB (reset), .CLK (clk), .DIN
       (_________28651), .QN (_________________9___18616));
  dffacs1 ____0________________9_(.CLRB (reset), .CLK (clk), .DIN
       (_________28665), .QN (____0____________9_));
  xor2s1 _______441410(.DIN1 (_____9___28697), .DIN2 (_____0__19966),
       .Q (______0__29571));
  xor2s1 _____0_441411(.DIN1 (_____0___28618), .DIN2 (______9__33247),
       .Q (_________28719));
  nor2s1 _______441412(.DIN1 (____0___23976), .DIN2 (_________28646),
       .Q (_________28718));
  or2s1 _______441413(.DIN1 (___0__9__27588), .DIN2 (_________28645),
       .Q (_________28717));
  and2s1 _______441414(.DIN1 (_________28715), .DIN2 (______9__28642),
       .Q (_________28716));
  nor2s1 _______441415(.DIN1 (___0_0__20743), .DIN2 (_________28645),
       .Q (______0__28714));
  nor2s1 ______441416(.DIN1 (____00__21260), .DIN2 (_________28645), .Q
       (_____09__28713));
  or2s1 ______441417(.DIN1 (_____0___28711), .DIN2 (_________28715), .Q
       (_____0___28712));
  and2s1 _______441418(.DIN1 (_________28715), .DIN2
       (_____________18905), .Q (_____0___28710));
  nnd2s1 _______441419(.DIN1 (_________28650), .DIN2 (_________28644),
       .Q (_____0___28709));
  nnd2s1 _______441420(.DIN1 (______0__28925), .DIN2 (________21126),
       .Q (_____0___28708));
  nor2s1 _______441421(.DIN1 (____9___23339), .DIN2 (_____0___28706),
       .Q (_____0___28707));
  nnd2s1 _____9_441422(.DIN1 (_____99__28704), .DIN2 (_________29585),
       .Q (_____00__28705));
  hi1s1 ______441423(.DIN (_____9___28702), .Q (_____9___28703));
  nnd2s1 _______441424(.DIN1 (_____9___28700), .DIN2 (_________28652),
       .Q (_____9___28701));
  or2s1 _______441425(.DIN1 (____09__19123), .DIN2 (_____9___28697), .Q
       (_____9___28698));
  nnd2s1 _____9_441426(.DIN1 (_________28694), .DIN2 (___0_99__27849),
       .Q (_____90__28696));
  nnd2s1 ______441427(.DIN1 (_________28694), .DIN2 (___0__9__27898),
       .Q (______9__28695));
  nor2s1 ______441428(.DIN1 (_________28692), .DIN2 (______0__29466),
       .Q (_________28693));
  nnd2s1 _______441429(.DIN1 (_________28694), .DIN2 (__9__0__26834),
       .Q (_________28691));
  xor2s1 _____0_441430(.DIN1 (_____99__28615), .DIN2 (_________28457),
       .Q (_________28690));
  nnd2s1 _______441431(.DIN1 (_________28694), .DIN2 (____0____28197),
       .Q (_________28689));
  nnd2s1 _______441432(.DIN1 (_________28694), .DIN2 (___0_0___27371),
       .Q (_________28688));
  xor2s1 _______441433(.DIN1 (_____9___28608), .DIN2 (_________33564),
       .Q (_________28744));
  and2s1 _______441434(.DIN1 (_________28687), .DIN2
       (_________________18749), .Q (_________28753));
  and2s1 _______441435(.DIN1 (______0__29466), .DIN2 (_________28692),
       .Q (_________28748));
  nor2s1 _______441436(.DIN1 (_________________18749), .DIN2
       (_________28687), .Q (_________28754));
  xor2s1 _______441437(.DIN1 (______9__28605), .DIN2 (_________33268),
       .Q (_________28757));
  nor2s1 _______441438(.DIN1 (________________18757), .DIN2
       (_________28670), .Q (______0__28686));
  nor2s1 ______441439(.DIN1 (_________28684), .DIN2 (_________28682),
       .Q (______9__28685));
  or2s1 _______441440(.DIN1 (_________28682), .DIN2 (_________28681),
       .Q (_________28683));
  xor2s1 _______441441(.DIN1 (outData[28]), .DIN2 (_________28649), .Q
       (_________28680));
  nnd2s1 _____9_441442(.DIN1 (_________28631), .DIN2 (________24503),
       .Q (_________28679));
  nnd2s1 _____0_441443(.DIN1 (_________28630), .DIN2 (____0____28162),
       .Q (_________28678));
  nnd2s1 _____0_441444(.DIN1 (_________28663), .DIN2 (_________28632),
       .Q (______0__28677));
  nnd2s1 _______441445(.DIN1 (_________28673), .DIN2 (__9_____27069),
       .Q (______9__28676));
  nor2s1 _______441446(.DIN1 (__9_0___26338), .DIN2 (_____09__28624),
       .Q (_________28675));
  nor2s1 _______441447(.DIN1 (_____9__23914), .DIN2 (______0__28625),
       .Q (_________28674));
  nor2s1 _______441448(.DIN1 (_________28671), .DIN2 (_____0___28623),
       .Q (_________28672));
  nor2s1 _______441449(.DIN1
       (_______________0____________________18829), .DIN2
       (_________28670), .Q (_____9___28702));
  nor2s1 _______441450(.DIN1 (_________34746), .DIN2 (_________34744),
       .Q (_____9___28699));
  nor2s1 ______441451(.DIN1 (_________28647), .DIN2 (_________28629),
       .Q (_________28930));
  nor2s1 ______441452(.DIN1 (________25582), .DIN2 (______9__28633), .Q
       (_________28669));
  or2s1 _______441453(.DIN1 (_________28667), .DIN2 (_________28635),
       .Q (______9__28668));
  nor2s1 _______441454(.DIN1 (____9___26144), .DIN2 (_____0___28622),
       .Q (_________28666));
  nnd2s1 _______441455(.DIN1 (_________28627), .DIN2 (___09____28074),
       .Q (_________28665));
  and2s1 _______441456(.DIN1 (_________28663), .DIN2 (______0__28634),
       .Q (_________28664));
  nor2s1 _____0_441457(.DIN1 (_________28661), .DIN2 (_____90__28606),
       .Q (_________28662));
  nor2s1 _____441458(.DIN1 (__9_____27013), .DIN2 (_____0___28619), .Q
       (_________28660));
  nor2s1 _______441459(.DIN1 (________23762), .DIN2 (_____0___28621),
       .Q (______0__28659));
  nor2s1 _______441460(.DIN1 (_________28636), .DIN2 (_________28656),
       .Q (______9__28658));
  nor2s1 ______441461(.DIN1 (___0__9__27286), .DIN2 (_________28656),
       .Q (_________28657));
  nnd2s1 _______441462(.DIN1 (_____9___28613), .DIN2 (___0____23449),
       .Q (_________28655));
  nor2s1 _______441463(.DIN1 (______0__28810), .DIN2 (_________28653),
       .Q (_________28654));
  nnd2s1 _____9_441464(.DIN1 (_____0___28620), .DIN2 (_________28537),
       .Q (_________28651));
  xor2s1 _______441465(.DIN1 (_________28583), .DIN2 (_________31164),
       .Q (_________28728));
  and2s1 _______441466(.DIN1 (_________34744), .DIN2 (_________34746),
       .Q (_________28726));
  or2s1 _____9_441467(.DIN1 (______0__28643), .DIN2 (_________28649),
       .Q (_________28650));
  nor2s1 _______441468(.DIN1 (_________28591), .DIN2 (_________28647),
       .Q (_________28648));
  nor2s1 _____441469(.DIN1 (_____9___30454), .DIN2 (_________28594), .Q
       (_________28646));
  hi1s1 _______441470(.DIN (_________28670), .Q (_________28645));
  nnd2s1 ______441471(.DIN1 (_________28600), .DIN2 (______0__28643),
       .Q (_________28644));
  nnd2s1 _______441472(.DIN1 (_________28649), .DIN2 (outData[29]), .Q
       (______9__28642));
  nnd2s1 _____441473(.DIN1 (_________28595), .DIN2 (_____0__23115), .Q
       (_____0___28706));
  or2s1 _______441474(.DIN1 (_________28604), .DIN2 (_________28649),
       .Q (_________28715));
  xnr2s1 _______441475(.DIN1 (_________28641), .DIN2 (_________28564),
       .Q (______0__28925));
  nor2s1 _______441476(.DIN1 (______9__28262), .DIN2 (_________28576),
       .Q (_________28640));
  nnd2s1 _______441477(.DIN1 (_________28574), .DIN2 (_____0___28526),
       .Q (_________28639));
  nor2s1 _____0_441478(.DIN1
       (______________________________________0___________), .DIN2
       (_________28637), .Q (_________28638));
  xor2s1 ______441479(.DIN1 (_________28548), .DIN2 (_________32644),
       .Q (_____99__28704));
  nor2s1 _______441480(.DIN1 (________19276), .DIN2 (_________28585),
       .Q (_____9___28697));
  or2s1 _____0_441481(.DIN1 (_______________18874), .DIN2
       (_________28637), .Q (_____9___28700));
  nnd2s1 _____0_441482(.DIN1 (_________28637), .DIN2
       (_______________18874), .Q (_________28652));
  nor2s1 _____441483(.DIN1 (______0__28542), .DIN2 (_________28582), .Q
       (_________28687));
  xor2s1 _______441484(.DIN1 (_____________18902), .DIN2
       (_____9___28611), .Q (____0____32826));
  dffacs1 _______________________441485(.CLRB (reset), .CLK (clk), .DIN
       (_________28575), .QN (_____________________18613));
  nor2s1 ______441486(.DIN1 (_________28636), .DIN2 (_________28573),
       .Q (_________28694));
  hi1s1 _____9_441487(.DIN (_________29472), .Q (______0__29466));
  dffacs1 _______________________441488(.CLRB (reset), .CLK (clk), .DIN
       (______0__28589), .QN (_____________________18609));
  nnd2s1 _______441489(.DIN1 (_________28561), .DIN2 (__99____27110),
       .Q (_________28635));
  nnd2s1 _____441490(.DIN1 (_________28566), .DIN2 (_________33444), .Q
       (______0__28634));
  nnd2s1 _____9_441491(.DIN1 (_________28563), .DIN2 (___00____27222),
       .Q (______9__28633));
  nnd2s1 ______441492(.DIN1 (______0__28569), .DIN2 (_________33444),
       .Q (_________28632));
  nnd2s1 _______441493(.DIN1 (______9__28568), .DIN2 (_________34966),
       .Q (_________28631));
  nor2s1 _______441494(.DIN1 (___0_____27911), .DIN2 (_________28570),
       .Q (_________28630));
  and2s1 ______441495(.DIN1 (_________28590), .DIN2 (_________28628),
       .Q (_________28629));
  and2s1 _______441496(.DIN1 (_________28562), .DIN2 (_________28626),
       .Q (_________28627));
  nnd2s1 _______441497(.DIN1 (_________28553), .DIN2 (_________28478),
       .Q (______0__28625));
  nnd2s1 ______441498(.DIN1 (_________28571), .DIN2 (____00__25948), .Q
       (_____09__28624));
  nnd2s1 ______441499(.DIN1 (_________28567), .DIN2 (____9___23167), .Q
       (_____0___28623));
  nnd2s1 _______441500(.DIN1 (_________28558), .DIN2 (________25704),
       .Q (_____0___28622));
  xor2s1 _____0_441501(.DIN1 (_________28535), .DIN2 (______0__29851),
       .Q (_________28681));
  xor2s1 _____0_441502(.DIN1 (_________28536), .DIN2 (_________29496),
       .Q (_________28682));
  nor2s1 _______441503(.DIN1 (_________28572), .DIN2 (_________28599),
       .Q (____0____30071));
  xor2s1 _______441504(.DIN1 (_________28540), .DIN2 (_________28737),
       .Q (_________28670));
  nnd2s1 _______441505(.DIN1 (_________28546), .DIN2 (________23197),
       .Q (_____0___28621));
  nor2s1 _______441506(.DIN1 (_________28497), .DIN2 (_________28544),
       .Q (_____0___28620));
  nor2s1 ______441507(.DIN1 (__99_9__27116), .DIN2 (_________28547), .Q
       (_____0___28619));
  and2s1 _______441508(.DIN1 (_____9___28609), .DIN2 (_____0___28617),
       .Q (_____0___28618));
  xor2s1 _______441509(.DIN1 (______0__28579), .DIN2
       (_______________18873), .Q (_____00__28616));
  xor2s1 ______441510(.DIN1 (_____00__28523), .DIN2 (_____0___31450),
       .Q (_____99__28615));
  nnd2s1 _______441511(.DIN1 (_____9___28607), .DIN2
       (_______________18873), .Q (_____9___28614));
  nnd2s1 _______441512(.DIN1 (_________28543), .DIN2 (___0_____27862),
       .Q (_____9___28613));
  nnd2s1 _______441513(.DIN1 (_____9___28611), .DIN2 (outData[29]), .Q
       (_____9___28612));
  nor2s1 _____0_441514(.DIN1 (_____0___28617), .DIN2 (_____9___28609),
       .Q (_____9___28610));
  nnd2s1 _______441515(.DIN1 (_____9___28607), .DIN2 (_________28603),
       .Q (_____9___28608));
  hi1s1 _______441516(.DIN (_________28637), .Q (_____90__28606));
  or2s1 _______441517(.DIN1 (_________28604), .DIN2 (_____9___28611),
       .Q (______9__28605));
  nor2s1 _______441518(.DIN1 (_________28603), .DIN2 (_____9___28607),
       .Q (_________28653));
  nnd2s1 _______441519(.DIN1 (_________28545), .DIN2 (_________28602),
       .Q (_________28656));
  nor2s1 _______441520(.DIN1 (________22146), .DIN2 (_________28552),
       .Q (_________28673));
  dffacs1 _______________________441521(.CLRB (reset), .CLK (clk), .DIN
       (_________28554), .QN (_____________________18598));
  xor2s1 _______441522(.DIN1 (_________28584), .DIN2 (_________28601),
       .Q (_________29472));
  and2s1 ______441523(.DIN1 (_________28599), .DIN2 (outData[27]), .Q
       (_________28600));
  nnd2s1 _______441524(.DIN1 (______0__28597), .DIN2 (_________28586),
       .Q (_________28598));
  nor2s1 _______441525(.DIN1 (________19475), .DIN2 (_________28599),
       .Q (______9__28596));
  xnr2s1 _______441526(.DIN1 (____0_9__30961), .DIN2 (______0__28504),
       .Q (_________28595));
  xor2s1 _______441527(.DIN1 (_________28512), .DIN2 (_________31983),
       .Q (_________28594));
  hi1s1 _____9_441528(.DIN (_________28590), .Q (_________28591));
  or2s1 ______441529(.DIN1 (______9__28588), .DIN2 (______0__28532), .Q
       (______0__28589));
  nor2s1 _______441530(.DIN1 (_________28586), .DIN2 (______0__28597),
       .Q (_________28587));
  nor2s1 ______441531(.DIN1 (________19275), .DIN2 (_________28584), .Q
       (_________28585));
  nnd2s1 _______441532(.DIN1 (_________28565), .DIN2 (_____99__31353),
       .Q (_________28663));
  nnd2s1 _______441533(.DIN1 (_________28599), .DIN2 (_________28581),
       .Q (_________28649));
  nor2s1 _______441534(.DIN1 (____0____28202), .DIN2 (_____0___28528),
       .Q (_________28583));
  nor2s1 ______441535(.DIN1 (_________28581), .DIN2 (_____0___28524),
       .Q (_________28582));
  nnd2s1 _______441536(.DIN1 (______0__28579), .DIN2 (______9__28578),
       .Q (_________28580));
  nor2s1 _______441537(.DIN1 (__9_0___26800), .DIN2 (_________29396),
       .Q (_________28577));
  xor2s1 _______441538(.DIN1 (_________28487), .DIN2 (____00___33677),
       .Q (_________28576));
  nnd2s1 _______441539(.DIN1 (_________28538), .DIN2 (________25049),
       .Q (_________28575));
  nnd2s1 _______441540(.DIN1 (_____99__28522), .DIN2 (____9_9__33643),
       .Q (_________28574));
  nor2s1 ______441541(.DIN1 (__9090), .DIN2 (_____9___28520), .Q
       (_________28573));
  dffacs1 ________________________441542(.CLRB (reset), .CLK (clk),
       .DIN (_____9___28521), .QN (______________________18617));
  hi1s1 _______441543(.DIN (_____9___28609), .Q (_________30587));
  dffacs1 ________________0_441544(.CLRB (reset), .CLK (clk), .DIN
       (_________28539), .Q (_________34472));
  dffacs1 _______________________441545(.CLRB (reset), .CLK (clk), .DIN
       (_____9___28518), .QN (_____________________18640));
  xor2s1 _______441546(.DIN1 (_________28451), .DIN2 (_________28488),
       .Q (_________28637));
  dffacs1 ____0__________________441547(.CLRB (reset), .CLK (clk), .DIN
       (_____0___28525), .QN (____0______________));
  nor2s1 _______441548(.DIN1 (_____________18901), .DIN2
       (_________28510), .Q (_________28572));
  nor2s1 ______441549(.DIN1 (___9_9__25202), .DIN2 (_________28501), .Q
       (_________28571));
  nnd2s1 _____9_441550(.DIN1 (_________28505), .DIN2 (___0_____27910),
       .Q (_________28570));
  xor2s1 _____0_441551(.DIN1 (_____0___28530), .DIN2 (_________29291),
       .Q (______0__28569));
  xor2s1 _____0_441552(.DIN1 (______0__34471), .DIN2 (_________28472),
       .Q (______9__28568));
  nor2s1 _______441553(.DIN1 (____0___23261), .DIN2 (______9__28484),
       .Q (_________28567));
  hi1s1 _______441554(.DIN (_________28565), .Q (_________28566));
  xor2s1 ______441555(.DIN1 (_____0___28529), .DIN2 (____0____28174),
       .Q (_________28564));
  nor2s1 _______441556(.DIN1 (__9_09__26995), .DIN2 (_________28502),
       .Q (_________28563));
  nor2s1 _______441557(.DIN1 (______9__28464), .DIN2 (_________28499),
       .Q (_________28562));
  nor2s1 _______441558(.DIN1 (_____00__28331), .DIN2 (_________28498),
       .Q (_________28561));
  nor2s1 ______441559(.DIN1 (__990___27088), .DIN2 (_____9___28514), .Q
       (_________28558));
  nor2s1 _______441560(.DIN1 (_________28556), .DIN2 (_________28557),
       .Q (_________28647));
  nnd2s1 _______441561(.DIN1 (_________28557), .DIN2 (_________28556),
       .Q (_________28590));
  nnd2s1 _______441562(.DIN1 (______9__28513), .DIN2 (_________28506),
       .Q (_________29784));
  nnd2s1 _______441563(.DIN1 (_________28495), .DIN2 (________23207),
       .Q (_________28555));
  nnd2s1 _______441564(.DIN1 (______9__28493), .DIN2 (________25113),
       .Q (_________28554));
  nor2s1 _______441565(.DIN1 (_________28483), .DIN2 (_________28500),
       .Q (_________28553));
  or2s1 _______441566(.DIN1 (______0__28551), .DIN2 (_________28508),
       .Q (_________28552));
  nor2s1 _______441567(.DIN1 (_________28549), .DIN2 (_____9___28515),
       .Q (_________28550));
  nor2s1 ______441568(.DIN1 (____09___28228), .DIN2 (_____0___28527),
       .Q (_________28548));
  nnd2s1 ____9_441569(.DIN1 (_________28480), .DIN2 (__9_____26623), .Q
       (_________28547));
  nor2s1 _____9_441570(.DIN1 (____0____28172), .DIN2 (______0__28485),
       .Q (_________28546));
  nor2s1 _____9_441571(.DIN1 (____0___23894), .DIN2 (_____9___28519),
       .Q (_________28545));
  nnd2s1 _____441572(.DIN1 (_________28486), .DIN2 (___0_____27902), .Q
       (_________28544));
  nor2s1 ____441573(.DIN1 (__9_9___26888), .DIN2 (_________28496), .Q
       (_________28543));
  nor2s1 ____9__441574(.DIN1 (___9____20680), .DIN2 (______9__28541),
       .Q (______0__28542));
  nor2s1 ____9__441575(.DIN1 (_________28458), .DIN2 (_________28482),
       .Q (_____9___28989));
  hi1s1 ____9__441576(.DIN (______0__28579), .Q (_____9___28607));
  xor2s1 _______441577(.DIN1 (_________28460), .DIN2
       (___________0___18872), .Q (_____9___28609));
  nnd2s1 ____90_441578(.DIN1 (______9__28541), .DIN2 (_________28581),
       .Q (_____9___28611));
  xnr2s1 _______441579(.DIN1 (______9__28503), .DIN2 (________23116),
       .Q (_________28540));
  nnd2s1 _______441580(.DIN1 (_________28469), .DIN2 (_________31303),
       .Q (_________28539));
  and2s1 _____9_441581(.DIN1 (_________28467), .DIN2 (_________28537),
       .Q (_________28538));
  nor2s1 _____0_441582(.DIN1 (_________28533), .DIN2 (_________28534),
       .Q (_________28536));
  nnd2s1 _______441583(.DIN1 (_________28534), .DIN2 (_________28533),
       .Q (_________28535));
  nnd2s1 _____9_441584(.DIN1 (_________28462), .DIN2 (_________28832),
       .Q (______0__28532));
  and2s1 _______441585(.DIN1 (_________29291), .DIN2 (_____0___28530),
       .Q (_____09__28531));
  nor2s1 ____90_441586(.DIN1 (________19427), .DIN2 (______9__28474),
       .Q (_________28584));
  nor2s1 _______441587(.DIN1 (_____0___28530), .DIN2 (_________29291),
       .Q (_________28565));
  nnd2s1 ______441588(.DIN1 (_____0___28529), .DIN2 (____0____28171),
       .Q (_________28592));
  nor2s1 _______441589(.DIN1 (outData[26]), .DIN2 (_________28509), .Q
       (_________28599));
  dffacs1 _______________________441590(.CLRB (reset), .CLK (clk), .DIN
       (_________28479), .QN (_____________________18614));
  dffacs1 ____0__________________441591(.CLRB (reset), .CLK (clk), .DIN
       (______0__28465), .QN (____0________________18595));
  hi1s1 ____9__441592(.DIN (_____0___28527), .Q (_____0___28528));
  nnd2s1 ____9_441593(.DIN1 (_________28452), .DIN2 (____0___21083), .Q
       (_____0___28526));
  nnd2s1 ____9__441594(.DIN1 (_________28463), .DIN2 (___0_0___27563),
       .Q (_____0___28525));
  or2s1 ____9__441595(.DIN1 (_________31154), .DIN2 (_____9___28516),
       .Q (_____0___28524));
  nnd2s1 ____9_441596(.DIN1 (_________28481), .DIN2 (_________28410),
       .Q (_____00__28523));
  nnd2s1 ____9__441597(.DIN1 (______9__28454), .DIN2 (____0___19303),
       .Q (_____99__28522));
  nnd2s1 ____9_441598(.DIN1 (_________28456), .DIN2 (___09_0__28051),
       .Q (_____9___28521));
  hi1s1 ____9_441599(.DIN (_____9___28519), .Q (_____9___28520));
  nnd2s1 ____9__441600(.DIN1 (______0__28455), .DIN2 (_____9___28517),
       .Q (_____9___28518));
  dffacs1 ______________0__0_(.CLRB (reset), .CLK (clk), .DIN
       (_________28470), .Q (__________0__0_));
  nnd2s1 ____90_441601(.DIN1 (_____9___28516), .DIN2 (_________28384),
       .Q (______0__28597));
  xor2s1 ____9_441602(.DIN1 (_____09__28434), .DIN2 (______0__31254),
       .Q (______0__28579));
  hi1s1 ____9__441603(.DIN (_____9___28515), .Q (_________29396));
  dffacs1 ____0__________________441604(.CLRB (reset), .CLK (clk), .DIN
       (_________28466), .QN (____0________________18591));
  nnd2s1 _______441605(.DIN1 (_________28507), .DIN2 (___0_____27327),
       .Q (_____9___28514));
  nnd2s1 _______441606(.DIN1 (_________28511), .DIN2 (____0____32823),
       .Q (______9__28513));
  nor2s1 _______441607(.DIN1 (______9__28405), .DIN2 (_________28511),
       .Q (_________28512));
  hi1s1 _______441608(.DIN (_________28509), .Q (_________28510));
  nnd2s1 ____9__441609(.DIN1 (_________28507), .DIN2 (________25836),
       .Q (_________28508));
  or2s1 _______441610(.DIN1 (____0____32823), .DIN2 (_________28448),
       .Q (_________28506));
  xor2s1 _______441611(.DIN1 (_____9___28419), .DIN2 (_____0___28427),
       .Q (_________28505));
  nor2s1 _______441612(.DIN1 (________23096), .DIN2 (______9__28503),
       .Q (______0__28504));
  nnd2s1 _____9_441613(.DIN1 (______0__28494), .DIN2 (____90__23074),
       .Q (_________28502));
  nnd2s1 _______441614(.DIN1 (_________28507), .DIN2 (__9_____27060),
       .Q (_________28501));
  nnd2s1 _______441615(.DIN1 (_________28439), .DIN2 (___09____28105),
       .Q (_________28500));
  nnd2s1 _____441616(.DIN1 (_________28450), .DIN2 (___0_____27720), .Q
       (_________28499));
  or2s1 _____9_441617(.DIN1 (_________28497), .DIN2 (_________28440),
       .Q (_________28498));
  hi1s1 _______441618(.DIN (_________28534), .Q (_________28557));
  xor2s1 _______441619(.DIN1 (_____________18900), .DIN2
       (_________28468), .Q (____9_0__29970));
  nnd2s1 ____90_441620(.DIN1 (_________28441), .DIN2 (_________28471),
       .Q (_________28559));
  dffacs1 _____________________9_441621(.CLRB (reset), .CLK (clk), .DIN
       (_________28446), .QN (_________________9___18669));
  nnd2s1 ____9_441622(.DIN1 (_____0___28433), .DIN2 (_________28294),
       .Q (_________28496));
  and2s1 ____9__441623(.DIN1 (______0__28494), .DIN2 (_________34772),
       .Q (_________28495));
  nor2s1 ____9__441624(.DIN1 (___9____26232), .DIN2 (_____0___28429),
       .Q (______9__28493));
  and2s1 ____9_441625(.DIN1 (_________28490), .DIN2 (_________28489),
       .Q (_________28491));
  xnr2s1 ____99_441626(.DIN1 (_________28737), .DIN2 (_________28453),
       .Q (_________28488));
  xor2s1 ____99_441627(.DIN1 (_________28413), .DIN2 (_________28269),
       .Q (_________28487));
  nor2s1 ____9__441628(.DIN1 (___0_____27284), .DIN2 (_____0___28428),
       .Q (_________28486));
  nnd2s1 ____9_441629(.DIN1 (_________28437), .DIN2 (___0_____27473),
       .Q (______0__28485));
  or2s1 ____9__441630(.DIN1 (_________28483), .DIN2 (_________28447),
       .Q (______9__28484));
  hi1s1 ____9_441631(.DIN (_________28481), .Q (_________28482));
  nor2s1 ____9__441632(.DIN1 (___0____23471), .DIN2 (_____0___28432),
       .Q (_________28480));
  nor2s1 ____99_441633(.DIN1 (___0_____27483), .DIN2 (_____0___28431),
       .Q (_____9___28519));
  hi1s1 ____9__441634(.DIN (_____9___28516), .Q (______9__28541));
  xor2s1 ____9__441635(.DIN1 (_________28473), .DIN2 (___0____19841),
       .Q (_____9___28515));
  nnd2s1 ____9__441636(.DIN1 (_________28436), .DIN2 (_________28459),
       .Q (_____0___28527));
  dffacs1 ______________________0_441637(.CLRB (reset), .CLK (clk),
       .DIN (______0__28445), .QN (__________________0_));
  dffacs1 ____0___________________441638(.CLRB (reset), .CLK (clk),
       .DIN (_____0___28430), .QN (____0_______________));
  nnd2s1 _____9_441639(.DIN1 (_____9___28421), .DIN2 (_________28478),
       .Q (_________28479));
  nor2s1 _______441640(.DIN1 (_________28476), .DIN2 (______0__28475),
       .Q (_________28477));
  nor2s1 ____9__441641(.DIN1 (________19426), .DIN2 (_________28473),
       .Q (______9__28474));
  xor2s1 ____9__441642(.DIN1 (_________28442), .DIN2 (_________28471),
       .Q (_________28472));
  nor2s1 ____9__441643(.DIN1 (_________34187), .DIN2 (_____00__28425),
       .Q (_________28470));
  nor2s1 _______441644(.DIN1 (____0___23978), .DIN2 (_____99__28424),
       .Q (_________28469));
  xor2s1 ____9__441645(.DIN1 (_________28388), .DIN2 (_____0___33866),
       .Q (_____0___28529));
  nnd2s1 _______441646(.DIN1 (_________28468), .DIN2
       (_____________18900), .Q (_________28509));
  or2s1 _______441647(.DIN1 (_________28368), .DIN2 (_________28468),
       .Q (_____9___29899));
  xor2s1 _______441648(.DIN1 (_________28403), .DIN2 (_________28313),
       .Q (_________28534));
  dffacs1 ______________________0_441649(.CLRB (reset), .CLK (clk),
       .DIN (_________28408), .Q (__________________0___18643));
  xor2s1 ____9__441650(.DIN1 (______0__28386), .DIN2 (_____0___29178),
       .Q (_________29291));
  nor2s1 ____9__441651(.DIN1 (_________28497), .DIN2 (_____9___28420),
       .Q (_________28467));
  nnd2s1 ____9__441652(.DIN1 (_____9___28422), .DIN2 (________23875),
       .Q (_________28466));
  or2s1 ____9__441653(.DIN1 (______9__28464), .DIN2 (_________28414),
       .Q (______0__28465));
  nor2s1 ____9__441654(.DIN1 (________23919), .DIN2 (______9__28415),
       .Q (_________28463));
  nor2s1 ____9__441655(.DIN1 (_________28461), .DIN2 (_____9___28418),
       .Q (_________28462));
  nnd2s1 ____441656(.DIN1 (______0__28435), .DIN2 (_________28459), .Q
       (_________28460));
  nor2s1 ____0__441657(.DIN1 (_________28457), .DIN2 (_________28411),
       .Q (_________28458));
  nor2s1 ____441658(.DIN1 (_________28461), .DIN2 (_____90__28416), .Q
       (_________28456));
  nor2s1 ____00_441659(.DIN1 (__9_____26659), .DIN2 (_________28412),
       .Q (______0__28455));
  nnd2s1 ____0_441660(.DIN1 (_________28453), .DIN2 (____0___19304), .Q
       (______9__28454));
  nor2s1 ____0__441661(.DIN1 (_________28451), .DIN2 (_________28453),
       .Q (_________28452));
  xor2s1 ____9__441662(.DIN1 (_________28387), .DIN2 (_____0___31450),
       .Q (_________28481));
  xor2s1 ____99_441663(.DIN1 (______0__28376), .DIN2 (_________32554),
       .Q (_____9___28516));
  dffacs2 ____0________________0_441664(.CLRB (reset), .CLK (clk), .DIN
       (_________28409), .Q (____0____________0_));
  nor2s1 ____9__441665(.DIN1 (_____0__26057), .DIN2 (_________28407),
       .Q (_________28450));
  xor2s1 _______441666(.DIN1 (_________28370), .DIN2 (_________32081),
       .Q (_________28449));
  nnd2s1 _____9_441667(.DIN1 (_________28438), .DIN2 (____0____28199),
       .Q (_________28448));
  nnd2s1 ____9__441668(.DIN1 (_________28393), .DIN2 (____0____28179),
       .Q (_________28447));
  nnd2s1 ____9__441669(.DIN1 (______0__28396), .DIN2 (__9__0__26394),
       .Q (_________28446));
  nnd2s1 ____9__441670(.DIN1 (_________28399), .DIN2 (______9__28444),
       .Q (______0__28445));
  and2s1 ____9__441671(.DIN1 (_________28442), .DIN2 (______0__34471),
       .Q (_________28443));
  or2s1 ____9__441672(.DIN1 (______0__34471), .DIN2 (_________28442),
       .Q (_________28441));
  or2s1 ____9_441673(.DIN1 (________24904), .DIN2 (_________28401), .Q
       (_________28440));
  nor2s1 ____9__441674(.DIN1 (___0_____27921), .DIN2 (_________28402),
       .Q (_________28439));
  nor2s1 ____90_441675(.DIN1 (___090___28045), .DIN2 (_________28438),
       .Q (_________28511));
  nor2s1 ____9__441676(.DIN1 (___0_____27778), .DIN2 (_________28398),
       .Q (______0__28494));
  nnd2s1 ____9__441677(.DIN1 (_________28404), .DIN2 (______0__34748),
       .Q (______9__28503));
  xor2s1 ____9_441678(.DIN1 (_________28362), .DIN2 (_________33144),
       .Q (_____0___29809));
  dffacs1 _______________________441679(.CLRB (reset), .CLK (clk), .DIN
       (_________28380), .QN (_____________________18615));
  nor2s1 ____00_441680(.DIN1 (___0_____27406), .DIN2 (_________28382),
       .Q (_________28437));
  nnd2s1 ____9__441681(.DIN1 (______0__28435), .DIN2 (____9___25551),
       .Q (_________28436));
  xor2s1 ____0__441682(.DIN1 (_________28345), .DIN2 (_________28939),
       .Q (_____09__28434));
  nor2s1 ____0__441683(.DIN1 (___0_____27804), .DIN2 (______9__28385),
       .Q (_____0___28433));
  nnd2s1 ____0__441684(.DIN1 (_________28377), .DIN2 (________21402),
       .Q (_____0___28432));
  nnd2s1 ____00_441685(.DIN1 (_________28391), .DIN2 (__9_____26496),
       .Q (_____0___28431));
  nnd2s1 ____441686(.DIN1 (_________28383), .DIN2 (_________28626), .Q
       (_____0___28430));
  nor2s1 ____9__441687(.DIN1 (__9_____26953), .DIN2 (_________28394),
       .Q (_____0___28429));
  nnd2s1 ____00_441688(.DIN1 (_________28378), .DIN2 (________23921),
       .Q (_____0___28428));
  nnd2s1 ____99_441689(.DIN1 (_________28442), .DIN2 (_____0___28426),
       .Q (_________28489));
  nnd2s1 ____9_441690(.DIN1 (_________28390), .DIN2 (_____0___28427),
       .Q (_________28492));
  or2s1 ____9__441691(.DIN1 (_____0___28426), .DIN2 (_________28442),
       .Q (_________28490));
  nnd2s1 ____99_441692(.DIN1 (______9__28395), .DIN2 (___0____25288),
       .Q (_________28507));
  nor2s1 ____0__441693(.DIN1 (_____9___28325), .DIN2 (_________28379),
       .Q (_________31306));
  dffacs1 ________________________441694(.CLRB (reset), .CLK (clk),
       .DIN (_________28397), .QN (____________________));
  xor2s1 ____9_441695(.DIN1 (_____9___28324), .DIN2 (_________28251),
       .Q (_____00__28425));
  nor2s1 ____9__441696(.DIN1 (_____9___30454), .DIN2 (_________28369),
       .Q (_____99__28424));
  xor2s1 ____9__441697(.DIN1 (___9_0__21608), .DIN2 (____0____32816),
       .Q (_____9___28423));
  nor2s1 ____0_441698(.DIN1 (______9__28464), .DIN2 (_________28354),
       .Q (_____9___28422));
  nor2s1 ____9__441699(.DIN1 (_________28667), .DIN2 (_________28372),
       .Q (_____9___28421));
  or2s1 ____00_441700(.DIN1 (___09____28066), .DIN2 (______0__28358),
       .Q (_____9___28420));
  xor2s1 ____99_441701(.DIN1 (_________28389), .DIN2 (_________28363),
       .Q (_____9___28419));
  nnd2s1 ____00_441702(.DIN1 (_________28352), .DIN2 (____0____28219),
       .Q (_____9___28418));
  hi1s1 ____9__441703(.DIN (_____9___28417), .Q (______0__28475));
  xnr2s1 ____9__441704(.DIN1 (_________33384), .DIN2 (_________28341),
       .Q (_________28468));
  nnd2s1 ____0_441705(.DIN1 (_________28350), .DIN2 (___09____28113),
       .Q (_____90__28416));
  nnd2s1 ____0__441706(.DIN1 (_________28351), .DIN2 (__9__9__27043),
       .Q (______9__28415));
  or2s1 ____0__441707(.DIN1 (___0_____27783), .DIN2 (_________28360),
       .Q (_________28414));
  nnd2s1 ____441708(.DIN1 (_________28349), .DIN2 (_________28268), .Q
       (_________28413));
  nnd2s1 ____09_441709(.DIN1 (_________28359), .DIN2 (__9_____26629),
       .Q (_________28412));
  hi1s1 ____0_441710(.DIN (_________28410), .Q (_________28411));
  nnd2s1 ____0__441711(.DIN1 (_________28355), .DIN2 (_________28353),
       .Q (_________28409));
  nnd2s1 ____0__441712(.DIN1 (_________28346), .DIN2 (__9_____26471),
       .Q (_________28408));
  xor2s1 ____0_441713(.DIN1 (_____9___28323), .DIN2 (______0__30607),
       .Q (_________28459));
  xor2s1 ____0_441714(.DIN1 (_________28312), .DIN2 (____0____32777),
       .Q (____9____32681));
  nor2s1 ____0__441715(.DIN1 (________19280), .DIN2 (______9__28357),
       .Q (_________28473));
  nnd2s1 _____0_441716(.DIN1 (______9__28347), .DIN2 (_________28344),
       .Q (_________28453));
  nnd2s1 ____0__441717(.DIN1 (_____0___28338), .DIN2 (_________28381),
       .Q (_________28407));
  and2s1 ____9__441718(.DIN1 (____0____32816), .DIN2 (_________34447),
       .Q (______0__28406));
  nor2s1 ____9__441719(.DIN1 (_________28392), .DIN2 (____0____28201),
       .Q (______9__28405));
  nnd2s1 ____9__441720(.DIN1 (_____0___28334), .DIN2 (_________31336),
       .Q (_________28404));
  xor2s1 ____99_441721(.DIN1 (_________28306), .DIN2 (____9____31798),
       .Q (_________28403));
  nnd2s1 ____00_441722(.DIN1 (_____0___28333), .DIN2 (___0_90__27938),
       .Q (_________28402));
  nnd2s1 ____0__441723(.DIN1 (_____9___28327), .DIN2 (____09___28232),
       .Q (_________28401));
  nor2s1 ____9__441724(.DIN1 (_________34447), .DIN2 (____0____32816),
       .Q (_________28400));
  nor2s1 ____0__441725(.DIN1 (________24121), .DIN2 (_____0___28336),
       .Q (_________28399));
  nnd2s1 ____0__441726(.DIN1 (_____09__28339), .DIN2 (____0___25470),
       .Q (_________28398));
  nnd2s1 ____0__441727(.DIN1 (_________28340), .DIN2 (______9__28444),
       .Q (_________28397));
  nor2s1 ____0_441728(.DIN1 (___00____27233), .DIN2 (_____0___28335),
       .Q (______0__28396));
  nor2s1 ____0__441729(.DIN1 (__9_9___26416), .DIN2 (_____9___28328),
       .Q (______9__28395));
  nnd2s1 ____0__441730(.DIN1 (_____99__28330), .DIN2 (________25905),
       .Q (_________28394));
  nor2s1 ____0_441731(.DIN1 (___0____25284), .DIN2 (_________28342), .Q
       (_________28393));
  xor2s1 ____9__441732(.DIN1 (____9_9__29949), .DIN2 (_________29500),
       .Q (_____9___28417));
  nnd2s1 ____9__441733(.DIN1 (____0____28200), .DIN2 (_________28392),
       .Q (_________28438));
  nor2s1 ____0__441734(.DIN1 (__90_9__26308), .DIN2 (_________28317),
       .Q (_________28391));
  nnd2s1 ____0__441735(.DIN1 (_________28389), .DIN2 (___09____28082),
       .Q (_________28390));
  nor2s1 ____0__441736(.DIN1 (___09____28122), .DIN2 (_________28314),
       .Q (_________28388));
  nor2s1 ____09_441737(.DIN1 (_________28373), .DIN2 (_________28374),
       .Q (_________28387));
  xor2s1 ____0__441738(.DIN1 (_________33264), .DIN2 (_________28356),
       .Q (______0__28386));
  nnd2s1 ____0__441739(.DIN1 (______0__28311), .DIN2 (_____9__22117),
       .Q (______9__28385));
  nnd2s1 ____0__441740(.DIN1 (______9__28375), .DIN2 (outData[26]), .Q
       (_________28384));
  nor2s1 ____0__441741(.DIN1 (______9__28301), .DIN2 (_____90__28321),
       .Q (_________28383));
  nnd2s1 ____0__441742(.DIN1 (_________28319), .DIN2 (_________28381),
       .Q (_________28382));
  nnd2s1 ____0_441743(.DIN1 (_____0___28332), .DIN2 (______9__28444),
       .Q (_________28380));
  nor2s1 ____0__441744(.DIN1 (_____________18900), .DIN2
       (_________28316), .Q (_________28379));
  nor2s1 ____0__441745(.DIN1 (________23120), .DIN2 (_____9___28322),
       .Q (_________28378));
  nor2s1 ____0__441746(.DIN1 (________26000), .DIN2 (_________28318),
       .Q (_________28377));
  nor2s1 ____0__441747(.DIN1 (outData[26]), .DIN2 (______9__28375), .Q
       (______0__28376));
  nnd2s1 _____0_441748(.DIN1 (_________28374), .DIN2 (_________28373),
       .Q (_________28410));
  xor2s1 ____0__441749(.DIN1 (_________28296), .DIN2 (_____9___33022),
       .Q (______0__28435));
  nor2s1 _____0_441750(.DIN1 (_________28270), .DIN2 (______0__28348),
       .Q (______0__28810));
  xnr2s1 ____0__441751(.DIN1 (_________29253), .DIN2 (_____9___34513),
       .Q (_________28442));
  nnd2s1 ____0__441752(.DIN1 (_________28309), .DIN2 (________24474),
       .Q (_________28372));
  nnd2s1 ____9__441753(.DIN1 (____9_9__29949), .DIN2
       (________________18756), .Q (_________28371));
  nnd2s1 ____9__441754(.DIN1 (____9_9__29949), .DIN2 (_________28476),
       .Q (_________28370));
  xor2s1 ____9__441755(.DIN1 (_________28285), .DIN2 (_________28289),
       .Q (_________28369));
  nor2s1 ____00_441756(.DIN1 (_____________18899), .DIN2
       (_________28361), .Q (_________28368));
  or2s1 ____9__441757(.DIN1 (________________18756), .DIN2
       (____9_9__29949), .Q (_________28367));
  nnd2s1 ____0__441758(.DIN1 (_____9___28326), .DIN2 (_________28363),
       .Q (_________28364));
  nor2s1 ____0__441759(.DIN1 (_________28286), .DIN2 (_________28361),
       .Q (_________28362));
  nnd2s1 ____0__441760(.DIN1 (______0__28302), .DIN2 (__9_____27041),
       .Q (_________28360));
  nnd2s1 _____0_441761(.DIN1 (_________28293), .DIN2 (___0____21654),
       .Q (_________28359));
  nnd2s1 ____0__441762(.DIN1 (_________28299), .DIN2 (_____9___34826),
       .Q (______0__28358));
  nor2s1 ____0__441763(.DIN1 (________19279), .DIN2 (_________28356),
       .Q (______9__28357));
  and2s1 ____0__441764(.DIN1 (_________28308), .DIN2 (_____9__25040),
       .Q (_________28355));
  nnd2s1 ____0__441765(.DIN1 (_________28307), .DIN2 (_________28353),
       .Q (_________28354));
  nor2s1 ____0__441766(.DIN1 (_____0___34930), .DIN2 (_________28297),
       .Q (_________28352));
  nor2s1 ____0_441767(.DIN1 (___0____22596), .DIN2 (_________28295), .Q
       (_________28351));
  nor2s1 _______441768(.DIN1 (___0_____27711), .DIN2 (______0__28292),
       .Q (_________28350));
  hi1s1 _______441769(.DIN (______0__28348), .Q (_________28349));
  nnd2s1 ______441770(.DIN1 (_________28343), .DIN2 (_________28939),
       .Q (______9__28347));
  nor2s1 _______441771(.DIN1 (__9_0___26519), .DIN2 (_________28300),
       .Q (_________28346));
  and2s1 _______441772(.DIN1 (_________28344), .DIN2 (_________28343),
       .Q (_________28345));
  nnd2s1 ____0_441773(.DIN1 (_________28280), .DIN2 (___0____24414), .Q
       (_________28342));
  nor2s1 ____0_441774(.DIN1 (outData[24]), .DIN2 (_________28304), .Q
       (_________28341));
  and2s1 ____09_441775(.DIN1 (_________28276), .DIN2 (_________28537),
       .Q (_________28340));
  nor2s1 ____09_441776(.DIN1 (__90____26265), .DIN2 (_____9___28329),
       .Q (_____09__28339));
  and2s1 ____0__441777(.DIN1 (______9__28282), .DIN2 (_____0___28337),
       .Q (_____0___28338));
  nnd2s1 ____0__441778(.DIN1 (_________28277), .DIN2 (____0_9__28185),
       .Q (_____0___28336));
  nnd2s1 ____0__441779(.DIN1 (_________28274), .DIN2 (___099__25366),
       .Q (_____0___28335));
  nnd2s1 ____441780(.DIN1 (_________28288), .DIN2 (________25410), .Q
       (_____0___28334));
  nor2s1 ____0__441781(.DIN1 (________24959), .DIN2 (_________28281),
       .Q (_____0___28333));
  nor2s1 ____0__441782(.DIN1 (_____00__28331), .DIN2 (_________28279),
       .Q (_____0___28332));
  nor2s1 ____0_441783(.DIN1 (___99___26240), .DIN2 (_____9___28329), .Q
       (_____99__28330));
  nnd2s1 ____0__441784(.DIN1 (______0__28273), .DIN2 (__9_____26389),
       .Q (_____9___28328));
  nor2s1 ____0__441785(.DIN1 (________24038), .DIN2 (______9__28291),
       .Q (_____9___28327));
  hi1s1 ____0__441786(.DIN (_____9___28326), .Q (_________28389));
  nnd2s1 ____0_441787(.DIN1 (_________28290), .DIN2 (_________28284),
       .Q (_________28392));
  hi1s1 ____0__441788(.DIN (______9__29651), .Q (____0____32816));
  nor2s1 _______441789(.DIN1 (____0___21818), .DIN2 (_________28315),
       .Q (_____9___28325));
  nor2s1 _____441790(.DIN1 (_________28252), .DIN2 (______9__28310), .Q
       (_____9___28324));
  nor2s1 ______441791(.DIN1 (___0__0__27762), .DIN2 (_________28260),
       .Q (_____9___28323));
  nnd2s1 _____441792(.DIN1 (_________28264), .DIN2 (________23576), .Q
       (_____9___28322));
  or2s1 _______441793(.DIN1 (______9__28320), .DIN2 (_________28261),
       .Q (_____90__28321));
  nor2s1 _______441794(.DIN1 (___0__9__27819), .DIN2 (_________28266),
       .Q (_________28319));
  nnd2s1 _______441795(.DIN1 (_________28265), .DIN2 (__9_____26489),
       .Q (_________28318));
  nnd2s1 ______441796(.DIN1 (_________28267), .DIN2 (___0_____27600),
       .Q (_________28317));
  nnd2s1 ______441797(.DIN1 (_________28315), .DIN2 (_________35086),
       .Q (_________28316));
  nor2s1 ____09_441798(.DIN1 (_________28313), .DIN2 (______9__28272),
       .Q (_________28314));
  or2s1 _______441799(.DIN1 (_____0___28236), .DIN2 (_________28315),
       .Q (_________28312));
  nor2s1 _______441800(.DIN1 (__9__0__26637), .DIN2 (_________28258),
       .Q (______0__28311));
  or2s1 _______441801(.DIN1 (_____0___28239), .DIN2 (_________28920),
       .Q (_________28373));
  xor2s1 _______441802(.DIN1 (____09___28229), .DIN2 (_________28365),
       .Q (______0__28348));
  nnd2s1 _______441803(.DIN1 (_________28315), .DIN2
       (_____________18900), .Q (______9__28375));
  nor2s1 _____0_441804(.DIN1 (______9__28253), .DIN2 (______9__28310),
       .Q (_________28684));
  dffacs1 _______________________441805(.CLRB (reset), .CLK (clk), .DIN
       (_________34750), .QN (_____________________18668));
  dffacs1 _______________________441806(.CLRB (reset), .CLK (clk), .DIN
       (_________28275), .QN (_____________________18665));
  nor2s1 ____0__441807(.DIN1 (______0__28263), .DIN2 (______0__28254),
       .Q (_________28309));
  nor2s1 ______441808(.DIN1 (________22796), .DIN2 (_____0___28242), .Q
       (_________28308));
  nor2s1 _____0_441809(.DIN1 (___0_____27968), .DIN2 (______0__28244),
       .Q (_________28307));
  nor2s1 ____09_441810(.DIN1 (_________28271), .DIN2 (_________28256),
       .Q (_________28306));
  xor2s1 _____0_441811(.DIN1 (____0_0__28206), .DIN2 (_________28305),
       .Q (_____9___28326));
  nor2s1 ____09_441812(.DIN1 (_________28305), .DIN2 (_________28255),
       .Q (_________28366));
  hi1s1 ____0_441813(.DIN (_________28304), .Q (_________28361));
  xor2s1 ____0__441814(.DIN1 (________25697), .DIN2 (_________28287),
       .Q (______9__29651));
  hi1s1 ____0__441815(.DIN (_________28303), .Q (______0__31456));
  nb1s1 ____0__441816(.DIN (_________28303), .Q (____9_9__29949));
  dffacs1 _______________________441817(.CLRB (reset), .CLK (clk), .DIN
       (_____09__28243), .QN (_____________________18664));
  nor2s1 _______441818(.DIN1 (______9__28301), .DIN2 (_____0___28237),
       .Q (______0__28302));
  nor2s1 _______441819(.DIN1 (___0_____27696), .DIN2 (____099__28234),
       .Q (_________28300));
  and2s1 _______441820(.DIN1 (_____0___28238), .DIN2 (_________28298),
       .Q (_________28299));
  nnd2s1 _______441821(.DIN1 (_________28247), .DIN2 (____0____28221),
       .Q (_________28297));
  nor2s1 _______441822(.DIN1 (___0_____27669), .DIN2 (_________28259),
       .Q (_________28296));
  nnd2s1 _______441823(.DIN1 (_____0___28240), .DIN2 (_________28294),
       .Q (_________28295));
  nor2s1 _______441824(.DIN1 (__9_____26660), .DIN2 (_____00__28235),
       .Q (_________28293));
  nnd2s1 _______441825(.DIN1 (____09___28233), .DIN2 (___9____25223),
       .Q (______0__28292));
  nnd2s1 _______441826(.DIN1 (____09___28231), .DIN2 (_________28661),
       .Q (_________28343));
  nor2s1 ______441827(.DIN1 (_________28245), .DIN2 (_________28250),
       .Q (_________28356));
  dffacs1 ____0__________________441828(.CLRB (reset), .CLK (clk), .DIN
       (_____0___28241), .QN (____0________________18594));
  nnd2s1 _______441829(.DIN1 (____09___28226), .DIN2 (____0___23713),
       .Q (______9__28291));
  nnd2s1 ____0_441830(.DIN1 (______0__28283), .DIN2 (_________28289),
       .Q (_________28290));
  nnd2s1 ____0__441831(.DIN1 (_________28287), .DIN2 (___0_0__25310),
       .Q (_________28288));
  xor2s1 ____0__441832(.DIN1 (____0_0__28196), .DIN2 (_________35086),
       .Q (_________28286));
  and2s1 ____09_441833(.DIN1 (_________28284), .DIN2 (______0__28283),
       .Q (_________28285));
  and2s1 _______441834(.DIN1 (____0____28217), .DIN2 (___0__0__27890),
       .Q (______9__28282));
  nnd2s1 _______441835(.DIN1 (____0_9__28214), .DIN2 (____9___25553),
       .Q (_________28281));
  nor2s1 _______441836(.DIN1 (___9____23417), .DIN2 (____0_9__28224),
       .Q (_________28280));
  nnd2s1 _______441837(.DIN1 (____0____28223), .DIN2 (_________28278),
       .Q (_________28279));
  and2s1 _______441838(.DIN1 (____0____28222), .DIN2 (___0_____27780),
       .Q (_________28277));
  and2s1 _______441839(.DIN1 (____0____28220), .DIN2 (_________28832),
       .Q (_________28276));
  nnd2s1 _______441840(.DIN1 (____09___28227), .DIN2 (___0_____27912),
       .Q (_________28275));
  nor2s1 _______441841(.DIN1 (___0__9__27520), .DIN2 (____0____28216),
       .Q (_________28274));
  xor2s1 ____0__441842(.DIN1 (____0____28198), .DIN2 (_________29253),
       .Q (_________28303));
  xor2s1 _____0_441843(.DIN1 (____0____28194), .DIN2 (_________35002),
       .Q (_________28304));
  nor2s1 _______441844(.DIN1 (________25148), .DIN2 (____0_0__28215),
       .Q (______0__28273));
  nor2s1 ______441845(.DIN1 (____0____28218), .DIN2 (_________28271),
       .Q (______9__28272));
  and2s1 _____0_441846(.DIN1 (_________28269), .DIN2 (_________28268),
       .Q (_________28270));
  nor2s1 _____441847(.DIN1 (___0_0__24362), .DIN2 (____0____28212), .Q
       (_________28267));
  nnd2s1 _______441848(.DIN1 (____0____28213), .DIN2 (________23110),
       .Q (_________28266));
  and2s1 ______441849(.DIN1 (____0____28207), .DIN2 (_________35074),
       .Q (_________28265));
  nor2s1 _______441850(.DIN1 (______0__28263), .DIN2 (____0_9__28205),
       .Q (_________28264));
  nnd2s1 _______441851(.DIN1 (____0____28204), .DIN2 (___09____28123),
       .Q (______9__28262));
  nnd2s1 _____441852(.DIN1 (____0____28211), .DIN2 (_____0__23656), .Q
       (_________28261));
  hi1s1 _____9_441853(.DIN (_________28259), .Q (_________28260));
  nnd2s1 _____9_441854(.DIN1 (____0____28203), .DIN2 (___9____25233),
       .Q (_________28258));
  nnd2s1 _______441855(.DIN1 (____09___28230), .DIN2
       (______________________________________0___________), .Q
       (_________28344));
  nor2s1 _______441856(.DIN1 (___9____26179), .DIN2 (____090__28225),
       .Q (_____9___28329));
  xor2s1 _______441857(.DIN1 (____0____28170), .DIN2 (____9____31746),
       .Q (______9__28310));
  nor2s1 ______441858(.DIN1 (____0____28210), .DIN2 (________25533), .Q
       (_________28920));
  nor2s1 _____9_441859(.DIN1 (outData[24]), .DIN2 (____0____28209), .Q
       (_________28315));
  xor2s1 ____0__441860(.DIN1 (______0__29502), .DIN2 (_________32644),
       .Q (_________28257));
  nor2s1 ______441861(.DIN1 (_________________0___18597), .DIN2
       (____0____28193), .Q (_________28256));
  xor2s1 _______441862(.DIN1 (___0999__28137), .DIN2 (____9____31798),
       .Q (_________28255));
  nnd2s1 _______441863(.DIN1 (____0____28192), .DIN2 (_________28537),
       .Q (______0__28254));
  nor2s1 _______441864(.DIN1 (_________28252), .DIN2 (_________28251),
       .Q (______9__28253));
  nor2s1 _______441865(.DIN1 (_________33278), .DIN2 (____0____28188),
       .Q (_________28250));
  nnd2s1 _______441866(.DIN1 (_________28248), .DIN2 (______0__34451),
       .Q (_________28249));
  and2s1 _______441867(.DIN1 (____0_0__28186), .DIN2 (_________28478),
       .Q (_________28247));
  or2s1 _______441868(.DIN1 (______0__34451), .DIN2 (_________28248),
       .Q (_________28246));
  nor2s1 _______441869(.DIN1 (________24923), .DIN2 (____0____28190),
       .Q (_________28245));
  nnd2s1 ______441870(.DIN1 (____0____28189), .DIN2 (____0____28183),
       .Q (______0__28244));
  or2s1 _______441871(.DIN1 (___0_____27698), .DIN2 (____0____28182),
       .Q (_____09__28243));
  nnd2s1 _______441872(.DIN1 (____0____28191), .DIN2 (____00__22989),
       .Q (_____0___28242));
  nnd2s1 _____9_441873(.DIN1 (____0____28184), .DIN2 (___09____28103),
       .Q (_____0___28241));
  nor2s1 _____9_441874(.DIN1 (________24833), .DIN2 (____0____28173),
       .Q (_____0___28240));
  nor2s1 _____0_441875(.DIN1 (_________18854), .DIN2 (________25534),
       .Q (_____0___28239));
  nor2s1 ______441876(.DIN1 (___0__0__28004), .DIN2 (____0____28180),
       .Q (_____0___28238));
  nnd2s1 _______441877(.DIN1 (____0____28178), .DIN2 (________25476),
       .Q (_____0___28237));
  nor2s1 _______441878(.DIN1 (_____________18899), .DIN2
       (____0____28208), .Q (_____0___28236));
  nnd2s1 _______441879(.DIN1 (____0_0__28168), .DIN2 (________25380),
       .Q (_____00__28235));
  nnd2s1 _______441880(.DIN1 (____0_9__28167), .DIN2 (___9____26235),
       .Q (____099__28234));
  and2s1 _______441881(.DIN1 (____0____28165), .DIN2 (____09___28232),
       .Q (____09___28233));
  hi1s1 _______441882(.DIN (____09___28230), .Q (____09___28231));
  nnd2s1 _____441883(.DIN1 (____09___28228), .DIN2
       (______________18867), .Q (____09___28229));
  nnd2s1 ______441884(.DIN1 (____0____28181), .DIN2 (___09____28127),
       .Q (_________28259));
  dffacs1 ____0_________________0_441885(.CLRB (reset), .CLK (clk),
       .DIN (____0____28187), .QN (____0_____________0_));
  nor2s1 _______441886(.DIN1 (___0_____27811), .DIN2 (____00___28144),
       .Q (____09___28227));
  nor2s1 _____0_441887(.DIN1 (___09_9__28080), .DIN2 (____0____28149),
       .Q (____09___28226));
  nnd2s1 _____0_441888(.DIN1 (____00___28142), .DIN2 (________21920),
       .Q (____090__28225));
  nnd2s1 _______441889(.DIN1 (____0_0__28148), .DIN2 (___9____25224),
       .Q (____0_9__28224));
  nor2s1 _______441890(.DIN1 (________23187), .DIN2 (____00___28146),
       .Q (____0____28223));
  and2s1 _______441891(.DIN1 (____0____28154), .DIN2 (____0____28221),
       .Q (____0____28222));
  and2s1 ______441892(.DIN1 (____00___28145), .DIN2 (____0____28219),
       .Q (____0____28220));
  nor2s1 _____0_441893(.DIN1 (_________________0___18597), .DIN2
       (____0____28152), .Q (____0____28218));
  nor2s1 _______441894(.DIN1 (________24929), .DIN2 (____0____28150),
       .Q (____0____28217));
  nnd2s1 _____9_441895(.DIN1 (____00___28140), .DIN2 (________24742),
       .Q (____0____28216));
  nnd2s1 _____0_441896(.DIN1 (___099___28132), .DIN2 (___99___25268),
       .Q (____0_0__28215));
  nor2s1 _____0_441897(.DIN1 (____0___23179), .DIN2 (____00___28141),
       .Q (____0_9__28214));
  xor2s1 _______441898(.DIN1 (___09_9__28119), .DIN2 (_____0___33866),
       .Q (______0__28283));
  xor2s1 ______441899(.DIN1 (___09_0__28120), .DIN2 (________19986), .Q
       (_________28284));
  nnd2s1 ______441900(.DIN1 (____0____28160), .DIN2 (__90____26256), .Q
       (_________28287));
  nor2s1 _______441901(.DIN1 (________23106), .DIN2 (___099___28133),
       .Q (____0____28213));
  nnd2s1 _______441902(.DIN1 (____00___28143), .DIN2 (__90____26310),
       .Q (____0____28212));
  nor2s1 _______441903(.DIN1 (________22929), .DIN2 (___0990__28128),
       .Q (____0____28211));
  hi1s1 _______441904(.DIN (_________18854), .Q (____0____28210));
  hi1s1 _______441905(.DIN (____0____28208), .Q (____0____28209));
  nor2s1 _______441906(.DIN1 (____90__26137), .DIN2 (___099___28131),
       .Q (____0____28207));
  xor2s1 _______441907(.DIN1 (____0____28169), .DIN2 (____000__28138),
       .Q (____0_0__28206));
  or2s1 _______441908(.DIN1 (___0_9___27940), .DIN2 (___099___28135),
       .Q (____0_9__28205));
  nor2s1 ______441909(.DIN1 (___0_____27930), .DIN2 (___099___28129),
       .Q (____0____28204));
  nor2s1 _______441910(.DIN1 (____09__24071), .DIN2 (___099___28134),
       .Q (____0____28203));
  xor2s1 _____9_441911(.DIN1 (___09____28108), .DIN2 (______0__35078),
       .Q (____09___28230));
  nnd2s1 _____9_441912(.DIN1 (____0____28202), .DIN2 (________26002),
       .Q (_________28268));
  nnd2s1 _______441913(.DIN1 (____0_9__28195), .DIN2 (____009__28147),
       .Q (_____9___29708));
  xor2s1 _______441914(.DIN1 (outData[23]), .DIN2 (____0____28163), .Q
       (____0____30938));
  and2s1 _______441915(.DIN1 (____0____28200), .DIN2 (____0____28199),
       .Q (____0____28201));
  xor2s1 _______441916(.DIN1 (____0____28159), .DIN2 (_________28866),
       .Q (____0____28198));
  nor2s1 ______441917(.DIN1 (__9__0__26346), .DIN2 (___09____28125), .Q
       (____0____28197));
  nnd2s1 _______441918(.DIN1 (____0_9__28195), .DIN2 (outData[23]), .Q
       (____0_0__28196));
  nor2s1 ______441919(.DIN1 (outData[23]), .DIN2 (____0_9__28195), .Q
       (____0____28194));
  xor2s1 _____0_441920(.DIN1 (____9_9__29072), .DIN2 (___09____28121),
       .Q (____0____28193));
  nor2s1 _____441921(.DIN1 (___0_____27877), .DIN2 (___09____28124), .Q
       (____0____28192));
  nor2s1 _______441922(.DIN1 (________24842), .DIN2 (___09____28115),
       .Q (____0____28191));
  nor2s1 _______441923(.DIN1 (___090___28048), .DIN2 (___09____28116),
       .Q (____0____28190));
  nor2s1 ______441924(.DIN1 (___9____24319), .DIN2 (___09____28102), .Q
       (____0____28189));
  nor2s1 ______441925(.DIN1 (___0_____28027), .DIN2 (___09____28112),
       .Q (____0____28188));
  nnd2s1 _______441926(.DIN1 (___09____28104), .DIN2 (_________28626),
       .Q (____0____28187));
  and2s1 _______441927(.DIN1 (___09____28099), .DIN2 (____0_9__28185),
       .Q (____0_0__28186));
  and2s1 _______441928(.DIN1 (___09_9__28100), .DIN2 (____0____28183),
       .Q (____0____28184));
  nnd2s1 _______441929(.DIN1 (___09_0__28101), .DIN2 (___0__9__27879),
       .Q (____0____28182));
  dffacs1 ________________0_441930(.CLRB (reset), .CLK (clk), .DIN
       (___09____28098), .QN (_________18854));
  nor2s1 _______441931(.DIN1 (_________32644), .DIN2 (____0____28151),
       .Q (_________28271));
  nnd2s1 _______441932(.DIN1 (____0_0__28177), .DIN2 (_________29253),
       .Q (____0____28181));
  nnd2s1 _______441933(.DIN1 (___09____28106), .DIN2 (____0____28179),
       .Q (____0____28180));
  nor2s1 _______441934(.DIN1 (___0_9___27459), .DIN2 (___09____28107),
       .Q (____0____28178));
  and2s1 ______441935(.DIN1 (____0____28175), .DIN2 (____0____28174),
       .Q (____0____28176));
  or2s1 _______441936(.DIN1 (____0____28172), .DIN2 (___09____28118),
       .Q (____0____28173));
  or2s1 _______441937(.DIN1 (____0____28174), .DIN2 (____0____28175),
       .Q (____0____28171));
  or2s1 _______441938(.DIN1 (____0____28164), .DIN2 (____0____28169),
       .Q (____0____28170));
  nor2s1 _____0_441939(.DIN1 (__9__9__26843), .DIN2 (____0____28166),
       .Q (____0_0__28168));
  nor2s1 _____0_441940(.DIN1 (__9_____26724), .DIN2 (____0____28166),
       .Q (____0_9__28167));
  nor2s1 _______441941(.DIN1 (____0___25370), .DIN2 (___09____28109),
       .Q (____0____28165));
  hi1s1 _______441942(.DIN (____0____28202), .Q (____09___28228));
  and2s1 _______441943(.DIN1 (____0____28169), .DIN2 (____0____28164),
       .Q (_________28252));
  nor2s1 _______441944(.DIN1 (outData[23]), .DIN2 (____0____28163), .Q
       (____0____28208));
  and2s1 ______441945(.DIN1 (____0____28163), .DIN2 (___09____28072),
       .Q (_________28248));
  dffacs1 _______________________441946(.CLRB (reset), .CLK (clk), .DIN
       (___09____28114), .QN (_____________________18608));
  xor2s1 _______441947(.DIN1 (___09_9__28060), .DIN2 (___09____28095),
       .Q (____0____28162));
  xor2s1 _______441948(.DIN1 (___09_0__28061), .DIN2 (_____0___30999),
       .Q (____0____28161));
  nnd2s1 _______441949(.DIN1 (____0____28159), .DIN2 (___9_9__26176),
       .Q (____0____28160));
  nnd2s1 _______441950(.DIN1 (____0_9__28157), .DIN2 (____0____28155),
       .Q (____0_0__28158));
  nor2s1 _______441951(.DIN1 (____0____28155), .DIN2 (____0_9__28157),
       .Q (____0____28156));
  and2s1 _______441952(.DIN1 (___09____28092), .DIN2 (____0____28153),
       .Q (____0____28154));
  hi1s1 _______441953(.DIN (____0____28151), .Q (____0____28152));
  nnd2s1 ______441954(.DIN1 (___09____28083), .DIN2 (____0___23626), .Q
       (____0____28150));
  nnd2s1 _______441955(.DIN1 (___09_0__28091), .DIN2 (___0_____27873),
       .Q (____0____28149));
  nor2s1 ______441956(.DIN1 (______0__28263), .DIN2 (___09____28088),
       .Q (____0_0__28148));
  nnd2s1 ______441957(.DIN1 (___09____28094), .DIN2 (outData[22]), .Q
       (____009__28147));
  nnd2s1 _______441958(.DIN1 (___09_0__28081), .DIN2 (___09____28078),
       .Q (____00___28146));
  nor2s1 _______441959(.DIN1 (________23644), .DIN2 (___09____28087),
       .Q (____00___28145));
  nnd2s1 _______441960(.DIN1 (___09____28085), .DIN2 (________24743),
       .Q (____00___28144));
  nnd2s1 _______441961(.DIN1 (___09_9__28090), .DIN2 (__9_____27009),
       .Q (_________28251));
  nnd2s1 _____441962(.DIN1 (___09____28096), .DIN2 (___0_____28018), .Q
       (_____0___28427));
  xor2s1 _______441963(.DIN1 (___09____28056), .DIN2 (____90___33582),
       .Q (______0__29502));
  nor2s1 _____441964(.DIN1 (_________28636), .DIN2 (___09____28073), .Q
       (____00___28143));
  nor2s1 ______441965(.DIN1 (_____9__25918), .DIN2 (___09____28086), .Q
       (____00___28142));
  nnd2s1 _______441966(.DIN1 (___09____28079), .DIN2 (____0___22898),
       .Q (____00___28141));
  nor2s1 _______441967(.DIN1 (_________34810), .DIN2 (___09____28084),
       .Q (____00___28140));
  or2s1 _______441968(.DIN1 (____000__28138), .DIN2 (___099___28136),
       .Q (____00___28139));
  nnd2s1 _______441969(.DIN1 (___099___28136), .DIN2 (____000__28138),
       .Q (___0999__28137));
  nnd2s1 _______441970(.DIN1 (___09____28067), .DIN2 (___0__9__27839),
       .Q (___099___28135));
  nnd2s1 _______441971(.DIN1 (___09____28069), .DIN2 (_________34884),
       .Q (___099___28134));
  nnd2s1 _____0_441972(.DIN1 (___09_0__28071), .DIN2 (________23160),
       .Q (___099___28133));
  nor2s1 _______441973(.DIN1 (___00___24334), .DIN2 (___09____28077),
       .Q (___099___28132));
  nnd2s1 _______441974(.DIN1 (___09____28097), .DIN2 (__9_____26870),
       .Q (___099___28131));
  nnd2s1 _______441975(.DIN1 (___09____28068), .DIN2 (____9___24979),
       .Q (___099___28130));
  nor2s1 _______441976(.DIN1 (___0_____27914), .DIN2 (___09_9__28070),
       .Q (___099___28129));
  nnd2s1 ______441977(.DIN1 (___09____28075), .DIN2 (________24029), .Q
       (___0990__28128));
  xor2s1 _____9_441978(.DIN1 (___0_____28025), .DIN2 (_________30693),
       .Q (_________28313));
  xor2s1 _____9_441979(.DIN1 (___0_____28024), .DIN2 (______9__32620),
       .Q (_________30667));
  xor2s1 _______441980(.DIN1 (______________18869), .DIN2
       (___0_99__28041), .Q (____0____28202));
  dffacs1 ________________________441981(.CLRB (reset), .CLK (clk),
       .DIN (___09____28089), .QN (______________________18671));
  nnd2s1 _______441982(.DIN1 (___09____28057), .DIN2 (inData[2]), .Q
       (___09____28126));
  nnd2s1 _______441983(.DIN1 (___09____28059), .DIN2 (___9____24323),
       .Q (___09____28125));
  nnd2s1 _______441984(.DIN1 (___09____28058), .DIN2 (_____9___34826),
       .Q (___09____28124));
  nor2s1 _______441985(.DIN1 (___0__0__27929), .DIN2 (___0__9__28031),
       .Q (___09____28123));
  nor2s1 ______441986(.DIN1 (___09____28121), .DIN2 (___09_9__28110),
       .Q (___09____28122));
  nnd2s1 _______441987(.DIN1 (_________34754), .DIN2 (_____00__28898),
       .Q (___09_0__28120));
  nor2s1 _____9_441988(.DIN1 (_____00__28898), .DIN2 (_________34754),
       .Q (___09_9__28119));
  or2s1 _______441989(.DIN1 (___09____28117), .DIN2 (___090___28049),
       .Q (___09____28118));
  and2s1 _____441990(.DIN1 (___09_0__28111), .DIN2 (outData[9]), .Q
       (___09____28116));
  nnd2s1 _____0_441991(.DIN1 (___0909__28050), .DIN2 (____99__24791),
       .Q (___09____28115));
  nnd2s1 _____0_441992(.DIN1 (___09____28052), .DIN2 (___09____28113),
       .Q (___09____28114));
  nor2s1 _______441993(.DIN1 (__909___26328), .DIN2 (___09_0__28111),
       .Q (___09____28112));
  nnd2s1 _____9_441994(.DIN1 (___09_9__28110), .DIN2 (___09____28121),
       .Q (____0____28151));
  xor2s1 _______441995(.DIN1 (___0__9__28013), .DIN2 (_________30693),
       .Q (____0____28200));
  nnd2s1 _______441996(.DIN1 (___09____28093), .DIN2 (________20899),
       .Q (____0_9__28195));
  nnd2s1 _______441997(.DIN1 (___0__9__28021), .DIN2 (___0_____27725),
       .Q (___09____28109));
  nnd2s1 _____441998(.DIN1 (___0_____28023), .DIN2 (___0_9___28040), .Q
       (___09____28108));
  nnd2s1 ______441999(.DIN1 (___0_9___28033), .DIN2 (_____9__23107), .Q
       (___09____28107));
  and2s1 _______442000(.DIN1 (___0_9___28035), .DIN2 (___09____28105),
       .Q (___09____28106));
  and2s1 _______442001(.DIN1 (___0_9___28037), .DIN2 (___09____28103),
       .Q (___09____28104));
  nnd2s1 _______442002(.DIN1 (___0_90__28032), .DIN2 (___900__24241),
       .Q (___09____28102));
  nor2s1 ______442003(.DIN1 (___0__0__27994), .DIN2 (___0_____28029),
       .Q (___09_0__28101));
  nor2s1 _______442004(.DIN1 (____9___22712), .DIN2 (___0900__28042),
       .Q (___09_9__28100));
  nor2s1 _______442005(.DIN1 (___0_9___28034), .DIN2 (___0_____28028),
       .Q (___09____28099));
  nnd2s1 _______442006(.DIN1 (___090___28043), .DIN2 (_________33279),
       .Q (___09____28098));
  hi1s1 _______442007(.DIN (___09____28097), .Q (____0____28166));
  nnd2s1 _______442008(.DIN1 (___0_9___28036), .DIN2 (___0__0__27984),
       .Q (_________28269));
  nnd2s1 _______442009(.DIN1 (___0_9___28039), .DIN2 (___0_____27495),
       .Q (____0_0__28177));
  xor2s1 _______442010(.DIN1 (___0__9__27983), .DIN2 (____0_0__31861),
       .Q (____0____28163));
  hi1s1 _______442011(.DIN (_________28641), .Q (____0____28175));
  hi1s1 _______442012(.DIN (___099___28136), .Q (____0____28169));
  nnd2s1 _______442013(.DIN1 (___09____28095), .DIN2 (___0_____27977),
       .Q (___09____28096));
  hi1s1 _______442014(.DIN (___09____28093), .Q (___09____28094));
  nor2s1 _______442015(.DIN1 (___0_____28002), .DIN2 (___0_____28012),
       .Q (___09____28092));
  nor2s1 _______442016(.DIN1 (___0_____27549), .DIN2 (___0_____28006),
       .Q (___09_0__28091));
  nor2s1 _______442017(.DIN1 (___0_____27615), .DIN2 (___0__0__28014),
       .Q (___09_9__28090));
  nnd2s1 ______442018(.DIN1 (___0_____27995), .DIN2 (___0_____27594),
       .Q (___09____28089));
  nnd2s1 ______442019(.DIN1 (___0__9__28003), .DIN2 (____0____28153),
       .Q (___09____28088));
  nnd2s1 _______442020(.DIN1 (___0_____27996), .DIN2 (___0_____27705),
       .Q (___09____28087));
  nnd2s1 _______442021(.DIN1 (_________34756), .DIN2 (________23270),
       .Q (___09____28086));
  nor2s1 _______442022(.DIN1 (____9___25073), .DIN2 (___0_____28010),
       .Q (___09____28085));
  nnd2s1 _______442023(.DIN1 (___0_____27987), .DIN2 (___0_____27709),
       .Q (___09____28084));
  nor2s1 _______442024(.DIN1 (________24628), .DIN2 (___0_____27997),
       .Q (___09____28083));
  nnd2s1 _______442025(.DIN1 (___0_____28019), .DIN2 (___0_____28011),
       .Q (____0____28159));
  hi1s1 _______442026(.DIN (___09____28082), .Q (_________28363));
  xor2s1 _____442027(.DIN1 (___9_9__21607), .DIN2 (___09____28055), .Q
       (____0_9__28157));
  hi1s1 _______442028(.DIN (___09_9__28110), .Q (____9_9__29072));
  nor2s1 _______442029(.DIN1 (___09_9__28080), .DIN2 (___0_____28020),
       .Q (___09_0__28081));
  and2s1 _______442030(.DIN1 (___0_____28005), .DIN2 (___09____28078),
       .Q (___09____28079));
  nnd2s1 _______442031(.DIN1 (___0__9__27993), .DIN2 (___9____26174),
       .Q (___09____28077));
  xor2s1 ______442032(.DIN1 (_____9___30449), .DIN2
       (_________________0___18633), .Q (___09____28076));
  and2s1 _______442033(.DIN1 (___0_____27999), .DIN2 (___09____28074),
       .Q (___09____28075));
  nnd2s1 _______442034(.DIN1 (___0_____27982), .DIN2 (___0_____27905),
       .Q (___09____28073));
  nnd2s1 _______442035(.DIN1 (___0_____27990), .DIN2 (outData[22]), .Q
       (___09____28072));
  nor2s1 _______442036(.DIN1 (_____0__22644), .DIN2 (___0_____27981),
       .Q (___09_0__28071));
  nnd2s1 _____9_442037(.DIN1 (___0_____27985), .DIN2 (___09____28065),
       .Q (___09_9__28070));
  nor2s1 _____9_442038(.DIN1 (________23330), .DIN2 (___0_____27986),
       .Q (___09____28069));
  nor2s1 _____442039(.DIN1 (________24741), .DIN2 (___0_____27980), .Q
       (___09____28068));
  nor2s1 _____0_442040(.DIN1 (___09____28066), .DIN2 (___0_____27991),
       .Q (___09____28067));
  nnd2s1 _____0_442041(.DIN1 (___0_____27988), .DIN2 (________22026),
       .Q (___09____28097));
  nnd2s1 _______442042(.DIN1 (___0_9___28038), .DIN2 (___09____28065),
       .Q (___09____28127));
  xor2s1 _______442043(.DIN1 (_________28979), .DIN2 (___090___28047),
       .Q (_________28641));
  xor2s1 _______442044(.DIN1 (___09____28064), .DIN2 (___0_____27956),
       .Q (___099___28136));
  dffacs1 ________________________442045(.CLRB (reset), .CLK (clk),
       .DIN (___0_____27992), .QN (______________________18672));
  nor2s1 _______442046(.DIN1 (___09____28062), .DIN2 (_________31252),
       .Q (___09____28063));
  nnd2s1 ______442047(.DIN1 (_________31252), .DIN2 (___09____28062),
       .Q (___09_0__28061));
  xor2s1 _____9_442048(.DIN1 (___0_____28017), .DIN2 (___0_____27976),
       .Q (___09_9__28060));
  nor2s1 _____0_442049(.DIN1 (________24814), .DIN2 (___0__9__27974),
       .Q (___09____28059));
  nor2s1 _______442050(.DIN1 (___99___23430), .DIN2 (___0_____27972),
       .Q (___09____28058));
  nor2s1 ______442051(.DIN1 (___0_____27978), .DIN2 (________24111), .Q
       (___09____28057));
  nnd2s1 _______442052(.DIN1 (___09____28055), .DIN2 (___0_____27875),
       .Q (___09____28056));
  or2s1 _____442053(.DIN1 (_________34452), .DIN2 (___09____28053), .Q
       (___09____28054));
  and2s1 _______442054(.DIN1 (___0_____27967), .DIN2 (___09_0__28051),
       .Q (___09____28052));
  nor2s1 _______442055(.DIN1 (_____0__24227), .DIN2 (___0_____27960),
       .Q (___0909__28050));
  or2s1 _______442056(.DIN1 (___0__0__27714), .DIN2 (___0_____27961),
       .Q (___090___28049));
  and2s1 _______442057(.DIN1 (___090___28047), .DIN2
       (____________18893), .Q (___090___28048));
  nnd2s1 ______442058(.DIN1 (___09____28053), .DIN2 (_________34452),
       .Q (___090___28046));
  hi1s1 _______442059(.DIN (___090___28045), .Q (____0____28199));
  xnr2s1 _____9_442060(.DIN1 (_________35012), .DIN2 (___0_9___27945),
       .Q (___09____28082));
  nor2s1 _______442061(.DIN1 (outData[21]), .DIN2 (___09____28055), .Q
       (___09____28093));
  xor2s1 ______442062(.DIN1 (___090___28044), .DIN2 (___0_____27926),
       .Q (___09_9__28110));
  nor2s1 _______442063(.DIN1 (___0_____27979), .DIN2 (_________28471),
       .Q (___090___28043));
  nnd2s1 _____9_442064(.DIN1 (___0_____27970), .DIN2 (________25154),
       .Q (___0900__28042));
  nnd2s1 _____0_442065(.DIN1 (___0__0__28022), .DIN2 (___0_9___28040),
       .Q (___0_99__28041));
  hi1s1 _____0_442066(.DIN (___0_9___28038), .Q (___0_9___28039));
  nor2s1 _______442067(.DIN1 (__9_____26671), .DIN2 (___0_____27969),
       .Q (___0_9___28037));
  xor2s1 _______442068(.DIN1 (___0_____28030), .DIN2 (_________33895),
       .Q (___0_9___28036));
  nor2s1 _______442069(.DIN1 (___0_9___28034), .DIN2 (___0__0__27965),
       .Q (___0_9___28035));
  nor2s1 ______442070(.DIN1 (________23735), .DIN2 (___0_____27963), .Q
       (___0_9___28033));
  nor2s1 _______442071(.DIN1 (_____9__23581), .DIN2 (___0_____27962),
       .Q (___0_90__28032));
  nor2s1 _____9_442072(.DIN1 (___0_____28030), .DIN2 (___0_____27957),
       .Q (___0__9__28031));
  nnd2s1 _______442073(.DIN1 (___0_____27958), .DIN2 (________25874),
       .Q (___0_____28029));
  nnd2s1 _______442074(.DIN1 (___0_____27975), .DIN2 (___0_____27915),
       .Q (___0_____28028));
  nor2s1 _______442075(.DIN1 (___0_____28026), .DIN2 (___090___28047),
       .Q (___0_____28027));
  nor2s1 _______442076(.DIN1 (___0__0__27955), .DIN2 (___0_____27959),
       .Q (___0_____28025));
  xor2s1 _______442077(.DIN1 (___0_____27989), .DIN2 (outData[21]), .Q
       (___0_____28024));
  nnd2s1 _______442078(.DIN1 (___0__0__28022), .DIN2 (_________28866),
       .Q (___0_____28023));
  nor2s1 _______442079(.DIN1 (________23157), .DIN2 (___0__9__27964),
       .Q (___0__9__28021));
  or2s1 _____442080(.DIN1 (____________18893), .DIN2 (___090___28047),
       .Q (___09_0__28111));
  dffacs1 _______________________442081(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27971), .QN (_____________________18663));
  nnd2s1 _______442082(.DIN1 (___0_____27931), .DIN2 (____0____28153),
       .Q (___0_____28020));
  nnd2s1 _____0_442083(.DIN1 (___0_0___27951), .DIN2
       (______________________________________0___________), .Q
       (___0_____28019));
  nnd2s1 ______442084(.DIN1 (___0_____28017), .DIN2 (___0__9__27908),
       .Q (___0_____28018));
  hi1s1 _______442085(.DIN (___0_____28015), .Q (___0_____28016));
  nnd2s1 ______442086(.DIN1 (___0_9___27946), .DIN2 (__9_____26835), .Q
       (___0__0__28014));
  nnd2s1 _______442087(.DIN1 (___0_____28000), .DIN2 (___0_____28001),
       .Q (___0__9__28013));
  or2s1 _______442088(.DIN1 (_____00__28331), .DIN2 (___0_9___27939),
       .Q (___0_____28012));
  nnd2s1 _____0_442089(.DIN1 (___0_0___27948), .DIN2
       (______________________________________0__________0), .Q
       (___0_____28011));
  nnd2s1 _______442090(.DIN1 (___0_9___27943), .DIN2 (________25046),
       .Q (___0_____28010));
  or2s1 _______442091(.DIN1 (_________________18709), .DIN2
       (___0_____28008), .Q (___0_____28009));
  and2s1 _______442092(.DIN1 (___0_____28008), .DIN2
       (_________________18709), .Q (___0_____28007));
  nnd2s1 _______442093(.DIN1 (___0_9___27942), .DIN2 (________24187),
       .Q (___0_____28006));
  nor2s1 _______442094(.DIN1 (___0__0__28004), .DIN2 (___0_9___27941),
       .Q (___0_____28005));
  nor2s1 _______442095(.DIN1 (___0_____28002), .DIN2 (___0_____27922),
       .Q (___0__9__28003));
  nor2s1 _______442096(.DIN1 (___0_____28001), .DIN2 (___0_____28000),
       .Q (___090___28045));
  nnd2s1 ______442097(.DIN1 (___0_99__27947), .DIN2 (___0__9__27742),
       .Q (___09____28095));
  and2s1 ______442098(.DIN1 (___0_____27924), .DIN2 (___0_____27998),
       .Q (___0_____27999));
  nnd2s1 _____9_442099(.DIN1 (___0_9___27944), .DIN2 (___0____25353),
       .Q (___0_____27997));
  nor2s1 _______442100(.DIN1 (____9___23166), .DIN2 (___0_____27932),
       .Q (___0_____27996));
  nor2s1 _______442101(.DIN1 (___0__0__27994), .DIN2 (___0_____27936),
       .Q (___0_____27995));
  nor2s1 _______442102(.DIN1 (___9_0__26167), .DIN2 (___0_____27927),
       .Q (___0__9__27993));
  nnd2s1 _______442103(.DIN1 (___0_____27935), .DIN2 (__9_____26812),
       .Q (___0_____27992));
  or2s1 _____9_442104(.DIN1 (___0_9___28034), .DIN2 (___0_____27916),
       .Q (___0_____27991));
  nnd2s1 _______442105(.DIN1 (___0_____27989), .DIN2
       (_____________18898), .Q (___0_____27990));
  nor2s1 ______442106(.DIN1 (________25033), .DIN2 (___0_____27925), .Q
       (___0_____27988));
  and2s1 _____9_442107(.DIN1 (___0__9__27937), .DIN2 (________24752),
       .Q (___0_____27987));
  nnd2s1 ______442108(.DIN1 (___0__9__27918), .DIN2 (_____0__23108), .Q
       (___0_____27986));
  nnd2s1 _______442109(.DIN1 (___0_____28030), .DIN2 (___0__0__27984),
       .Q (___0_____27985));
  nor2s1 _______442110(.DIN1 (outData[21]), .DIN2 (___0_____27920), .Q
       (___0__9__27983));
  and2s1 _______442111(.DIN1 (___0_____27923), .DIN2 (___0_____27973),
       .Q (___0_____27982));
  nnd2s1 _______442112(.DIN1 (___0__0__27919), .DIN2 (___09____28074),
       .Q (___0_____27981));
  nnd2s1 _______442113(.DIN1 (___0_____27917), .DIN2 (___9____25243),
       .Q (___0_____27980));
  xor2s1 _______442114(.DIN1 (___0_____27893), .DIN2 (____99___31805),
       .Q (___0_9___28038));
  dffacs1 ________________________442115(.CLRB (reset), .CLK (clk),
       .DIN (___0_0___27952), .QN (______________________18632));
  nor2s1 _______442116(.DIN1 (__0), .DIN2 (_________28374), .Q
       (___0_____27979));
  xor2s1 _______442117(.DIN1 (_________________18718), .DIN2
       (____________0___18704), .Q (___0_____27978));
  nnd2s1 _______442118(.DIN1 (___0_____27934), .DIN2 (___0_____27976),
       .Q (___0_____27977));
  nor2s1 _______442119(.DIN1 (___0_____27966), .DIN2 (___0__9__27889),
       .Q (___0_____27975));
  nnd2s1 ______442120(.DIN1 (___0_____27906), .DIN2 (___0_____27973),
       .Q (___0__9__27974));
  nnd2s1 _______442121(.DIN1 (___0_____27907), .DIN2 (___0____23462),
       .Q (___0_____27972));
  nnd2s1 _______442122(.DIN1 (___0_____27886), .DIN2 (___0_0___27755),
       .Q (___0_____27971));
  nor2s1 _______442123(.DIN1 (________23573), .DIN2 (___0_____27888),
       .Q (___0_____27970));
  or2s1 _______442124(.DIN1 (___0_____27968), .DIN2 (___0_____27891),
       .Q (___0_____27969));
  nor2s1 _______442125(.DIN1 (___0_____27966), .DIN2 (___0_____27903),
       .Q (___0_____27967));
  xor2s1 ______442126(.DIN1 (___0_____27868), .DIN2 (___0_0___27857),
       .Q (___0_____28015));
  xor2s1 _______442127(.DIN1 (___0_0___27852), .DIN2 (____9_9__33643),
       .Q (___09____28055));
  xnr2s1 ______442128(.DIN1 (___0_0___27950), .DIN2 (________26005), .Q
       (_________31252));
  nnd2s1 _____9_442129(.DIN1 (___0_____27885), .DIN2 (___0_____27825),
       .Q (___0__0__27965));
  or2s1 _______442130(.DIN1 (_________28483), .DIN2 (___0_____27884),
       .Q (___0__9__27964));
  nnd2s1 ______442131(.DIN1 (___0_____27887), .DIN2 (________23586), .Q
       (___0_____27963));
  nnd2s1 _______442132(.DIN1 (___0__0__27909), .DIN2 (________21999),
       .Q (___0_____27962));
  nnd2s1 _______442133(.DIN1 (___0_____27904), .DIN2 (___0__9__27324),
       .Q (___0_____27961));
  nnd2s1 _______442134(.DIN1 (___0_____27895), .DIN2 (___0__0__27609),
       .Q (___0_____27960));
  nor2s1 _____442135(.DIN1 (___09____28064), .DIN2 (___0_09__27954), .Q
       (___0_____27959));
  nor2s1 _______442136(.DIN1 (________24967), .DIN2 (___0_____27901),
       .Q (___0_____27958));
  nnd2s1 _____0_442137(.DIN1 (___0__0__27984), .DIN2 (___0_9___27846),
       .Q (___0_____27957));
  nor2s1 _____0_442138(.DIN1 (___0__0__27955), .DIN2 (___0_09__27954),
       .Q (___0_____27956));
  nnd2s1 _______442139(.DIN1 (___0_____27883), .DIN2 (_________28603),
       .Q (___0__0__28022));
  xor2s1 _____0_442140(.DIN1 (___0_0___27953), .DIN2 (outData[20]), .Q
       (___09____28053));
  and2s1 _______442141(.DIN1 (___0_0___27953), .DIN2 (___0_____27892),
       .Q (_____9___30449));
  nnd2s1 _______442142(.DIN1 (___0_____27900), .DIN2 (________19286),
       .Q (___090___28047));
  dffacs1 _______________________442143(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27913), .QN (_____________________18662));
  nnd2s1 _______442144(.DIN1 (___0_____27864), .DIN2 (________25767),
       .Q (___0_0___27952));
  nnd2s1 ______442145(.DIN1 (___0_0___27950), .DIN2 (________20337), .Q
       (___0_0___27951));
  nnd2s1 ______442146(.DIN1 (___0_0___27950), .DIN2 (_____9__25060), .Q
       (___0_0___27948));
  nnd2s1 ______442147(.DIN1 (___0__9__27869), .DIN2 (___0_____27832),
       .Q (___0_99__27947));
  nor2s1 _______442148(.DIN1 (__99_0__27154), .DIN2 (___0_____27872),
       .Q (___0_9___27946));
  nor2s1 _______442149(.DIN1 (___0_____27823), .DIN2 (___0_____27871),
       .Q (___0_9___27945));
  nor2s1 _______442150(.DIN1 (__9_____26953), .DIN2 (___0_____27863),
       .Q (___0_9___27944));
  nor2s1 _______442151(.DIN1 (________24839), .DIN2 (___0_____27876),
       .Q (___0_9___27943));
  nor2s1 _______442152(.DIN1 (________22911), .DIN2 (___0_____27861),
       .Q (___0_9___27942));
  or2s1 _______442153(.DIN1 (___0_9___27940), .DIN2 (___0_____27878),
       .Q (___0_9___27941));
  nnd2s1 _______442154(.DIN1 (___0_____27874), .DIN2 (___0_90__27938),
       .Q (___0_9___27939));
  nor2s1 ______442155(.DIN1 (____99__25463), .DIN2 (___0__0__27880), .Q
       (___0__9__27937));
  nnd2s1 _______442156(.DIN1 (___0__0__27860), .DIN2 (___0_____27536),
       .Q (___0_____27936));
  nor2s1 _______442157(.DIN1 (___0_____27539), .DIN2 (___0_____27866),
       .Q (___0_____27935));
  hi1s1 _____0_442158(.DIN (___0_____27934), .Q (___0_____28017));
  nor2s1 ______442159(.DIN1 (_________34472), .DIN2 (___0_____27881),
       .Q (_________28471));
  nor2s1 _______442160(.DIN1 (___0_____27774), .DIN2 (___0_____27867),
       .Q (___0_____28008));
  nnd2s1 _______442161(.DIN1 (___0_____27933), .DIN2
       (____________0___18704), .Q (___0_____28001));
  nnd2s1 ______442162(.DIN1 (___0_0___27855), .DIN2 (________25877), .Q
       (___0_____27932));
  nor2s1 _______442163(.DIN1 (___0_____27767), .DIN2 (___0_90__27840),
       .Q (___0_____27931));
  nor2s1 _____9_442164(.DIN1 (_________31154), .DIN2 (___0__9__27928),
       .Q (___0_____27930));
  and2s1 _____9_442165(.DIN1 (___0__9__27928), .DIN2 (_________31154),
       .Q (___0__0__27929));
  nnd2s1 _____9_442166(.DIN1 (___0_0___27854), .DIN2 (__9__0__26664),
       .Q (___0_____27927));
  xor2s1 _____0_442167(.DIN1 (___0__0__27899), .DIN2 (_____0___30999),
       .Q (___0_____27926));
  nnd2s1 _______442168(.DIN1 (___0_9___27841), .DIN2 (________25866),
       .Q (___0_____27925));
  and2s1 ______442169(.DIN1 (___0_____27836), .DIN2 (____0___25656), .Q
       (___0_____27924));
  nor2s1 _______442170(.DIN1 (________26092), .DIN2 (___0_0___27856),
       .Q (___0_____27923));
  or2s1 _______442171(.DIN1 (___0_____27921), .DIN2 (___0_0___27858),
       .Q (___0_____27922));
  or2s1 _______442172(.DIN1 (________22684), .DIN2 (___0_0___27953), .Q
       (___0_____27920));
  nor2s1 _______442173(.DIN1 (__90____26275), .DIN2 (___0_____27835),
       .Q (___0__0__27919));
  nor2s1 _______442174(.DIN1 (_____0__23950), .DIN2 (___0_____27837),
       .Q (___0__9__27918));
  nor2s1 _______442175(.DIN1 (_____0__24676), .DIN2 (___0_9___27845),
       .Q (___0_____27917));
  nnd2s1 ______442176(.DIN1 (___0_00__27850), .DIN2 (___0_____27915),
       .Q (___0_____27916));
  nor2s1 _______442177(.DIN1 (outData[20]), .DIN2 (___0_0___27953), .Q
       (___0_____27989));
  nnd2s1 _______442178(.DIN1 (___0_____27882), .DIN2
       (______________18868), .Q (___0_9___28040));
  nor2s1 _______442179(.DIN1 (___0_____27914), .DIN2 (___0_9___27847),
       .Q (___0_____28030));
  dffacs1 ____0__________________442180(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27865), .QN (____0________________18590));
  dffacs1 _______________________442181(.CLRB (reset), .CLK (clk), .DIN
       (___0_09__27859), .QN (_____________________18666));
  nnd2s1 _______442182(.DIN1 (___0_____27813), .DIN2 (___0_____27912),
       .Q (___0_____27913));
  nnd2s1 _______442183(.DIN1 (___0_____27831), .DIN2 (___0_____27545),
       .Q (___0_____27911));
  nor2s1 ______442184(.DIN1 (___0_____27546), .DIN2 (___0_____27833),
       .Q (___0_____27910));
  nor2s1 _______442185(.DIN1 (___0_____27894), .DIN2 (___0_____27814),
       .Q (___0__0__27909));
  hi1s1 _______442186(.DIN (___0_____27976), .Q (___0__9__27908));
  nor2s1 _______442187(.DIN1 (___0_____27730), .DIN2 (___0_____27826),
       .Q (___0_____27907));
  and2s1 _____9_442188(.DIN1 (___0_____27824), .DIN2 (___0_____27905),
       .Q (___0_____27906));
  nor2s1 _____0_442189(.DIN1 (________23660), .DIN2 (___0_____27817),
       .Q (___0_____27904));
  nnd2s1 _______442190(.DIN1 (___0_____27821), .DIN2 (___0_____27902),
       .Q (___0_____27903));
  or2s1 _______442191(.DIN1 (________24443), .DIN2 (___0_____27815), .Q
       (___0_____27901));
  nnd2s1 ______442192(.DIN1 (___0__0__27899), .DIN2 (________19285), .Q
       (___0_____27900));
  and2s1 ______442193(.DIN1 (___0_____27806), .DIN2 (___0_____27897),
       .Q (___0__9__27898));
  xor2s1 ______442194(.DIN1 (___0__0__27870), .DIN2 (_____0__24044), .Q
       (___0_____27934));
  xor2s1 ______442195(.DIN1 (___0__9__27791), .DIN2 (___0_____27896),
       .Q (_________29746));
  nor2s1 _______442196(.DIN1 (___0_____27894), .DIN2 (___0_____27805),
       .Q (___0_____27895));
  nor2s1 _______442197(.DIN1 (___0__0__27511), .DIN2 (___0__0__27810),
       .Q (___0_____27893));
  nnd2s1 _______442198(.DIN1 (___0_____27809), .DIN2 (outData[19]), .Q
       (___0_____27892));
  nnd2s1 _______442199(.DIN1 (___0__0__27820), .DIN2 (___0__0__27890),
       .Q (___0_____27891));
  nnd2s1 _______442200(.DIN1 (___0_____27818), .DIN2 (________23920),
       .Q (___0__9__27889));
  nnd2s1 ______442201(.DIN1 (___0_____27803), .DIN2 (________24194), .Q
       (___0_____27888));
  and2s1 _______442202(.DIN1 (___0__9__27801), .DIN2 (___09____28074),
       .Q (___0_____27887));
  nor2s1 _______442203(.DIN1 (___0_____27477), .DIN2 (___0_____27812),
       .Q (___0_____27886));
  nor2s1 _______442204(.DIN1 (____0___23715), .DIN2 (___0_____27822),
       .Q (___0_____27885));
  nnd2s1 _____0_442205(.DIN1 (___0_____27799), .DIN2 (___09____28105),
       .Q (___0_____27884));
  hi1s1 _______442206(.DIN (___0_____27882), .Q (___0_____27883));
  nor2s1 _______442207(.DIN1 (________24466), .DIN2 (___0_____27807),
       .Q (___0_09__27954));
  hi1s1 _______442208(.DIN (___0_____27881), .Q (_________28374));
  xor2s1 _______442209(.DIN1 (___0_____27763), .DIN2 (_________33895),
       .Q (___0__0__27984));
  dffacs1 ____0__________________442210(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27834), .QN (____0________________18652));
  nnd2s1 _______442211(.DIN1 (___0_____27769), .DIN2 (___0__9__27879),
       .Q (___0__0__27880));
  or2s1 _______442212(.DIN1 (___0_____27877), .DIN2 (___0_____27764),
       .Q (___0_____27878));
  nnd2s1 _______442213(.DIN1 (___0_____27797), .DIN2 (_____0__24473),
       .Q (___0_____27876));
  nnd2s1 ______442214(.DIN1 (___0_0___27851), .DIN2 (outData[20]), .Q
       (___0_____27875));
  and2s1 _______442215(.DIN1 (___0_____27766), .DIN2 (___0_____27873),
       .Q (___0_____27874));
  xor2s1 ______442216(.DIN1 (___0_9___27745), .DIN2 (_________33385),
       .Q (___0_____27872));
  nor2s1 _____9_442217(.DIN1 (_____0___33866), .DIN2 (___0__0__27870),
       .Q (___0_____27871));
  xor2s1 _____9_442218(.DIN1 (___0_____27740), .DIN2 (_________32624),
       .Q (___0__9__27869));
  xor2s1 _____0_442219(.DIN1 (_____0__23092), .DIN2 (_____99__29445),
       .Q (___0_____27868));
  nor2s1 _____0_442220(.DIN1 (_________9_), .DIN2 (___0_____27776), .Q
       (___0_____27867));
  nnd2s1 ______442221(.DIN1 (___0_____27777), .DIN2 (__9_____27019), .Q
       (___0_____27866));
  nnd2s1 _______442222(.DIN1 (___0_____27793), .DIN2 (___0_____27816),
       .Q (___0_____27865));
  nor2s1 _______442223(.DIN1 (__9_____26404), .DIN2 (___0__0__27772),
       .Q (___0_____27864));
  nnd2s1 _______442224(.DIN1 (___0_____27784), .DIN2 (___0_____27862),
       .Q (___0_____27863));
  nnd2s1 ______442225(.DIN1 (___0__0__27782), .DIN2 (____9___23338), .Q
       (___0_____27861));
  nor2s1 _______442226(.DIN1 (____0___24430), .DIN2 (___0_____27786),
       .Q (___0__0__27860));
  or2s1 _______442227(.DIN1 (__9__0__27035), .DIN2 (___0_____27787), .Q
       (___0_09__27859));
  nnd2s1 _______442228(.DIN1 (___0__9__27781), .DIN2 (___9____24304),
       .Q (___0_0___27858));
  nnd2s1 _______442229(.DIN1 (___0_____27795), .DIN2 (___0_0___27857),
       .Q (___0_0___27949));
  nor2s1 ______442230(.DIN1 (___9____21595), .DIN2 (___0_____27789), .Q
       (___0_0___27950));
  nnd2s1 _______442231(.DIN1 (___0_____27796), .DIN2 (___0_____27580),
       .Q (___0_____27976));
  dffacs1 ________________0_442232(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27794), .Q (____________0___18704));
  or2s1 _____9_442233(.DIN1 (___0090__27257), .DIN2 (___0_0___27759),
       .Q (___0_0___27856));
  nor2s1 ______442234(.DIN1 (___0__0__28004), .DIN2 (___0_____27768),
       .Q (___0_0___27855));
  nor2s1 _______442235(.DIN1 (__9_____26831), .DIN2 (___0_0___27757),
       .Q (___0_0___27854));
  and2s1 _______442236(.DIN1 (___0_____27779), .DIN2 (_________28837),
       .Q (___0_0___27853));
  nor2s1 ______442237(.DIN1 (outData[20]), .DIN2 (___0_0___27851), .Q
       (___0_0___27852));
  nor2s1 ______442238(.DIN1 (___0_____27798), .DIN2 (___0_09__27761),
       .Q (___0_00__27850));
  nor2s1 _______442239(.DIN1 (___0_9___27848), .DIN2 (___0_____27770),
       .Q (___0_99__27849));
  nnd2s1 ______442240(.DIN1 (___0_9___27846), .DIN2 (___09____28065),
       .Q (___0_9___27847));
  nnd2s1 ______442241(.DIN1 (___0_0___27756), .DIN2 (________24449), .Q
       (___0_9___27845));
  and2s1 _______442242(.DIN1 (___0_9___27843), .DIN2 (___0_9___27842),
       .Q (___0_9___27844));
  nor2s1 _____442243(.DIN1 (_____9___34926), .DIN2 (___0_0___27760), .Q
       (___0_9___27841));
  nnd2s1 _______442244(.DIN1 (___0_____27765), .DIN2 (___0__9__27839),
       .Q (___0_90__27840));
  nor2s1 _____9_442245(.DIN1 (___0_9___27842), .DIN2 (___0_9___27843),
       .Q (___0_____27838));
  nor2s1 _______442246(.DIN1 (____99__22894), .DIN2 (___0_0___27758),
       .Q (___0_____27837));
  nor2s1 _______442247(.DIN1 (____9___22715), .DIN2 (___0_0___27754),
       .Q (___0_____27836));
  nnd2s1 _______442248(.DIN1 (___0_00__27753), .DIN2 (___00____27213),
       .Q (___0_____27835));
  nnd2s1 _____442249(.DIN1 (______0__34758), .DIN2 (___0_____27672), .Q
       (___0_____27882));
  xor2s1 _______442250(.DIN1 (___0_____27513), .DIN2 (_________34762),
       .Q (___0_____27881));
  nor2s1 _______442251(.DIN1 (________24467), .DIN2 (_________34760),
       .Q (___0__0__27955));
  nor2s1 ______442252(.DIN1 (___0__9__27392), .DIN2 (___0_____27775),
       .Q (___0__9__27928));
  nnd2s1 _______442253(.DIN1 (___0_____27808), .DIN2 (_________9_), .Q
       (___0_0___27953));
  dffacs1 ____0________________9_442254(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27788), .QN (____0____________9___18654));
  nnd2s1 _____0_442255(.DIN1 (___0_____27728), .DIN2 (____9____29042),
       .Q (___0_____27834));
  and2s1 _____442256(.DIN1 (___0__0__27830), .DIN2 (___0_____27832), .Q
       (___0_____27833));
  or2s1 _____442257(.DIN1 (___0_____27832), .DIN2 (___0__0__27830), .Q
       (___0_____27831));
  nnd2s1 _______442258(.DIN1 (___0_____27828), .DIN2 (_________34479),
       .Q (___0__9__27829));
  or2s1 _______442259(.DIN1 (_________34479), .DIN2 (___0_____27828),
       .Q (___0_____27827));
  nnd2s1 _______442260(.DIN1 (___0_9___27747), .DIN2 (___0_____27825),
       .Q (___0_____27826));
  nor2s1 _______442261(.DIN1 (_____0__26127), .DIN2 (___0_9___27749),
       .Q (___0_____27824));
  nnd2s1 _______442262(.DIN1 (___0_____27741), .DIN2 (________23959),
       .Q (___0_____27823));
  nnd2s1 ______442263(.DIN1 (___0__0__27733), .DIN2 (________24093), .Q
       (___0_____27822));
  nor2s1 _______442264(.DIN1 (_____0__24936), .DIN2 (___0_____27726),
       .Q (___0_____27821));
  nor2s1 _______442265(.DIN1 (___0__9__27819), .DIN2 (___0_____27734),
       .Q (___0__0__27820));
  nor2s1 ______442266(.DIN1 (________23826), .DIN2 (___0_____27718), .Q
       (___0_____27818));
  nnd2s1 _____442267(.DIN1 (___0_____27722), .DIN2 (___0_____27816), .Q
       (___0_____27817));
  dffacs1 ____0__________________442268(.CLRB (reset), .CLK (clk), .DIN
       (___0_9___27746), .QN (____0________________18650));
  nnd2s1 ______442269(.DIN1 (___0_____27727), .DIN2 (___0_____27690),
       .Q (___0_____27815));
  nnd2s1 _____0_442270(.DIN1 (___0_9___27750), .DIN2 (_____9___35026),
       .Q (___0_____27814));
  nor2s1 _____0_442271(.DIN1 (____9___25462), .DIN2 (___0_____27719),
       .Q (___0_____27813));
  or2s1 _____0_442272(.DIN1 (___0_____27811), .DIN2 (___0__9__27732),
       .Q (___0_____27812));
  nor2s1 _____0_442273(.DIN1 (_________34762), .DIN2 (___0_____27512),
       .Q (___0__0__27810));
  hi1s1 _______442274(.DIN (___0_____27808), .Q (___0_____27809));
  hi1s1 _______442275(.DIN (_________34760), .Q (___0_____27807));
  and2s1 _____0_442276(.DIN1 (___0_____27737), .DIN2 (__9_____26447),
       .Q (___0_____27806));
  or2s1 _______442277(.DIN1 (___0_____27804), .DIN2 (___0_____27721),
       .Q (___0_____27805));
  and2s1 _______442278(.DIN1 (___0__9__27723), .DIN2 (___0__0__27802),
       .Q (___0_____27803));
  and2s1 _______442279(.DIN1 (___0__0__27724), .DIN2 (___0_____27800),
       .Q (___0__9__27801));
  nor2s1 _______442280(.DIN1 (___0_____27798), .DIN2 (___0_____27731),
       .Q (___0_____27799));
  xor2s1 _______442281(.DIN1 (___0__0__27676), .DIN2 (____9____29052),
       .Q (_________28533));
  nnd2s1 _______442282(.DIN1 (___0_____27736), .DIN2 (___0_90__27743),
       .Q (___0__0__27899));
  xor2s1 _______442283(.DIN1 (___0_99__27752), .DIN2 (outData[18]), .Q
       (_________32535));
  nor2s1 _______442284(.DIN1 (____90__24598), .DIN2 (___0_____27691),
       .Q (___0_____27797));
  nnd2s1 _______442285(.DIN1 (___0__9__27713), .DIN2 (___0____22547),
       .Q (___0_____27796));
  or2s1 _______442286(.DIN1 (_________34437), .DIN2 (_________29594),
       .Q (___0_____27795));
  nnd2s1 _______442287(.DIN1 (___0_____27702), .DIN2 (___0____24397),
       .Q (___0_____27794));
  and2s1 _______442288(.DIN1 (___0_____27715), .DIN2 (___0__0__27792),
       .Q (___0_____27793));
  nor2s1 _______442289(.DIN1 (___0_____27494), .DIN2 (___0_____27716),
       .Q (___0__9__27791));
  xnr2s1 _______442290(.DIN1 (_________35066), .DIN2 (______9__28944),
       .Q (___0_____27790));
  xor2s1 _______442291(.DIN1 (___0_____27668), .DIN2 (_________30131),
       .Q (___0_____27789));
  nnd2s1 _______442292(.DIN1 (___0__0__27704), .DIN2 (_________28942),
       .Q (___0_____27788));
  nnd2s1 _______442293(.DIN1 (___0_____27701), .DIN2 (___0_____27527),
       .Q (___0_____27787));
  nnd2s1 _______442294(.DIN1 (___0_____27717), .DIN2 (___00___24339),
       .Q (___0_____27786));
  and2s1 _____442295(.DIN1 (_________29594), .DIN2 (_________34437), .Q
       (___0_____27785));
  nor2s1 _______442296(.DIN1 (___0_____27783), .DIN2 (___0_____27700),
       .Q (___0_____27784));
  nor2s1 _____9_442297(.DIN1 (___0_____28002), .DIN2 (___0_____27695),
       .Q (___0__0__27782));
  and2s1 _____9_442298(.DIN1 (___0_____27707), .DIN2 (___0_____27780),
       .Q (___0__9__27781));
  nor2s1 _____0_442299(.DIN1 (___0_____27778), .DIN2 (___0__9__27703),
       .Q (___0_____27779));
  nor2s1 _______442300(.DIN1 (___9____25258), .DIN2 (___0_____27710),
       .Q (___0_____27777));
  nnd2s1 ______442301(.DIN1 (___0_____27773), .DIN2 (_________32624),
       .Q (___0_____27776));
  xor2s1 _______442302(.DIN1 (___0_____27639), .DIN2 (___0_____27914),
       .Q (___0_____27775));
  nor2s1 _______442303(.DIN1 (____9___23341), .DIN2 (___0_____27773),
       .Q (___0_____27774));
  nor2s1 _______442304(.DIN1 (___0__9__27771), .DIN2 (___0_____27697),
       .Q (___0__0__27772));
  xor2s1 _______442305(.DIN1 (___0_9___27744), .DIN2 (_____0__23958),
       .Q (___0__0__27870));
  nnd2s1 ______442306(.DIN1 (___0_____27677), .DIN2 (______0__35038),
       .Q (___0_____27770));
  nor2s1 _______442307(.DIN1 (________24593), .DIN2 (___0_____27699),
       .Q (___0_____27769));
  or2s1 _______442308(.DIN1 (___0_____27767), .DIN2 (___0_____27712),
       .Q (___0_____27768));
  nor2s1 ______442309(.DIN1 (___0__0__27637), .DIN2 (___0__0__27694),
       .Q (___0_____27766));
  and2s1 _______442310(.DIN1 (___0_____27706), .DIN2 (___0_90__27938),
       .Q (___0_____27765));
  nnd2s1 _______442311(.DIN1 (___0__9__27693), .DIN2 (_____9__24625),
       .Q (___0_____27764));
  nor2s1 _______442312(.DIN1 (___0_9___27751), .DIN2 (___0__0__27762),
       .Q (___0_____27763));
  nnd2s1 _______442313(.DIN1 (___0_____27678), .DIN2 (___0_____27573),
       .Q (___0_09__27761));
  nnd2s1 _______442314(.DIN1 (___0_____27680), .DIN2 (____0___24704),
       .Q (___0_0___27760));
  nnd2s1 ______442315(.DIN1 (___0_____27679), .DIN2 (____99__23801), .Q
       (___0_0___27759));
  nnd2s1 _______442316(.DIN1 (___0_____27688), .DIN2 (__9_____26846),
       .Q (___0_0___27758));
  nnd2s1 _______442317(.DIN1 (___0_____27692), .DIN2 (___0____25333),
       .Q (___0_0___27757));
  and2s1 _______442318(.DIN1 (___0_____27687), .DIN2 (___0_0___27755),
       .Q (___0_0___27756));
  nnd2s1 _____0_442319(.DIN1 (___0_____27682), .DIN2 (________24744),
       .Q (___0_0___27754));
  nor2s1 _____0_442320(.DIN1 (___00___25273), .DIN2 (___0_____27689),
       .Q (___0_00__27753));
  nor2s1 _______442321(.DIN1 (outData[18]), .DIN2 (___0_99__27752), .Q
       (___0_____27808));
  nnd2s1 _______442322(.DIN1 (___0_____27681), .DIN2 (___0_____27674),
       .Q (_________29468));
  nnd2s1 _______442323(.DIN1 (___0__0__27762), .DIN2 (___0_9___27751),
       .Q (___0_9___27846));
  nnd2s1 _______442324(.DIN1 (___0_____27773), .DIN2 (_________9_), .Q
       (___0_0___27851));
  and2s1 _______442325(.DIN1 (___0_99__27752), .DIN2 (___0_____27673),
       .Q (___0_9___27843));
  dffacs1 ____0___________________442326(.CLRB (reset), .CLK (clk),
       .DIN (___0_____27708), .QN (____0_________________18596));
  nor2s1 _______442327(.DIN1 (___0____22605), .DIN2 (___0_9___27652),
       .Q (___0_9___27750));
  or2s1 _____9_442328(.DIN1 (___0_9___27748), .DIN2 (___0_0___27664),
       .Q (___0_9___27749));
  nor2s1 _____9_442329(.DIN1 (___0_9___27557), .DIN2 (___0_0___27662),
       .Q (___0_9___27747));
  nnd2s1 _____442330(.DIN1 (___0_0___27661), .DIN2 (____9____29042), .Q
       (___0_9___27746));
  nnd2s1 ______442331(.DIN1 (___0_9___27744), .DIN2 (___99___20691), .Q
       (___0_9___27745));
  nnd2s1 _______442332(.DIN1 (___0_____27643), .DIN2 (_________31134),
       .Q (___0_90__27743));
  nnd2s1 ______442333(.DIN1 (___0_____27738), .DIN2 (___0_____27739),
       .Q (___0__9__27742));
  nnd2s1 _______442334(.DIN1 (___0_9___27744), .DIN2 (________24045),
       .Q (___0_____27741));
  nor2s1 _______442335(.DIN1 (___0_____27739), .DIN2 (___0_____27738),
       .Q (___0_____27740));
  nor2s1 _______442336(.DIN1 (__9_____26535), .DIN2 (___0__0__27666),
       .Q (___0_____27737));
  nnd2s1 _______442337(.DIN1 (___0_9___27647), .DIN2 (___0_____27735),
       .Q (___0_____27736));
  or2s1 _______442338(.DIN1 (________24553), .DIN2 (___0_0___27658), .Q
       (___0_____27734));
  and2s1 _______442339(.DIN1 (___0_____27644), .DIN2 (________23282),
       .Q (___0__0__27733));
  xor2s1 _______442340(.DIN1 (___0_9___27654), .DIN2 (___0_____27739),
       .Q (___0__0__27830));
  xor2s1 ______442341(.DIN1 (___0_____27671), .DIN2 (outData[18]), .Q
       (___0_____27828));
  hi1s1 _______442342(.DIN (_________29594), .Q (_____99__29445));
  or2s1 ______442343(.DIN1 (__99____27128), .DIN2 (___0_9___27650), .Q
       (___0__9__27732));
  or2s1 ______442344(.DIN1 (___0_____27730), .DIN2 (___0_____27638), .Q
       (___0_____27731));
  nor2s1 _____9_442345(.DIN1 (________25676), .DIN2 (___0_90__27646),
       .Q (___0_____27728));
  nor2s1 _____9_442346(.DIN1 (___9____25216), .DIN2 (___0_____27640),
       .Q (___0_____27727));
  nnd2s1 _____9_442347(.DIN1 (___0_00__27656), .DIN2 (___0_____27725),
       .Q (___0_____27726));
  nor2s1 _____9_442348(.DIN1 (___9____24322), .DIN2 (___0_99__27655),
       .Q (___0__0__27724));
  nor2s1 _____9_442349(.DIN1 (___0_____27783), .DIN2 (___0_9___27649),
       .Q (___0__9__27723));
  nor2s1 _____442350(.DIN1 (___0_9___27648), .DIN2 (___0_9___27653), .Q
       (___0_____27722));
  nnd2s1 _____442351(.DIN1 (___0_____27642), .DIN2 (___0_____27720), .Q
       (___0_____27721));
  nnd2s1 _______442352(.DIN1 (___0_9___27651), .DIN2 (___0_____27612),
       .Q (___0_____27719));
  nnd2s1 _______442353(.DIN1 (___0_____27641), .DIN2 (____09__23180),
       .Q (___0_____27718));
  dffacs1 ____0___________________442354(.CLRB (reset), .CLK (clk),
       .DIN (___0_0___27660), .QN (____0_________________18657));
  dffacs1 _______________________442355(.CLRB (reset), .CLK (clk), .DIN
       (___0_0___27657), .QN (_____________________18600));
  dffacs1 ____0__________________442356(.CLRB (reset), .CLK (clk), .DIN
       (___0_0___27663), .QN (____0________________18647));
  dffacs1 ________________9_442357(.CLRB (reset), .CLK (clk), .DIN
       (___0__9__27645), .QN
       (______________________________________0_____________18891));
  nor2s1 _______442358(.DIN1 (___0_____27281), .DIN2 (___0_____27620),
       .Q (___0_____27717));
  and2s1 _____9_442359(.DIN1 (___0_____27635), .DIN2 (_________34485),
       .Q (___0_____27716));
  nor2s1 _____9_442360(.DIN1 (___0__0__27714), .DIN2 (___0_____27625),
       .Q (___0_____27715));
  xor2s1 _______442361(.DIN1 (___0_____27577), .DIN2 (_________33174),
       .Q (___0__9__27713));
  or2s1 _____442362(.DIN1 (___0_____27711), .DIN2 (___0__9__27636), .Q
       (___0_____27712));
  nnd2s1 _______442363(.DIN1 (___0_____27633), .DIN2 (___0_____27709),
       .Q (___0_____27710));
  nnd2s1 _______442364(.DIN1 (___0_____27630), .DIN2 (________23109),
       .Q (___0_____27708));
  nor2s1 _______442365(.DIN1 (___099__24428), .DIN2 (___0_____27629),
       .Q (___0_____27707));
  and2s1 _______442366(.DIN1 (___0__9__27627), .DIN2 (___0_____27705),
       .Q (___0_____27706));
  nor2s1 ______442367(.DIN1 (___90___26149), .DIN2 (___0_____27626), .Q
       (___0__0__27704));
  nnd2s1 _______442368(.DIN1 (___0_____27619), .DIN2 (__9_____26370),
       .Q (___0__9__27703));
  and2s1 _______442369(.DIN1 (___0_____27634), .DIN2 (_____0__25012),
       .Q (___0_____27702));
  nor2s1 ______442370(.DIN1 (___0_____27631), .DIN2 (___0_____27613),
       .Q (___0_____27701));
  nnd2s1 _____0_442371(.DIN1 (___0_____27611), .DIN2 (___0_____27998),
       .Q (___0_____27700));
  or2s1 _____9_442372(.DIN1 (___0_____27698), .DIN2 (___0_____27632),
       .Q (___0_____27699));
  nor2s1 _____0_442373(.DIN1 (___0_____27696), .DIN2 (___0__0__27618),
       .Q (___0_____27697));
  or2s1 _____0_442374(.DIN1 (___0_____27767), .DIN2 (___0_____27623),
       .Q (___0_____27695));
  nnd2s1 _____0_442375(.DIN1 (___0_____27621), .DIN2 (________24040),
       .Q (___0__0__27694));
  nor2s1 _____0_442376(.DIN1 (____0___24611), .DIN2 (___0_____27616),
       .Q (___0__9__27693));
  nor2s1 _____0_442377(.DIN1 (____90__25165), .DIN2 (___0_____27624),
       .Q (___0_____27692));
  hi1s1 _____9_442378(.DIN (_____0___28807), .Q (___09____28064));
  xor2s1 _______442379(.DIN1 (_____99__34517), .DIN2 (___0_____27667),
       .Q (_________29594));
  nnd2s1 ______442380(.DIN1 (___0__9__27617), .DIN2 (___0_____27690),
       .Q (___0_____27691));
  nnd2s1 _____9_442381(.DIN1 (___0_____27603), .DIN2 (________23701),
       .Q (___0_____27689));
  nor2s1 ______442382(.DIN1 (________23932), .DIN2 (___0_____27610), .Q
       (___0_____27688));
  nor2s1 _______442383(.DIN1 (________24954), .DIN2 (___0_____27595),
       .Q (___0_____27687));
  and2s1 _______442384(.DIN1 (___0__0__27685), .DIN2 (___0_____27683),
       .Q (___0_____27686));
  nor2s1 _______442385(.DIN1 (___0_____27683), .DIN2 (___0__0__27685),
       .Q (___0__9__27684));
  nor2s1 ______442386(.DIN1 (________23869), .DIN2 (___0_____27604), .Q
       (___0_____27682));
  nnd2s1 ______442387(.DIN1 (___0__9__27675), .DIN2 (____9____29052),
       .Q (___0_____27681));
  nor2s1 _______442388(.DIN1 (________24662), .DIN2 (___0__9__27598),
       .Q (___0_____27680));
  nor2s1 _______442389(.DIN1 (___0_0___27370), .DIN2 (___0_____27602),
       .Q (___0_____27679));
  and2s1 _______442390(.DIN1 (___0_____27596), .DIN2 (___0_____27524),
       .Q (___0_____27678));
  nor2s1 _______442391(.DIN1 (________24902), .DIN2 (___0_____27601),
       .Q (___0_____27677));
  nnd2s1 _______442392(.DIN1 (___0__9__27675), .DIN2 (___0_____27674),
       .Q (___0__0__27676));
  nnd2s1 ______442393(.DIN1 (___0_____27670), .DIN2 (outData[17]), .Q
       (___0_____27673));
  nnd2s1 _______442394(.DIN1 (___0__9__27608), .DIN2 (_________31505),
       .Q (___0_____27672));
  and2s1 _______442395(.DIN1 (___0_____27671), .DIN2 (___0_____27622),
       .Q (___0_____27729));
  or2s1 _______442396(.DIN1 (outData[17]), .DIN2 (___0_____27670), .Q
       (___0_99__27752));
  hi1s1 ______442397(.DIN (___0_____27669), .Q (___0__0__27762));
  nor2s1 ______442398(.DIN1 (outData[18]), .DIN2 (___0_____27671), .Q
       (___0_____27773));
  dffacs1 _______________________442399(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27605), .QN (_____________________18638));
  dffacs1 _______________________442400(.CLRB (reset), .CLK (clk), .DIN
       (___0__0__27628), .QN (_____________________18619));
  or2s1 ______442401(.DIN1 (________21039), .DIN2 (___0_____27667), .Q
       (___0_____27668));
  nnd2s1 _______442402(.DIN1 (___0_0___27565), .DIN2 (___0_09__27665),
       .Q (___0__0__27666));
  nnd2s1 ______442403(.DIN1 (___0__0__27579), .DIN2 (___0____25329), .Q
       (___0_0___27664));
  nnd2s1 _______442404(.DIN1 (___0_____27586), .DIN2 (___0_0___27659),
       .Q (___0_0___27663));
  nnd2s1 _______442405(.DIN1 (___0_____27585), .DIN2 (____0___23624),
       .Q (___0_0___27662));
  nor2s1 _______442406(.DIN1 (____9___25846), .DIN2 (___0_____27584),
       .Q (___0_0___27661));
  nnd2s1 _______442407(.DIN1 (___0_____27583), .DIN2 (___0_0___27659),
       .Q (___0_0___27660));
  nnd2s1 _______442408(.DIN1 (___0_9___27554), .DIN2 (________22041),
       .Q (___0_0___27658));
  nnd2s1 _______442409(.DIN1 (___0_____27572), .DIN2 (___0_____27318),
       .Q (___0_0___27657));
  and2s1 _______442410(.DIN1 (___0_____27574), .DIN2 (___09____28078),
       .Q (___0_00__27656));
  nnd2s1 _______442411(.DIN1 (___0_9___27552), .DIN2 (____9___25167),
       .Q (___0_99__27655));
  xor2s1 _______442412(.DIN1 (___0__0__27541), .DIN2 (_________33564),
       .Q (___0_____28000));
  nnd2s1 _______442413(.DIN1 (___0_____27582), .DIN2 (___0_____27479),
       .Q (___0_0___27857));
  hi1s1 _____442414(.DIN (___0_9___27654), .Q (___0_____27738));
  xor2s1 _______442415(.DIN1 (___0_____27507), .DIN2 (___0_____27496),
       .Q (___0_9___27744));
  nnd2s1 _______442416(.DIN1 (___0__9__27578), .DIN2 (___0_____27390),
       .Q (___0_____27832));
  xor2s1 _______442417(.DIN1 (___0_____27509), .DIN2 (______0__30607),
       .Q (______9__28944));
  xor2s1 ______442418(.DIN1 (___0_____27542), .DIN2 (___0_____27581),
       .Q (_________28953));
  xor2s1 _______442419(.DIN1 (___0_____27514), .DIN2 (________20212),
       .Q (_____0___28807));
  nnd2s1 _______442420(.DIN1 (___0_0___27562), .DIN2 (_________28353),
       .Q (___0_9___27653));
  nnd2s1 _______442421(.DIN1 (___0_90__27551), .DIN2 (___999__26246),
       .Q (___0_9___27652));
  nor2s1 _______442422(.DIN1 (________24827), .DIN2 (___0_____27576),
       .Q (___0_9___27651));
  nnd2s1 _______442423(.DIN1 (___0_____27575), .DIN2 (________25043),
       .Q (___0_9___27650));
  or2s1 _______442424(.DIN1 (___0_9___27648), .DIN2 (___0_9___27555),
       .Q (___0_9___27649));
  nnd2s1 _______442425(.DIN1 (___0_____27570), .DIN2 (___0__9__27452),
       .Q (___0_9___27647));
  nnd2s1 _______442426(.DIN1 (___0_0___27566), .DIN2 (__9_____26348),
       .Q (___0_90__27646));
  nnd2s1 _______442427(.DIN1 (___0_0___27567), .DIN2 (____0___25758),
       .Q (___0__9__27645));
  nor2s1 _______442428(.DIN1 (___0_9___27940), .DIN2 (___0_9___27553),
       .Q (___0_____27644));
  nnd2s1 ______442429(.DIN1 (___0_____27571), .DIN2 (___0_9___27457),
       .Q (___0_____27643));
  nor2s1 _______442430(.DIN1 (___0_____27446), .DIN2 (___0_0___27560),
       .Q (___0_____27642));
  nor2s1 _____442431(.DIN1 (___9____23419), .DIN2 (___0_9___27558), .Q
       (___0_____27641));
  nnd2s1 _____9_442432(.DIN1 (___0_9___27556), .DIN2 (________25067),
       .Q (___0_____27640));
  xor2s1 _____0_442433(.DIN1 (___09____28065), .DIN2 (_________33564),
       .Q (___0_____27639));
  or2s1 _______442434(.DIN1 (___0__0__27637), .DIN2 (___0__9__27550),
       .Q (___0_____27638));
  xor2s1 _____442435(.DIN1 (___0_____27607), .DIN2 (___0_____27606), .Q
       (___0_____27669));
  xor2s1 ______442436(.DIN1 (outData[16]), .DIN2 (___0_____27593), .Q
       (_________30122));
  dffacs1 ____0__________________442437(.CLRB (reset), .CLK (clk), .DIN
       (___0_0___27564), .QN (____0________________18593));
  or2s1 _______442438(.DIN1 (___09____28066), .DIN2 (___0__9__27530),
       .Q (___0__9__27636));
  xor2s1 _____9_442439(.DIN1 (___0_____27476), .DIN2 (_____9___30624),
       .Q (___0_____27635));
  or2s1 _______442440(.DIN1 (_________32158), .DIN2 (___0_____27547),
       .Q (___0_____27634));
  nor2s1 _______442441(.DIN1 (________24211), .DIN2 (___0_____27528),
       .Q (___0_____27633));
  or2s1 ______442442(.DIN1 (___0_____27631), .DIN2 (___0__9__27540), .Q
       (___0_____27632));
  nor2s1 _______442443(.DIN1 (___9____24290), .DIN2 (___0_____27534),
       .Q (___0_____27630));
  nnd2s1 _______442444(.DIN1 (___0_____27548), .DIN2 (________23159),
       .Q (___0_____27629));
  nnd2s1 _______442445(.DIN1 (___0_____27535), .DIN2 (___00____27215),
       .Q (___0__0__27628));
  and2s1 _______442446(.DIN1 (___0__0__27531), .DIN2 (__90____26284),
       .Q (___0__9__27627));
  or2s1 _______442447(.DIN1 (___0____25350), .DIN2 (___0_____27522), .Q
       (___0_____27626));
  nnd2s1 _______442448(.DIN1 (___0_____27532), .DIN2 (________24627),
       .Q (___0_____27625));
  nnd2s1 _______442449(.DIN1 (___0_____27526), .DIN2 (___09___25358),
       .Q (___0_____27624));
  or2s1 _______442450(.DIN1 (___0_____27877), .DIN2 (___0_____27525),
       .Q (___0_____27623));
  nnd2s1 _______442451(.DIN1 (___0_____27591), .DIN2 (outData[17]), .Q
       (___0_____27622));
  nor2s1 _______442452(.DIN1 (________24048), .DIN2 (___0_____27516),
       .Q (___0_____27621));
  or2s1 _______442453(.DIN1 (___0_____27811), .DIN2 (___0__0__27521),
       .Q (___0_____27620));
  nor2s1 _______442454(.DIN1 (________25782), .DIN2 (___0_____27533),
       .Q (___0_____27619));
  nnd2s1 ______442455(.DIN1 (___0_____27499), .DIN2 (_____0__25770), .Q
       (___0__0__27618));
  nor2s1 _____9_442456(.DIN1 (___0_____27505), .DIN2 (___0_____27537),
       .Q (___0__9__27617));
  nnd2s1 _____9_442457(.DIN1 (___0_____27517), .DIN2 (________23946),
       .Q (___0_____27616));
  xor2s1 _______442458(.DIN1 (___9____23390), .DIN2 (___0_____27615),
       .Q (___0_9___27654));
  nnd2s1 _____0_442459(.DIN1 (___0_____27538), .DIN2 (___0_____27612),
       .Q (___0_____27613));
  nor2s1 _____442460(.DIN1 (____0____28172), .DIN2 (___0_____27518), .Q
       (___0_____27611));
  nnd2s1 _______442461(.DIN1 (___0_____27515), .DIN2 (___0__0__27609),
       .Q (___0_____27610));
  nor2s1 _______442462(.DIN1 (___0_____27607), .DIN2 (___0_____27606),
       .Q (___0__9__27608));
  nnd2s1 _______442463(.DIN1 (___0_____27504), .DIN2 (__9__9__26691),
       .Q (___0_____27605));
  nnd2s1 ______442464(.DIN1 (___0_____27503), .DIN2 (___0__0__27802),
       .Q (___0_____27604));
  nor2s1 _______442465(.DIN1 (________23184), .DIN2 (___0_____27502),
       .Q (___0_____27603));
  nnd2s1 _______442466(.DIN1 (___0_____27498), .DIN2 (___0_____27289),
       .Q (___0_____27602));
  nnd2s1 _______442467(.DIN1 (___0__9__27500), .DIN2 (___0_____27600),
       .Q (___0_____27601));
  xor2s1 ____442468(.DIN1 (___0_____27450), .DIN2 (_________35086), .Q
       (___0__0__27599));
  nnd2s1 ______442469(.DIN1 (___0__9__27510), .DIN2 (_____9___34924),
       .Q (___0__9__27598));
  nnd2s1 ______442470(.DIN1 (___0_____27606), .DIN2 (___9____26228), .Q
       (___0_____27597));
  nor2s1 _______442471(.DIN1 (___0_____27529), .DIN2 (___0__0__27501),
       .Q (___0_____27596));
  nnd2s1 _______442472(.DIN1 (___0_____27506), .DIN2 (___0_____27594),
       .Q (___0_____27595));
  or2s1 _____442473(.DIN1 (outData[16]), .DIN2 (___0_____27593), .Q
       (___0_____27670));
  nnd2s1 _______442474(.DIN1 (___0_____27592), .DIN2 (_________18851),
       .Q (___0_____27674));
  or2s1 _______442475(.DIN1 (_________18851), .DIN2 (___0_____27592),
       .Q (___0__9__27675));
  or2s1 _______442476(.DIN1 (outData[17]), .DIN2 (___0_____27591), .Q
       (___0_____27671));
  and2s1 ____90_442477(.DIN1 (___0_____27593), .DIN2 (___0_____27351),
       .Q (___0__0__27685));
  dffacs1 _______________________442478(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27523), .QN (_____________________18625));
  dffacs1 _______________________442479(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27519), .QN (_____________________18667));
  dffacs1 _______________________442480(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27497), .QN (_____________________18626));
  or2s1 _______442481(.DIN1 (________________18706), .DIN2
       (___0__0__27589), .Q (___0_____27590));
  and2s1 _______442482(.DIN1 (___0__0__27589), .DIN2
       (________________18706), .Q (___0__9__27588));
  nnd2s1 _______442483(.DIN1 (___0_____27493), .DIN2 (__9__0__27005),
       .Q (___0_____27587));
  and2s1 ______442484(.DIN1 (___0__9__27490), .DIN2 (____90___28999),
       .Q (___0_____27586));
  nor2s1 ______442485(.DIN1 (________24123), .DIN2 (___0_____27489), .Q
       (___0_____27585));
  nnd2s1 _______442486(.DIN1 (___0_____27488), .DIN2 (__9_____27006),
       .Q (___0_____27584));
  nor2s1 _______442487(.DIN1 (___0_0__25328), .DIN2 (___0_____27487),
       .Q (___0_____27583));
  or2s1 _______442488(.DIN1 (___0_____27581), .DIN2 (___0_____27482),
       .Q (___0_____27582));
  or2s1 _____9_442489(.DIN1 (_____0__22310), .DIN2 (___0_____27615), .Q
       (___0_____27580));
  nor2s1 _____9_442490(.DIN1 (________22686), .DIN2 (___0_____27492),
       .Q (___0__0__27579));
  nnd2s1 _____0_442491(.DIN1 (___0__9__27480), .DIN2 (___0_0___27369),
       .Q (___0__9__27578));
  and2s1 _____0_442492(.DIN1 (___0_____27615), .DIN2 (___9____23389),
       .Q (___0_____27577));
  nnd2s1 _______442493(.DIN1 (___0_0___27467), .DIN2 (_____9__24738),
       .Q (___0_____27576));
  nor2s1 _______442494(.DIN1 (________24454), .DIN2 (___0_0___27465),
       .Q (___0_____27575));
  and2s1 _______442495(.DIN1 (___0_0___27468), .DIN2 (___0_____27573),
       .Q (___0_____27574));
  nor2s1 _______442496(.DIN1 (___909__25183), .DIN2 (___0_00__27461),
       .Q (___0_____27572));
  or2s1 _______442497(.DIN1 (outData[5]), .DIN2 (___0__0__27569), .Q
       (___0_____27571));
  nnd2s1 _______442498(.DIN1 (___0__0__27569), .DIN2 (___9____25205),
       .Q (___0_____27570));
  xor2s1 _____0_442499(.DIN1 (___0_____27415), .DIN2 (___0_09__27568),
       .Q (___0_____27667));
  xor2s1 _______442500(.DIN1 (outData[16]), .DIN2 (___0_____27508), .Q
       (____0____29106));
  nor2s1 ______442501(.DIN1 (___0_____27451), .DIN2 (________22795), .Q
       (___0_0___27567));
  or2s1 _______442502(.DIN1 (_____0___28805), .DIN2 (___0_____27484),
       .Q (___0_0___27566));
  nor2s1 _______442503(.DIN1 (___0_____27303), .DIN2 (___0_____27472),
       .Q (___0_0___27565));
  nnd2s1 _______442504(.DIN1 (___0_0___27463), .DIN2 (___0_0___27563),
       .Q (___0_0___27564));
  nor2s1 _______442505(.DIN1 (___0_0___27561), .DIN2 (___0_0___27466),
       .Q (___0_0___27562));
  nnd2s1 _______442506(.DIN1 (___0_99__27460), .DIN2 (___0_____27800),
       .Q (___0_0___27560));
  or2s1 _______442507(.DIN1 (___0_9___27557), .DIN2 (___0_90__27453),
       .Q (___0_9___27558));
  nor2s1 ______442508(.DIN1 (________24677), .DIN2 (___0__0__27471), .Q
       (___0_9___27556));
  nnd2s1 ______442509(.DIN1 (___0_____27474), .DIN2 (________26123), .Q
       (___0_9___27555));
  nor2s1 _______442510(.DIN1 (_____0__22914), .DIN2 (___0_09__27470),
       .Q (___0_9___27554));
  or2s1 _______442511(.DIN1 (___0_____27921), .DIN2 (___0_9___27458),
       .Q (___0_9___27553));
  nor2s1 _______442512(.DIN1 (________24716), .DIN2 (___0_9___27454),
       .Q (___0_9___27552));
  and2s1 _______442513(.DIN1 (___0_9___27455), .DIN2 (___0__0__27802),
       .Q (___0_90__27551));
  or2s1 ____9__442514(.DIN1 (___0_____27549), .DIN2 (___0_0___27462),
       .Q (___0__9__27550));
  xor2s1 _____9_442515(.DIN1 (___0_____27400), .DIN2 (_________28939),
       .Q (____0____28164));
  dffacs1 _______________________442516(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27486), .QN (_____________________18605));
  dffacs1 _______________________442517(.CLRB (reset), .CLK (clk), .DIN
       (___0_0___27469), .QN (_____________________18635));
  dffacs1 ______________________0_442518(.CLRB (reset), .CLK (clk),
       .DIN (___0_____27478), .QN (__________________0___18670));
  dffacs1 _______________________442519(.CLRB (reset), .CLK (clk), .DIN
       (___0_0___27464), .QN (_____________________18621));
  nnd2s1 _______442520(.DIN1 (___0__9__27442), .DIN2 (________21469),
       .Q (___0_____27548));
  xnr2s1 ______442521(.DIN1 (____________0___18686), .DIN2
       (_________29326), .Q (___0_____27547));
  nor2s1 _______442522(.DIN1 (___0_____27543), .DIN2 (___0_____27544),
       .Q (___0_____27546));
  nnd2s1 _____0_442523(.DIN1 (___0_____27544), .DIN2 (___0_____27543),
       .Q (___0_____27545));
  xor2s1 _____0_442524(.DIN1 (____________0___18769), .DIN2
       (_________29326), .Q (___0_____27542));
  xor2s1 _____0_442525(.DIN1 (__9_____26482), .DIN2 (_________29326),
       .Q (___0__0__27541));
  or2s1 _______442526(.DIN1 (___0_____27539), .DIN2 (___0__9__27432),
       .Q (___0__9__27540));
  nor2s1 _______442527(.DIN1 (____9___24976), .DIN2 (___0_____27436),
       .Q (___0_____27538));
  nnd2s1 ______442528(.DIN1 (___0_____27437), .DIN2 (___0_____27536),
       .Q (___0_____27537));
  and2s1 ______442529(.DIN1 (___0__0__27423), .DIN2 (____09__25956), .Q
       (___0_____27535));
  nnd2s1 _______442530(.DIN1 (___0__0__27443), .DIN2 (___0_9___27357),
       .Q (___0_____27534));
  nnd2s1 _______442531(.DIN1 (___0_____27438), .DIN2 (____0___25560),
       .Q (___0_____27533));
  and2s1 _______442532(.DIN1 (___0_____27434), .DIN2 (________25971),
       .Q (___0_____27532));
  nor2s1 _______442533(.DIN1 (________23025), .DIN2 (___0_____27441),
       .Q (___0__0__27531));
  or2s1 _______442534(.DIN1 (___0_____27529), .DIN2 (___0_____27427),
       .Q (___0__9__27530));
  nnd2s1 _______442535(.DIN1 (___0_____27428), .DIN2 (___0_____27527),
       .Q (___0_____27528));
  nor2s1 _______442536(.DIN1 (_____9__23637), .DIN2 (___0_____27448),
       .Q (___0_____27526));
  nnd2s1 _______442537(.DIN1 (___0__9__27422), .DIN2 (___0_____27524),
       .Q (___0_____27525));
  nnd2s1 _______442538(.DIN1 (___0_____27429), .DIN2 (__9_____26377),
       .Q (___0_____27523));
  nor2s1 ______442539(.DIN1 (_____0___28805), .DIN2 (___0_____27431),
       .Q (___0_____27522));
  or2s1 _______442540(.DIN1 (___0__9__27520), .DIN2 (___0_____27425),
       .Q (___0__0__27521));
  nnd2s1 _______442541(.DIN1 (___0_____27426), .DIN2 (___0_____27912),
       .Q (___0_____27519));
  or2s1 _______442542(.DIN1 (___09____28117), .DIN2 (___0_____27447),
       .Q (___0_____27518));
  nor2s1 _______442543(.DIN1 (___0____23503), .DIN2 (___0_____27435),
       .Q (___0_____27517));
  nnd2s1 _______442544(.DIN1 (___0_____27439), .DIN2 (________25055),
       .Q (___0_____27516));
  nor2s1 ____9__442545(.DIN1 (__9_____26773), .DIN2 (___0__9__27412),
       .Q (___0_____27515));
  xor2s1 _____442546(.DIN1 (___0_9___27456), .DIN2 (_________35086), .Q
       (___0_____27514));
  nor2s1 _____9_442547(.DIN1 (___0_____27512), .DIN2 (___0__0__27511),
       .Q (___0_____27513));
  nor2s1 ____9__442548(.DIN1 (__9_____26964), .DIN2 (___0__0__27413),
       .Q (___0__9__27510));
  nor2s1 _____9_442549(.DIN1 (___0_____27445), .DIN2 (___0_____27508),
       .Q (___0_____27509));
  xor2s1 _____9_442550(.DIN1 (_________28692), .DIN2 (________24042),
       .Q (___0_____27507));
  nor2s1 ____9__442551(.DIN1 (___0_____27505), .DIN2 (___0__0__27393),
       .Q (___0_____27506));
  nor2s1 ____9__442552(.DIN1 (___0_____27405), .DIN2 (___0_____27280),
       .Q (___0_____27504));
  and2s1 ____9__442553(.DIN1 (___0_____27407), .DIN2 (__9_____26722),
       .Q (___0_____27503));
  nnd2s1 ____9__442554(.DIN1 (___0_____27414), .DIN2 (_____9__24745),
       .Q (___0_____27502));
  nnd2s1 ____9__442555(.DIN1 (___0_____27401), .DIN2 (________23913),
       .Q (___0__0__27501));
  nor2s1 ____9__442556(.DIN1 (________25831), .DIN2 (___0_____27411),
       .Q (___0__9__27500));
  nor2s1 _______442557(.DIN1 (________23752), .DIN2 (___0_____27424),
       .Q (___0_____27499));
  nor2s1 ____9_442558(.DIN1 (________23233), .DIN2 (___0_____27404), .Q
       (___0_____27498));
  nnd2s1 ____9__442559(.DIN1 (___0_____27395), .DIN2 (__9_____26360),
       .Q (___0_____27497));
  nnd2s1 ____9__442560(.DIN1 (___0_____27409), .DIN2 (___0_____27399),
       .Q (___0_____27592));
  nnd2s1 _____9_442561(.DIN1 (___0_____27508), .DIN2 (________19231),
       .Q (___0_____27591));
  nor2s1 _____9_442562(.DIN1 (___0_____27496), .DIN2 (___0_____27418),
       .Q (___0_____27614));
  xor2s1 ____9__442563(.DIN1 (___0_____27350), .DIN2 (______0__30283),
       .Q (___0_____27593));
  dffacs1 _____________________9_442564(.CLRB (reset), .CLK (clk), .DIN
       (___0__0__27433), .QN (_________________9___18627));
  nnd2s1 ____9_442565(.DIN1 (___0_____27397), .DIN2 (__9_0___26610), .Q
       (___0_____27606));
  dffacs1 _______________________442566(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27394), .QN (_____________________18634));
  hi1s1 ____9__442567(.DIN (___0_____27495), .Q (___09____28065));
  dffacs1 ________________________442568(.CLRB (reset), .CLK (clk),
       .DIN (___0_____27444), .QN (______________________18629));
  dffacs1 ____0__________________442569(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27440), .QN (____0________________18651));
  and2s1 _______442570(.DIN1 (___0_____27475), .DIN2 (_________29326),
       .Q (___0_____27494));
  nnd2s1 _______442571(.DIN1 (___0__0__27491), .DIN2 (________22243),
       .Q (___0_____27493));
  nnd2s1 _______442572(.DIN1 (___0__0__27491), .DIN2 (____99__26046),
       .Q (___0_____27492));
  and2s1 _______442573(.DIN1 (___0_____27379), .DIN2 (________25824),
       .Q (___0__9__27490));
  nnd2s1 ______442574(.DIN1 (___0_____27382), .DIN2 (____00__23618), .Q
       (___0_____27489));
  nnd2s1 ______442575(.DIN1 (___0_____27388), .DIN2 (___0_____27386),
       .Q (___0_____27488));
  nnd2s1 _______442576(.DIN1 (___0_____27387), .DIN2 (________25822),
       .Q (___0_____27487));
  nnd2s1 ____9__442577(.DIN1 (___0_____27378), .DIN2 (___0_____27485),
       .Q (___0_____27486));
  nor2s1 ____9__442578(.DIN1 (___0_____27483), .DIN2 (___0_____27375),
       .Q (___0_____27484));
  nor2s1 ______442579(.DIN1 (___0__0__27481), .DIN2 (_________29326),
       .Q (___0_____27482));
  xor2s1 _______442580(.DIN1 (___0_____27391), .DIN2 (___0_09__27568),
       .Q (___0__9__27480));
  nnd2s1 _______442581(.DIN1 (_________29326), .DIN2 (___0__0__27481),
       .Q (___0_____27479));
  or2s1 _______442582(.DIN1 (___0_____27477), .DIN2 (___0_____27385),
       .Q (___0_____27478));
  nor2s1 _____9_442583(.DIN1 (_________29326), .DIN2 (___0_____27475),
       .Q (___0_____27476));
  and2s1 ____9_442584(.DIN1 (___0_0___27365), .DIN2 (___0_____27473),
       .Q (___0_____27474));
  nnd2s1 ____90_442585(.DIN1 (___0_0___27372), .DIN2 (_____0__24666),
       .Q (___0_____27472));
  nor2s1 ____90_442586(.DIN1 (___00____27202), .DIN2 (___0__0__27374),
       .Q (___0__0__27471));
  nnd2s1 ____90_442587(.DIN1 (___0_9___27355), .DIN2 (__99____27150),
       .Q (___0_09__27470));
  nnd2s1 ____90_442588(.DIN1 (___0_9___27360), .DIN2 (___0_0___27272),
       .Q (___0_0___27469));
  nnd2s1 ______442589(.DIN1 (___0__9__27383), .DIN2 (___0_0___27368),
       .Q (___0__0__27589));
  or2s1 ______442590(.DIN1 (____________0___18686), .DIN2
       (_________29326), .Q (_________29287));
  xor2s1 ____90_442591(.DIN1 (___0_____27312), .DIN2 (_________32554),
       .Q (___0_____27615));
  nor2s1 ____9__442592(.DIN1 (_____0__24534), .DIN2 (___0_____27377),
       .Q (___0_0___27468));
  nor2s1 ____9_442593(.DIN1 (________25631), .DIN2 (___0_____27380), .Q
       (___0_0___27467));
  or2s1 ____9_442594(.DIN1 (__99_0__27144), .DIN2 (___0_9___27358), .Q
       (___0_0___27466));
  or2s1 ____9__442595(.DIN1 (__999___27167), .DIN2 (___0_09__27373), .Q
       (___0_0___27465));
  or2s1 ____9__442596(.DIN1 (__9_____26391), .DIN2 (___0_____27389), .Q
       (___0_0___27464));
  and2s1 ____9__442597(.DIN1 (___0_0___27366), .DIN2 (________23733),
       .Q (___0_0___27463));
  nnd2s1 ____0__442598(.DIN1 (___0_____27347), .DIN2 (____9___24513),
       .Q (___0_0___27462));
  nor2s1 ____9__442599(.DIN1 (__9_____26621), .DIN2 (___0_9___27362),
       .Q (___0_00__27461));
  nor2s1 ____9__442600(.DIN1 (___0_9___27459), .DIN2 (___0_9___27361),
       .Q (___0_99__27460));
  nnd2s1 ____9_442601(.DIN1 (___0_0___27367), .DIN2 (____0___23806), .Q
       (___0_9___27458));
  nnd2s1 ____9__442602(.DIN1 (___0_9___27456), .DIN2 (outData[7]), .Q
       (___0_9___27457));
  and2s1 ____9__442603(.DIN1 (___0_____27376), .DIN2 (________22677),
       .Q (___0_9___27455));
  nnd2s1 ____9__442604(.DIN1 (___0_9___27359), .DIN2 (________21886),
       .Q (___0_9___27454));
  nnd2s1 ____9__442605(.DIN1 (___0_90__27354), .DIN2 (________23702),
       .Q (___0_90__27453));
  or2s1 ____9__442606(.DIN1 (________19440), .DIN2 (___0_9___27456), .Q
       (___0__9__27452));
  nor2s1 ____9_442607(.DIN1 (___0_00__27364), .DIN2 (___9____25213), .Q
       (___0_____27451));
  and2s1 ____0_442608(.DIN1 (___0_____27449), .DIN2 (___00_0__27247),
       .Q (___0_____27450));
  nor2s1 ____9__442609(.DIN1 (____9____29052), .DIN2 (___0__9__27353),
       .Q (___0_9___27559));
  xor2s1 ____9_442610(.DIN1 (__9_____26715), .DIN2 (___0_____27396), .Q
       (___0_____27495));
  nor2s1 ____9_442611(.DIN1 (outData[7]), .DIN2 (___0_9___27456), .Q
       (___0__0__27569));
  dffacs1 _____________________9_442612(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27346), .Q (_________________9___18642));
  dffacs1 _______________________442613(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27352), .QN (_____________________18603));
  nnd2s1 ____9__442614(.DIN1 (___0__0__27316), .DIN2 (_____9__24569),
       .Q (___0_____27448));
  or2s1 ____90_442615(.DIN1 (___0_____27446), .DIN2 (___0_____27321),
       .Q (___0_____27447));
  nor2s1 ____90_442616(.DIN1 (_____________18896), .DIN2
       (___0_____27421), .Q (___0_____27445));
  nnd2s1 ____442617(.DIN1 (___0__0__27335), .DIN2 (__9_____26913), .Q
       (___0_____27444));
  nor2s1 ____9__442618(.DIN1 (____00__23802), .DIN2 (___0__0__27325),
       .Q (___0__0__27443));
  nnd2s1 ____9__442619(.DIN1 (___0_____27333), .DIN2 (___0_0__23500),
       .Q (___0__9__27442));
  nor2s1 ____9_442620(.DIN1 (________21758), .DIN2 (___0_____27332), .Q
       (___0_____27441));
  nnd2s1 ____9__442621(.DIN1 (___0_____27331), .DIN2 (_________28942),
       .Q (___0_____27440));
  nor2s1 ____9__442622(.DIN1 (____9___25647), .DIN2 (___0__0__27345),
       .Q (___0_____27439));
  nor2s1 ____9__442623(.DIN1 (___9_0__22472), .DIN2 (___0_____27328),
       .Q (___0_____27438));
  nor2s1 ____9__442624(.DIN1 (____9___25075), .DIN2 (___0_____27337),
       .Q (___0_____27437));
  nnd2s1 ____9__442625(.DIN1 (___0_____27323), .DIN2 (________24451),
       .Q (___0_____27436));
  nnd2s1 ____9__442626(.DIN1 (___0_____27313), .DIN2 (________23148),
       .Q (___0_____27435));
  nor2s1 ______442627(.DIN1 (___0____22574), .DIN2 (___0_____27343), .Q
       (___0_____27434));
  nnd2s1 ____9__442628(.DIN1 (___0__9__27334), .DIN2 (__9_____26552),
       .Q (___0__0__27433));
  nnd2s1 ____9_442629(.DIN1 (___0__9__27315), .DIN2 (________24463), .Q
       (___0__9__27432));
  nor2s1 ____9_442630(.DIN1 (___0_____27430), .DIN2 (___0_____27320),
       .Q (___0_____27431));
  nor2s1 ____9__442631(.DIN1 (__9_____26690), .DIN2 (___0_____27326),
       .Q (___0_____27429));
  nor2s1 ____9__442632(.DIN1 (________25541), .DIN2 (___0_____27340),
       .Q (___0_____27428));
  nnd2s1 ____9__442633(.DIN1 (___0_____27319), .DIN2 (____0___23719),
       .Q (___0_____27427));
  and2s1 ____9_442634(.DIN1 (___0_____27338), .DIN2 (___0_0___27755),
       .Q (___0_____27426));
  nnd2s1 ____9_442635(.DIN1 (___0_____27339), .DIN2 (___9____25253), .Q
       (___0_____27425));
  nnd2s1 ____9__442636(.DIN1 (___0_____27301), .DIN2 (__9_____26358),
       .Q (___0_____27424));
  nnd2s1 ____9__442637(.DIN1 (___0_____27317), .DIN2 (___00____27211),
       .Q (___0__0__27423));
  nor2s1 ____9__442638(.DIN1 (__9_____26959), .DIN2 (___0__9__27344),
       .Q (___0__9__27422));
  and2s1 ____9__442639(.DIN1 (___0_____27421), .DIN2
       (_____________18896), .Q (___0_____27508));
  nnd2s1 ____0__442640(.DIN1 (___0_____27419), .DIN2
       (_________________18741), .Q (___0_____27420));
  nor2s1 ____9__442641(.DIN1 (outData[0]), .DIN2 (___0__9__27402), .Q
       (___0_____27418));
  nor2s1 ____0__442642(.DIN1 (___0_____27416), .DIN2 (___0_____27348),
       .Q (___0_____27417));
  nor2s1 ____9__442643(.DIN1 (__90____26267), .DIN2 (___0_____27330),
       .Q (___0_____27415));
  and2s1 ____0_442644(.DIN1 (___0_____27299), .DIN2 (___0_____27862),
       .Q (___0_____27414));
  nnd2s1 ____0_442645(.DIN1 (___0_____27295), .DIN2 (__99____27157), .Q
       (___0__0__27413));
  nnd2s1 ____99_442646(.DIN1 (___0__0__27307), .DIN2 (__9_00), .Q
       (___0__9__27412));
  nnd2s1 ____99_442647(.DIN1 (___0_____27298), .DIN2 (___0_____27410),
       .Q (___0_____27411));
  nnd2s1 ____99_442648(.DIN1 (___0_____27398), .DIN2 (_________28939),
       .Q (___0_____27409));
  or2s1 ____00_442649(.DIN1 (_________________18741), .DIN2
       (___0_____27419), .Q (___0_____27408));
  nor2s1 ____00_442650(.DIN1 (___0_____27406), .DIN2 (___0_____27308),
       .Q (___0_____27407));
  nnd2s1 ____442651(.DIN1 (___0_____27305), .DIN2 (__90_9__26327), .Q
       (___0_____27405));
  nnd2s1 ____0__442652(.DIN1 (___0_____27304), .DIN2 (___90___26151),
       .Q (___0_____27404));
  nnd2s1 ____9_442653(.DIN1 (___0__9__27402), .DIN2 (outData[0]), .Q
       (___0__0__27403));
  and2s1 ____0_442654(.DIN1 (___0_____27302), .DIN2 (___9____24279), .Q
       (___0_____27401));
  and2s1 ____0__442655(.DIN1 (___0_____27399), .DIN2 (___0_____27398),
       .Q (___0_____27400));
  nnd2s1 ____0__442656(.DIN1 (___0_____27396), .DIN2 (__9_0___26611),
       .Q (___0_____27397));
  nor2s1 ____0__442657(.DIN1 (__9_0___26994), .DIN2 (___0__9__27296),
       .Q (___0_____27395));
  nnd2s1 ____0__442658(.DIN1 (___0__9__27306), .DIN2 (__99____27100),
       .Q (___0_____27394));
  nnd2s1 ____0__442659(.DIN1 (___0__0__27297), .DIN2 (___9____25254),
       .Q (___0__0__27393));
  and2s1 ____9__442660(.DIN1 (___0__9__27392), .DIN2
       (______________________________________0__________0), .Q
       (___0__0__27511));
  and2s1 ____9__442661(.DIN1 (___0_____27391), .DIN2 (___0_____27390),
       .Q (___0_____27544));
  nor2s1 ____9__442662(.DIN1
       (______________________________________0__________0), .DIN2
       (___0__9__27392), .Q (___0_____27512));
  dffacs1 ____0__________________442663(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27314), .QN (____0________________18648));
  dffacs1 _______________________442664(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27341), .QN (_____________________18622));
  dffacs1 _______________________442665(.CLRB (reset), .CLK (clk), .DIN
       (___0_____27322), .QN (_____________________18601));
  nnd2s1 ____99_442666(.DIN1 (___0_0___27275), .DIN2 (________25933),
       .Q (___0_____27389));
  nnd2s1 ____9_442667(.DIN1 (___0_____27292), .DIN2 (___0__0__27287),
       .Q (___0_____27388));
  nnd2s1 ____9__442668(.DIN1 (___0_____27288), .DIN2 (___0_____27386),
       .Q (___0_____27387));
  nnd2s1 ____9__442669(.DIN1 (___0_____27282), .DIN2 (___0_____27536),
       .Q (___0_____27385));
  xor2s1 ____9__442670(.DIN1 (_____9___29527), .DIN2 (____9____30874),
       .Q (___0__0__27384));
  xnr2s1 ____9__442671(.DIN1 (____0____30981), .DIN2 (___00____27194),
       .Q (___0__9__27383));
  and2s1 ____9__442672(.DIN1 (___0_____27285), .DIN2 (___0_____27873),
       .Q (___0_____27382));
  nor2s1 ____9__442673(.DIN1 (________22146), .DIN2 (___0_____27283),
       .Q (___0_____27381));
  nnd2s1 ____0__442674(.DIN1 (___009___27263), .DIN2 (_____9__26116),
       .Q (___0_____27380));
  nor2s1 ____9__442675(.DIN1 (____99__25849), .DIN2 (___0_____27279),
       .Q (___0_____27379));
  and2s1 ____00_442676(.DIN1 (___0_0___27274), .DIN2 (__9_9___26987),
       .Q (___0_____27378));
  nnd2s1 ____00_442677(.DIN1 (___0_0___27271), .DIN2 (___999__23436),
       .Q (___0_____27377));
  nor2s1 ____00_442678(.DIN1 (________23562), .DIN2 (___00____27255),
       .Q (___0_____27376));
  nnd2s1 ____00_442679(.DIN1 (___0099__27266), .DIN2 (__9__9__27014),
       .Q (___0_____27375));
  nor2s1 ____00_442680(.DIN1 (_____9__24719), .DIN2 (___009___27260),
       .Q (___0__0__27374));
  nnd2s1 ____0__442681(.DIN1 (___009___27261), .DIN2 (___0_____27336),
       .Q (___0_09__27373));
  nor2s1 ____0__442682(.DIN1 (___0____24406), .DIN2 (___009___27264),
       .Q (___0_0___27372));
  nor2s1 ____0__442683(.DIN1 (___0_0___27370), .DIN2 (___0_09__27276),
       .Q (___0_0___27371));
  xor2s1 _____9_442684(.DIN1 (___0_0___27369), .DIN2
       (_________________0___18618), .Q (___0_____27543));
  nnd2s1 ____0_442685(.DIN1 (___000___27173), .DIN2 (_____00__28898),
       .Q (___0_____27581));
  nor2s1 ____9__442686(.DIN1 (___0_____27430), .DIN2 (___0_____27290),
       .Q (___0__0__27491));
  xor2s1 ____9__442687(.DIN1 (_____________18895), .DIN2
       (___0_0___27368), .Q (_____9___30268));
  hi1s1 ____0__442688(.DIN (___0__9__27402), .Q (_________28692));
  xnr2s1 ____442689(.DIN1 (__90____26269), .DIN2 (___0_____27329), .Q
       (_________29326));
  nor2s1 ____0__442690(.DIN1 (________23986), .DIN2 (___00_9__27256),
       .Q (___0_0___27367));
  nor2s1 ____0__442691(.DIN1 (______9__28464), .DIN2 (___00____27251),
       .Q (___0_0___27366));
  and2s1 ____0__442692(.DIN1 (___00____27254), .DIN2 (________24000),
       .Q (___0_0___27365));
  xor2s1 ____0__442693(.DIN1 (___0_99__27363), .DIN2 (__90_9__26270),
       .Q (___0_00__27364));
  nor2s1 ____0__442694(.DIN1 (________21758), .DIN2 (___009___27259),
       .Q (___0_9___27362));
  nnd2s1 ____0_442695(.DIN1 (___0_____27293), .DIN2 (________24485), .Q
       (___0_9___27361));
  nor2s1 ____0__442696(.DIN1 (___09___23521), .DIN2 (___0_0___27270),
       .Q (___0_9___27360));
  nor2s1 ____0__442697(.DIN1 (____00__23528), .DIN2 (___009___27262),
       .Q (___0_9___27359));
  nnd2s1 ____0__442698(.DIN1 (___009___27265), .DIN2 (___0_9___27357),
       .Q (___0_9___27358));
  nnd2s1 ____0__442699(.DIN1 (___009___27258), .DIN2 (_____9___28891),
       .Q (___0_9___27356));
  nor2s1 ____0_442700(.DIN1 (__90____26262), .DIN2 (___00____27252), .Q
       (___0_9___27355));
  nor2s1 ____0__442701(.DIN1 (________23726), .DIN2 (___0_0___27269),
       .Q (___0_90__27354));
  xor2s1 ____0__442702(.DIN1 (___0009__27178), .DIN2 (______0__33107),
       .Q (___0__9__27353));
  nnd2s1 _____9_442703(.DIN1 (___00____27249), .DIN2 (___0_____27485),
       .Q (___0_____27352));
  or2s1 ____442704(.DIN1 (_____________18896), .DIN2 (___0_____27349),
       .Q (___0_____27351));
  and2s1 ______442705(.DIN1 (___0_____27349), .DIN2
       (_____________18896), .Q (___0_____27350));
  nor2s1 _______442706(.DIN1 (___9____23415), .DIN2 (___00____27243),
       .Q (___0_____27347));
  nnd2s1 _______442707(.DIN1 (___00_9__27246), .DIN2 (___9____25236),
       .Q (___0_____27346));
  xnr2s1 _____9_442708(.DIN1 (___0____21656), .DIN2 (___00____27192),
       .Q (___0_____27449));
  dffacs1 _________________0_442709(.CLRB (reset), .CLK (clk), .DIN
       (___00____27245), .QN (_____________0___18679));
  dffacs1 _______________________442710(.CLRB (reset), .CLK (clk), .DIN
       (___0_0___27273), .QN (_____________________18637));
  nnd2s1 ____09_442711(.DIN1 (___0_0___27268), .DIN2 (________22872),
       .Q (___0_9___27456));
  dffacs1 _______________________442712(.CLRB (reset), .CLK (clk), .DIN
       (___00____27253), .QN (_____________________18620));
  dffacs1 _______________________442713(.CLRB (reset), .CLK (clk), .DIN
       (___00____27250), .QN (_____________________18661));
  nnd2s1 ____0_442714(.DIN1 (___00____27224), .DIN2 (__9__0__26816), .Q
       (___0__0__27345));
  nnd2s1 ____0__442715(.DIN1 (___00____27240), .DIN2 (___9____23414),
       .Q (___0__9__27344));
  nnd2s1 ____9__442716(.DIN1 (___00____27241), .DIN2 (___9____26220),
       .Q (___0_____27343));
  xor2s1 ____9__442717(.DIN1 (__99____27155), .DIN2 (____0____30977),
       .Q (___0_____27342));
  nnd2s1 ____99_442718(.DIN1 (__999___27169), .DIN2 (___00____27212),
       .Q (___0_____27341));
  nnd2s1 ____99_442719(.DIN1 (___00____27239), .DIN2 (___0____24401),
       .Q (___0_____27340));
  nor2s1 ____99_442720(.DIN1 (________24687), .DIN2 (___00_0__27238),
       .Q (___0_____27339));
  nor2s1 ____442721(.DIN1 (___0_____27477), .DIN2 (___00____27234), .Q
       (___0_____27338));
  nnd2s1 ____442722(.DIN1 (___00____27210), .DIN2 (___0_____27336), .Q
       (___0_____27337));
  nor2s1 ____00_442723(.DIN1 (__9_____26475), .DIN2 (___00____27205),
       .Q (___0__0__27335));
  nor2s1 ____0_442724(.DIN1 (__9_____26649), .DIN2 (___00_0__27199), .Q
       (___0__9__27334));
  nor2s1 ____0__442725(.DIN1 (__9_____26784), .DIN2 (___00_0__27228),
       .Q (___0_____27333));
  nor2s1 ____0__442726(.DIN1 (__9_____26655), .DIN2 (___00____27226),
       .Q (___0_____27332));
  nor2s1 ____0__442727(.DIN1 (__990___27085), .DIN2 (___00____27206),
       .Q (___0_____27331));
  nor2s1 ____0__442728(.DIN1 (__90____26268), .DIN2 (___0_____27329),
       .Q (___0_____27330));
  nnd2s1 ____0__442729(.DIN1 (___00____27223), .DIN2 (__9_____26631),
       .Q (___0_____27328));
  nor2s1 ____0__442730(.DIN1 (________22657), .DIN2 (___00_9__27227),
       .Q (___0_____27327));
  nor2s1 ____0__442731(.DIN1 (___0__9__27771), .DIN2 (___00_9__27237),
       .Q (___0_____27326));
  nnd2s1 ____0__442732(.DIN1 (___00____27184), .DIN2 (___0__9__27324),
       .Q (___0__0__27325));
  nor2s1 ____0_442733(.DIN1 (__9_____26907), .DIN2 (___00____27231), .Q
       (___0_____27323));
  nnd2s1 ____0_442734(.DIN1 (___00____27236), .DIN2 (___0_____27485),
       .Q (___0_____27322));
  nnd2s1 ____0__442735(.DIN1 (___00____27214), .DIN2 (________22960),
       .Q (___0_____27321));
  nnd2s1 ____0__442736(.DIN1 (___00____27197), .DIN2 (__9_0___26517),
       .Q (___0_____27320));
  nor2s1 ____0__442737(.DIN1 (___0____23487), .DIN2 (___00_0__27208),
       .Q (___0_____27319));
  nnd2s1 ____0_442738(.DIN1 (___00____27207), .DIN2 (________21886), .Q
       (___0_____27318));
  nnd2s1 ____0__442739(.DIN1 (___00____27221), .DIN2 (__9_____26387),
       .Q (___0_____27317));
  nor2s1 ____0__442740(.DIN1 (outData[14]), .DIN2 (___0_0___27368), .Q
       (___0_____27421));
  dffacs1 _______________________442741(.CLRB (reset), .CLK (clk), .DIN
       (___00____27232), .QN (_____________________18636));
  dffacs1 __________________442742(.CLRB (reset), .CLK (clk), .DIN
       (___00____27229), .QN
       (______________________________________0_____________18890));
  nor2s1 ____0__442743(.DIN1 (__9__0__26356), .DIN2 (___00____27201),
       .Q (___0__0__27316));
  nor2s1 ____0__442744(.DIN1 (_____9__24472), .DIN2 (___00____27203),
       .Q (___0__9__27315));
  nnd2s1 ____0__442745(.DIN1 (___00_9__27198), .DIN2 (_________28942),
       .Q (___0_____27314));
  nnd2s1 ____0__442746(.DIN1 (___00____27195), .DIN2 (________21469),
       .Q (___0_____27313));
  nnd2s1 ____0__442747(.DIN1 (___00____27209), .DIN2 (___0_____27496),
       .Q (___0_____27312));
  nor2s1 ______442748(.DIN1 (___0_____27310), .DIN2 (___0_____27309),
       .Q (___0_____27311));
  nnd2s1 ____09_442749(.DIN1 (___00____27186), .DIN2 (________23952),
       .Q (___0_____27308));
  nor2s1 ____09_442750(.DIN1 (__9_____26647), .DIN2 (___00_0__27179),
       .Q (___0__0__27307));
  nor2s1 _____0_442751(.DIN1 (________25878), .DIN2 (___00____27190),
       .Q (___0__9__27306));
  nnd2s1 _______442752(.DIN1 (___00_0__27189), .DIN2 (__9_____27045),
       .Q (___0_____27305));
  nor2s1 _______442753(.DIN1 (___0_____27303), .DIN2 (___00____27204),
       .Q (___0_____27304));
  nnd2s1 _______442754(.DIN1 (___00____27183), .DIN2 (________21469),
       .Q (___0_____27302));
  nor2s1 ____0__442755(.DIN1 (__9__0__26749), .DIN2 (___00____27225),
       .Q (___0_____27301));
  nnd2s1 _____9_442756(.DIN1 (___0__0__27277), .DIN2 (___000___27176),
       .Q (___0_____27300));
  nor2s1 _______442757(.DIN1 (________24908), .DIN2 (___000___27175),
       .Q (___0_____27299));
  nor2s1 _______442758(.DIN1 (________24722), .DIN2 (___000___27177),
       .Q (___0_____27298));
  nor2s1 ______442759(.DIN1 (_____0__24209), .DIN2 (___00____27181), .Q
       (___0__0__27297));
  nor2s1 _______442760(.DIN1 (________22146), .DIN2 (___00____27180),
       .Q (___0__9__27296));
  nor2s1 ______442761(.DIN1 (__9_____26487), .DIN2 (___000___27174), .Q
       (___0_____27295));
  nnd2s1 _______442762(.DIN1 (___0_____27294), .DIN2
       (___________________________________), .Q (___0_____27398));
  xnr2s1 _____442763(.DIN1 (_________32901), .DIN2 (__99____27130), .Q
       (___0_____27348));
  nnd2s1 ______442764(.DIN1 (___00____27185), .DIN2 (__9_____26454), .Q
       (___0_____27396));
  or2s1 _______442765(.DIN1 (___________________________________),
       .DIN2 (___0_____27294), .Q (___0_____27399));
  nnd2s1 ____0_442766(.DIN1 (___00____27219), .DIN2 (__9_____26999), .Q
       (___0_____27391));
  dffacs1 _______________0_(.CLRB (reset), .CLK (clk), .DIN
       (___00_9__27188), .QN
       (______________0______________________18828));
  xor2s1 _____0_442767(.DIN1 (_____________18895), .DIN2
       (___00____27242), .Q (___0_____27419));
  xor2s1 ____442768(.DIN1 (__99____27120), .DIN2 (__9_0___26703), .Q
       (___0__9__27392));
  xor2s1 ____09_442769(.DIN1 (________22873), .DIN2 (___0_00__27267),
       .Q (___0__9__27402));
  dffacs2 _________________(.CLRB (reset), .CLK (clk), .DIN
       (___00____27230), .Q
       (______________________________________0__________0));
  dffacs1 _________________442770(.CLRB (reset), .CLK (clk), .DIN
       (___00____27187), .QN (______________18868));
  nor2s1 ______442771(.DIN1 (________23201), .DIN2 (__99____27156), .Q
       (___0_____27293));
  nor2s1 ____99_442772(.DIN1 (___0_____27291), .DIN2 (__9990), .Q
       (___0_____27292));
  nnd2s1 ____0__442773(.DIN1 (__999_), .DIN2 (___0_____27289), .Q
       (___0_____27290));
  nnd2s1 ____0__442774(.DIN1 (__999___27165), .DIN2 (___0__0__27287),
       .Q (___0_____27288));
  nnd2s1 ____0__442775(.DIN1 (__999___27164), .DIN2 (____9___24057), .Q
       (___0__9__27286));
  nor2s1 ____0__442776(.DIN1 (___0_____27284), .DIN2 (__99____27160),
       .Q (___0_____27285));
  nor2s1 ____0__442777(.DIN1 (___00____27200), .DIN2 (_________34766),
       .Q (___0_____27283));
  nor2s1 ____0__442778(.DIN1 (___0_____27281), .DIN2 (__999___27168),
       .Q (___0_____27282));
  nor2s1 ____0__442779(.DIN1 (___0_____27696), .DIN2 (__99____27158),
       .Q (___0_____27280));
  nor2s1 ____0_442780(.DIN1 (_____0___28805), .DIN2 (__99____27159), .Q
       (___0_____27279));
  nnd2s1 ____0__442781(.DIN1 (___0__0__27277), .DIN2 (___000___27172),
       .Q (___0_____27278));
  or2s1 ______442782(.DIN1 (_________35060), .DIN2 (__99____27127), .Q
       (___0_09__27276));
  nnd2s1 ____09_442783(.DIN1 (__99_9__27133), .DIN2 (__9_____27061), .Q
       (___0_0___27275));
  nor2s1 _____0_442784(.DIN1 (__9_____26437), .DIN2 (__99____27131), .Q
       (___0_0___27274));
  nnd2s1 _____0_442785(.DIN1 (__99____27147), .DIN2 (___0_0___27272),
       .Q (___0_0___27273));
  nor2s1 _____0_442786(.DIN1 (__99____27123), .DIN2 (__9_____26662), .Q
       (___0_0___27271));
  nnd2s1 _____0_442787(.DIN1 (__99____27146), .DIN2 (__9_____27046), .Q
       (___0_0___27270));
  nnd2s1 _______442788(.DIN1 (__99____27149), .DIN2 (________23597), .Q
       (___0_0___27269));
  or2s1 _______442789(.DIN1 (________22788), .DIN2 (___0_00__27267), .Q
       (___0_0___27268));
  nor2s1 ______442790(.DIN1 (__9_____26548), .DIN2 (__99____27142), .Q
       (___0099__27266));
  nor2s1 _______442791(.DIN1 (___099__23527), .DIN2 (__99_9__27153), .Q
       (___009___27265));
  nnd2s1 _______442792(.DIN1 (__99____27152), .DIN2 (_________34906),
       .Q (___009___27264));
  nnd2s1 ____0__442793(.DIN1 (___00_0__27218), .DIN2 (__9_____27000),
       .Q (___0_____27390));
  dffacs1 _______________________442794(.CLRB (reset), .CLK (clk), .DIN
       (__999___27163), .QN (_____________________18639));
  dffacs1 __________________442795(.CLRB (reset), .CLK (clk), .DIN
       (__999___27166), .QN
       (______________________________________0__________0__18892));
  nnd2s1 _____9_442796(.DIN1 (__99____27124), .DIN2 (________22673), .Q
       (___009___27263));
  nnd2s1 _______442797(.DIN1 (__99____27148), .DIN2 (___00___23444), .Q
       (___009___27262));
  nor2s1 _______442798(.DIN1 (________25680), .DIN2 (__99____27137), .Q
       (___009___27261));
  nnd2s1 _______442799(.DIN1 (__99____27135), .DIN2 (__9_____26354), .Q
       (___009___27260));
  nnd2s1 _______442800(.DIN1 (__99_0__27134), .DIN2 (_____0__25790), .Q
       (___009___27259));
  or2s1 _______442801(.DIN1 (___0090__27257), .DIN2 (__99____27122), .Q
       (___009___27258));
  nnd2s1 _______442802(.DIN1 (__99_9__27143), .DIN2 (____09__23091), .Q
       (___00_9__27256));
  or2s1 _______442803(.DIN1 (___0_9___27648), .DIN2 (__99____27151), .Q
       (___00____27255));
  nor2s1 ______442804(.DIN1 (________23943), .DIN2 (___0000__27170), .Q
       (___00____27254));
  nnd2s1 _______442805(.DIN1 (__99_9__27125), .DIN2 (________25907), .Q
       (___00____27253));
  or2s1 _____442806(.DIN1 (___0_____27446), .DIN2 (__99____27145), .Q
       (___00____27252));
  nnd2s1 _____9_442807(.DIN1 (__99____27132), .DIN2 (__9__9__26476), .Q
       (___00____27251));
  or2s1 _______442808(.DIN1 (___0_____27505), .DIN2 (__99____27129), .Q
       (___00____27250));
  nor2s1 _______442809(.DIN1 (___00____27235), .DIN2 (__99____27121),
       .Q (___00____27249));
  or2s1 _______442810(.DIN1 (___00_0__27247), .DIN2 (________21955), .Q
       (___00____27248));
  nor2s1 _______442811(.DIN1 (________26112), .DIN2 (__99_0__27117), .Q
       (___00_9__27246));
  nnd2s1 ______442812(.DIN1 (________22295), .DIN2 (__99____27119), .Q
       (___00____27245));
  nnd2s1 _______442813(.DIN1 (__99____27114), .DIN2 (_________34770),
       .Q (___00____27244));
  nnd2s1 _____0_442814(.DIN1 (__99____27111), .DIN2 (________22912), .Q
       (___00____27243));
  nnd2s1 _______442815(.DIN1 (_________34764), .DIN2
       (______________18870), .Q (_________28457));
  nor2s1 _______442816(.DIN1 (outData[14]), .DIN2 (___00____27242), .Q
       (___0_____27349));
  nnd2s1 _______442817(.DIN1 (___00____27242), .DIN2 (__9_____27050),
       .Q (_________32427));
  dffacs2 _____________________0_442818(.CLRB (reset), .CLK (clk), .DIN
       (__99____27115), .QN (_________________0___18607));
  xor2s1 _____0_442819(.DIN1 (____0____34552), .DIN2 (__9_0___26805),
       .Q (_____00__28898));
  dffacs1 _______________________442820(.CLRB (reset), .CLK (clk), .DIN
       (__99_0__27126), .QN (_____________________18602));
  nor2s1 ____0__442821(.DIN1 (________22424), .DIN2 (__99____27102), .Q
       (___00____27241));
  nor2s1 _______442822(.DIN1 (____9___22892), .DIN2 (__9_9___27075), .Q
       (___00____27240));
  nnd2s1 ____09_442823(.DIN1 (__9900), .DIN2 (________22673), .Q
       (___00____27239));
  nnd2s1 ____09_442824(.DIN1 (__9909), .DIN2 (________24740), .Q
       (___00_0__27238));
  nor2s1 _____442825(.DIN1 (__90_0__26318), .DIN2 (__99____27094), .Q
       (___00_9__27237));
  nor2s1 _____0_442826(.DIN1 (___00____27235), .DIN2 (__99__), .Q
       (___00____27236));
  or2s1 _____0_442827(.DIN1 (___00____27233), .DIN2 (__99____27108), .Q
       (___00____27234));
  nnd2s1 _____442828(.DIN1 (__99____27101), .DIN2 (_____9___28517), .Q
       (___00____27232));
  nnd2s1 ______442829(.DIN1 (__99_0__27097), .DIN2 (___9____24262), .Q
       (___00____27231));
  or2s1 _______442830(.DIN1 (_____9__23684), .DIN2 (__9__0__27064), .Q
       (___00____27230));
  nnd2s1 _______442831(.DIN1 (__9_____27067), .DIN2 (___9____23361), .Q
       (___00____27229));
  nnd2s1 _______442832(.DIN1 (__99_9), .DIN2 (_____9__22884), .Q
       (___00_0__27228));
  nnd2s1 _______442833(.DIN1 (___00____27216), .DIN2 (__9_____26635),
       .Q (___00_9__27227));
  nnd2s1 _______442834(.DIN1 (__99____27096), .DIN2 (___00____27182),
       .Q (___00____27226));
  nnd2s1 _______442835(.DIN1 (__99____27093), .DIN2 (_____90__34918),
       .Q (___00____27225));
  nor2s1 _______442836(.DIN1 (___9____25237), .DIN2 (__9_____27071), .Q
       (___00____27224));
  and2s1 _______442837(.DIN1 (__99____27095), .DIN2 (___00____27222),
       .Q (___00____27223));
  and2s1 _______442838(.DIN1 (__9_90__27074), .DIN2 (___00____27220),
       .Q (___00____27221));
  hi1s1 ______442839(.DIN (___00_0__27218), .Q (___00____27219));
  or2s1 _______442840(.DIN1 (___0__9__27771), .DIN2 (___00____27216),
       .Q (___00_9__27217));
  nnd2s1 _______442841(.DIN1 (__99____27092), .DIN2 (____9___21899), .Q
       (___00____27215));
  and2s1 _______442842(.DIN1 (__990___27087), .DIN2 (___00____27213),
       .Q (___00____27214));
  nnd2s1 _______442843(.DIN1 (__9_9___27079), .DIN2 (___00____27211),
       .Q (___00____27212));
  nor2s1 ______442844(.DIN1 (_____9__24597), .DIN2 (__9_____27058), .Q
       (___00____27210));
  xor2s1 _______442845(.DIN1 (__9_____26971), .DIN2 (_________34362),
       .Q (___00____27209));
  nor2s1 _______442846(.DIN1 (________21758), .DIN2 (__9_9___27077), .Q
       (___00_0__27208));
  nnd2s1 _______442847(.DIN1 (__9_____27072), .DIN2 (__90_0__26271), .Q
       (___00____27207));
  nnd2s1 ______442848(.DIN1 (__9_____27070), .DIN2 (__9_____26927), .Q
       (___00____27206));
  nor2s1 _______442849(.DIN1 (___0__9__27771), .DIN2 (__9_____27056),
       .Q (___00____27205));
  xor2s1 ____0__442850(.DIN1 (__9_____27003), .DIN2 (_________30472),
       .Q (___0_0___27369));
  nnd2s1 _______442851(.DIN1 (__990___27083), .DIN2 (__99____27109), .Q
       (___0_0___27368));
  nnd2s1 _______442852(.DIN1 (__9_9___27076), .DIN2 (__9_____26401), .Q
       (___00____27204));
  nor2s1 _______442853(.DIN1 (___00____27202), .DIN2 (__99_0), .Q
       (___00____27203));
  or2s1 _______442854(.DIN1 (___00____27200), .DIN2 (__990___27089), .Q
       (___00____27201));
  nor2s1 _______442855(.DIN1 (___0__9__27771), .DIN2 (__9_____27059),
       .Q (___00_0__27199));
  nor2s1 _______442856(.DIN1 (__9_____26933), .DIN2 (__9_____27065), .Q
       (___00_9__27198));
  and2s1 ______442857(.DIN1 (__9_____27066), .DIN2 (___00____27196), .Q
       (___00____27197));
  nor2s1 _____9_442858(.DIN1 (________24921), .DIN2 (__9_9___27081), .Q
       (___00____27195));
  nor2s1 _____442859(.DIN1 (___00___19777), .DIN2 (__9_9___27080), .Q
       (___00____27194));
  nor2s1 ______442860(.DIN1 (____9_0__29047), .DIN2 (_____9___30627),
       .Q (___00____27193));
  nnd2s1 _____0_442861(.DIN1 (____9_0__29047), .DIN2 (___00____27191),
       .Q (___00____27192));
  nnd2s1 _______442862(.DIN1 (__9__0__27054), .DIN2 (___0_0___27272),
       .Q (___00____27190));
  nnd2s1 _______442863(.DIN1 (__9__9__27053), .DIN2 (__9_____26717), .Q
       (___00_0__27189));
  nnd2s1 ______442864(.DIN1 (__99_0__27107), .DIN2 (_________32356), .Q
       (___00_9__27188));
  nnd2s1 ______442865(.DIN1 (__9_____27057), .DIN2 (_____9__24533), .Q
       (___00____27187));
  nor2s1 _______442866(.DIN1 (__990___27086), .DIN2 (__99_9__27106), .Q
       (___00____27186));
  nor2s1 _______442867(.DIN1 (________25999), .DIN2 (__99____27105), .Q
       (___00____27185));
  nor2s1 _______442868(.DIN1 (________23206), .DIN2 (__99____27098), .Q
       (___00____27184));
  nnd2s1 _______442869(.DIN1 (__9_____27049), .DIN2 (___00____27182),
       .Q (___00____27183));
  nor2s1 _______442870(.DIN1 (___00____27202), .DIN2 (__99____27090),
       .Q (___00____27181));
  nor2s1 _______442871(.DIN1 (___9____23399), .DIN2 (__99____27103), .Q
       (___00____27180));
  nnd2s1 _______442872(.DIN1 (__9_____27055), .DIN2 (________26059), .Q
       (___00_0__27179));
  nnd2s1 _______442873(.DIN1 (__99____27113), .DIN2 (__9__9__26968), .Q
       (___0009__27178));
  nnd2s1 _______442874(.DIN1 (__9_____27047), .DIN2 (________23773), .Q
       (___000___27177));
  nnd2s1 _______442875(.DIN1 (___000___27171), .DIN2 (__9_____27052),
       .Q (___000___27176));
  nnd2s1 ______442876(.DIN1 (__9__0__27044), .DIN2 (__90____26273), .Q
       (___000___27175));
  nnd2s1 ______442877(.DIN1 (__9_____27048), .DIN2 (__9__9__26540), .Q
       (___000___27174));
  xor2s1 _______442878(.DIN1 (_______________18876), .DIN2
       (_____9___30627), .Q (___0_99__27363));
  xor2s1 _____0_442879(.DIN1 (__9_____26972), .DIN2 (_________35050),
       .Q (___0_____27329));
  and2s1 _______442880(.DIN1 (___000___27173), .DIN2
       (______________18869), .Q (___0_____27294));
  nor2s1 _______442881(.DIN1 (____9_0__29047), .DIN2
       (_______________18873), .Q (___0_____27310));
  xor2s1 _____0_442882(.DIN1 (__9_____26975), .DIN2 (outData[12]), .Q
       (_____9___29527));
  dffacs1 __________________442883(.CLRB (reset), .CLK (clk), .DIN
       (__99____27099), .QN
       (______________________________________0_____________18889));
  nnd2s1 _____9_442884(.DIN1 (___000___27171), .DIN2 (__9_____27012),
       .Q (___000___27172));
  nnd2s1 _______442885(.DIN1 (__9_0___26993), .DIN2 (_____9__22643), .Q
       (___0000__27170));
  and2s1 ____09_442886(.DIN1 (__9_____27017), .DIN2 (___9_9__26226), .Q
       (__999___27169));
  or2s1 _____0_442887(.DIN1 (__999___27167), .DIN2 (__9_____27020), .Q
       (__999___27168));
  nnd2s1 _______442888(.DIN1 (__9_____27028), .DIN2 (___9_9__23385), .Q
       (__999___27166));
  nor2s1 _______442889(.DIN1 (___0_____27291), .DIN2 (__9_____27022),
       .Q (__999___27165));
  nor2s1 _______442890(.DIN1 (___0_9__25356), .DIN2 (__99____27161), .Q
       (__999___27164));
  nnd2s1 _______442891(.DIN1 (__9_____27016), .DIN2 (_____9___28517),
       .Q (__999___27163));
  and2s1 _______442892(.DIN1 (__9__0__27015), .DIN2 (___00____27196),
       .Q (__999_));
  nnd2s1 _______442893(.DIN1 (__9_____27011), .DIN2 (__99____27141), .Q
       (__9990));
  nnd2s1 _______442894(.DIN1 (__99____27161), .DIN2 (___0_____27386),
       .Q (__99_9__27162));
  nnd2s1 ______442895(.DIN1 (__9_____27008), .DIN2 (____0___23805), .Q
       (__99____27160));
  nor2s1 _______442896(.DIN1 (________23911), .DIN2 (__9__9__27024), .Q
       (__99____27159));
  and2s1 _______442897(.DIN1 (__9_____27010), .DIN2 (__99____27157), .Q
       (__99____27158));
  or2s1 _______442898(.DIN1 (____09__23535), .DIN2 (__9_____26976), .Q
       (__99____27156));
  or2s1 _____0_442899(.DIN1 (__99_0__27154), .DIN2 (__9_____27007), .Q
       (__99____27155));
  nnd2s1 _______442900(.DIN1 (__9_9___26983), .DIN2 (___9_0__24276), .Q
       (__99_9__27153));
  nor2s1 _______442901(.DIN1 (____0___24159), .DIN2 (__9_____26970), .Q
       (__99____27152));
  nnd2s1 _____0_442902(.DIN1 (__9_____26998), .DIN2 (__99____27150), .Q
       (__99____27151));
  nor2s1 _____442903(.DIN1 (_____0__23268), .DIN2 (__9_90__26979), .Q
       (__99____27149));
  nor2s1 ______442904(.DIN1 (____09__23983), .DIN2 (__9_9___26980), .Q
       (__99____27148));
  and2s1 _______442905(.DIN1 (__9_____26977), .DIN2 (__9_____26383), .Q
       (__99____27147));
  nor2s1 _______442906(.DIN1 (__9_0___26614), .DIN2 (__9_____27001), .Q
       (__99____27146));
  or2s1 _______442907(.DIN1 (__99_0__27144), .DIN2 (__9_____27030), .Q
       (__99____27145));
  nor2s1 _______442908(.DIN1 (________23281), .DIN2 (__9__9__26978), .Q
       (__99_9__27143));
  nnd2s1 _______442909(.DIN1 (__9_____27039), .DIN2 (__99____27141), .Q
       (__99____27142));
  xor2s1 _____0_442910(.DIN1 (outData[2]), .DIN2 (__9_____26909), .Q
       (___00_0__27218));
  xor2s1 _____0_442911(.DIN1 (__990_), .DIN2 (outData[12]), .Q
       (____9____29964));
  dffacs1 ___________________442912(.CLRB (reset), .CLK (clk), .DIN
       (__9_____27018), .Q (______________0____________________));
  dffacs1 __________________442913(.CLRB (reset), .CLK (clk), .DIN
       (__9_____27026), .QN
       (______________________________________0_____________18885));
  nor2s1 _______442914(.DIN1 (__99____27139), .DIN2 (__99____27138), .Q
       (__99____27140));
  nnd2s1 _______442915(.DIN1 (__9_____27036), .DIN2 (____09__24524), .Q
       (__99____27137));
  nor2s1 _______442916(.DIN1 (__9_0___26335), .DIN2 (__9__0__26996), .Q
       (__99____27136));
  nor2s1 _______442917(.DIN1 (________24845), .DIN2 (__9_____27004), .Q
       (__99____27135));
  nor2s1 ______442918(.DIN1 (__9_____26472), .DIN2 (__9_____26997), .Q
       (__99_0__27134));
  nnd2s1 _______442919(.DIN1 (__9_____27033), .DIN2 (__9__0__26739), .Q
       (__99_9__27133));
  nor2s1 ______442920(.DIN1 (________23552), .DIN2 (__9_____27042), .Q
       (__99____27132));
  nor2s1 _______442921(.DIN1 (__9_____26953), .DIN2 (__9_____26973), .Q
       (__99____27131));
  nnd2s1 _______442922(.DIN1 (_________33835), .DIN2
       (_______________18876), .Q (__99____27130));
  or2s1 _______442923(.DIN1 (__99____27128), .DIN2 (__9_____27032), .Q
       (__99____27129));
  nnd2s1 ______442924(.DIN1 (______0__34768), .DIN2 (__90____26306), .Q
       (__99____27127));
  nnd2s1 _______442925(.DIN1 (__9_99__26988), .DIN2 (___0_____27485),
       .Q (__99_0__27126));
  nor2s1 _____9_442926(.DIN1 (__9_9___26984), .DIN2 (__9_____26914), .Q
       (__99_9__27125));
  nnd2s1 _______442927(.DIN1 (__9__9__27034), .DIN2 (________24195), .Q
       (__99____27124));
  nor2s1 _______442928(.DIN1 (________21758), .DIN2 (__9_9___26981), .Q
       (__99____27123));
  nnd2s1 _______442929(.DIN1 (__9_____27038), .DIN2 (________25672), .Q
       (__99____27122));
  nnd2s1 _______442930(.DIN1 (__9_____26963), .DIN2 (__9_____26759), .Q
       (__99____27121));
  xor2s1 _______442931(.DIN1 (__99____27104), .DIN2 (_________32901),
       .Q (__99____27120));
  nnd2s1 _______442932(.DIN1 (__99____27118), .DIN2
       (_______________18876), .Q (__99____27119));
  nor2s1 _____9_442933(.DIN1 (__99_9__27116), .DIN2 (__9_____26965), .Q
       (__99_0__27117));
  nnd2s1 ______442934(.DIN1 (__9__0__26961), .DIN2 (________23954), .Q
       (__99____27115));
  hi1s1 _______442935(.DIN (__99____27113), .Q (__99____27114));
  nor2s1 _______442936(.DIN1 (_______________18876), .DIN2
       (______________________________________0_____________18888), .Q
       (__99____27112));
  and2s1 _______442937(.DIN1 (__9__9__26960), .DIN2 (__99____27110), .Q
       (__99____27111));
  nnd2s1 _______442938(.DIN1 (_____90__31526), .DIN2 (__9_____27051),
       .Q (___0__0__27277));
  nor2s1 _______442939(.DIN1 (_______________18876), .DIN2
       (______9__28578), .Q (___0_____27309));
  nor2s1 ______442940(.DIN1 (__9_____26820), .DIN2 (__9_9___26982), .Q
       (___0_00__27267));
  nor2s1 _______442941(.DIN1 (_______________18876), .DIN2
       (_________33835), .Q (___0_____27416));
  nnd2s1 _____0_442942(.DIN1 (_______________18876), .DIN2
       (_________9___0_), .Q (___00_0__27247));
  nnd2s1 _______442943(.DIN1 (__9_____26967), .DIN2 (__99____27109), .Q
       (___00____27242));
  nor2s1 _______442944(.DIN1 (__9_____26974), .DIN2 (__9_0___26990), .Q
       (_________29457));
  nnd2s1 ______442945(.DIN1 (__9_____26957), .DIN2 (____90__25645), .Q
       (__99____27108));
  nor2s1 _______442946(.DIN1 (___9_0__24257), .DIN2 (__9_____26880), .Q
       (__99_0__27107));
  nnd2s1 ______442947(.DIN1 (__9_9___26889), .DIN2 (____9___22893), .Q
       (__99_9__27106));
  and2s1 _______442948(.DIN1 (__99____27104), .DIN2 (________26003), .Q
       (__99____27105));
  nnd2s1 _______442949(.DIN1 (__9_0___26898), .DIN2 (__9_9___26604), .Q
       (__99____27103));
  nnd2s1 ______442950(.DIN1 (__9_____26947), .DIN2 (___0__0__27609), .Q
       (__99____27102));
  and2s1 _______442951(.DIN1 (__9_____26944), .DIN2 (__99____27100), .Q
       (__99____27101));
  nnd2s1 _______442952(.DIN1 (__9__0__27025), .DIN2 (__9__9__26950), .Q
       (__99____27099));
  nnd2s1 _______442953(.DIN1 (__9_____26954), .DIN2 (__9_____26723), .Q
       (__99____27098));
  nnd2s1 _______442954(.DIN1 (__9_99__26891), .DIN2 (________22673), .Q
       (__99_0__27097));
  nor2s1 ______442955(.DIN1 (________22146), .DIN2 (__9_____26952), .Q
       (__99_9));
  nor2s1 _______442956(.DIN1 (__9__9__26921), .DIN2 (__9_____26938), .Q
       (__99____27096));
  and2s1 ______442957(.DIN1 (__9_____26904), .DIN2 (________24854), .Q
       (__99____27095));
  nnd2s1 ______442958(.DIN1 (__9_____26948), .DIN2 (___0____22610), .Q
       (__99____27094));
  and2s1 _______442959(.DIN1 (__9_____26906), .DIN2 (__9_____26840), .Q
       (__99____27093));
  nnd2s1 _______442960(.DIN1 (__9_____26946), .DIN2 (__99____27091), .Q
       (__99____27092));
  nor2s1 _______442961(.DIN1 (__9_____26572), .DIN2 (__9_0___26895), .Q
       (__99____27090));
  or2s1 _______442962(.DIN1 (________24753), .DIN2 (__9__0__26951), .Q
       (__99__));
  nor2s1 _______442963(.DIN1 (________23248), .DIN2 (__9_____26932), .Q
       (__99_0));
  nor2s1 _______442964(.DIN1 (________24919), .DIN2 (__9_____26945), .Q
       (__9909));
  or2s1 _____9_442965(.DIN1 (__990___27088), .DIN2 (__9__9__26930), .Q
       (__990___27089));
  nor2s1 _____442966(.DIN1 (__990___27086), .DIN2 (__9_____26925), .Q
       (__990___27087));
  nor2s1 _______442967(.DIN1 (__990___27084), .DIN2 (__9_____26929), .Q
       (__990___27085));
  nor2s1 _______442968(.DIN1 (outData[12]), .DIN2 (__990_), .Q
       (__990___27083));
  nnd2s1 _______442969(.DIN1 (__9_____26928), .DIN2 (________24557), .Q
       (__9900));
  nnd2s1 ______442970(.DIN1 (__9_____27068), .DIN2 (___00____27211), .Q
       (__9_99__27082));
  nnd2s1 _______442971(.DIN1 (__9_____26949), .DIN2 (_________34900),
       .Q (__9_9___27081));
  and2s1 _______442972(.DIN1 (__990_), .DIN2 (outData[13]), .Q
       (__9_9___27080));
  nnd2s1 _______442973(.DIN1 (__9_____26956), .DIN2 (__9_____26779), .Q
       (__9_9___27079));
  nor2s1 _______442974(.DIN1 (___0_9__22581), .DIN2 (__9_0___26992), .Q
       (__9_9___27078));
  nor2s1 ______442975(.DIN1 (________22146), .DIN2 (__9_____26910), .Q
       (__9_9___27077));
  nor2s1 _______442976(.DIN1 (__9_____26381), .DIN2 (__9_____26955), .Q
       (___00____27216));
  nnd2s1 _______442977(.DIN1 (__990_), .DIN2 (__9_____26666), .Q
       (_________28476));
  nor2s1 _______442978(.DIN1 (________25722), .DIN2 (__9_90__26883), .Q
       (__9_9___27076));
  nor2s1 _____9_442979(.DIN1 (________21758), .DIN2 (__9__0__26922), .Q
       (__9_9___27075));
  nor2s1 _____9_442980(.DIN1 (__9__9__27073), .DIN2 (__9__0__26941), .Q
       (__9_90__27074));
  nor2s1 _____9_442981(.DIN1 (________25064), .DIN2 (__9__0__26931), .Q
       (__9_____27072));
  nnd2s1 _____442982(.DIN1 (__9_____26926), .DIN2 (________22910), .Q
       (__9_____27071));
  nnd2s1 _____442983(.DIN1 (__9_____26939), .DIN2 (_____9___28891), .Q
       (__9_____27070));
  nor2s1 _____0_442984(.DIN1 (__9_____27068), .DIN2 (__9_____27062), .Q
       (__9_____27069));
  nnd2s1 _____0_442985(.DIN1 (__9_____26915), .DIN2 (__9_____27027), .Q
       (__9_____27067));
  nor2s1 _____0_442986(.DIN1 (________25739), .DIN2 (__9_____26920), .Q
       (__9_____27066));
  nor2s1 _____0_442987(.DIN1 (_____0___28805), .DIN2 (__9_____26936),
       .Q (__9_____27065));
  nor2s1 _______442988(.DIN1 (________23683), .DIN2 (__9__9__26940), .Q
       (__9__0__27064));
  nnd2s1 _______442989(.DIN1 (__9_____27062), .DIN2 (__9_____27061), .Q
       (__9__9__27063));
  nor2s1 _______442990(.DIN1 (___0_0__24352), .DIN2 (__9_____26924), .Q
       (__9_____27060));
  nor2s1 _______442991(.DIN1 (___0_____27696), .DIN2 (__9_____26919),
       .Q (__9_____27059));
  nnd2s1 ______442992(.DIN1 (__9_____26916), .DIN2 (________24439), .Q
       (__9_____27058));
  nnd2s1 ______442993(.DIN1 (____9___24784), .DIN2 (__9_0___26899), .Q
       (__9_____27057));
  nor2s1 _____9_442994(.DIN1 (___00____27200), .DIN2 (__9_____26923),
       .Q (__9_____27056));
  nor2s1 _____9_442995(.DIN1 (________25881), .DIN2 (__9_0___26894), .Q
       (__9_____27055));
  nor2s1 _____9_442996(.DIN1 (__9_0___26709), .DIN2 (__9_9___26887), .Q
       (__9__0__27054));
  nor2s1 _______442997(.DIN1 (__9_0___26422), .DIN2 (__9_0___26900), .Q
       (__9__9__27053));
  hi1s1 ______442998(.DIN (__9_____27051), .Q (__9_____27052));
  nnd2s1 _______442999(.DIN1 (__9_____26966), .DIN2 (outData[13]), .Q
       (__9_____27050));
  nor2s1 _______443000(.DIN1 (__9_____26553), .DIN2 (__9_0___26893), .Q
       (__9_____27049));
  nor2s1 ______443001(.DIN1 (________26125), .DIN2 (__9_____26903), .Q
       (__9_____27048));
  nor2s1 _______443002(.DIN1 (____9___24884), .DIN2 (__9_0___26896), .Q
       (__9_____27047));
  nnd2s1 _______443003(.DIN1 (__9_09__26901), .DIN2 (__9_____27045), .Q
       (__9_____27046));
  and2s1 _______443004(.DIN1 (__9_9___26886), .DIN2 (__9__9__27043), .Q
       (__9__0__27044));
  nor2s1 _____0_443005(.DIN1 (__9_0___26801), .DIN2 (__99____27104), .Q
       (___000___27173));
  nnd2s1 _______443006(.DIN1 (__9__0__26902), .DIN2
       (______________18870), .Q (__99____27113));
  dffacs1 ___________________443007(.CLRB (reset), .CLK (clk), .DIN
       (__9_00__26892), .Q (______________0___________________));
  hi1s1 _____9_443008(.DIN (_______________18876), .Q (____9_0__29047));
  dffacs1 ________________________443009(.CLRB (reset), .CLK (clk),
       .DIN (__9_____26943), .QN (______________________18631));
  nnd2s1 _______443010(.DIN1 (__9_____26845), .DIN2 (__9_____27041), .Q
       (__9_____27042));
  or2s1 _______443011(.DIN1 (_____0___28805), .DIN2 (__9__0__26969), .Q
       (__9_____27040));
  nor2s1 _______443012(.DIN1 (___0____21669), .DIN2 (__9_____26830), .Q
       (__9_____27039));
  nor2s1 ______443013(.DIN1 (__9_____27037), .DIN2 (__9_____26839), .Q
       (__9_____27038));
  nor2s1 _______443014(.DIN1 (__9__0__27035), .DIN2 (__9_____26813), .Q
       (__9_____27036));
  nor2s1 _______443015(.DIN1 (_____0__25156), .DIN2 (__9_____26836), .Q
       (__9__9__27034));
  nor2s1 _______443016(.DIN1 (__9_____26583), .DIN2 (__9_____26832), .Q
       (__9_____27033));
  nnd2s1 _______443017(.DIN1 (__9_____27031), .DIN2 (____9___25646), .Q
       (__9_____27032));
  or2s1 _______443018(.DIN1 (____0___23264), .DIN2 (__9_____26823), .Q
       (__9_____27030));
  xor2s1 _____9_443019(.DIN1 (__9_99__26797), .DIN2 (_________31290),
       .Q (__9_____27029));
  nnd2s1 _______443020(.DIN1 (__9_____26827), .DIN2 (__9_____27027), .Q
       (__9_____27028));
  nnd2s1 _______443021(.DIN1 (__9__0__27025), .DIN2 (__9_____26865), .Q
       (__9_____27026));
  or2s1 _______443022(.DIN1 (__9_____27023), .DIN2 (__9__0__26873), .Q
       (__9__9__27024));
  nnd2s1 _______443023(.DIN1 (__9_____26874), .DIN2 (__9_____27021), .Q
       (__9_____27022));
  nnd2s1 _______443024(.DIN1 (__9_____26866), .DIN2 (__9_____27019), .Q
       (__9_____27020));
  or2s1 _______443025(.DIN1 (_________31949), .DIN2 (__9_____26867), .Q
       (__9_____27018));
  nnd2s1 _______443026(.DIN1 (__9__9__26863), .DIN2 (__9_____27061), .Q
       (__9_____27017));
  nor2s1 _______443027(.DIN1 (_____9__25789), .DIN2 (__9_____26859), .Q
       (__9_____27016));
  and2s1 _______443028(.DIN1 (__9_____26876), .DIN2 (__9__9__27014), .Q
       (__9__0__27015));
  nnd2s1 _______443029(.DIN1 (__9_____26851), .DIN2 (________25629), .Q
       (__9_____27013));
  xor2s1 _____9_443030(.DIN1
       (______________________________________0__________0__18892),
       .DIN2 (_______________18875), .Q (__9_____27012));
  nor2s1 _____9_443031(.DIN1 (______0__28751), .DIN2 (__9_____26857),
       .Q (__9_____27011));
  nor2s1 _____0_443032(.DIN1 (__9_0___26521), .DIN2 (__9_____26858), .Q
       (__9_____27010));
  xor2s1 _____0_443033(.DIN1 (__9__0__26729), .DIN2 (____9___19200), .Q
       (__9_____27009));
  nor2s1 _____0_443034(.DIN1 (___0____23485), .DIN2 (__9_____26856), .Q
       (__9_____27008));
  nnd2s1 _____443035(.DIN1 (__9_____27002), .DIN2 (___99___24328), .Q
       (__9_____27007));
  nnd2s1 _______443036(.DIN1 (__9_____26855), .DIN2 (__9__0__27005), .Q
       (__9_____27006));
  nnd2s1 _______443037(.DIN1 (__9_____26849), .DIN2 (________23003), .Q
       (__9_____27004));
  nnd2s1 _______443038(.DIN1 (__9_____27002), .DIN2 (_____0__25820), .Q
       (__9_____27003));
  nor2s1 _______443039(.DIN1 (___0_____27696), .DIN2 (__9__0__26844),
       .Q (__9_____27001));
  hi1s1 _______443040(.DIN (__9_____26999), .Q (__9_____27000));
  nor2s1 _______443041(.DIN1 (_____9__22280), .DIN2 (__9_____26837), .Q
       (__9_____26998));
  nnd2s1 _______443042(.DIN1 (__9_____26860), .DIN2 (__9_____27021), .Q
       (__99____27161));
  nor2s1 _______443043(.DIN1 (__9_____26908), .DIN2 (__9_____26869), .Q
       (___0_____27739));
  nnd2s1 _______443044(.DIN1 (__9__9__26853), .DIN2 (________25864), .Q
       (__9_____26997));
  and2s1 _______443045(.DIN1 (__9_09__26995), .DIN2 (__9_____26576), .Q
       (__9__0__26996));
  and2s1 _______443046(.DIN1 (__9_____26841), .DIN2 (__9_____27061), .Q
       (__9_0___26994));
  nor2s1 ______443047(.DIN1 (________23225), .DIN2 (__9_____26842), .Q
       (__9_0___26993));
  xor2s1 _______443048(.DIN1 (__9_____26716), .DIN2 (__9_00__26989), .Q
       (__9_0___26990));
  and2s1 _______443049(.DIN1 (__9_____26822), .DIN2 (__9_9___26987), .Q
       (__9_99__26988));
  nor2s1 _______443050(.DIN1 (__990___27084), .DIN2 (__9_9___26985), .Q
       (__9_9___26986));
  nor2s1 _______443051(.DIN1 (___0__9__27771), .DIN2 (__9_____26818),
       .Q (__9_9___26984));
  nor2s1 _______443052(.DIN1 (________22701), .DIN2 (__9_____26847), .Q
       (__9_9___26983));
  nor2s1 _______443053(.DIN1 (_________30166), .DIN2 (__9_____26814),
       .Q (__9_9___26982));
  nor2s1 _______443054(.DIN1 (________22146), .DIN2 (__9_____26819), .Q
       (__9_9___26981));
  nnd2s1 ______443055(.DIN1 (__9_____26821), .DIN2 (______0__35048), .Q
       (__9_9___26980));
  nnd2s1 _______443056(.DIN1 (__9_____26817), .DIN2 (________24012), .Q
       (__9_90__26979));
  nor2s1 _______443057(.DIN1 (________21758), .DIN2 (__9_____26829), .Q
       (__9__9__26978));
  nor2s1 _______443058(.DIN1 (________25667), .DIN2 (__9__9__26815), .Q
       (__9_____26977));
  nnd2s1 _______443059(.DIN1 (__9_____26848), .DIN2 (___9____25195), .Q
       (__9_____26976));
  xor2s1 ______443060(.DIN1 (______9__32620), .DIN2 (__9_____26974), .Q
       (__9_____26975));
  nor2s1 _______443061(.DIN1 (________21758), .DIN2 (__9__9__26872), .Q
       (__9_____26973));
  nor2s1 _______443062(.DIN1 (__9_0___26806), .DIN2 (__9_9___26890), .Q
       (__9_____26972));
  nor2s1 ______443063(.DIN1 (__9_____26958), .DIN2 (_________28549), .Q
       (__9_____26971));
  nnd2s1 _______443064(.DIN1 (__9__0__26969), .DIN2 (________26103), .Q
       (__9_____26970));
  hi1s1 ______443065(.DIN (_________34770), .Q (__9__9__26968));
  hi1s1 _____443066(.DIN (__9_____26966), .Q (__9_____26967));
  nor2s1 _____0_443067(.DIN1 (__9_____26964), .DIN2 (__9_0___26803), .Q
       (__9_____26965));
  nnd2s1 _______443068(.DIN1 (__9__9__26824), .DIN2 (__9_____26962), .Q
       (__9_____26963));
  nor2s1 _______443069(.DIN1 (________22878), .DIN2 (__9_0___26802), .Q
       (__9__0__26961));
  nor2s1 _____0_443070(.DIN1 (__9_____26959), .DIN2 (__9_____26811), .Q
       (__9__9__26960));
  nor2s1 _______443071(.DIN1 (_____0___30458), .DIN2 (____09___30086),
       .Q (__99____27139));
  nor2s1 _______443072(.DIN1 (_________29585), .DIN2 (____09___30086),
       .Q (__9_____27051));
  nnd2s1 _______443073(.DIN1 (_________28549), .DIN2 (__9_____26958),
       .Q (___0_____27496));
  dffacs2 __________________443074(.CLRB (reset), .CLK (clk), .DIN
       (__9_0___26804), .Q (_______________18876));
  nor2s1 ______443075(.DIN1 (____9___24975), .DIN2 (__9_9___26793), .Q
       (__9_____26957));
  nor2s1 _______443076(.DIN1 (________25478), .DIN2 (__9_0___26799), .Q
       (__9_____26956));
  nnd2s1 _______443077(.DIN1 (__9__9__26787), .DIN2 (__9_00__26419), .Q
       (__9_____26955));
  nor2s1 _______443078(.DIN1 (__9_____26953), .DIN2 (__9_9___26792), .Q
       (__9_____26954));
  nnd2s1 _______443079(.DIN1 (__9_9___26789), .DIN2 (__9_____26937), .Q
       (__9_____26952));
  nnd2s1 ______443080(.DIN1 (__9_____26776), .DIN2 (_____9__25769), .Q
       (__9__0__26951));
  nor2s1 _______443081(.DIN1 (________23681), .DIN2 (__9_____26770), .Q
       (__9__9__26950));
  nnd2s1 _______443082(.DIN1 (__9_9___26790), .DIN2 (___99___23429), .Q
       (__9_____26949));
  nor2s1 ______443083(.DIN1 (__9_____26754), .DIN2 (__9_____26772), .Q
       (__9_____26948));
  nor2s1 ______443084(.DIN1 (________24205), .DIN2 (__9_____26774), .Q
       (__9_____26947));
  nor2s1 _______443085(.DIN1 (___00____27200), .DIN2 (__9_____26780),
       .Q (__9_____26946));
  nnd2s1 _______443086(.DIN1 (__9_____26742), .DIN2 (________24751), .Q
       (__9_____26945));
  nor2s1 ______443087(.DIN1 (________22637), .DIN2 (__9_____26783), .Q
       (__9_____26944));
  nnd2s1 _____443088(.DIN1 (__9_____26771), .DIN2 (__9__0__26467), .Q
       (__9_____26943));
  nnd2s1 _____9_443089(.DIN1 (__9_90__26788), .DIN2 (_____9___28891),
       .Q (__9_____26942));
  nnd2s1 _____9_443090(.DIN1 (__9__0__26768), .DIN2 (__9__0__26494), .Q
       (__9__0__26941));
  nor2s1 _____443091(.DIN1 (_____0___31003), .DIN2 (__9_9___26794), .Q
       (__9__9__26940));
  nnd2s1 _____443092(.DIN1 (__9_____26766), .DIN2 (__9_____27021), .Q
       (__9_____26939));
  nnd2s1 _____0_443093(.DIN1 (__9_____26756), .DIN2 (__9_____26937), .Q
       (__9_____26938));
  nor2s1 _______443094(.DIN1 (__9_____26935), .DIN2 (__9_____26737), .Q
       (__9_____26936));
  nnd2s1 _______443095(.DIN1 (__99____27118), .DIN2
       (_______________18875), .Q (__9_____26934));
  nnd2s1 _______443096(.DIN1 (__9_____26760), .DIN2 (________25575), .Q
       (__9_____26933));
  nnd2s1 ______443097(.DIN1 (__9_____26775), .DIN2 (_____0__24588), .Q
       (__9_____26932));
  nnd2s1 _______443098(.DIN1 (__9__0__26778), .DIN2 (________25044), .Q
       (__9__0__26931));
  nnd2s1 _______443099(.DIN1 (__9_____26755), .DIN2 (___9____23398), .Q
       (__9__9__26930));
  nor2s1 _______443100(.DIN1 (___0_____27430), .DIN2 (__9_____26752),
       .Q (__9_____26929));
  nor2s1 _______443101(.DIN1 (__9_____26764), .DIN2 (__9_____26745), .Q
       (__9_____26928));
  nnd2s1 ______443102(.DIN1 (__9__0__26720), .DIN2 (___0_____27386), .Q
       (__9_____26927));
  nnd2s1 _______443103(.DIN1 (__9_____26751), .DIN2 (________21469), .Q
       (__9_____26926));
  nnd2s1 _______443104(.DIN1 (__9_9___26795), .DIN2 (________23819), .Q
       (__9_____26925));
  nnd2s1 _______443105(.DIN1 (_________34774), .DIN2 (_____9__22416),
       .Q (__9_____26924));
  nnd2s1 _______443106(.DIN1 (__9__0__26758), .DIN2 (__9_____26862), .Q
       (__9_____26923));
  nor2s1 _______443107(.DIN1 (__9__9__26921), .DIN2 (__9_____26741), .Q
       (__9__0__26922));
  nnd2s1 _______443108(.DIN1 (__9_____26786), .DIN2 (________26121), .Q
       (__9_____26920));
  nnd2s1 _______443109(.DIN1 (__9__9__26767), .DIN2 (__9_____26917), .Q
       (__9_____26919));
  nor2s1 _______443110(.DIN1 (_______________18875), .DIN2
       (________21243), .Q (__9_____26918));
  nnd2s1 _____0_443111(.DIN1 (__9_____26750), .DIN2 (__9_____26917), .Q
       (__9_____27068));
  nnd2s1 _____0_443112(.DIN1 (__9_9___26796), .DIN2 (________24488), .Q
       (__9_____26999));
  nor2s1 _______443113(.DIN1 (___0_____27698), .DIN2 (__9_____26735),
       .Q (__9_____26916));
  nnd2s1 _______443114(.DIN1 (__9_____26677), .DIN2
       (_______________18875), .Q (__9_____26915));
  nor2s1 _______443115(.DIN1 (___0_9__22581), .DIN2 (__9_____26744), .Q
       (__9_____26914));
  nnd2s1 _______443116(.DIN1 (__9_____26769), .DIN2 (____9___21899), .Q
       (__9_____26913));
  nnd2s1 _______443117(.DIN1 (__9_____26762), .DIN2 (__9__9__26911), .Q
       (__9__0__26912));
  nnd2s1 _______443118(.DIN1 (__9_____26785), .DIN2 (__9_____26828), .Q
       (__9_____26910));
  or2s1 ______443119(.DIN1 (__9_____26868), .DIN2 (__9_____26908), .Q
       (__9_____26909));
  nnd2s1 _______443120(.DIN1 (__9__9__26777), .DIN2 (___0_____27690),
       .Q (__9_____26907));
  nor2s1 _______443121(.DIN1 (__9_____26905), .DIN2 (__9_____26781), .Q
       (__9_____26906));
  nor2s1 ______443122(.DIN1 (____00__22626), .DIN2 (__9_____26782), .Q
       (__9_____26904));
  nnd2s1 _____9_443123(.DIN1 (__9_0___26705), .DIN2 (________25817), .Q
       (__9_____26903));
  nnd2s1 _____9_443124(.DIN1 (__9_09__26807), .DIN2 (___0_____27914),
       .Q (__9__0__26902));
  nnd2s1 _____443125(.DIN1 (__9_____26718), .DIN2 (________24651), .Q
       (__9_09__26901));
  nnd2s1 _____0_443126(.DIN1 (__9_____26725), .DIN2 (__9_0___26424), .Q
       (__9_0___26900));
  nnd2s1 _____0_443127(.DIN1 (__9_0___26704), .DIN2 (__9__0__26532), .Q
       (__9_0___26899));
  nor2s1 _____0_443128(.DIN1 (__9_0___26897), .DIN2 (__9_____26714), .Q
       (__9_0___26898));
  nnd2s1 ______443129(.DIN1 (__9_9___26884), .DIN2 (___0____24407), .Q
       (__9_0___26896));
  nnd2s1 _______443130(.DIN1 (__9_____26721), .DIN2 (________25399), .Q
       (__9_0___26895));
  nnd2s1 _______443131(.DIN1 (__9__0__26712), .DIN2 (___0____24386), .Q
       (__9_0___26894));
  nnd2s1 _______443132(.DIN1 (__9__9__26719), .DIN2 (__900_), .Q
       (__9_0___26893));
  or2s1 _____0_443133(.DIN1 (____9____30867), .DIN2 (__9_____26726), .Q
       (__9_00__26892));
  nnd2s1 _______443134(.DIN1 (__9_____26765), .DIN2 (____99__25750), .Q
       (__9_99__26891));
  nor2s1 _______443135(.DIN1 (__9_9___26888), .DIN2 (__9_09__26711), .Q
       (__9_9___26889));
  and2s1 _______443136(.DIN1 (__9_0___26708), .DIN2 (__9_____27045), .Q
       (__9_9___26887));
  nor2s1 _______443137(.DIN1 (_____0__22962), .DIN2 (__9_0___26710), .Q
       (__9_9___26886));
  or2s1 _____9_443138(.DIN1 (_____0___28805), .DIN2 (__9_9___26884), .Q
       (__9_9___26885));
  nnd2s1 _____0_443139(.DIN1 (__9__9__26748), .DIN2 (_________28602),
       .Q (__9_90__26883));
  nnd2s1 _______443140(.DIN1 (__9_____26881), .DIN2 (__9_____27061), .Q
       (__9__9__26882));
  nor2s1 ______443141(.DIN1 (__9_0___26706), .DIN2 (_________32344), .Q
       (__9_____26880));
  nnd2s1 _______443142(.DIN1 (__9_____26879), .DIN2 (__9_____26878), .Q
       (__9_0___26991));
  nnd2s1 _______443143(.DIN1 (__9_____26974), .DIN2
       (_____________18894), .Q (__9_____26966));
  nnd2s1 ______443144(.DIN1 (__9_____26740), .DIN2 (__9_____26877), .Q
       (__9_____27062));
  nor2s1 _______443145(.DIN1 (___0_____27696), .DIN2 (__9_____26747),
       .Q (__9_0___26992));
  nor2s1 _______443146(.DIN1 (_______________18875), .DIN2
       (_________34409), .Q (__99____27138));
  xnr2s1 ______443147(.DIN1 (__9_____26809), .DIN2 (____99___31805), .Q
       (__99____27104));
  xor2s1 ______443148(.DIN1 (__9__9__26644), .DIN2 (_________31478), .Q
       (__990_));
  and2s1 ______443149(.DIN1 (__9__0__26683), .DIN2 (__9_____26875), .Q
       (__9_____26876));
  nor2s1 _______443150(.DIN1 (____0___25853), .DIN2 (__9_9___26699), .Q
       (__9_____26874));
  or2s1 _______443151(.DIN1 (__9_____26736), .DIN2 (__9_____26689), .Q
       (__9__0__26873));
  nnd2s1 _______443152(.DIN1 (_________34776), .DIN2 (__9_____26871),
       .Q (__9__9__26872));
  nor2s1 ______443153(.DIN1 (___9____25186), .DIN2 (__9_____26850), .Q
       (__9_____26870));
  nor2s1 _______443154(.DIN1 (___9____24300), .DIN2 (__9_____26868), .Q
       (__9_____26869));
  nnd2s1 _______443155(.DIN1 (__9__0__26674), .DIN2 (___9____24283), .Q
       (__9_____26867));
  nor2s1 _____9_443156(.DIN1 (_________34810), .DIN2 (__9_9___26693),
       .Q (__9_____26866));
  nor2s1 _____9_443157(.DIN1 (___9____23370), .DIN2 (__9_____26676), .Q
       (__9_____26865));
  nor2s1 _______443158(.DIN1 (_____9__21884), .DIN2 (__9_9___26696), .Q
       (__9__0__26864));
  nnd2s1 ______443159(.DIN1 (__9_____26687), .DIN2 (__9_____26862), .Q
       (__9__9__26863));
  and2s1 _______443160(.DIN1 (__9__9__26833), .DIN2 (__9__0__27005), .Q
       (__9_____26861));
  nor2s1 _______443161(.DIN1 (_____0__25967), .DIN2 (__9_____26685), .Q
       (__9_____26860));
  nnd2s1 _______443162(.DIN1 (__9_____26680), .DIN2 (__9__0__26439), .Q
       (__9_____26859));
  nnd2s1 ______443163(.DIN1 (__9__9__26682), .DIN2 (_____9__25928), .Q
       (__9_____26858));
  nnd2s1 _______443164(.DIN1 (__9_9___26697), .DIN2 (________26099), .Q
       (__9_____26857));
  nnd2s1 _______443165(.DIN1 (__9_____26688), .DIN2 (___0_9__23517), .Q
       (__9_____26856));
  nnd2s1 ______443166(.DIN1 (__9_____26684), .DIN2 (__9__0__26854), .Q
       (__9_____26855));
  nor2s1 _______443167(.DIN1 (__9_____26440), .DIN2 (__9_____26651), .Q
       (__9__9__26853));
  nnd2s1 _______443168(.DIN1 (__9_____26679), .DIN2 (___0____23469), .Q
       (__9_____26852));
  nnd2s1 _______443169(.DIN1 (__9_____26850), .DIN2 (__9_____27045), .Q
       (__9_____26851));
  and2s1 _______443170(.DIN1 (__9_____26652), .DIN2 (________24682), .Q
       (__9_____26849));
  nor2s1 _______443171(.DIN1 (___90___23347), .DIN2 (__9__9__26653), .Q
       (__9_____26848));
  nnd2s1 _____9_443172(.DIN1 (__9_____26638), .DIN2 (__9_____26846), .Q
       (__9_____26847));
  nor2s1 _____9_443173(.DIN1 (________25801), .DIN2 (__9_____26646), .Q
       (__9_____26845));
  nor2s1 _____443174(.DIN1 (________26130), .DIN2 (__9_____26661), .Q
       (__9__0__26844));
  nnd2s1 _____0_443175(.DIN1 (__9_____26658), .DIN2 (_____9__21800), .Q
       (__9__9__26843));
  nnd2s1 ______443176(.DIN1 (__9_____26667), .DIN2 (__9_9___26791), .Q
       (__9_____26842));
  nnd2s1 _______443177(.DIN1 (__9__0__26645), .DIN2 (__9_____26840), .Q
       (__9_____26841));
  or2s1 _______443178(.DIN1 (__9_____26838), .DIN2 (__9_____26634), .Q
       (__9_____26839));
  nnd2s1 _______443179(.DIN1 (__9_____26672), .DIN2 (______0__34968),
       .Q (__9_____26837));
  or2s1 _______443180(.DIN1 (____0___23622), .DIN2 (__9__9__26627), .Q
       (__9_____26836));
  xor2s1 _______443181(.DIN1 (________24547), .DIN2 (__9_____26835), .Q
       (__9_____27002));
  dffacs1 ________________0_443182(.CLRB (reset), .CLK (clk), .DIN
       (__9__9__26673), .QN (___________0___18877));
  hi1s1 _____9_443183(.DIN (_______________18875), .Q (____09___30086));
  dffacs1 _______________________443184(.CLRB (reset), .CLK (clk), .DIN
       (__9_9___26694), .QN (_____________________18599));
  nor2s1 ______443185(.DIN1 (________26072), .DIN2 (__9__9__26833), .Q
       (__9__0__26834));
  or2s1 _______443186(.DIN1 (__9_____26831), .DIN2 (__9_____26665), .Q
       (__9_____26832));
  nnd2s1 _______443187(.DIN1 (__9_____26630), .DIN2 (_________34982),
       .Q (__9_____26830));
  and2s1 _______443188(.DIN1 (__9_____26656), .DIN2 (__9_____26828), .Q
       (__9_____26829));
  nnd2s1 _______443189(.DIN1 (__9_____26678), .DIN2 (inData[18]), .Q
       (__9_____26827));
  xor2s1 _____443190(.DIN1 (__9_____26547), .DIN2 (____0____30965), .Q
       (__9_____26826));
  nor2s1 _______443191(.DIN1 (__9_0___26615), .DIN2 (__9_____26730), .Q
       (__9__0__26825));
  nnd2s1 _______443192(.DIN1 (__9_0___26609), .DIN2 (________25035), .Q
       (__9__9__26824));
  nnd2s1 _______443193(.DIN1 (__9_0___26616), .DIN2 (________23898), .Q
       (__9_____26823));
  nor2s1 _______443194(.DIN1 (__9_____26622), .DIN2 (__9_____26501), .Q
       (__9_____26822));
  nor2s1 _______443195(.DIN1 (________22859), .DIN2 (__9_____26648), .Q
       (__9_____26821));
  and2s1 _______443196(.DIN1 (__9_____26620), .DIN2 (_________30166),
       .Q (__9_____26820));
  nnd2s1 _____9_443197(.DIN1 (__9_____26640), .DIN2 (___00____27182),
       .Q (__9_____26819));
  nor2s1 _____0_443198(.DIN1 (___9_0__25184), .DIN2 (__9__9__26663), .Q
       (__9_____26818));
  and2s1 ______443199(.DIN1 (__9__0__26654), .DIN2 (__9__0__26816), .Q
       (__9_____26817));
  nor2s1 _______443200(.DIN1 (__99_9__27116), .DIN2 (__9_____26624), .Q
       (__9__9__26815));
  nor2s1 _______443201(.DIN1 (________19132), .DIN2 (__9_09__26617), .Q
       (__9_____26814));
  nnd2s1 _______443202(.DIN1 (__9_____26670), .DIN2 (__9_____26812), .Q
       (__9_____26813));
  nnd2s1 _______443203(.DIN1 (__9_99__26608), .DIN2 (________22926), .Q
       (__9_____26811));
  nnd2s1 _______443204(.DIN1 (____0____31872), .DIN2 (__9_____26809),
       .Q (__9_____26810));
  or2s1 _______443205(.DIN1 (__9_____26809), .DIN2 (____0____31872), .Q
       (__9_____26808));
  nor2s1 ______443206(.DIN1 (__9_____26728), .DIN2 (__9_0___26805), .Q
       (__9_0___26806));
  nnd2s1 _______443207(.DIN1 (__9_9___26607), .DIN2 (________22827), .Q
       (__9_0___26804));
  nnd2s1 _______443208(.DIN1 (__9_0___26612), .DIN2 (__9_0___26707), .Q
       (__9_0___26803));
  nor2s1 ______443209(.DIN1 (________21758), .DIN2 (__9_0___26613), .Q
       (__9_0___26802));
  nor2s1 ______443210(.DIN1 (___9____26182), .DIN2 (__9_____26668), .Q
       (__9__0__26969));
  xnr2s1 _______443211(.DIN1 (__9_00__26702), .DIN2 (______0__33107),
       .Q (__9_9___26890));
  and2s1 _______443212(.DIN1 (__9_____26625), .DIN2 (__9__0__26854), .Q
       (__9_9___26985));
  nor2s1 _______443213(.DIN1 (__9_____26809), .DIN2 (__9_0___26801), .Q
       (_________28289));
  xor2s1 _______443214(.DIN1 (__9_____26543), .DIN2 (_________31431),
       .Q (_________32304));
  nor2s1 ______443215(.DIN1 (_____0__24819), .DIN2 (__9_____26669), .Q
       (__9_____27031));
  or2s1 _______443216(.DIN1 (___9____26215), .DIN2 (__9_____26633), .Q
       (__9_09__26995));
  hi1s1 _______443217(.DIN (__9_0___26800), .Q (_________28549));
  dffacs1 _______________________443218(.CLRB (reset), .CLK (clk), .DIN
       (__9_90__26692), .QN (_____________________18641));
  nnd2s1 _______443219(.DIN1 (__9_____26578), .DIN2 (__9_00__26798), .Q
       (__9_0___26799));
  xor2s1 _______443220(.DIN1 (_______________18881), .DIN2
       (_________33007), .Q (__9_99__26797));
  nnd2s1 _____9_443221(.DIN1 (__9_____26835), .DIN2 (________23778), .Q
       (__9_9___26796));
  nor2s1 _____9_443222(.DIN1 (________22401), .DIN2 (__9_9___26603), .Q
       (__9_9___26795));
  nnd2s1 _____0_443223(.DIN1 (________23692), .DIN2 (__9_9___26601), .Q
       (__9_9___26794));
  nnd2s1 _____0_443224(.DIN1 (__9_____26561), .DIN2 (________24754), .Q
       (__9_9___26793));
  nnd2s1 _____443225(.DIN1 (__9_____26558), .DIN2 (__9_9___26791), .Q
       (__9_9___26792));
  nor2s1 _______443226(.DIN1 (___99___23432), .DIN2 (__9_90__26599), .Q
       (__9_9___26790));
  nor2s1 _______443227(.DIN1 (_____9__24828), .DIN2 (__9_____26568), .Q
       (__9_9___26789));
  nnd2s1 _______443228(.DIN1 (__9_____26594), .DIN2 (_________35006),
       .Q (__9_90__26788));
  nor2s1 _______443229(.DIN1 (__9_____26905), .DIN2 (__9_____26592), .Q
       (__9__9__26787));
  nor2s1 _______443230(.DIN1 (____9___25945), .DIN2 (__9__9__26588), .Q
       (__9_____26786));
  nor2s1 _______443231(.DIN1 (__9_____26784), .DIN2 (__9_____26587), .Q
       (__9_____26785));
  nnd2s1 _______443232(.DIN1 (__9_____26565), .DIN2 (________25692), .Q
       (__9_____26783));
  nnd2s1 _______443233(.DIN1 (__9_____26586), .DIN2 (___0____22566), .Q
       (__9_____26782));
  nnd2s1 _______443234(.DIN1 (__9_____26585), .DIN2 (__9_____26555), .Q
       (__9_____26781));
  nnd2s1 ______443235(.DIN1 (__9_____26596), .DIN2 (__9_____26779), .Q
       (__9_____26780));
  nor2s1 ______443236(.DIN1 (________24132), .DIN2 (__9_____26582), .Q
       (__9__0__26778));
  nor2s1 _______443237(.DIN1 (____99__24607), .DIN2 (__9__9__26569), .Q
       (__9__9__26777));
  nnd2s1 _______443238(.DIN1 (__9_____26580), .DIN2 (__9_____26962), .Q
       (__9_____26776));
  nor2s1 _______443239(.DIN1 (_____0___35036), .DIN2 (__9__9__26579),
       .Q (__9_____26775));
  or2s1 _______443240(.DIN1 (__9_____26773), .DIN2 (__9_9___26606), .Q
       (__9_____26774));
  nnd2s1 _______443241(.DIN1 (__9_____26574), .DIN2 (________24089), .Q
       (__9_____26772));
  nor2s1 _______443242(.DIN1 (__9_____26590), .DIN2 (__9_____26575), .Q
       (__9_____26771));
  nor2s1 _______443243(.DIN1 (__9__0__26570), .DIN2 (__9_____26675), .Q
       (__9_____26770));
  nnd2s1 ______443244(.DIN1 (__9_9___26602), .DIN2 (__9_____26686), .Q
       (__9_____26769));
  nor2s1 ______443245(.DIN1 (__9_9___26414), .DIN2 (__9_____26556), .Q
       (__9__0__26768));
  nor2s1 _______443246(.DIN1 (__9_____26499), .DIN2 (__9_____26584), .Q
       (__9__9__26767));
  nor2s1 _______443247(.DIN1 (__90_0), .DIN2 (__9__0__26589), .Q
       (__9_____26766));
  nor2s1 _______443248(.DIN1 (__9_____26764), .DIN2 (__9_____26573), .Q
       (__9_____26765));
  nnd2s1 _______443249(.DIN1 (_________31290), .DIN2 (_________31940),
       .Q (__9_____26763));
  hi1s1 _______443250(.DIN (__9_____26761), .Q (__9_____26762));
  nnd2s1 ______443251(.DIN1 (__9_____26567), .DIN2 (__9__0__27005), .Q
       (__9_____26760));
  nor2s1 ______443252(.DIN1 (_____9__26076), .DIN2 (__9__0__26560), .Q
       (__9_____26759));
  nor2s1 _______443253(.DIN1 (__9__9__26757), .DIN2 (__9_____26566), .Q
       (__9__0__26758));
  nor2s1 _______443254(.DIN1 (________22688), .DIN2 (__9_____26593), .Q
       (__9_____26756));
  nor2s1 _______443255(.DIN1 (__9_____26754), .DIN2 (__9_____26564), .Q
       (__9_____26755));
  nor2s1 _______443256(.DIN1 (_________31940), .DIN2 (_____0___35109),
       .Q (__9_____26753));
  nnd2s1 _______443257(.DIN1 (__9_____26549), .DIN2 (__9__9__27014), .Q
       (__9_____26752));
  nnd2s1 _______443258(.DIN1 (__9_____26571), .DIN2 (__9_____26937), .Q
       (__9_____26751));
  nor2s1 _______443259(.DIN1 (__9__0__26749), .DIN2 (__9__0__26551), .Q
       (__9_____26750));
  dffacs2 __________________443260(.CLRB (reset), .CLK (clk), .DIN
       (__9_9___26600), .Q (_______________18875));
  nor2s1 _______443261(.DIN1 (________25095), .DIN2 (______0__34778),
       .Q (__9__9__26748));
  nnd2s1 _____9_443262(.DIN1 (__9_9___26605), .DIN2 (__99____27091), .Q
       (__9_____26747));
  nnd2s1 _____9_443263(.DIN1 (_________31940), .DIN2 (_________31281),
       .Q (__9_____26746));
  nnd2s1 _____443264(.DIN1 (__9__9__26550), .DIN2 (________26084), .Q
       (__9_____26745));
  nor2s1 _____443265(.DIN1 (__9_____26743), .DIN2 (__9__9__26559), .Q
       (__9_____26744));
  nnd2s1 _____0_443266(.DIN1 (__9_____26563), .DIN2 (________22673), .Q
       (__9_____26742));
  nnd2s1 _____0_443267(.DIN1 (__9_____26554), .DIN2 (__9_____26639), .Q
       (__9_____26741));
  and2s1 _____0_443268(.DIN1 (__9_____26557), .DIN2 (__9__0__26739), .Q
       (__9_____26740));
  nnd2s1 _____443269(.DIN1 (__9_____26641), .DIN2 (__9__0__27005), .Q
       (__9__9__26738));
  or2s1 _______443270(.DIN1 (__9_____26736), .DIN2 (__9_____26595), .Q
       (__9_____26737));
  nnd2s1 ______443271(.DIN1 (__9_____26581), .DIN2 (__9_____26734), .Q
       (__9_____26735));
  nor2s1 _______443272(.DIN1 (__9_____26732), .DIN2 (__9_____26642), .Q
       (__9_____26733));
  nor2s1 ____9__443273(.DIN1 (__9_____26457), .DIN2 (__9_____26730), .Q
       (__9_____26731));
  nor2s1 _______443274(.DIN1 (outData[0]), .DIN2 (__9_99__26701), .Q
       (__9__0__26729));
  xor2s1 _______443275(.DIN1 (__9_____26433), .DIN2 (_________32901),
       .Q (__9_____26727));
  nnd2s1 _______443276(.DIN1 (__9_____26544), .DIN2 (________19536), .Q
       (__9_____26726));
  nor2s1 ______443277(.DIN1 (____0___26053), .DIN2 (__9_____26529), .Q
       (__9_____26725));
  nnd2s1 ______443278(.DIN1 (__9_____26536), .DIN2 (________25007), .Q
       (__9_____26724));
  and2s1 ______443279(.DIN1 (__9_____26530), .DIN2 (__9_____26722), .Q
       (__9_____26723));
  nor2s1 _______443280(.DIN1 (___9____24277), .DIN2 (__9_____26533), .Q
       (__9_____26721));
  or2s1 _____9_443281(.DIN1 (__9_9___26695), .DIN2 (__9__9__26598), .Q
       (__9__0__26720));
  nor2s1 _______443282(.DIN1 (________25437), .DIN2 (__9_____26539), .Q
       (__9__9__26719));
  and2s1 _____9_443283(.DIN1 (__9_____26538), .DIN2 (__9_____26717), .Q
       (__9_____26718));
  nnd2s1 _______443284(.DIN1 (__9_9___26700), .DIN2 (outData[11]), .Q
       (__9_____26716));
  xor2s1 _____9_443285(.DIN1 (____0___21076), .DIN2 (___0_9___27751),
       .Q (__9_____26715));
  or2s1 _______443286(.DIN1 (__9_____26713), .DIN2 (__9_____26534), .Q
       (__9_____26714));
  nor2s1 _______443287(.DIN1 (________23066), .DIN2 (__9__0__26523), .Q
       (__9__0__26712));
  nnd2s1 ______443288(.DIN1 (__9_0___26520), .DIN2 (__9_9___26791), .Q
       (__9_09__26711));
  nnd2s1 _______443289(.DIN1 (__9_____26524), .DIN2 (________23770), .Q
       (__9_0___26710));
  nor2s1 _______443290(.DIN1 (__99_9__27116), .DIN2 (__9_09__26522), .Q
       (__9_0___26709));
  nnd2s1 _______443291(.DIN1 (__9__0__26541), .DIN2 (__9_0___26707), .Q
       (__9_0___26708));
  xnr2s1 _______443292(.DIN1 (__9__9__26531), .DIN2 (___0_9___27751),
       .Q (__9_0___26706));
  nor2s1 _______443293(.DIN1 (_____0__24173), .DIN2 (__9_____26537), .Q
       (__9_0___26705));
  nnd2s1 _______443294(.DIN1 (__9_0___26703), .DIN2 (__9_____26527), .Q
       (__9_0___26704));
  nnd2s1 ______443295(.DIN1
       (______________________________________0_____________18887),
       .DIN2 (_________31940), .Q (__9_____26879));
  nor2s1 _____9_443296(.DIN1 (__90_9), .DIN2 (__9_____26526), .Q
       (__9_9___26884));
  nnd2s1 _____9_443297(.DIN1 (__9_____26528), .DIN2 (__9__0__26739), .Q
       (__9_____26881));
  nnd2s1 _______443298(.DIN1 (___99___26238), .DIN2 (__9_00__26702), .Q
       (__9_09__26807));
  xor2s1 ______443299(.DIN1 (__9_____26619), .DIN2 (__9__0__26618), .Q
       (__9_0___26800));
  nor2s1 _______443300(.DIN1 (________19609), .DIN2 (__9_99__26701), .Q
       (__9_____26908));
  nor2s1 _______443301(.DIN1 (outData[11]), .DIN2 (__9_9___26700), .Q
       (__9_____26974));
  or2s1 _______443302(.DIN1 (__9_9___26698), .DIN2 (__9_9___26509), .Q
       (__9_9___26699));
  nor2s1 _______443303(.DIN1 (__9_9___26505), .DIN2 (__9_9___26510), .Q
       (__9_9___26697));
  nor2s1 ______443304(.DIN1 (__9_9___26695), .DIN2 (__9_9___26508), .Q
       (__9_9___26696));
  nnd2s1 _______443305(.DIN1 (__9__9__26503), .DIN2 (____0___25858), .Q
       (__9_9___26694));
  nnd2s1 _______443306(.DIN1 (__900___26250), .DIN2 (__9__9__26493), .Q
       (__9_9___26693));
  nnd2s1 _______443307(.DIN1 (__9_99__26513), .DIN2 (__9__9__26691), .Q
       (__9_90__26692));
  nor2s1 _______443308(.DIN1 (___0_9__22581), .DIN2 (__9_____26502), .Q
       (__9_____26690));
  nnd2s1 _______443309(.DIN1 (__9_9___26512), .DIN2 (_________34982),
       .Q (__9_____26689));
  nor2s1 ______443310(.DIN1 (____9___22887), .DIN2 (__9_____26492), .Q
       (__9_____26688));
  and2s1 ______443311(.DIN1 (__9_____26500), .DIN2 (__9_____26686), .Q
       (__9_____26687));
  nnd2s1 ______443312(.DIN1 (__9_9___26506), .DIN2 (______0__35038), .Q
       (__9_____26685));
  and2s1 _____443313(.DIN1 (__9_____26497), .DIN2 (__9__9__27014), .Q
       (__9_____26684));
  nor2s1 _____9_443314(.DIN1 (_____9__23868), .DIN2 (__9_____26491), .Q
       (__9__0__26683));
  nor2s1 _____9_443315(.DIN1 (____00__24886), .DIN2 (__9_____26490), .Q
       (__9__9__26682));
  nnd2s1 _____9_443316(.DIN1
       (______________________________________0_____________18889),
       .DIN2 (_______________18881), .Q (__9_____26681));
  nnd2s1 _____0_443317(.DIN1 (__9_____26488), .DIN2 (___0____21654), .Q
       (__9_____26680));
  and2s1 _______443318(.DIN1 (__9_____26495), .DIN2 (__9_____26862), .Q
       (__9_____26679));
  and2s1 _______443319(.DIN1 (__9_____26677), .DIN2 (__9_0___26515), .Q
       (__9_____26678));
  nor2s1 _______443320(.DIN1 (_______________18881), .DIN2
       (__9_____26675), .Q (__9_____26676));
  or2s1 _______443321(.DIN1 (_______________18881), .DIN2
       (______0__32006), .Q (__9__0__26674));
  nnd2s1 _____0_443322(.DIN1 (_________34780), .DIN2 (_____9__22838),
       .Q (__9__9__26673));
  nor2s1 ______443323(.DIN1 (__9_____26671), .DIN2 (__9_____26478), .Q
       (__9_____26672));
  nor2s1 _______443324(.DIN1 (____0___24703), .DIN2 (__9_____26464), .Q
       (__9_____26670));
  nor2s1 _______443325(.DIN1 (___00____27202), .DIN2 (__9_____26626),
       .Q (__9_____26669));
  nnd2s1 ______443326(.DIN1 (__9_____26481), .DIN2 (__9_____26445), .Q
       (__9_____26668));
  nor2s1 _______443327(.DIN1 (________25983), .DIN2 (__9_____26466), .Q
       (__9_____26667));
  nnd2s1 _______443328(.DIN1 (__9_____26643), .DIN2 (outData[11]), .Q
       (__9_____26666));
  nnd2s1 _______443329(.DIN1 (__9_____26444), .DIN2 (__9__0__26664), .Q
       (__9_____26665));
  nnd2s1 _______443330(.DIN1 (__9_____26460), .DIN2 (____90__25840), .Q
       (__9__9__26663));
  nnd2s1 _______443331(.DIN1 (__9_____26474), .DIN2 (_________28478),
       .Q (__9_____26662));
  or2s1 _______443332(.DIN1 (__9_____26660), .DIN2 (__9_____26461), .Q
       (__9_____26661));
  and2s1 _______443333(.DIN1 (__9_____26657), .DIN2 (__9_____27045), .Q
       (__9_____26659));
  nor2s1 _______443334(.DIN1 (__9_____26657), .DIN2 (__9__0__26628), .Q
       (__9_____26658));
  nor2s1 _______443335(.DIN1 (__9_____26655), .DIN2 (__9_____26451), .Q
       (__9_____26656));
  nnd2s1 _______443336(.DIN1 (__9_____26483), .DIN2 (________21891), .Q
       (__9_____26850));
  nor2s1 _______443337(.DIN1 (____0___25857), .DIN2 (__9_____26562), .Q
       (__9_____26868));
  nnd2s1 _______443338(.DIN1 (__9_____26486), .DIN2 (__9_____26372), .Q
       (__9__9__26833));
  nnd2s1 ______443339(.DIN1 (_______________18881), .DIN2
       (_________31926), .Q (__9_____26878));
  nor2s1 _______443340(.DIN1 (_______________18881), .DIN2
       (______________________________________0_____________18886), .Q
       (__9_____26761));
  nnd2s1 _______443341(.DIN1
       (______________________________________0_____________18886),
       .DIN2 (_______________18881), .Q (__9__9__26911));
  nor2s1 _______443342(.DIN1 (___0____23491), .DIN2 (__9_____26443), .Q
       (__9__0__26654));
  nnd2s1 _____9_443343(.DIN1 (__9_____26465), .DIN2 (________22938), .Q
       (__9__9__26653));
  nor2s1 _____9_443344(.DIN1 (___0_0__24343), .DIN2 (__9_____26463), .Q
       (__9_____26652));
  or2s1 _____443345(.DIN1 (__9_____26650), .DIN2 (__9_____26462), .Q
       (__9_____26651));
  nor2s1 _____0_443346(.DIN1 (___0_9__22581), .DIN2 (__9_____26450), .Q
       (__9_____26649));
  or2s1 _____0_443347(.DIN1 (__9_____26647), .DIN2 (__9_____26498), .Q
       (__9_____26648));
  nnd2s1 _______443348(.DIN1 (__9_____26479), .DIN2 (____9___22713), .Q
       (__9_____26646));
  nor2s1 _______443349(.DIN1 (________25715), .DIN2 (__9_____26468), .Q
       (__9__0__26645));
  nor2s1 _______443350(.DIN1 (outData[11]), .DIN2 (__9_____26643), .Q
       (__9__9__26644));
  and2s1 _______443351(.DIN1 (__9_____26442), .DIN2 (__9_____26639), .Q
       (__9_____26640));
  nor2s1 _______443352(.DIN1 (__9__0__26637), .DIN2 (__9__0__26477), .Q
       (__9_____26638));
  nor2s1 _______443353(.DIN1 (___0_9__22581), .DIN2 (__9_____26635), .Q
       (__9__9__26636));
  nnd2s1 _______443354(.DIN1 (__9_____26453), .DIN2 (____9___23800), .Q
       (__9_____26634));
  or2s1 _______443355(.DIN1 (__9_____26632), .DIN2 (__9_____26473), .Q
       (__9_____26633));
  nor2s1 ______443356(.DIN1 (___9____25200), .DIN2 (__9__9__26448), .Q
       (__9_____26630));
  nnd2s1 _______443357(.DIN1 (__9__0__26628), .DIN2 (__9_____26469), .Q
       (__9_____26629));
  nnd2s1 _____9_443358(.DIN1 (__9_____26626), .DIN2 (________24074), .Q
       (__9__9__26627));
  nor2s1 _______443359(.DIN1 (__9_9___26695), .DIN2 (__9_____26446), .Q
       (__9_____26625));
  and2s1 ______443360(.DIN1 (__9_____26436), .DIN2 (__9_____26623), .Q
       (__9_____26624));
  nor2s1 ______443361(.DIN1 (__9_____26621), .DIN2 (__9_____26441), .Q
       (__9_____26622));
  and2s1 _______443362(.DIN1 (__9_____26619), .DIN2 (__9__0__26618), .Q
       (__9_____26620));
  nor2s1 _______443363(.DIN1 (____0___19121), .DIN2 (__9_____26619), .Q
       (__9_09__26617));
  nor2s1 _______443364(.DIN1 (________22278), .DIN2 (__9__9__26438), .Q
       (__9_0___26616));
  nor2s1 ____9__443365(.DIN1 (____9____34518), .DIN2 (__9_____26456),
       .Q (__9_0___26615));
  nor2s1 _______443366(.DIN1 (__99_9__27116), .DIN2 (__9_0___26425), .Q
       (__9_0___26614));
  nor2s1 _______443367(.DIN1 (________22393), .DIN2 (__9_0___26426), .Q
       (__9_0___26613));
  nor2s1 _______443368(.DIN1 (________26094), .DIN2 (__9_____26434), .Q
       (__9_0___26612));
  or2s1 ______443369(.DIN1 (_________28603), .DIN2 (___0_9___27751), .Q
       (__9_0___26611));
  nnd2s1 _______443370(.DIN1 (___0_9___27751), .DIN2 (_________28603),
       .Q (__9_0___26610));
  nor2s1 ______443371(.DIN1 (____90__23704), .DIN2 (__9_09__26428), .Q
       (__9_0___26609));
  nnd2s1 ____9__443372(.DIN1 (__9_____26455), .DIN2 (________21469), .Q
       (__9_99__26608));
  nnd2s1 ____443373(.DIN1 (________25142), .DIN2 (__9_____26430), .Q
       (__9_9___26607));
  nor2s1 ____9__443374(.DIN1 (___0_9___27751), .DIN2
       (______________18869), .Q (__9_____26728));
  xnr2s1 _____443375(.DIN1 (outData[10]), .DIN2 (__9_____26542), .Q
       (_________29406));
  nnd2s1 _______443376(.DIN1 (___0_9___27751), .DIN2 (___0_____27914),
       .Q (__9_____26809));
  or2s1 ______443377(.DIN1 (________25728), .DIN2 (__9_99), .Q
       (__9_9___26606));
  and2s1 _______443378(.DIN1 (__9_____26388), .DIN2 (__9_9___26604), .Q
       (__9_9___26605));
  nnd2s1 _______443379(.DIN1 (__9__9__26375), .DIN2 (________21759), .Q
       (__9_9___26603));
  nor2s1 _______443380(.DIN1 (____0___26055), .DIN2 (__9_____26411), .Q
       (__9_9___26602));
  nor2s1 _______443381(.DIN1 (___9_9__26166), .DIN2 (__9_____26385), .Q
       (__9_9___26601));
  nnd2s1 _______443382(.DIN1 (__9__9__26412), .DIN2 (________23678), .Q
       (__9_9___26600));
  nnd2s1 _______443383(.DIN1 (__9_____26410), .DIN2 (___99___26242), .Q
       (__9_90__26599));
  or2s1 _______443384(.DIN1 (__9_____26597), .DIN2 (__9_____26407), .Q
       (__9__9__26598));
  nor2s1 _______443385(.DIN1 (__9__0__26449), .DIN2 (__9_0___26420), .Q
       (__9_____26596));
  nnd2s1 ______443386(.DIN1 (__9_____26363), .DIN2 (________23243), .Q
       (__9_____26595));
  nor2s1 _______443387(.DIN1 (___0090__27257), .DIN2 (__9_____26409),
       .Q (__9_____26594));
  nnd2s1 _______443388(.DIN1 (__9_____26408), .DIN2 (___9____26159), .Q
       (__9_____26593));
  nnd2s1 _______443389(.DIN1 (__9_9___26417), .DIN2 (__9_____26591), .Q
       (__9_____26592));
  nor2s1 _______443390(.DIN1 (________22146), .DIN2 (__9_____26382), .Q
       (__9_____26590));
  nnd2s1 _______443391(.DIN1 (__9_____26405), .DIN2 (________25774), .Q
       (__9__0__26589));
  or2s1 ______443392(.DIN1 (________25872), .DIN2 (__9_____26402), .Q
       (__9__9__26588));
  nnd2s1 _______443393(.DIN1 (__9_____26374), .DIN2 (___00____27182),
       .Q (__9_____26587));
  nor2s1 _______443394(.DIN1 (____0___25368), .DIN2 (__9_____26398), .Q
       (__9_____26586));
  nor2s1 _____443395(.DIN1 (________25593), .DIN2 (__9_____26400), .Q
       (__9_____26585));
  or2s1 _____9_443396(.DIN1 (__9_____26583), .DIN2 (__9__0__26403), .Q
       (__9_____26584));
  nnd2s1 _____9_443397(.DIN1 (__9_____26371), .DIN2 (________25452), .Q
       (__9_____26582));
  nor2s1 _____9_443398(.DIN1 (________24691), .DIN2 (__9_____26396), .Q
       (__9_____26581));
  nnd2s1 _____0_443399(.DIN1 (__9__0__26366), .DIN2 (___900__26147), .Q
       (__9_____26580));
  nnd2s1 _____0_443400(.DIN1 (__9_____26392), .DIN2 (________23652), .Q
       (__9__9__26579));
  nor2s1 _____0_443401(.DIN1 (____90__21345), .DIN2 (__9_____26390), .Q
       (__9_____26578));
  nnd2s1 ______443402(.DIN1 (__9_____26480), .DIN2 (__9_____26576), .Q
       (__9_____26577));
  nor2s1 _______443403(.DIN1 (___0_9__22581), .DIN2 (__9__9__26365), .Q
       (__9_____26575));
  nor2s1 _______443404(.DIN1 (____90__25939), .DIN2 (__9_90), .Q
       (__9_____26574));
  or2s1 _______443405(.DIN1 (__9_____26572), .DIN2 (__9_____26380), .Q
       (__9_____26573));
  nor2s1 ______443406(.DIN1 (___9_0__26157), .DIN2 (__9_____26379), .Q
       (__9_____26571));
  nor2s1 ______443407(.DIN1 (____0___24155), .DIN2 (__9_____26369), .Q
       (__9__0__26570));
  nnd2s1 _______443408(.DIN1 (__9_____26395), .DIN2 (________25643), .Q
       (__9__9__26569));
  nnd2s1 _______443409(.DIN1 (__9__0__26376), .DIN2 (___0____23502), .Q
       (__9_____26568));
  nnd2s1 _______443410(.DIN1 (__9_____26373), .DIN2 (___0__0__27287),
       .Q (__9_____26567));
  nnd2s1 _______443411(.DIN1 (__9_____26351), .DIN2 (__9_____26840), .Q
       (__9_____26566));
  nor2s1 _______443412(.DIN1 (________25536), .DIN2 (__9_9_), .Q
       (__9_____26565));
  nnd2s1 _______443413(.DIN1 (__9_____26397), .DIN2 (________22879), .Q
       (__9_____26564));
  nnd2s1 ______443414(.DIN1 (__9_____26367), .DIN2 (___9____26163), .Q
       (__9_____26563));
  hi1s1 _______443415(.DIN (__9_____26562), .Q (__9_99__26701));
  hi1s1 _______443416(.DIN (_______________18881), .Q (_________31940));
  nor2s1 _______443417(.DIN1 (__9_____26386), .DIN2 (__9__9__26393), .Q
       (__9_____26561));
  nor2s1 _______443418(.DIN1 (__90____26312), .DIN2 (__9_____26349), .Q
       (__9__0__26560));
  nnd2s1 ______443419(.DIN1 (__9_____26359), .DIN2 (___00____27220), .Q
       (__9__9__26559));
  nor2s1 _______443420(.DIN1 (________22425), .DIN2 (__9_9___26413), .Q
       (__9_____26558));
  and2s1 _______443421(.DIN1 (__9_9___26415), .DIN2 (______0__28974),
       .Q (__9_____26557));
  nnd2s1 ______443422(.DIN1 (__9_____26357), .DIN2 (__9_____26555), .Q
       (__9_____26556));
  nor2s1 ______443423(.DIN1 (__9_____26553), .DIN2 (__9_____26353), .Q
       (__9_____26554));
  nnd2s1 _______443424(.DIN1 (__9_____26361), .DIN2 (____9___21899), .Q
       (__9_____26552));
  nnd2s1 _______443425(.DIN1 (__9_____26399), .DIN2 (_____0__22337), .Q
       (__9__0__26551));
  nor2s1 _______443426(.DIN1 (____9___26142), .DIN2 (__9__9__26355), .Q
       (__9__9__26550));
  nor2s1 _______443427(.DIN1 (__9_____26548), .DIN2 (__9_____26347), .Q
       (__9_____26549));
  or2s1 _______443428(.DIN1 (__9_____26546), .DIN2 (__9_____26545), .Q
       (__9_____26547));
  nor2s1 ____0__443429(.DIN1 (________19083), .DIN2 (__9_____26345), .Q
       (__9_____26544));
  and2s1 ____9__443430(.DIN1 (__9_____26542), .DIN2 (__90____26260), .Q
       (__9_____26543));
  and2s1 ____9__443431(.DIN1 (__909___26331), .DIN2 (__9__9__26540), .Q
       (__9__0__26541));
  nnd2s1 _____0_443432(.DIN1 (__9_0___26340), .DIN2 (________25726), .Q
       (__9_____26539));
  nor2s1 _______443433(.DIN1 (___0____22597), .DIN2 (__9_____26341), .Q
       (__9_____26538));
  nnd2s1 _______443434(.DIN1 (__9__0), .DIN2 (__90_0__26291), .Q
       (__9_____26537));
  nor2s1 _______443435(.DIN1 (__9_0___26518), .DIN2 (__9_____26470), .Q
       (__9_____26536));
  nnd2s1 _______443436(.DIN1 (__9_0___26339), .DIN2 (________25451), .Q
       (__9_____26534));
  nnd2s1 _______443437(.DIN1 (__909___26332), .DIN2 (____9___23794), .Q
       (__9_____26533));
  nnd2s1 ______443438(.DIN1 (__9__9__26531), .DIN2 (____________), .Q
       (__9__0__26532));
  and2s1 _____9_443439(.DIN1 (__9_09), .DIN2 (__99____27150), .Q
       (__9_____26530));
  nnd2s1 ____90_443440(.DIN1 (__909___26333), .DIN2 (___0____25307), .Q
       (__9_____26529));
  and2s1 ____90_443441(.DIN1 (__9_0___26336), .DIN2 (_________35010),
       .Q (__9_____26528));
  nnd2s1 ____9__443442(.DIN1 (____________), .DIN2
       (______________18867), .Q (__9_____26527));
  nnd2s1 ____9__443443(.DIN1 (__9099), .DIN2 (__9_____26525), .Q
       (__9_____26526));
  nor2s1 ____9__443444(.DIN1 (____0___22812), .DIN2 (__9_0_), .Q
       (__9_____26524));
  nnd2s1 ____9_443445(.DIN1 (__9_0___26337), .DIN2 (____99__25654), .Q
       (__9__0__26523));
  nor2s1 ____9__443446(.DIN1 (__9_0___26521), .DIN2 (__9___), .Q
       (__9_09__26522));
  nor2s1 ____9__443447(.DIN1 (____9___22078), .DIN2 (__9_0___26334), .Q
       (__9_0___26520));
  and2s1 ____9_443448(.DIN1 (__9_0___26518), .DIN2 (__9_____27045), .Q
       (__9_0___26519));
  nnd2s1 _____9_443449(.DIN1 (__9_____26352), .DIN2 (__9_0___26517), .Q
       (__9_____26641));
  or2s1 ____9__443450(.DIN1 (outData[10]), .DIN2 (__9_____26542), .Q
       (__9_9___26700));
  nor2s1 ____9__443451(.DIN1 (____________), .DIN2 (_________28866), .Q
       (__9_00__26702));
  xor2s1 _____9_443452(.DIN1 (____9___19200), .DIN2 (___99___26239), .Q
       (__9_____26642));
  nor2s1 _______443453(.DIN1 (__9__0__26459), .DIN2 (__9_0___26516), .Q
       (_____9___30175));
  nor2s1 _______443454(.DIN1 (__9_____26344), .DIN2 (_________33174),
       .Q (__9_____26730));
  nor2s1 _____443455(.DIN1 (____99__26146), .DIN2 (__9_____26364), .Q
       (__9_____26835));
  xor2s1 _____9_443456(.DIN1 (outData[10]), .DIN2 (__9_0___26423), .Q
       (___09____28062));
  xor2s1 _______443457(.DIN1 (__9__9__26384), .DIN2 (__9_00__26514), .Q
       (__9_0___26515));
  nor2s1 _______443458(.DIN1 (________25620), .DIN2 (__90____26326), .Q
       (__9_99__26513));
  nor2s1 ______443459(.DIN1 (__9_9___26511), .DIN2 (__90____26323), .Q
       (__9_9___26512));
  or2s1 _______443460(.DIN1 (__9_____26452), .DIN2 (__90____26321), .Q
       (__9_9___26510));
  nnd2s1 _______443461(.DIN1 (__90____26311), .DIN2 (_____0__22952), .Q
       (__9_9___26509));
  nnd2s1 _______443462(.DIN1 (__90____26320), .DIN2 (__9_9___26507), .Q
       (__9_9___26508));
  nor2s1 _______443463(.DIN1 (__9_9___26505), .DIN2 (__90____26307), .Q
       (__9_9___26506));
  nnd2s1 _______443464(.DIN1 (__9_9___26418), .DIN2 (___00____27211),
       .Q (__9_90__26504));
  nor2s1 _____9_443465(.DIN1 (________25797), .DIN2 (__90____26313), .Q
       (__9__9__26503));
  and2s1 _____443466(.DIN1 (__90_0__26300), .DIN2 (_________35010), .Q
       (__9_____26502));
  nnd2s1 _____0_443467(.DIN1 (__90____26305), .DIN2 (________25017), .Q
       (__9_____26501));
  nor2s1 _____443468(.DIN1 (__9_____26499), .DIN2 (__90____26319), .Q
       (__9_____26500));
  or2s1 _______443469(.DIN1 (________25424), .DIN2 (__90____26277), .Q
       (__9_____26498));
  and2s1 _______443470(.DIN1 (__90_0__26309), .DIN2 (__9_____26496), .Q
       (__9_____26497));
  and2s1 _______443471(.DIN1 (__90____26322), .DIN2 (__9__0__26494), .Q
       (__9_____26495));
  nnd2s1 _______443472(.DIN1 (__90_9__26317), .DIN2 (________22673), .Q
       (__9__9__26493));
  nnd2s1 ______443473(.DIN1 (__90_9__26299), .DIN2 (________23112), .Q
       (__9_____26492));
  or2s1 _______443474(.DIN1 (______0__28751), .DIN2 (__90____26301), .Q
       (__9_____26491));
  nnd2s1 _______443475(.DIN1 (__90____26302), .DIN2 (__9_____26489), .Q
       (__9_____26490));
  or2s1 _______443476(.DIN1 (__9_____26487), .DIN2 (__90____26298), .Q
       (__9_____26488));
  nor2s1 _______443477(.DIN1 (__9__0__26485), .DIN2 (__90____26304), .Q
       (__9_____26486));
  nor2s1 _______443478(.DIN1 (_____9__21884), .DIN2 (__909_), .Q
       (__9__9__26484));
  nor2s1 _______443479(.DIN1 (__9_____26435), .DIN2 (__90____26303), .Q
       (__9_____26483));
  xor2s1 _____9_443480(.DIN1 (_________34485), .DIN2 (___0_____27475),
       .Q (__9_____26482));
  nor2s1 _______443481(.DIN1 (___0090__27257), .DIN2 (__90_0__26261),
       .Q (__9_____26481));
  and2s1 _____443482(.DIN1 (__90____26263), .DIN2 (___0____22575), .Q
       (__9_____26479));
  nnd2s1 ______443483(.DIN1 (__90____26254), .DIN2 (________25509), .Q
       (__9_____26478));
  nnd2s1 _______443484(.DIN1 (__90____26276), .DIN2 (__9__9__26476), .Q
       (__9__0__26477));
  nor2s1 _______443485(.DIN1 (___0_9__22581), .DIN2 (__90____26324), .Q
       (__9_____26475));
  nor2s1 _______443486(.DIN1 (___0__0__28004), .DIN2 (__90____26293),
       .Q (__9_____26474));
  or2s1 _______443487(.DIN1 (__9_____26472), .DIN2 (__90____26272), .Q
       (__9_____26473));
  nnd2s1 _______443488(.DIN1 (__9_____26470), .DIN2 (__9_____26469), .Q
       (__9_____26471));
  nnd2s1 _______443489(.DIN1 (__90____26257), .DIN2 (________25991), .Q
       (__9_____26468));
  or2s1 _______443490(.DIN1 (___0__9__27771), .DIN2 (__90____26285), .Q
       (__9__0__26467));
  nnd2s1 _______443491(.DIN1 (__9000), .DIN2 (___0____24393), .Q
       (__9_____26466));
  xor2s1 _____9_443492(.DIN1 (_____0___28530), .DIN2 (__909___26329),
       .Q (__9_____26562));
  dffacs2 __________________443493(.CLRB (reset), .CLK (clk), .DIN
       (__90____26325), .Q (_______________18881));
  nor2s1 _______443494(.DIN1 (________22965), .DIN2 (__90_9__26280), .Q
       (__9_____26465));
  or2s1 _______443495(.DIN1 (___9_0__24267), .DIN2 (__900___26251), .Q
       (__9_____26464));
  nnd2s1 ______443496(.DIN1 (__90____26279), .DIN2 (________23738), .Q
       (__9_____26463));
  nnd2s1 _______443497(.DIN1 (__90____26278), .DIN2 (___00____27222),
       .Q (__9_____26462));
  or2s1 _______443498(.DIN1 (________25887), .DIN2 (__90____26294), .Q
       (__9_____26461));
  and2s1 _______443499(.DIN1 (__90____26283), .DIN2 (________25926), .Q
       (__9_____26460));
  nor2s1 _______443500(.DIN1 (_______________18878), .DIN2
       (__90____26264), .Q (__9__9__26458));
  nor2s1 ______443501(.DIN1 (__9_____26343), .DIN2 (__9_____26456), .Q
       (__9_____26457));
  nnd2s1 _______443502(.DIN1 (___9____26233), .DIN2 (____9___22886), .Q
       (__9_____26455));
  or2s1 _____0_443503(.DIN1 (__9_0___26703), .DIN2 (_________32049), .Q
       (__9_____26454));
  nor2s1 ____90_443504(.DIN1 (__9_____26452), .DIN2 (__90__), .Q
       (__9_____26453));
  nnd2s1 ____90_443505(.DIN1 (__90____26259), .DIN2 (________23119), .Q
       (__9_____26451));
  nor2s1 ____443506(.DIN1 (__9__0__26449), .DIN2 (__9009), .Q
       (__9_____26450));
  nnd2s1 ____9_443507(.DIN1 (__90____26314), .DIN2 (__9_____26447), .Q
       (__9__9__26448));
  nnd2s1 ____9__443508(.DIN1 (__90____26288), .DIN2 (__9_____26445), .Q
       (__9_____26446));
  nor2s1 ____9_443509(.DIN1 (___9____26213), .DIN2 (__90____26295), .Q
       (__9_____26444));
  nor2s1 ____9__443510(.DIN1 (________21758), .DIN2 (__900___26247), .Q
       (__9_____26443));
  nor2s1 ____9__443511(.DIN1 (__9_____26784), .DIN2 (___99___26243), .Q
       (__9_____26442));
  nor2s1 ____9__443512(.DIN1 (__9_____26440), .DIN2 (__900___26248), .Q
       (__9_____26441));
  nnd2s1 ____9__443513(.DIN1 (__90____26292), .DIN2 (__9_____27045), .Q
       (__9__0__26439));
  nnd2s1 ____9__443514(.DIN1 (__90____26274), .DIN2 (_____0__22653), .Q
       (__9__9__26438));
  nnd2s1 ____9__443515(.DIN1 (___99___26245), .DIN2 (___99___26241), .Q
       (__9_____26437));
  nor2s1 ____9__443516(.DIN1 (__9_____26435), .DIN2 (__900___26249), .Q
       (__9_____26436));
  or2s1 ____09_443517(.DIN1 (__90_0__26281), .DIN2 (___9_9__26236), .Q
       (__9_____26434));
  nor2s1 ____9__443518(.DIN1 (__9_____26432), .DIN2 (__9_____26431), .Q
       (__9_____26433));
  xor2s1 ____09_443519(.DIN1 (_____0___30458), .DIN2 (_____9___30627),
       .Q (__9_____26430));
  xor2s1 ____09_443520(.DIN1 (_________31058), .DIN2 (_____0___30458),
       .Q (__9__0__26429));
  or2s1 ____0__443521(.DIN1 (__9_0___26427), .DIN2 (__90____26266), .Q
       (__9_09__26428));
  nnd2s1 ____99_443522(.DIN1 (___9____26234), .DIN2 (________24660), .Q
       (__9_0___26426));
  nor2s1 ____9__443523(.DIN1 (___9____26171), .DIN2 (___990__26237), .Q
       (__9_0___26425));
  nnd2s1 _______443524(.DIN1 (__90____26282), .DIN2 (__9_0___26424), .Q
       (__9_____26657));
  nor2s1 ____9_443525(.DIN1 (__90____26289), .DIN2 (__9_0___26423), .Q
       (_________29637));
  and2s1 ____9__443526(.DIN1 (__90____26255), .DIN2 (__99____27091), .Q
       (__9_____26635));
  or2s1 ____9_443527(.DIN1 (__9_0___26422), .DIN2 (__90_9__26290), .Q
       (__9__0__26628));
  dffacs1 __________________443528(.CLRB (reset), .CLK (clk), .DIN
       (___99___26244), .Q (________________18675));
  nor2s1 _______443529(.DIN1 (__9_____26342), .DIN2 (__9_0___26421), .Q
       (_________29592));
  nnd2s1 _______443530(.DIN1 (__9_0___26423), .DIN2 (____99__19113), .Q
       (__9_____26643));
  nor2s1 _______443531(.DIN1 (__9_____26572), .DIN2 (__90____26296), .Q
       (__9_____26626));
  xor2s1 ____9__443532(.DIN1 (________26111), .DIN2 (______0__33107),
       .Q (__9_____26619));
  hi1s1 ____9__443533(.DIN (____________), .Q (___0_9___27751));
  nnd2s1 _______443534(.DIN1 (___9____26198), .DIN2 (__9_00__26419), .Q
       (__9_0___26420));
  nnd2s1 _______443535(.DIN1 (___9____26225), .DIN2 (___99___22533), .Q
       (__9_99));
  nor2s1 _____0_443536(.DIN1 (__9_9___26416), .DIN2 (___9_9__26186), .Q
       (__9_9___26417));
  nor2s1 _____0_443537(.DIN1 (__9_9___26414), .DIN2 (___9____26219), .Q
       (__9_9___26415));
  nnd2s1 _____0_443538(.DIN1 (___9____26208), .DIN2 (________22706), .Q
       (__9_9___26413));
  and2s1 _____0_443539(.DIN1 (___9____26212), .DIN2 (__9_____26469), .Q
       (__9_9_));
  nnd2s1 _______443540(.DIN1 (___9____26188), .DIN2 (__9_00__26419), .Q
       (__9_90));
  nnd2s1 _______443541(.DIN1 (___9____26169), .DIN2 (inData[30]), .Q
       (__9__9__26412));
  or2s1 ______443542(.DIN1 (___9____23391), .DIN2 (___909__26156), .Q
       (__9_____26411));
  nor2s1 ______443543(.DIN1 (________25901), .DIN2 (___9____26204), .Q
       (__9_____26410));
  nnd2s1 _______443544(.DIN1 (___9____26165), .DIN2 (_____9__25596), .Q
       (__9_____26409));
  nor2s1 _______443545(.DIN1 (________23101), .DIN2 (___9____26203), .Q
       (__9_____26408));
  nnd2s1 _______443546(.DIN1 (___9____26202), .DIN2 (__9_____26406), .Q
       (__9_____26407));
  and2s1 _______443547(.DIN1 (___9____26183), .DIN2 (________25392), .Q
       (__9_____26405));
  nor2s1 _______443548(.DIN1 (___0_9__22581), .DIN2 (___9____26201), .Q
       (__9_____26404));
  nnd2s1 _______443549(.DIN1 (___9_0__26187), .DIN2 (_____90__34918),
       .Q (__9__0__26403));
  nnd2s1 _______443550(.DIN1 (___90___26152), .DIN2 (__9_____26401), .Q
       (__9_____26402));
  nnd2s1 _______443551(.DIN1 (___9____26222), .DIN2 (________25641), .Q
       (__9_____26400));
  nor2s1 _______443552(.DIN1 (________25989), .DIN2 (___9____26214), .Q
       (__9_____26399));
  nnd2s1 _______443553(.DIN1 (__90____26297), .DIN2 (_____0__24916), .Q
       (__9_____26398));
  nor2s1 ____9__443554(.DIN1 (________23328), .DIN2 (___9____26189), .Q
       (__9_____26397));
  nor2s1 ______443555(.DIN1 (___00____27202), .DIN2 (___9____26224), .Q
       (__9_____26396));
  and2s1 _______443556(.DIN1 (___9_0__26197), .DIN2 (__9__0__26394), .Q
       (__9_____26395));
  nnd2s1 _______443557(.DIN1 (___9____26205), .DIN2 (___0_____27594),
       .Q (__9__9__26393));
  nor2s1 _______443558(.DIN1 (_____9__23554), .DIN2 (___9_9__26196), .Q
       (__9_____26392));
  nor2s1 ______443559(.DIN1 (___0_9__22581), .DIN2 (___9____26195), .Q
       (__9_____26391));
  nnd2s1 _______443560(.DIN1 (___9____26168), .DIN2 (__9_____26389), .Q
       (__9_____26390));
  and2s1 _______443561(.DIN1 (___9____26190), .DIN2 (__9_____26387), .Q
       (__9_____26388));
  nor2s1 ____9_443562(.DIN1 (___00____27202), .DIN2 (___9____26178), .Q
       (__9_____26386));
  nor2s1 _______443563(.DIN1
       (______________________________________0__________0), .DIN2
       (__9__9__26384), .Q (__9_____26385));
  nnd2s1 ______443564(.DIN1 (___9____26172), .DIN2 (__9_____27045), .Q
       (__9_____26383));
  nor2s1 _____443565(.DIN1 (__9_____26381), .DIN2 (___9____26173), .Q
       (__9_____26382));
  nnd2s1 _____9_443566(.DIN1 (____9___26143), .DIN2 (______0__34998),
       .Q (__9_____26380));
  nnd2s1 _____9_443567(.DIN1 (___9____26160), .DIN2 (________26018), .Q
       (__9_____26379));
  nor2s1 _____9_443568(.DIN1 (________23221), .DIN2 (___9____26184), .Q
       (__9_____26378));
  nnd2s1 _____9_443569(.DIN1 (___9_0__26217), .DIN2 (____9___21899), .Q
       (__9_____26377));
  nor2s1 _____9_443570(.DIN1 (__90____26258), .DIN2 (___9____26191), .Q
       (__9__0__26376));
  nor2s1 _____443571(.DIN1 (___0____22579), .DIN2 (___9____26221), .Q
       (__9__9__26375));
  nor2s1 ____90_443572(.DIN1 (________25524), .DIN2 (___9____26192), .Q
       (__9_____26374));
  and2s1 ____90_443573(.DIN1 (________26128), .DIN2 (__9_____26372), .Q
       (__9_____26373));
  nor2s1 ____90_443574(.DIN1 (____9___24060), .DIN2 (___9____26180), .Q
       (__9_____26371));
  nnd2s1 _______443575(.DIN1 (___9_9__26216), .DIN2 (__9_____26370), .Q
       (__9_____26480));
  dffacs1 ___________________443576(.CLRB (reset), .CLK (clk), .DIN
       (___9____26193), .Q (_________________18680));
  dffacs1 _____________________0_443577(.CLRB (reset), .CLK (clk), .DIN
       (___9____26170), .QN (_________________0___18597));
  xor2s1 ____9__443578(.DIN1 (__9_____26368), .DIN2 (_____0__26007), .Q
       (__9_____26369));
  nor2s1 ____9__443579(.DIN1 (___9____24318), .DIN2 (___9____26211), .Q
       (__9_____26367));
  nor2s1 ____9__443580(.DIN1 (________26101), .DIN2 (___90___26155), .Q
       (__9__0__26366));
  nor2s1 ____9__443581(.DIN1 (___09___23520), .DIN2 (___9____26175), .Q
       (__9__9__26365));
  nor2s1 ____9__443582(.DIN1 (______9__33856), .DIN2 (____9___26140),
       .Q (__9_____26364));
  and2s1 ____9__443583(.DIN1 (___9____26185), .DIN2 (__9_____26362), .Q
       (__9_____26363));
  or2s1 ____9__443584(.DIN1 (__9_____26381), .DIN2 (___9_9__26206), .Q
       (__9_____26361));
  nnd2s1 ____9__443585(.DIN1 (___90___26150), .DIN2 (___00____27211),
       .Q (__9_____26360));
  and2s1 ____9__443586(.DIN1 (___9____26199), .DIN2 (__9_____26358), .Q
       (__9_____26359));
  nor2s1 ____9_443587(.DIN1 (__9__0__26356), .DIN2 (___9____26210), .Q
       (__9_____26357));
  nnd2s1 ____9__443588(.DIN1 (___9____26164), .DIN2 (__9_____26354), .Q
       (__9__9__26355));
  nnd2s1 ____9__443589(.DIN1 (___9____26158), .DIN2 (________23917), .Q
       (__9_____26353));
  nor2s1 ____9__443590(.DIN1 (___90___22450), .DIN2 (___90___26153), .Q
       (__9_____26352));
  nor2s1 ____9_443591(.DIN1 (__9_____26350), .DIN2 (____9___26145), .Q
       (__9_____26351));
  nor2s1 ____9__443592(.DIN1 (________21758), .DIN2 (___90___26148), .Q
       (__9_____26349));
  nnd2s1 ____9__443593(.DIN1 (____9___26141), .DIN2 (__9__0__27005), .Q
       (__9_____26348));
  or2s1 ____9__443594(.DIN1 (__9__0__26346), .DIN2 (___9____26161), .Q
       (__9_____26347));
  nnd2s1 ____9__443595(.DIN1 (________26024), .DIN2 (____9___26139), .Q
       (__9__9));
  nor2s1 ______443596(.DIN1 (_____0___30458), .DIN2
       (_____________________18662), .Q (__9_____26345));
  hi1s1 _______443597(.DIN (__9_____26343), .Q (__9_____26344));
  nnd2s1 ____9__443598(.DIN1 (________26132), .DIN2 (________25604), .Q
       (__9_____26341));
  nnd2s1 ____9__443599(.DIN1 (________26118), .DIN2 (___009__25280), .Q
       (__9___));
  and2s1 ____99_443600(.DIN1 (____9___26138), .DIN2 (________26079), .Q
       (__9__0));
  and2s1 ____00_443601(.DIN1 (________26124), .DIN2 (___09____28103),
       .Q (__9_09));
  nor2s1 ____0__443602(.DIN1 (____0___24888), .DIN2 (________26120), .Q
       (__9_0___26340));
  nor2s1 ____0__443603(.DIN1 (__9_0___26338), .DIN2 (________26115), .Q
       (__9_0___26339));
  nor2s1 ____0__443604(.DIN1 (____9___25746), .DIN2 (________26114), .Q
       (__9_0___26337));
  nor2s1 ____0__443605(.DIN1 (________23238), .DIN2 (________26119), .Q
       (__9_0___26336));
  and2s1 ____0__443606(.DIN1 (________26113), .DIN2 (________21886), .Q
       (__9_0___26335));
  nnd2s1 _______443607(.DIN1 (________26110), .DIN2 (________26020), .Q
       (__9_0___26334));
  nnd2s1 _____0_443608(.DIN1 (________26135), .DIN2 (__9_00), .Q
       (__9_0_));
  nor2s1 ____0__443609(.DIN1 (___0_0___27370), .DIN2 (________26122),
       .Q (__9099));
  nor2s1 ____0_443610(.DIN1 (________24749), .DIN2 (___9____26162), .Q
       (__909___26333));
  nor2s1 ____0__443611(.DIN1 (________25710), .DIN2 (________26134), .Q
       (__909___26332));
  and2s1 ____09_443612(.DIN1 (________26131), .DIN2 (__9_0___26424), .Q
       (__909___26331));
  nnd2s1 ____09_443613(.DIN1 (________26133), .DIN2 (_____9___28891),
       .Q (__909___26330));
  and2s1 ____9__443614(.DIN1 (__909___26329), .DIN2 (_____9__26106), .Q
       (__9_____26958));
  nor2s1 ______443615(.DIN1 (______9__30537), .DIN2 (_____0___30458),
       .Q (__9__0__26459));
  nnd2s1 ____0_443616(.DIN1 (_____9__26126), .DIN2 (__9_0___26424), .Q
       (__9_0___26518));
  nor2s1 _______443617(.DIN1 (_______________18874), .DIN2
       (_____0___30458), .Q (__9_____26546));
  nor2s1 ____9_443618(.DIN1 (_____0__26107), .DIN2 (___9____26181), .Q
       (____9_9__30888));
  nnd2s1 _______443619(.DIN1 (________26109), .DIN2 (__909___26328), .Q
       (__9_____26542));
  dffacs1 _________________443620(.CLRB (reset), .CLK (clk), .DIN
       (________26129), .Q (____________));
  nor2s1 ____9__443621(.DIN1 (__9090), .DIN2 (________26073), .Q
       (__909_));
  nnd2s1 _______443622(.DIN1 (________26098), .DIN2 (__9_____26469), .Q
       (__90_9__26327));
  nnd2s1 ______443623(.DIN1 (_____9__26096), .DIN2 (____9___25555), .Q
       (__90____26326));
  nnd2s1 ______443624(.DIN1 (_____0__26097), .DIN2 (___9____23358), .Q
       (__90____26325));
  nor2s1 ____0__443625(.DIN1 (__9_____26381), .DIN2 (____9___26038), .Q
       (__90____26324));
  nnd2s1 _______443626(.DIN1 (________26091), .DIN2 (________25923), .Q
       (__90____26323));
  nor2s1 ______443627(.DIN1 (_____0__25694), .DIN2 (________26082), .Q
       (__90____26322));
  nnd2s1 ______443628(.DIN1 (________26075), .DIN2 (________24865), .Q
       (__90____26321));
  nor2s1 ______443629(.DIN1 (________25913), .DIN2 (________26100), .Q
       (__90____26320));
  or2s1 _______443630(.DIN1 (__90_0__26318), .DIN2 (________26083), .Q
       (__90____26319));
  nnd2s1 _______443631(.DIN1 (________26085), .DIN2 (___9____26223), .Q
       (__90_9__26317));
  nor2s1 _______443632(.DIN1 (__9_____26621), .DIN2 (__90____26315), .Q
       (__90____26316));
  nor2s1 ____0_443633(.DIN1 (__9_____26452), .DIN2 (_____9__26036), .Q
       (__90____26314));
  nor2s1 _____9_443634(.DIN1 (__90____26312), .DIN2 (________26105), .Q
       (__90____26313));
  and2s1 _____9_443635(.DIN1 (________26090), .DIN2 (__90____26310), .Q
       (__90____26311));
  nor2s1 ____9__443636(.DIN1 (__90_9__26308), .DIN2 (________26078), .Q
       (__90_0__26309));
  nnd2s1 ____9_443637(.DIN1 (________26088), .DIN2 (__90____26306), .Q
       (__90____26307));
  nnd2s1 ____9__443638(.DIN1 (________26102), .DIN2 (________21886), .Q
       (__90____26305));
  nnd2s1 ____9__443639(.DIN1 (_____0__26067), .DIN2 (________24726), .Q
       (__90____26304));
  nnd2s1 ____9__443640(.DIN1 (________26095), .DIN2 (____9___25742), .Q
       (__90____26303));
  and2s1 ____9__443641(.DIN1 (________26069), .DIN2 (_________35074),
       .Q (__90____26302));
  nnd2s1 ____9_443642(.DIN1 (________26093), .DIN2 (________26074), .Q
       (__90____26301));
  nor2s1 _______443643(.DIN1 (________24171), .DIN2 (_____0__26087), .Q
       (__90_0__26300));
  nnd2s1 ____9__443644(.DIN1 (_____9__26066), .DIN2 (________21469), .Q
       (__90_9__26299));
  nnd2s1 ____9_443645(.DIN1 (________26065), .DIN2 (__9__9__26540), .Q
       (__90____26298));
  nnd2s1 ____9__443646(.DIN1 (_____9__26026), .DIN2 (________25627), .Q
       (__90____26296));
  nnd2s1 ____9__443647(.DIN1 (_____0__26027), .DIN2 (________25419), .Q
       (__90____26295));
  nnd2s1 ____9_443648(.DIN1 (____0___26054), .DIN2 (________26068), .Q
       (__90____26294));
  nnd2s1 ____99_443649(.DIN1 (____0___26052), .DIN2 (___0__9__27839),
       .Q (__90____26293));
  nnd2s1 ____99_443650(.DIN1 (____0___26051), .DIN2 (__90_0__26291), .Q
       (__90____26292));
  nnd2s1 ____99_443651(.DIN1 (________26022), .DIN2 (____0___25661), .Q
       (__90_9__26290));
  and2s1 ____00_443652(.DIN1 (___9_0__26227), .DIN2 (outData[9]), .Q
       (__90____26289));
  nor2s1 ____0_443653(.DIN1 (________23700), .DIN2 (____9___26045), .Q
       (__90____26288));
  nor2s1 ____0__443654(.DIN1 (__990___27084), .DIN2 (__90____26286), .Q
       (__90____26287));
  nor2s1 ____0__443655(.DIN1 (__9_____26499), .DIN2 (________26035), .Q
       (__90____26285));
  nor2s1 ____0__443656(.DIN1 (________23185), .DIN2 (________26061), .Q
       (__90____26284));
  nor2s1 ____0__443657(.DIN1 (________25812), .DIN2 (_____0__26017), .Q
       (__90____26283));
  nor2s1 ____0__443658(.DIN1 (__90_0__26281), .DIN2 (________26080), .Q
       (__90____26282));
  or2s1 ____0__443659(.DIN1 (__9_____26647), .DIN2 (____9___26040), .Q
       (__90_9__26280));
  nor2s1 ____0_443660(.DIN1 (_____9__24847), .DIN2 (________26015), .Q
       (__90____26279));
  nor2s1 ____0_443661(.DIN1 (________24563), .DIN2 (____9___26039), .Q
       (__90____26278));
  nnd2s1 ____0__443662(.DIN1 (________26060), .DIN2 (___9____22495), .Q
       (__90____26277));
  nor2s1 ____0_443663(.DIN1 (__90____26275), .DIN2 (________26058), .Q
       (__90____26276));
  nnd2s1 ______443664(.DIN1 (_____9__26086), .DIN2 (__9_____26389), .Q
       (__9_9___26418));
  dffacs1 _________________443665(.CLRB (reset), .CLK (clk), .DIN
       (____0___26050), .QN (______________18871));
  and2s1 _______443666(.DIN1 (________26021), .DIN2 (__90____26273), .Q
       (__90____26274));
  nnd2s1 ____0__443667(.DIN1 (_____9__26016), .DIN2 (__90_0__26271), .Q
       (__90____26272));
  nor2s1 _______443668(.DIN1 (_________34409), .DIN2 (______9__30537),
       .Q (__90_9__26270));
  nor2s1 _______443669(.DIN1 (__90____26268), .DIN2 (__90____26267), .Q
       (__90____26269));
  or2s1 ______443670(.DIN1 (__90____26265), .DIN2 (________26033), .Q
       (__90____26266));
  nnd2s1 _______443671(.DIN1 (_________33174), .DIN2 (_________34409),
       .Q (__90____26264));
  nor2s1 ____0__443672(.DIN1 (__90____26262), .DIN2 (____0___26048), .Q
       (__90____26263));
  or2s1 ____0__443673(.DIN1 (__90_9), .DIN2 (________26034), .Q
       (__90_0__26261));
  nnd2s1 ____0__443674(.DIN1 (________26108), .DIN2 (outData[9]), .Q
       (__90____26260));
  nor2s1 ____0__443675(.DIN1 (__90____26258), .DIN2 (____9___26044), .Q
       (__90____26259));
  nor2s1 ____0_443676(.DIN1 (________25137), .DIN2 (____09__26056), .Q
       (__90____26257));
  nnd2s1 ____0__443677(.DIN1 (_________29253), .DIN2
       (______________18869), .Q (__90____26256));
  nor2s1 ____0__443678(.DIN1 (___9____26194), .DIN2 (________26023), .Q
       (__90____26255));
  nor2s1 ____09_443679(.DIN1 (___9_9__23404), .DIN2 (________26011), .Q
       (__90____26254));
  or2s1 ____443680(.DIN1 (__90_0), .DIN2 (________26030), .Q (__90__));
  nnd2s1 _____443681(.DIN1 (________26029), .DIN2 (________22946), .Q
       (__9009));
  nnd2s1 _____0_443682(.DIN1
       (______________________________________0__________0__18892),
       .DIN2 (_________29253), .Q (__900___26253));
  nor2s1 _____0_443683(.DIN1
       (______________________________________0__________0__18892),
       .DIN2 (_________29253), .Q (__900___26252));
  nor2s1 _______443684(.DIN1 (___00____27202), .DIN2 (____90__26037),
       .Q (__900___26251));
  nor2s1 ______443685(.DIN1 (_____9__24446), .DIN2 (________26025), .Q
       (__900___26250));
  or2s1 _______443686(.DIN1 (__9_____26487), .DIN2 (________26013), .Q
       (__900___26249));
  nnd2s1 _______443687(.DIN1 (____9___26041), .DIN2 (____0___25752), .Q
       (__900___26248));
  and2s1 _______443688(.DIN1 (________26010), .DIN2 (__900_), .Q
       (__900___26247));
  and2s1 ____0__443689(.DIN1 (____9___26042), .DIN2 (___999__26246), .Q
       (__9000));
  nnd2s1 _______443690(.DIN1 (________26012), .DIN2 (__9_____26576), .Q
       (___99___26245));
  nor2s1 ______443691(.DIN1 (_________29253), .DIN2
       (_________________0___18660), .Q (___99___26244));
  nnd2s1 _______443692(.DIN1 (________26019), .DIN2 (___99___26242), .Q
       (___99___26243));
  nnd2s1 _______443693(.DIN1 (________26009), .DIN2 (__9_____26962), .Q
       (___99___26241));
  nnd2s1 _______443694(.DIN1 (___9____26231), .DIN2 (________25112), .Q
       (___99___26240));
  nor2s1 _______443695(.DIN1 (____0____30075), .DIN2 (_________29253),
       .Q (___99___26239));
  hi1s1 _______443696(.DIN (__9_0___26801), .Q (___99___26238));
  nnd2s1 _______443697(.DIN1 (________26001), .DIN2 (___9____26230), .Q
       (___990__26237));
  nnd2s1 _____9_443698(.DIN1 (________25998), .DIN2 (___9____26235), .Q
       (___9_9__26236));
  nor2s1 _____443699(.DIN1 (____0___21992), .DIN2 (________26004), .Q
       (___9____26234));
  nor2s1 _____9_443700(.DIN1 (________24855), .DIN2 (________26031), .Q
       (___9____26233));
  nor2s1 _______443701(.DIN1 (__9_____26621), .DIN2 (___9____26231), .Q
       (___9____26232));
  nnd2s1 ____0__443702(.DIN1 (____0___26049), .DIN2 (___9____26230), .Q
       (__9_____26470));
  nnd2s1 _______443703(.DIN1 (________26028), .DIN2 (________25762), .Q
       (___0_____27933));
  nor2s1 ____0_443704(.DIN1 (_________9______18799), .DIN2
       (_________29253), .Q (__9_____26342));
  nor2s1 _______443705(.DIN1 (_________34409), .DIN2 (_________31058),
       .Q (__9_____26343));
  and2s1 ____0__443706(.DIN1 (_________29253), .DIN2
       (_________9______18799), .Q (__9_0___26421));
  nor2s1 _______443707(.DIN1 (____9____29052), .DIN2 (_________29253),
       .Q (__9_____26432));
  nor2s1 _______443708(.DIN1 (_________34409), .DIN2
       (______________________________________0_____________18891), .Q
       (__9_0___26516));
  nor2s1 _______443709(.DIN1 (_________34409), .DIN2 (____0____30075),
       .Q (__9_____26545));
  nnd2s1 _______443710(.DIN1 (___9____26229), .DIN2 (___9____26228), .Q
       (___0_____27607));
  nor2s1 _______443711(.DIN1 (_____9__25879), .DIN2 (__9__9__26531), .Q
       (__9_0___26703));
  nor2s1 ____0__443712(.DIN1 (outData[9]), .DIN2 (___9_0__26227), .Q
       (__9_0___26423));
  nnd2s1 ____0__443713(.DIN1 (____0___25952), .DIN2 (____9___21899), .Q
       (___9_9__26226));
  nor2s1 _______443714(.DIN1 (___9_0__26207), .DIN2 (_____0__25957), .Q
       (___9____26225));
  and2s1 ____9__443715(.DIN1 (________25930), .DIN2 (___9____26223), .Q
       (___9____26224));
  nor2s1 ____9_443716(.DIN1 (________25985), .DIN2 (________25992), .Q
       (___9____26222));
  nnd2s1 ____9_443717(.DIN1 (________25984), .DIN2 (___9____26220), .Q
       (___9____26221));
  nnd2s1 ____9__443718(.DIN1 (____0___25951), .DIN2 (___9____26218), .Q
       (___9____26219));
  or2s1 ____9__443719(.DIN1 (______0__28551), .DIN2 (____0___25950), .Q
       (___9_0__26217));
  nor2s1 ____9__443720(.DIN1 (___9____26215), .DIN2 (________25988), .Q
       (___9_9__26216));
  or2s1 ____9__443721(.DIN1 (___9____26213), .DIN2 (____9___25941), .Q
       (___9____26214));
  nnd2s1 ____99_443722(.DIN1 (________25981), .DIN2 (__9_____26623), .Q
       (___9____26212));
  nnd2s1 ____443723(.DIN1 (________25993), .DIN2 (________25394), .Q
       (___9____26211));
  or2s1 ____00_443724(.DIN1 (___9____26209), .DIN2 (____9___25944), .Q
       (___9____26210));
  nor2s1 ____00_443725(.DIN1 (___9_0__26207), .DIN2 (_____9__25908), .Q
       (___9____26208));
  nnd2s1 ____00_443726(.DIN1 (________25979), .DIN2 (________25132), .Q
       (___9_9__26206));
  and2s1 ____00_443727(.DIN1 (________25917), .DIN2 (________25162), .Q
       (___9____26205));
  nnd2s1 ____443728(.DIN1 (________25936), .DIN2 (________22739), .Q
       (___9____26204));
  nnd2s1 ____0__443729(.DIN1 (________25969), .DIN2 (________25973), .Q
       (___9____26203));
  nor2s1 ____0__443730(.DIN1 (__9_____27023), .DIN2 (________25968), .Q
       (___9____26202));
  and2s1 ____0__443731(.DIN1 (________25965), .DIN2 (___9____26200), .Q
       (___9____26201));
  nor2s1 ____0__443732(.DIN1 (__90_0__26318), .DIN2 (____9___25942), .Q
       (___9____26199));
  nor2s1 ____0__443733(.DIN1 (________25910), .DIN2 (________25994), .Q
       (___9____26198));
  and2s1 ____0__443734(.DIN1 (____0___25955), .DIN2 (________24502), .Q
       (___9_0__26197));
  nnd2s1 ____0__443735(.DIN1 (________25975), .DIN2 (___9_0__26177), .Q
       (___9_9__26196));
  nor2s1 ____0__443736(.DIN1 (___9____26194), .DIN2 (____0___25954), .Q
       (___9____26195));
  nnd2s1 ____0_443737(.DIN1 (________20193), .DIN2 (_____0__25909), .Q
       (___9____26193));
  nnd2s1 _______443738(.DIN1 (________25920), .DIN2 (____9___26043), .Q
       (___9____26192));
  nnd2s1 ____0__443739(.DIN1 (________25974), .DIN2 (________23140), .Q
       (___9____26191));
  nor2s1 ____0__443740(.DIN1 (_____9__25684), .DIN2 (________25990), .Q
       (___9____26190));
  nnd2s1 ____0__443741(.DIN1 (________25765), .DIN2 (________25962), .Q
       (___9____26189));
  nor2s1 ____0__443742(.DIN1 (__9_0___26897), .DIN2 (_____0__25987), .Q
       (___9____26188));
  and2s1 ____0_443743(.DIN1 (____0___25949), .DIN2 (__9_____26840), .Q
       (___9_0__26187));
  nnd2s1 ____0__443744(.DIN1 (_____9__25986), .DIN2 (________25861), .Q
       (___9_9__26186));
  nor2s1 ____0__443745(.DIN1 (_____0__23860), .DIN2 (____9___25946), .Q
       (___9____26185));
  nor2s1 _______443746(.DIN1 (________22146), .DIN2 (____9___25940), .Q
       (___9____26184));
  nor2s1 ____0__443747(.DIN1 (___9____26182), .DIN2 (_____9__25966), .Q
       (___9____26183));
  xor2s1 ____0__443748(.DIN1 (________25792), .DIN2 (_________31667),
       .Q (___9____26181));
  or2s1 ____0__443749(.DIN1 (___9____26179), .DIN2 (_____0__25919), .Q
       (___9____26180));
  and2s1 ____0__443750(.DIN1 (________25912), .DIN2 (___9_0__26177), .Q
       (___9____26178));
  nnd2s1 ____0__443751(.DIN1 (__________9_), .DIN2 (_________28866), .Q
       (___9_9__26176));
  nnd2s1 ____0_443752(.DIN1 (____99__25947), .DIN2 (___9____26174), .Q
       (___9____26175));
  nnd2s1 ____443753(.DIN1 (________25982), .DIN2 (__9_____26877), .Q
       (___9____26173));
  or2s1 ____09_443754(.DIN1 (___9____26171), .DIN2 (_____0__25929), .Q
       (___9____26172));
  nnd2s1 ____09_443755(.DIN1 (________25906), .DIN2 (____9___25552), .Q
       (___9____26170));
  nnd2s1 _____0_443756(.DIN1 (___0____25302), .DIN2 (________25925), .Q
       (___9____26169));
  nor2s1 _____443757(.DIN1 (___9_0__26167), .DIN2 (________25927), .Q
       (___9____26168));
  nor2s1 ______443758(.DIN1 (__________9_), .DIN2 (________25489), .Q
       (___9_9__26166));
  nor2s1 _______443759(.DIN1 (____0___22992), .DIN2 (________25972), .Q
       (___9____26165));
  and2s1 _______443760(.DIN1 (____0___25953), .DIN2 (___9____26163), .Q
       (___9____26164));
  nor2s1 ____0__443761(.DIN1 (__9_____26632), .DIN2 (________25961), .Q
       (__90____26297));
  dffacs1 __________________443762(.CLRB (reset), .CLK (clk), .DIN
       (_____9__25976), .QN (_______________18873));
  nnd2s1 _______443763(.DIN1 (_____9__25889), .DIN2 (____0___25754), .Q
       (___9____26162));
  or2s1 ______443764(.DIN1 (__9_____26838), .DIN2 (________25924), .Q
       (___9____26161));
  and2s1 _______443765(.DIN1 (________25902), .DIN2 (___9____26159), .Q
       (___9____26160));
  nor2s1 _______443766(.DIN1 (___9_0__26157), .DIN2 (________25937), .Q
       (___9____26158));
  nnd2s1 _______443767(.DIN1 (________25970), .DIN2 (________25444), .Q
       (___909__26156));
  or2s1 _______443768(.DIN1 (___90___26154), .DIN2 (________25900), .Q
       (___90___26155));
  nnd2s1 _______443769(.DIN1 (________25964), .DIN2 (_____0__26077), .Q
       (___90___26153));
  and2s1 ______443770(.DIN1 (________25903), .DIN2 (___90___26151), .Q
       (___90___26152));
  nnd2s1 _______443771(.DIN1 (________25911), .DIN2 (__9_____26862), .Q
       (___90___26150));
  nor2s1 _______443772(.DIN1 (_____9__21884), .DIN2 (________25904), .Q
       (___90___26149));
  nnd2s1 _______443773(.DIN1 (________25915), .DIN2 (___900__26147), .Q
       (___90___26148));
  and2s1 _______443774(.DIN1 (____0____28174), .DIN2 (________25423),
       .Q (____99__26146));
  or2s1 _______443775(.DIN1 (____9___26144), .DIN2 (________25916), .Q
       (____9___26145));
  nor2s1 _______443776(.DIN1 (____9___26142), .DIN2 (_____0__25899), .Q
       (____9___26143));
  or2s1 _______443777(.DIN1 (___0_____27430), .DIN2 (_________34782),
       .Q (____9___26141));
  or2s1 _______443778(.DIN1 (________25422), .DIN2 (____0____28174), .Q
       (____9___26140));
  nnd2s1 _______443779(.DIN1 (________25931), .DIN2
       (______________________________________0_____________18886), .Q
       (____9___26139));
  nor2s1 ______443780(.DIN1 (____90__26137), .DIN2 (_____0__25890), .Q
       (____9___26138));
  nor2s1 _______443781(.DIN1 (___9____25226), .DIN2 (_____0__25860), .Q
       (_____9__26136));
  nor2s1 _______443782(.DIN1 (___0____22571), .DIN2 (________25882), .Q
       (________26135));
  nnd2s1 _____0_443783(.DIN1 (________25868), .DIN2 (_____9__25674), .Q
       (________26134));
  nnd2s1 _____9_443784(.DIN1 (________25863), .DIN2 (__9_____26525), .Q
       (________26133));
  nor2s1 _______443785(.DIN1 (_____0__26117), .DIN2 (____09__25859), .Q
       (________26132));
  nor2s1 _______443786(.DIN1 (________26130), .DIN2 (________25891), .Q
       (________26131));
  nnd2s1 _______443787(.DIN1 (________25893), .DIN2 (________24532), .Q
       (________26129));
  nor2s1 _______443788(.DIN1 (_____0__26127), .DIN2 (________25914), .Q
       (________26128));
  nor2s1 _____9_443789(.DIN1 (________26125), .DIN2 (________25867), .Q
       (_____9__26126));
  and2s1 _____443790(.DIN1 (________25884), .DIN2 (________26123), .Q
       (________26124));
  nnd2s1 _____443791(.DIN1 (________25873), .DIN2 (________26121), .Q
       (________26122));
  nnd2s1 _______443792(.DIN1 (_____9__25869), .DIN2 (_____9__25528), .Q
       (________26120));
  nnd2s1 _______443793(.DIN1 (________25862), .DIN2 (___9____26218), .Q
       (________26119));
  nor2s1 _______443794(.DIN1 (_____0__26117), .DIN2 (________25892), .Q
       (________26118));
  nor2s1 _______443795(.DIN1 (___0_____27698), .DIN2 (________25875),
       .Q (_____9__26116));
  or2s1 _______443796(.DIN1 (________26081), .DIN2 (_____0__25880), .Q
       (________26115));
  nnd2s1 _______443797(.DIN1 (________25876), .DIN2 (________25806), .Q
       (________26114));
  nnd2s1 _______443798(.DIN1 (________25865), .DIN2 (__9_____26370), .Q
       (________26113));
  and2s1 _______443799(.DIN1 (________25888), .DIN2 (__9_____27045), .Q
       (________26112));
  nnd2s1 _______443800(.DIN1 (________25871), .DIN2 (________22870), .Q
       (________26111));
  nor2s1 _______443801(.DIN1 (____9___22440), .DIN2 (________25886), .Q
       (________26110));
  hi1s1 _______443802(.DIN (________26108), .Q (________26109));
  nor2s1 ______443803(.DIN1 (__________9_), .DIN2
       (_______________18874), .Q (__9_____26732));
  nor2s1 _______443804(.DIN1 (__________9_), .DIN2
       (______________18871), .Q (__9_____26431));
  nor2s1 ______443805(.DIN1 (________25107), .DIN2 (____0____28174), .Q
       (__909___26329));
  nnd2s1 ______443806(.DIN1 (__________9_), .DIN2
       (___________0___18872), .Q (__9__9__26384));
  xnr2s1 _______443807(.DIN1 (outData[8]), .DIN2 (_____9__25996), .Q
       (___0_____27475));
  nnd2s1 _______443808(.DIN1 (________25883), .DIN2
       (______________________________________0___________), .Q
       (__9_0___26801));
  xor2s1 _______443809(.DIN1 (outData[8]), .DIN2 (_____0__26107), .Q
       (____9____29056));
  hi1s1 ______443810(.DIN (_____9__26106), .Q (_____0___28530));
  dffacs1 __________________443811(.CLRB (reset), .CLK (clk), .DIN
       (_____0__25977), .QN (_______________18880));
  hi1s1 ______443812(.DIN (_________34409), .Q (_____0___30458));
  and2s1 _____0_443813(.DIN1 (____0___25856), .DIN2 (__9_____26631), .Q
       (________26105));
  nor2s1 ____9__443814(.DIN1 (__990___27084), .DIN2 (________26103), .Q
       (________26104));
  or2s1 ____9__443815(.DIN1 (________26101), .DIN2 (________25834), .Q
       (________26102));
  nnd2s1 ____443816(.DIN1 (____9___25844), .DIN2 (________26099), .Q
       (________26100));
  nnd2s1 ____99_443817(.DIN1 (____0___25852), .DIN2 (_____9___28891),
       .Q (________26098));
  nnd2s1 ____99_443818(.DIN1 (________25827), .DIN2 (inData[18]), .Q
       (_____0__26097));
  nnd2s1 ____443819(.DIN1 (____00__25850), .DIN2 (___0____21654), .Q
       (_____9__26096));
  nor2s1 ____00_443820(.DIN1 (________26094), .DIN2 (________25825), .Q
       (________26095));
  nor2s1 ____00_443821(.DIN1 (________26092), .DIN2 (________25826), .Q
       (________26093));
  nor2s1 ____0__443822(.DIN1 (___0_9___27848), .DIN2 (____9___25848),
       .Q (________26091));
  and2s1 ____0_443823(.DIN1 (____9___25845), .DIN2 (________26089), .Q
       (________26090));
  nor2s1 ____0_443824(.DIN1 (___9_0__25241), .DIN2 (____9___25843), .Q
       (________26088));
  nnd2s1 ____0__443825(.DIN1 (____9___25842), .DIN2 (__9_____26877), .Q
       (_____0__26087));
  nor2s1 ____0__443826(.DIN1 (________25513), .DIN2 (____9___25841), .Q
       (_____9__26086));
  and2s1 ____0__443827(.DIN1 (_____9__25839), .DIN2 (________26084), .Q
       (________26085));
  or2s1 ____0__443828(.DIN1 (__9_____26905), .DIN2 (________25837), .Q
       (________26083));
  or2s1 ____0__443829(.DIN1 (________26081), .DIN2 (____0___25855), .Q
       (________26082));
  nnd2s1 _______443830(.DIN1 (________25805), .DIN2 (________26079), .Q
       (________26080));
  nnd2s1 ____0_443831(.DIN1 (________25832), .DIN2 (_____0__26077), .Q
       (________26078));
  nor2s1 ____0_443832(.DIN1 (__9_____26953), .DIN2 (________25838), .Q
       (_____9__26076));
  and2s1 ____0__443833(.DIN1 (________25833), .DIN2 (________26074), .Q
       (________26075));
  or2s1 ____0__443834(.DIN1 (________26072), .DIN2 (____0___25854), .Q
       (________26073));
  xor2s1 _____0_443835(.DIN1 (________26070), .DIN2
       (_______________18878), .Q (________26071));
  dffacs2 _____________________0_443836(.CLRB (reset), .CLK (clk), .DIN
       (________25821), .QN (_________________0___18633));
  and2s1 _____0_443837(.DIN1 (________25823), .DIN2 (________26068), .Q
       (________26069));
  and2s1 _______443838(.DIN1 (_____0__25830), .DIN2 (__90____26310), .Q
       (_____0__26067));
  or2s1 _______443839(.DIN1 (__90____26258), .DIN2 (____9___25847), .Q
       (_____9__26066));
  nor2s1 _______443840(.DIN1 (________25980), .DIN2 (____0___25851), .Q
       (________26065));
  xor2s1 ______443841(.DIN1
       (______________________________________0_____________18889),
       .DIN2 (_______________18878), .Q (________26064));
  xnr2s1 _______443842(.DIN1 (________26062), .DIN2 (______0__29851),
       .Q (________26063));
  nnd2s1 _______443843(.DIN1 (________25802), .DIN2 (____0___22997), .Q
       (________26061));
  and2s1 ______443844(.DIN1 (________25816), .DIN2 (________26059), .Q
       (________26060));
  or2s1 _______443845(.DIN1 (_____0__26057), .DIN2 (________25811), .Q
       (________26058));
  or2s1 _______443846(.DIN1 (____0___26055), .DIN2 (________25794), .Q
       (____09__26056));
  nor2s1 ______443847(.DIN1 (____0___26053), .DIN2 (_____9__25809), .Q
       (____0___26054));
  nor2s1 _______443848(.DIN1 (___0_____27711), .DIN2 (________25808),
       .Q (____0___26052));
  and2s1 _______443849(.DIN1 (_____0__25810), .DIN2 (________23295), .Q
       (____0___26051));
  nnd2s1 _____443850(.DIN1 (________25788), .DIN2 (________23650), .Q
       (____0___26050));
  nor2s1 _____9_443851(.DIN1 (___0____25354), .DIN2 (________25818), .Q
       (____0___26049));
  nnd2s1 _____9_443852(.DIN1 (________25815), .DIN2 (____0___23529), .Q
       (____0___26048));
  nor2s1 _____9_443853(.DIN1 (_____0___28805), .DIN2 (____99__26046),
       .Q (____00__26047));
  nnd2s1 _____0_443854(.DIN1 (_____9__25819), .DIN2 (_____0__22108), .Q
       (____9___26045));
  nnd2s1 _____0_443855(.DIN1 (________25828), .DIN2 (____9___26043), .Q
       (____9___26044));
  and2s1 _______443856(.DIN1 (________25777), .DIN2 (_____0__23811), .Q
       (____9___26042));
  nor2s1 ____0__443857(.DIN1 (_____0__25997), .DIN2 (________25835), .Q
       (__90____26315));
  hi1s1 _______443858(.DIN (__________9_), .Q (_________29253));
  nor2s1 _______443859(.DIN1 (___990__25261), .DIN2 (________25763), .Q
       (____9___26041));
  or2s1 _______443860(.DIN1 (________23318), .DIN2 (________25795), .Q
       (____9___26040));
  or2s1 ______443861(.DIN1 (________26008), .DIN2 (________25783), .Q
       (____9___26039));
  nnd2s1 _______443862(.DIN1 (________25813), .DIN2 (__9__0__26739), .Q
       (____9___26038));
  nor2s1 ______443863(.DIN1 (________23556), .DIN2 (________25796), .Q
       (____90__26037));
  or2s1 _______443864(.DIN1 (_____9__25001), .DIN2 (_____9__25799), .Q
       (_____9__26036));
  nnd2s1 _______443865(.DIN1 (_____0__25780), .DIN2 (_____90__34918),
       .Q (________26035));
  nnd2s1 ______443866(.DIN1 (_____0__25800), .DIN2 (________26121), .Q
       (________26034));
  or2s1 _______443867(.DIN1 (________26032), .DIN2 (________25791), .Q
       (________26033));
  nnd2s1 _______443868(.DIN1 (____00__25751), .DIN2 (___0____23484), .Q
       (________26031));
  nnd2s1 _______443869(.DIN1 (________25786), .DIN2 (_____0__25520), .Q
       (________26030));
  nor2s1 _______443870(.DIN1 (________25793), .DIN2 (________25773), .Q
       (________26029));
  nnd2s1 _______443871(.DIN1 (________25766), .DIN2 (outData[7]), .Q
       (________26028));
  nor2s1 _______443872(.DIN1 (________25978), .DIN2 (________25781), .Q
       (_____0__26027));
  and2s1 _______443873(.DIN1 (________26014), .DIN2 (____99__23345), .Q
       (_____9__26026));
  nnd2s1 _______443874(.DIN1 (________25778), .DIN2 (___0_____27527),
       .Q (________26025));
  nnd2s1 _____9_443875(.DIN1 (________25934), .DIN2 (_________31058),
       .Q (________26024));
  nnd2s1 _____9_443876(.DIN1 (_____9__25779), .DIN2 (__9_____26389), .Q
       (________26023));
  nor2s1 _____443877(.DIN1 (________23104), .DIN2 (________25804), .Q
       (________26022));
  and2s1 _____0_443878(.DIN1 (________25807), .DIN2 (________26020), .Q
       (________26021));
  and2s1 _______443879(.DIN1 (________25776), .DIN2 (________26018), .Q
       (________26019));
  or2s1 _______443880(.DIN1 (__9_____26499), .DIN2 (________25771), .Q
       (_____0__26017));
  nor2s1 _______443881(.DIN1 (___0____24412), .DIN2 (________25787), .Q
       (_____9__26016));
  nnd2s1 _______443882(.DIN1 (________26014), .DIN2 (_____9__25606), .Q
       (________26015));
  or2s1 _______443883(.DIN1 (________26130), .DIN2 (________25785), .Q
       (________26013));
  nnd2s1 ______443884(.DIN1 (________25768), .DIN2 (___900__26147), .Q
       (________26012));
  nnd2s1 _______443885(.DIN1 (________25764), .DIN2 (________22647), .Q
       (________26011));
  nor2s1 _______443886(.DIN1 (_____0__23591), .DIN2 (________25784), .Q
       (________26010));
  or2s1 ______443887(.DIN1 (________26008), .DIN2 (____0___25753), .Q
       (________26009));
  nor2s1 _______443888(.DIN1 (_____9__26006), .DIN2 (_________31058),
       .Q (_____0__26007));
  xor2s1 _______443889(.DIN1 (_____9___34515), .DIN2 (_________31060),
       .Q (________26005));
  nnd2s1 _______443890(.DIN1 (____0___25757), .DIN2 (________22954), .Q
       (________26004));
  nnd2s1 _______443891(.DIN1
       (______________0______________________18828), .DIN2
       (________26002), .Q (________26003));
  nor2s1 _____443892(.DIN1 (________26000), .DIN2 (____0___25756), .Q
       (________26001));
  nor2s1 _____0_443893(.DIN1 (________26002), .DIN2 (____0___22994), .Q
       (________25999));
  and2s1 _______443894(.DIN1 (____0___25755), .DIN2 (__90_0__26291), .Q
       (________25998));
  nnd2s1 _______443895(.DIN1 (_________28661), .DIN2 (________26002),
       .Q (___9____26229));
  xnr2s1 ______443896(.DIN1 (_____0__25870), .DIN2 (________22871), .Q
       (_____9__26106));
  nnd2s1 _______443897(.DIN1 (_____0__26107), .DIN2 (________25995), .Q
       (________26108));
  nor2s1 _______443898(.DIN1 (__9__0__26485), .DIN2 (________25775), .Q
       (__90____26286));
  nor2s1 _______443899(.DIN1 (_____0__25997), .DIN2 (_________34784),
       .Q (___9____26231));
  nor2s1 ______443900(.DIN1 (________26002), .DIN2
       (______________18870), .Q (__90____26268));
  nnd2s1 _______443901(.DIN1 (_____9__25996), .DIN2 (________25995), .Q
       (___9_0__26227));
  xor2s1 _______443902(.DIN1 (________25681), .DIN2 (_________30166),
       .Q (_____0___28617));
  nor2s1 _______443903(.DIN1 (___0_____27914), .DIN2 (________26002),
       .Q (__9__9__26531));
  dffacs2 __________________443904(.CLRB (reset), .CLK (clk), .DIN
       (____0___25759), .Q (_________34409));
  nnd2s1 _______443905(.DIN1 (________25716), .DIN2 (__9_____26389), .Q
       (________25994));
  nor2s1 _______443906(.DIN1 (____9___25458), .DIN2 (_____0__25675), .Q
       (________25993));
  nnd2s1 _______443907(.DIN1 (_____9__25730), .DIN2 (________25991), .Q
       (________25992));
  or2s1 _______443908(.DIN1 (________25989), .DIN2 (________25705), .Q
       (________25990));
  nnd2s1 ______443909(.DIN1 (_____9__25702), .DIN2 (____00__24792), .Q
       (________25988));
  nnd2s1 _______443910(.DIN1 (____9___25744), .DIN2 (___0_9__21666), .Q
       (_____0__25987));
  nor2s1 _______443911(.DIN1 (________25985), .DIN2 (________25738), .Q
       (_____9__25986));
  nor2s1 ______443912(.DIN1 (________25983), .DIN2 (________25737), .Q
       (________25984));
  nor2s1 _______443913(.DIN1 (__9_____26743), .DIN2 (________25735), .Q
       (________25982));
  nor2s1 _______443914(.DIN1 (________25980), .DIN2 (________25733), .Q
       (________25981));
  nor2s1 _______443915(.DIN1 (________25978), .DIN2 (____9___25745), .Q
       (________25979));
  nnd2s1 _____9_443916(.DIN1 (________25688), .DIN2 (___9_0__23366), .Q
       (_____0__25977));
  nnd2s1 _____9_443917(.DIN1 (_____0__25731), .DIN2 (_________34800),
       .Q (_____9__25976));
  nor2s1 _____0_443918(.DIN1 (____9___23255), .DIN2 (________25708), .Q
       (________25975));
  and2s1 _____0_443919(.DIN1 (________25727), .DIN2 (________25973), .Q
       (________25974));
  nnd2s1 _____0_443920(.DIN1 (_____9__25740), .DIN2 (________22955), .Q
       (________25972));
  nor2s1 ______443921(.DIN1 (________25725), .DIN2 (____0___25657), .Q
       (________25971));
  nor2s1 _______443922(.DIN1 (____0____34554), .DIN2 (________25736),
       .Q (________25970));
  nor2s1 _______443923(.DIN1 (_____9__25145), .DIN2 (________25724), .Q
       (________25969));
  or2s1 _______443924(.DIN1 (_____0__25967), .DIN2 (_____0__25721), .Q
       (________25968));
  or2s1 _______443925(.DIN1 (________26072), .DIN2 (_____9__25720), .Q
       (_____9__25966));
  and2s1 ______443926(.DIN1 (________25695), .DIN2 (____0___23173), .Q
       (________25965));
  nor2s1 _______443927(.DIN1 (________25963), .DIN2 (________25719), .Q
       (________25964));
  and2s1 _______443928(.DIN1 (______0__34788), .DIN2 (_____9__24007),
       .Q (________25962));
  nnd2s1 ______443929(.DIN1 (________25698), .DIN2 (__90_0__26271), .Q
       (________25961));
  and2s1 ______443930(.DIN1 (________25959), .DIN2 (_________28788), .Q
       (________25960));
  nor2s1 _______443931(.DIN1 (_________28788), .DIN2 (________25959),
       .Q (________25958));
  nnd2s1 ______443932(.DIN1 (____9___25747), .DIN2 (___9____22463), .Q
       (_____0__25957));
  nnd2s1 _______443933(.DIN1 (________25714), .DIN2 (__9_____27061), .Q
       (____09__25956));
  nor2s1 ______443934(.DIN1 (________24501), .DIN2 (________25617), .Q
       (____0___25955));
  nnd2s1 _______443935(.DIN1 (_________34786), .DIN2 (________22945),
       .Q (____0___25954));
  nor2s1 _______443936(.DIN1 (____9___23163), .DIN2 (________25706), .Q
       (____0___25953));
  nnd2s1 _______443937(.DIN1 (_____0__25703), .DIN2 (__9__0__26494), .Q
       (____0___25952));
  nor2s1 _______443938(.DIN1 (____9___26144), .DIN2 (________25718), .Q
       (____0___25951));
  nnd2s1 _______443939(.DIN1 (______0__34788), .DIN2 (___009__24342),
       .Q (____0___25950));
  and2s1 _______443940(.DIN1 (________25701), .DIN2 (____00__25948), .Q
       (____0___25949));
  nor2s1 _______443941(.DIN1 (____0____34554), .DIN2 (____90__25741),
       .Q (____99__25947));
  or2s1 ______443942(.DIN1 (____9___25945), .DIN2 (_____0__25635), .Q
       (____9___25946));
  or2s1 _____0_443943(.DIN1 (____9___25943), .DIN2 (________25686), .Q
       (____9___25944));
  or2s1 _______443944(.DIN1 (__9_____26831), .DIN2 (________25690), .Q
       (____9___25942));
  nnd2s1 _______443945(.DIN1 (________25669), .DIN2 (________25707), .Q
       (____9___25941));
  nor2s1 ______443946(.DIN1 (____90__25939), .DIN2 (________25691), .Q
       (____9___25940));
  nnd2s1 _______443947(.DIN1 (________25417), .DIN2
       (_______________18878), .Q (_____9__25938));
  nnd2s1 _______443948(.DIN1 (________25682), .DIN2 (___9____23416), .Q
       (________25937));
  nor2s1 ______443949(.DIN1 (___9____25249), .DIN2 (________25671), .Q
       (________25936));
  nor2s1 _____443950(.DIN1 (_______________18878), .DIN2
       (________25934), .Q (________25935));
  nnd2s1 _____9_443951(.DIN1 (________25699), .DIN2 (____9___21899), .Q
       (________25933));
  nnd2s1 _____9_443952(.DIN1 (________25490), .DIN2
       (_______________18878), .Q (________25932));
  and2s1 _____9_443953(.DIN1 (____0____32762), .DIN2
       (_______________18878), .Q (________25931));
  and2s1 _____443954(.DIN1 (________25700), .DIN2 (___9_0__26177), .Q
       (________25930));
  nnd2s1 _____0_443955(.DIN1 (____9___25743), .DIN2 (_____9__25928), .Q
       (_____0__25929));
  nnd2s1 _____0_443956(.DIN1 (________25668), .DIN2 (________25926), .Q
       (________25927));
  nnd2s1 _____0_443957(.DIN1 (________23900), .DIN2 (____9___25748), .Q
       (________25925));
  dffacs1 _______________9_(.CLRB (reset), .CLK (clk), .DIN
       (________25732), .Q (__________9_));
  dffacs1 ________________0_443958(.CLRB (reset), .CLK (clk), .DIN
       (________25633), .QN (___________0___18883));
  nnd2s1 _____0_443959(.DIN1 (________25723), .DIN2 (________25923), .Q
       (________25924));
  nnd2s1 _______443960(.DIN1 (_______________18878), .DIN2
       (_________31281), .Q (________25922));
  nor2s1 _______443961(.DIN1 (_______________18878), .DIN2
       (_________31281), .Q (________25921));
  nor2s1 _______443962(.DIN1 (_____9__23161), .DIN2 (________25678), .Q
       (________25920));
  or2s1 _______443963(.DIN1 (_____9__25918), .DIN2 (________25713), .Q
       (_____0__25919));
  nor2s1 ______443964(.DIN1 (___0_____27698), .DIN2 (________25679), .Q
       (________25917));
  or2s1 ______443965(.DIN1 (__9_9___26416), .DIN2 (________25666), .Q
       (________25916));
  nor2s1 _______443966(.DIN1 (___9____26215), .DIN2 (________25683), .Q
       (________25915));
  or2s1 _______443967(.DIN1 (________25913), .DIN2 (_____9__25693), .Q
       (________25914));
  nor2s1 _______443968(.DIN1 (___0_9__25318), .DIN2 (________25677), .Q
       (________25912));
  nor2s1 _______443969(.DIN1 (________25910), .DIN2 (_____0__25685), .Q
       (________25911));
  nnd2s1 _______443970(.DIN1 (__99____27118), .DIN2
       (_______________18878), .Q (_____0__25909));
  or2s1 _______443971(.DIN1 (__9_____26647), .DIN2 (________25729), .Q
       (_____9__25908));
  nnd2s1 _______443972(.DIN1 (________25689), .DIN2 (____9___21899), .Q
       (________25907));
  or2s1 _______443973(.DIN1 (__9_____26953), .DIN2 (________25905), .Q
       (________25906));
  nor2s1 ______443974(.DIN1 (__9_9___26695), .DIN2 (________25673), .Q
       (________25904));
  nor2s1 _______443975(.DIN1 (_____9__25829), .DIN2 (________25696), .Q
       (________25903));
  nor2s1 _______443976(.DIN1 (________25901), .DIN2 (________25670), .Q
       (________25902));
  nnd2s1 _______443977(.DIN1 (________25709), .DIN2 (____9___23707), .Q
       (________25900));
  nnd2s1 _______443978(.DIN1 (_____9__25711), .DIN2 (________24230), .Q
       (_____0__25899));
  nor2s1 ______443979(.DIN1 (________25897), .DIN2 (________25896), .Q
       (________25898));
  xor2s1 _______443980(.DIN1 (________25508), .DIN2 (_________35066),
       .Q (________25895));
  nnd2s1 _______443981(.DIN1 (____9___25651), .DIN2 (clk), .Q
       (________25894));
  nnd2s1 _______443982(.DIN1 (____9___24783), .DIN2
       (______________18867), .Q (________25893));
  nnd2s1 _______443983(.DIN1 (____0___25663), .DIN2 (_________35074),
       .Q (________25892));
  or2s1 _______443984(.DIN1 (________26094), .DIN2 (____0___25662), .Q
       (________25891));
  nnd2s1 _____9_443985(.DIN1 (____0___25659), .DIN2 (_____0__25090), .Q
       (_____0__25890));
  and2s1 _____9_443986(.DIN1 (________25632), .DIN2 (____90__23792), .Q
       (_____9__25889));
  or2s1 _____0_443987(.DIN1 (________25887), .DIN2 (____0___25658), .Q
       (________25888));
  nnd2s1 _____0_443988(.DIN1 (____00__25655), .DIN2 (___0____23508), .Q
       (________25886));
  nnd2s1 _____443989(.DIN1 (______0__32006), .DIN2 (________25638), .Q
       (________25885));
  nor2s1 _______443990(.DIN1 (________25814), .DIN2 (________25626), .Q
       (________25884));
  nor2s1 _______443991(.DIN1 (_________28603), .DIN2
       (______________18867), .Q (________25883));
  or2s1 _______443992(.DIN1 (________25881), .DIN2 (____9___25650), .Q
       (________25882));
  nnd2s1 _______443993(.DIN1 (________25642), .DIN2 (_____9__24655), .Q
       (_____0__25880));
  nor2s1 _______443994(.DIN1 (______________18867), .DIN2
       (______________0______________________18828), .Q
       (_____9__25879));
  nor2s1 _______443995(.DIN1 (___0_____27696), .DIN2 (____09__25664),
       .Q (________25878));
  nor2s1 _______443996(.DIN1 (___0_____27730), .DIN2 (____9___25648),
       .Q (________25877));
  nor2s1 _______443997(.DIN1 (____0___24522), .DIN2 (_____9__25624), .Q
       (________25876));
  nnd2s1 _______443998(.DIN1 (_____9__25644), .DIN2 (________25874), .Q
       (________25875));
  nor2s1 _______443999(.DIN1 (________25872), .DIN2 (____9___25653), .Q
       (________25873));
  nnd2s1 _____9_444000(.DIN1 (_____0__25870), .DIN2 (________22869), .Q
       (________25871));
  nor2s1 _____0_444001(.DIN1 (________24083), .DIN2 (________25630), .Q
       (_____9__25869));
  nor2s1 _______444002(.DIN1 (___9_0__24316), .DIN2 (________25628), .Q
       (________25868));
  nnd2s1 _______444003(.DIN1 (________25623), .DIN2 (________25866), .Q
       (________25867));
  and2s1 _______444004(.DIN1 (________25640), .DIN2 (________25864), .Q
       (________25865));
  nor2s1 _______444005(.DIN1 (___9____23381), .DIN2 (________25619), .Q
       (________25863));
  and2s1 _______444006(.DIN1 (________25621), .DIN2 (________25861), .Q
       (________25862));
  nnd2s1 _______444007(.DIN1 (____9___25649), .DIN2 (____0___22632), .Q
       (_____0__25860));
  nnd2s1 ______444008(.DIN1 (____0___25660), .DIN2 (_________35062), .Q
       (____09__25859));
  nnd2s1 ______444009(.DIN1 (________25618), .DIN2 (________21886), .Q
       (____0___25858));
  nor2s1 _______444010(.DIN1 (______________18867), .DIN2
       (_________28939), .Q (__90____26267));
  nnd2s1 _______444011(.DIN1
       (______________________________________0___________), .DIN2
       (______________18867), .Q (___9____26228));
  xor2s1 _______444012(.DIN1 (________25502), .DIN2 (____0___25857), .Q
       (____0____28174));
  and2s1 _______444013(.DIN1 (________25586), .DIN2 (___00____27222),
       .Q (____0___25856));
  nnd2s1 _______444014(.DIN1 (________25594), .DIN2 (________25158), .Q
       (____0___25855));
  or2s1 _______444015(.DIN1 (____0___25853), .DIN2 (________25570), .Q
       (____0___25854));
  nor2s1 _______444016(.DIN1 (________25389), .DIN2 (________25605), .Q
       (____0___25852));
  nnd2s1 ______444017(.DIN1 (________25585), .DIN2 (___9____26235), .Q
       (____0___25851));
  nnd2s1 _____9_444018(.DIN1 (________25590), .DIN2 (___09___23526), .Q
       (____00__25850));
  nor2s1 _____0_444019(.DIN1 (__990___27084), .DIN2 (________25602), .Q
       (____99__25849));
  nnd2s1 _____0_444020(.DIN1 (_____0__25588), .DIN2 (________26121), .Q
       (____9___25848));
  nnd2s1 _____0_444021(.DIN1 (________25601), .DIN2 (____0___22814), .Q
       (____9___25847));
  nor2s1 _______444022(.DIN1 (_____9__21884), .DIN2 (________25569), .Q
       (____9___25846));
  nor2s1 ______444023(.DIN1 (________23961), .DIN2 (________25598), .Q
       (____9___25845));
  nor2s1 _______444024(.DIN1 (___0____22559), .DIN2 (_____0__25597), .Q
       (____9___25844));
  or2s1 _______444025(.DIN1 (________25123), .DIN2 (________25595), .Q
       (____9___25843));
  nor2s1 _______444026(.DIN1 (________25772), .DIN2 (________25592), .Q
       (____9___25842));
  nnd2s1 _______444027(.DIN1 (________25576), .DIN2 (____90__25840), .Q
       (____9___25841));
  nor2s1 _______444028(.DIN1 (___9____24263), .DIN2 (_____0__25607), .Q
       (_____9__25839));
  nor2s1 _______444029(.DIN1 (________22132), .DIN2 (________25591), .Q
       (________25838));
  nnd2s1 _______444030(.DIN1 (________25589), .DIN2 (________25836), .Q
       (________25837));
  nnd2s1 ______444031(.DIN1 (________25581), .DIN2 (________24632), .Q
       (________25835));
  or2s1 ______444032(.DIN1 (_____0__25997), .DIN2 (________25583), .Q
       (________25834));
  nor2s1 _______444033(.DIN1 (____9___23973), .DIN2 (________25600), .Q
       (________25833));
  nor2s1 _______444034(.DIN1 (________25831), .DIN2 (________25572), .Q
       (________25832));
  nor2s1 ______444035(.DIN1 (_____9__25829), .DIN2 (________25599), .Q
       (_____0__25830));
  nor2s1 _______444036(.DIN1 (________23284), .DIN2 (_____0__25529), .Q
       (________25828));
  nor2s1 _______444037(.DIN1 (________25580), .DIN2 (________25687), .Q
       (________25827));
  or2s1 _____9_444038(.DIN1 (___9____26182), .DIN2 (________25571), .Q
       (________25826));
  or2s1 _____444039(.DIN1 (__90_0__26281), .DIN2 (_____9__25587), .Q
       (________25825));
  nnd2s1 ______444040(.DIN1 (________25603), .DIN2 (_____9___28891), .Q
       (________25824));
  nor2s1 _______444041(.DIN1 (________25499), .DIN2 (_____0__25578), .Q
       (________25823));
  nnd2s1 _______444042(.DIN1 (_____9__25577), .DIN2 (_____9___28891),
       .Q (________25822));
  nnd2s1 ______444043(.DIN1 (________25574), .DIN2 (________23559), .Q
       (________25821));
  or2s1 _______444044(.DIN1 (________24546), .DIN2 (__99_0__27154), .Q
       (_____0__25820));
  nor2s1 _______444045(.DIN1 (__9__0__26485), .DIN2 (_____0__25568), .Q
       (_____9__25819));
  nnd2s1 _____0_444046(.DIN1 (________25517), .DIN2 (________25817), .Q
       (________25818));
  and2s1 _______444047(.DIN1 (____0___25565), .DIN2 (___9____23397), .Q
       (________25816));
  nor2s1 _______444048(.DIN1 (________25814), .DIN2 (________25537), .Q
       (________25815));
  nor2s1 _______444049(.DIN1 (________25812), .DIN2 (____0___25562), .Q
       (________25813));
  nnd2s1 _______444050(.DIN1 (_____9__25510), .DIN2 (___00____27213),
       .Q (________25811));
  nor2s1 _______444051(.DIN1 (________22001), .DIN2 (____00__25558), .Q
       (_____0__25810));
  nnd2s1 _______444052(.DIN1 (_________34792), .DIN2 (________25803),
       .Q (_____9__25809));
  nnd2s1 _____9_444053(.DIN1 (_____9__25519), .DIN2 (___0_____27915),
       .Q (________25808));
  and2s1 _____9_444054(.DIN1 (____0___25559), .DIN2 (________25806), .Q
       (________25807));
  and2s1 _____444055(.DIN1 (____99__25557), .DIN2 (________25866), .Q
       (________25805));
  nnd2s1 _____444056(.DIN1 (____9___25556), .DIN2 (________25803), .Q
       (________25804));
  nor2s1 _______444057(.DIN1 (__9090), .DIN2 (________25584), .Q
       (________26103));
  dffacs1 _________________9_444058(.CLRB (reset), .CLK (clk), .DIN
       (_____0__25539), .Q
       (______________0______________________18825));
  hi1s1 _______444059(.DIN (_______________18878), .Q (_________31058));
  and2s1 _______444060(.DIN1 (_____0__25501), .DIN2 (___0_____27780),
       .Q (________25802));
  nnd2s1 _______444061(.DIN1 (_____9__25538), .DIN2 (________23780), .Q
       (________25801));
  nor2s1 _______444062(.DIN1 (__9_9___26698), .DIN2 (____0___25564), .Q
       (_____0__25800));
  nnd2s1 ______444063(.DIN1 (________25521), .DIN2 (________25798), .Q
       (_____9__25799));
  nor2s1 _______444064(.DIN1 (__9_____26621), .DIN2 (________25547), .Q
       (________25797));
  nnd2s1 _______444065(.DIN1 (________25546), .DIN2 (___90___24242), .Q
       (________25796));
  nnd2s1 ______444066(.DIN1 (________25545), .DIN2 (___90___25180), .Q
       (________25795));
  or2s1 _______444067(.DIN1 (________25793), .DIN2 (____09__25567), .Q
       (________25794));
  nor2s1 _______444068(.DIN1 (____________18893), .DIN2
       (____9___25749), .Q (________25792));
  nnd2s1 _______444069(.DIN1 (_____9__25491), .DIN2 (_____0__25790), .Q
       (________25791));
  nor2s1 _______444070(.DIN1 (__99_9__27116), .DIN2 (_____0__25492), .Q
       (_____9__25789));
  nnd2s1 ______444071(.DIN1 (________25518), .DIN2 (inData[20]), .Q
       (________25788));
  nnd2s1 ______444072(.DIN1 (____0___25561), .DIN2 (________24822), .Q
       (________25787));
  nor2s1 _______444073(.DIN1 (____0___24520), .DIN2 (________25530), .Q
       (________25786));
  nnd2s1 ______444074(.DIN1 (________25526), .DIN2 (___0____22598), .Q
       (________25785));
  nnd2s1 _____9_444075(.DIN1 (________25523), .DIN2 (____9___25168), .Q
       (________25784));
  or2s1 _____9_444076(.DIN1 (________25782), .DIN2 (________25527), .Q
       (________25783));
  nnd2s1 _____9_444077(.DIN1 (________25540), .DIN2 (_____0__23326), .Q
       (________25781));
  nor2s1 _____9_444078(.DIN1 (__9_____26831), .DIN2 (____90__25549), .Q
       (_____0__25780));
  nor2s1 _____9_444079(.DIN1 (________25989), .DIN2 (________25532), .Q
       (_____9__25779));
  and2s1 _____0_444080(.DIN1 (________25542), .DIN2 (__9_____26812), .Q
       (________25778));
  nor2s1 _____0_444081(.DIN1 (___90___22447), .DIN2 (____0___25563), .Q
       (________25777));
  nor2s1 _______444082(.DIN1 (___9_9__23395), .DIN2 (________25525), .Q
       (________25776));
  nnd2s1 _______444083(.DIN1 (________25608), .DIN2 (________25774), .Q
       (________25775));
  or2s1 _______444084(.DIN1 (________25772), .DIN2 (________25543), .Q
       (________25773));
  nnd2s1 ______444085(.DIN1 (________25514), .DIN2 (_____0__25770), .Q
       (________25771));
  nnd2s1 _______444086(.DIN1 (________25512), .DIN2 (__9_____26576), .Q
       (_____9__25769));
  nor2s1 _______444087(.DIN1 (________26101), .DIN2 (_____0__25511), .Q
       (________25768));
  nnd2s1 _______444088(.DIN1 (____9___25550), .DIN2 (____9___21899), .Q
       (________25767));
  nor2s1 _______444089(.DIN1 (_________31505), .DIN2 (________25761),
       .Q (________25766));
  nor2s1 _______444090(.DIN1 (________23754), .DIN2 (_________34790),
       .Q (________25765));
  nor2s1 _______444091(.DIN1 (____0___23717), .DIN2 (_____9__25548), .Q
       (________25764));
  nnd2s1 ______444092(.DIN1 (________25515), .DIN2 (____9___23885), .Q
       (________25763));
  nnd2s1 _______444093(.DIN1 (________25761), .DIN2 (____00__21166), .Q
       (________25762));
  xor2s1 _______444094(.DIN1 (_________________18699), .DIN2
       (_________________18685), .Q (____09__25760));
  nnd2s1 _______444095(.DIN1 (________25498), .DIN2 (____0___25758), .Q
       (____0___25759));
  nor2s1 _______444096(.DIN1 (_____0__24447), .DIN2 (________25496), .Q
       (____0___25757));
  nnd2s1 _____9_444097(.DIN1 (________25497), .DIN2 (__90_0__26291), .Q
       (____0___25756));
  and2s1 _____0_444098(.DIN1 (_____9__25500), .DIN2 (____0___25754), .Q
       (____0___25755));
  nnd2s1 _______444099(.DIN1 (________25493), .DIN2 (____0___25752), .Q
       (____0___25753));
  nor2s1 _______444100(.DIN1 (____9___23169), .DIN2 (________25495), .Q
       (____00__25751));
  and2s1 ______444101(.DIN1 (________25522), .DIN2 (____99__25750), .Q
       (________26014));
  nor2s1 ______444102(.DIN1 (outData[7]), .DIN2 (________25761), .Q
       (_____9__25996));
  and2s1 _______444103(.DIN1 (____9___25554), .DIN2 (__9__0__26854), .Q
       (____99__26046));
  and2s1 _______444104(.DIN1 (____9___25749), .DIN2
       (____________18893), .Q (_____0__26107));
  hi1s1 _______444105(.DIN (______________18867), .Q (________26002));
  nor2s1 _______444106(.DIN1 (________25440), .DIN2 (___0____22549), .Q
       (____9___25748));
  nor2s1 _____0_444107(.DIN1 (____9___25746), .DIN2 (________25488), .Q
       (____9___25747));
  nnd2s1 _______444108(.DIN1 (_____9__25445), .DIN2 (___9____24298), .Q
       (____9___25745));
  and2s1 _______444109(.DIN1 (________25441), .DIN2 (_____0__25770), .Q
       (____9___25744));
  and2s1 _______444110(.DIN1 (_____0__25446), .DIN2 (____9___25742), .Q
       (____9___25743));
  nnd2s1 _______444111(.DIN1 (________25449), .DIN2 (________25717), .Q
       (____90__25741));
  nor2s1 ______444112(.DIN1 (________25739), .DIN2 (________25448), .Q
       (_____9__25740));
  nnd2s1 ______444113(.DIN1 (________25411), .DIN2 (________25991), .Q
       (________25738));
  nnd2s1 _____9_444114(.DIN1 (________25485), .DIN2 (________22229), .Q
       (________25737));
  nnd2s1 _____9_444115(.DIN1 (________25486), .DIN2 (________24824), .Q
       (________25736));
  nnd2s1 _____9_444116(.DIN1 (________25473), .DIN2 (________25734), .Q
       (________25735));
  nnd2s1 _____9_444117(.DIN1 (________25450), .DIN2 (________25378), .Q
       (________25733));
  nnd2s1 _____0_444118(.DIN1 (_____0__25482), .DIN2 (________23664), .Q
       (________25732));
  and2s1 _____0_444119(.DIN1 (________25398), .DIN2 (________23677), .Q
       (_____0__25731));
  nor2s1 _____0_444120(.DIN1 (________25812), .DIN2 (_________34796),
       .Q (_____9__25730));
  or2s1 ______444121(.DIN1 (________25728), .DIN2 (_____9__25425), .Q
       (________25729));
  and2s1 _______444122(.DIN1 (________25480), .DIN2 (________25726), .Q
       (________25727));
  nnd2s1 _______444123(.DIN1 (________25477), .DIN2 (_____0__25625), .Q
       (________25725));
  nnd2s1 _______444124(.DIN1 (_____0__25436), .DIN2 (________22289), .Q
       (________25724));
  nor2s1 _______444125(.DIN1 (________25722), .DIN2 (________25475), .Q
       (________25723));
  nnd2s1 ______444126(.DIN1 (________25474), .DIN2 (______0__35038), .Q
       (_____0__25721));
  or2s1 ______444127(.DIN1 (____9___25652), .DIN2 (_____0__25472), .Q
       (_____9__25720));
  or2s1 _______444128(.DIN1 (________24024), .DIN2 (_____9__25405), .Q
       (________25719));
  nnd2s1 _______444129(.DIN1 (________25404), .DIN2 (________25717), .Q
       (________25718));
  nor2s1 _______444130(.DIN1 (________25715), .DIN2 (____0___25469), .Q
       (________25716));
  nnd2s1 _______444131(.DIN1 (____0___25468), .DIN2 (_____90__34918),
       .Q (________25714));
  or2s1 ______444132(.DIN1 (_____0__25712), .DIN2 (____0___25467), .Q
       (________25713));
  nor2s1 _______444133(.DIN1 (________25710), .DIN2 (____0___25466), .Q
       (_____9__25711));
  nor2s1 _______444134(.DIN1 (___0____24368), .DIN2 (____9___25461), .Q
       (________25709));
  nnd2s1 _______444135(.DIN1 (____9___25459), .DIN2 (____0___25465), .Q
       (________25708));
  nnd2s1 _______444136(.DIN1 (____9___25456), .DIN2 (_________35046),
       .Q (________25706));
  nnd2s1 _______444137(.DIN1 (________25428), .DIN2 (________25704), .Q
       (________25705));
  nor2s1 ______444138(.DIN1 (________24483), .DIN2 (_____9__25454), .Q
       (_____0__25703));
  nor2s1 _______444139(.DIN1 (________24183), .DIN2 (________25453), .Q
       (_____9__25702));
  and2s1 ______444140(.DIN1 (_____0__25416), .DIN2 (________25836), .Q
       (________25701));
  nor2s1 _______444141(.DIN1 (___9____24313), .DIN2 (________25487), .Q
       (________25700));
  or2s1 _______444142(.DIN1 (______0__28551), .DIN2 (________25431), .Q
       (________25699));
  nor2s1 _______444143(.DIN1 (________25639), .DIN2 (____0___25471), .Q
       (________25698));
  nnd2s1 _______444144(.DIN1 (________25427), .DIN2 (_________34956),
       .Q (________25696));
  nor2s1 _______444145(.DIN1 (_____0__25694), .DIN2 (________25420), .Q
       (________25695));
  nnd2s1 _______444146(.DIN1 (________25439), .DIN2 (_________35064),
       .Q (_____9__25693));
  nnd2s1 _______444147(.DIN1 (________25432), .DIN2 (___0____21654), .Q
       (________25692));
  nnd2s1 _____444148(.DIN1 (________25429), .DIN2 (________24939), .Q
       (________25691));
  nnd2s1 _____9_444149(.DIN1 (________25479), .DIN2 (___9____26200), .Q
       (________25690));
  nnd2s1 _____444150(.DIN1 (________25430), .DIN2 (__9_____26387), .Q
       (________25689));
  or2s1 _____444151(.DIN1 (________25418), .DIN2 (________25687), .Q
       (________25688));
  nnd2s1 _____0_444152(.DIN1 (_____0__25426), .DIN2 (_____0__25665), .Q
       (________25686));
  or2s1 _____0_444153(.DIN1 (_____9__25684), .DIN2 (_____0__25406), .Q
       (_____0__25685));
  nnd2s1 _____0_444154(.DIN1 (________25421), .DIN2 (________25864), .Q
       (________25683));
  nor2s1 _____444155(.DIN1 (________25901), .DIN2 (________25438), .Q
       (________25682));
  dffacs1 __________________444156(.CLRB (reset), .CLK (clk), .DIN
       (____0___25374), .QN (________________18678));
  dffacs1 __________________444157(.CLRB (reset), .CLK (clk), .DIN
       (_____9__25396), .Q (________________18676));
  dffacs1 ___________________444158(.CLRB (reset), .CLK (clk), .DIN
       (___09___25363), .Q (______________0___________________9));
  dffacs2 __________________444159(.CLRB (reset), .CLK (clk), .DIN
       (_____9__25481), .Q (_______________18878));
  nnd2s1 _____0_444160(.DIN1 (________25609), .DIN2 (________25383), .Q
       (________25681));
  nor2s1 _______444161(.DIN1 (_____0__25616), .DIN2 (________25395), .Q
       (________25680));
  or2s1 _______444162(.DIN1 (___0_____27281), .DIN2 (____00__25464), .Q
       (________25679));
  nnd2s1 ______444163(.DIN1 (_____0__25397), .DIN2 (________25726), .Q
       (________25678));
  nnd2s1 _______444164(.DIN1 (________25443), .DIN2 (________24804), .Q
       (________25677));
  nor2s1 _______444165(.DIN1 (_____9__21884), .DIN2 (________25433), .Q
       (________25676));
  nnd2s1 ______444166(.DIN1 (____9___25457), .DIN2 (_____9__25674), .Q
       (_____0__25675));
  nnd2s1 _______444167(.DIN1 (________25393), .DIN2 (________25672), .Q
       (________25673));
  nnd2s1 _______444168(.DIN1 (________25407), .DIN2 (________24944), .Q
       (________25671));
  nnd2s1 _______444169(.DIN1 (________25402), .DIN2 (________22882), .Q
       (________25670));
  nor2s1 _______444170(.DIN1 (________25531), .DIN2 (________25434), .Q
       (________25669));
  nor2s1 _______444171(.DIN1 (_____9__25415), .DIN2 (______0__34798),
       .Q (________25668));
  nor2s1 _______444172(.DIN1 (___0_____27696), .DIN2 (________25484),
       .Q (________25667));
  nnd2s1 ______444173(.DIN1 (________25414), .DIN2 (_____0__25665), .Q
       (________25666));
  nor2s1 _______444174(.DIN1 (___9____25206), .DIN2 (________25381), .Q
       (____09__25664));
  nor2s1 _______444175(.DIN1 (________23273), .DIN2 (________25379), .Q
       (____0___25663));
  nnd2s1 ______444176(.DIN1 (___0____25349), .DIN2 (____0___25661), .Q
       (____0___25662));
  and2s1 _____444177(.DIN1 (_____0__25377), .DIN2 (________26079), .Q
       (____0___25660));
  and2s1 _____0_444178(.DIN1 (________25382), .DIN2 (________24629), .Q
       (____0___25659));
  or2s1 _____0_444179(.DIN1 (________24105), .DIN2 (____09__25376), .Q
       (____0___25658));
  nnd2s1 _____0_444180(.DIN1 (___0____25345), .DIN2 (____0___25656), .Q
       (____0___25657));
  and2s1 _____444181(.DIN1 (____0___25369), .DIN2 (____99__25654), .Q
       (____00__25655));
  or2s1 ______444182(.DIN1 (____9___25652), .DIN2 (____0___25372), .Q
       (____9___25653));
  nor2s1 _______444183(.DIN1 (________23996), .DIN2 (____0___25375), .Q
       (____9___25651));
  or2s1 _______444184(.DIN1 (________23288), .DIN2 (________25385), .Q
       (____9___25650));
  nor2s1 ______444185(.DIN1 (____09__23896), .DIN2 (____0___25373), .Q
       (____9___25649));
  or2s1 ______444186(.DIN1 (____9___25647), .DIN2 (____0___25371), .Q
       (____9___25648));
  and2s1 _______444187(.DIN1 (___0____25352), .DIN2 (____90__25645), .Q
       (____9___25646));
  and2s1 _______444188(.DIN1 (___09___25365), .DIN2 (________25643), .Q
       (_____9__25644));
  and2s1 ______444189(.DIN1 (___09___25362), .DIN2 (________25641), .Q
       (________25642));
  nor2s1 _______444190(.DIN1 (________25639), .DIN2 (_____9__25386), .Q
       (________25640));
  or2s1 _______444191(.DIN1 (_____0___31003), .DIN2
       (_________________18685), .Q (________25638));
  nnd2s1 _____9_444192(.DIN1 (________25636), .DIN2 (________25105), .Q
       (________25637));
  nnd2s1 _______444193(.DIN1 (_____9__25435), .DIN2 (_____9__25634), .Q
       (_____0__25635));
  nnd2s1 _____444194(.DIN1 (________25384), .DIN2 (___9____21591), .Q
       (________25633));
  nor2s1 _____0_444195(.DIN1 (________25622), .DIN2 (_____0__25387), .Q
       (________25632));
  nnd2s1 ______444196(.DIN1 (____00__25367), .DIN2 (___0_____27594), .Q
       (________25631));
  nnd2s1 _______444197(.DIN1 (___0____25348), .DIN2 (________23063), .Q
       (________25630));
  nnd2s1 _______444198(.DIN1 (___0____25355), .DIN2 (___0____21654), .Q
       (________25629));
  nnd2s1 _______444199(.DIN1 (________25388), .DIN2 (________25627), .Q
       (________25628));
  nnd2s1 ______444200(.DIN1 (________25412), .DIN2 (_____0__25625), .Q
       (________25626));
  nnd2s1 ______444201(.DIN1 (___09___25364), .DIN2 (________23307), .Q
       (_____9__25624));
  nor2s1 ______444202(.DIN1 (________25622), .DIN2 (___09___25360), .Q
       (________25623));
  and2s1 _______444203(.DIN1 (___09___25359), .DIN2 (____0___25566), .Q
       (________25621));
  nor2s1 _______444204(.DIN1 (________25535), .DIN2 (________25390), .Q
       (________25620));
  nnd2s1 ______444205(.DIN1 (________25391), .DIN2 (________23226), .Q
       (________25619));
  nnd2s1 _______444206(.DIN1 (___0____25344), .DIN2 (________23222), .Q
       (________25618));
  nor2s1 _______444207(.DIN1 (_____0__25616), .DIN2 (________25400), .Q
       (________25617));
  nor2s1 _______444208(.DIN1 (_____9__25615), .DIN2 (________25614), .Q
       (__9_00__26514));
  nor2s1 _______444209(.DIN1 (__9_____26632), .DIN2 (________25403), .Q
       (________25905));
  xor2s1 _______444210(.DIN1 (___9____25218), .DIN2 (_________31431),
       .Q (________25896));
  nnd2s1 _______444211(.DIN1 (________25613), .DIN2 (________25612), .Q
       (________26062));
  nnd2s1 _______444212(.DIN1 (________25611), .DIN2 (________25610), .Q
       (____0____29150));
  nnd2s1 _____0_444213(.DIN1 (___0_0__25347), .DIN2 (________19454), .Q
       (_____0__25870));
  xor2s1 ______444214(.DIN1 (________25609), .DIN2 (outData[6]), .Q
       (________25959));
  dffacs1 ___________________444215(.CLRB (reset), .CLK (clk), .DIN
       (____90__25455), .QN (_________________18681));
  dffacs1 _________________444216(.CLRB (reset), .CLK (clk), .DIN
       (___0____25351), .Q (______________18867));
  and2s1 _______444217(.DIN1 (___0_9__25299), .DIN2 (________25923), .Q
       (________25608));
  nnd2s1 ______444218(.DIN1 (___0_0__25319), .DIN2 (_____9__25606), .Q
       (_____0__25607));
  nnd2s1 _____0_444219(.DIN1 (___0____25340), .DIN2 (________25604), .Q
       (________25605));
  or2s1 ______444220(.DIN1 (____9___25945), .DIN2 (___0____25320), .Q
       (________25603));
  nor2s1 ______444221(.DIN1 (___0_____27483), .DIN2 (___0_9__25337), .Q
       (________25602));
  nor2s1 _______444222(.DIN1 (_____0__22924), .DIN2 (___0____25335), .Q
       (________25601));
  or2s1 _______444223(.DIN1 (________26092), .DIN2 (___0____25331), .Q
       (________25600));
  nnd2s1 _______444224(.DIN1 (___0____25330), .DIN2 (________22682), .Q
       (________25599));
  nnd2s1 _______444225(.DIN1 (___0_9__25327), .DIN2 (________23021), .Q
       (________25598));
  nnd2s1 _______444226(.DIN1 (___0____25326), .DIN2 (_____9__25596), .Q
       (_____0__25597));
  nnd2s1 ______444227(.DIN1 (___0____25325), .DIN2 (_____9__23544), .Q
       (________25595));
  nor2s1 _______444228(.DIN1 (________25593), .DIN2 (___0____25339), .Q
       (________25594));
  nnd2s1 _______444229(.DIN1 (___0_9__25309), .DIN2 (___09___25361), .Q
       (________25592));
  or2s1 ______444230(.DIN1 (________24100), .DIN2 (___0____25322), .Q
       (________25591));
  nor2s1 _______444231(.DIN1 (_____9___34926), .DIN2 (___0____25315),
       .Q (________25590));
  nor2s1 _______444232(.DIN1 (________25413), .DIN2 (___0____25341), .Q
       (________25589));
  nor2s1 _______444233(.DIN1 (___0____25303), .DIN2 (___0____25317), .Q
       (_____0__25588));
  nnd2s1 _______444234(.DIN1 (___0____25308), .DIN2 (________26079), .Q
       (_____9__25587));
  nor2s1 _____9_444235(.DIN1 (___0_0__25290), .DIN2 (___0____25313), .Q
       (________25586));
  nor2s1 _____0_444236(.DIN1 (_____9__24490), .DIN2 (________25573), .Q
       (________25585));
  nnd2s1 _____0_444237(.DIN1 (___0_0__25300), .DIN2 (__9_0___26517), .Q
       (________25584));
  or2s1 ______444238(.DIN1 (________25582), .DIN2 (___0____25314), .Q
       (________25583));
  nor2s1 _______444239(.DIN1 (________26008), .DIN2 (___0____25321), .Q
       (________25581));
  xor2s1 _______444240(.DIN1 (________25579), .DIN2 (________25104), .Q
       (________25580));
  nnd2s1 _______444241(.DIN1 (___0____25316), .DIN2 (________24216), .Q
       (_____0__25578));
  nnd2s1 _______444242(.DIN1 (___0_0__25338), .DIN2 (________24735), .Q
       (_____9__25577));
  nor2s1 ______444243(.DIN1 (___9_0__26167), .DIN2 (___0____25334), .Q
       (________25576));
  nnd2s1 _______444244(.DIN1 (___0____25312), .DIN2 (_____9___28891),
       .Q (________25575));
  nnd2s1 _______444245(.DIN1 (________25573), .DIN2 (___0____21654), .Q
       (________25574));
  nnd2s1 _______444246(.DIN1 (___0____25304), .DIN2 (_____0__24551), .Q
       (________25572));
  nnd2s1 _______444247(.DIN1 (___0____25311), .DIN2 (___0_____27600),
       .Q (________25571));
  nnd2s1 _______444248(.DIN1 (___0____25342), .DIN2 (_____0__26077), .Q
       (________25570));
  nor2s1 _______444249(.DIN1 (___9____23387), .DIN2 (___0____25332), .Q
       (________25569));
  nnd2s1 _______444250(.DIN1 (___0____25294), .DIN2 (________25447), .Q
       (_____0__25568));
  nnd2s1 _______444251(.DIN1 (___0_9__25289), .DIN2 (____0___25566), .Q
       (____09__25567));
  nor2s1 _______444252(.DIN1 (________22727), .DIN2 (___9____25257), .Q
       (____0___25565));
  or2s1 _______444253(.DIN1 (__9_9___26505), .DIN2 (___9____25227), .Q
       (____0___25564));
  nnd2s1 _____9_444254(.DIN1 (___9____25259), .DIN2 (___909__24248), .Q
       (____0___25563));
  nnd2s1 _____9_444255(.DIN1 (___0____25286), .DIN2 (_____9__24838), .Q
       (____0___25562));
  and2s1 _____9_444256(.DIN1 (___0____25291), .DIN2 (____0___25560), .Q
       (____0___25561));
  and2s1 _____444257(.DIN1 (___0____25283), .DIN2 (___0_____27816), .Q
       (____0___25559));
  nnd2s1 _____0_444258(.DIN1 (___0_0__25281), .DIN2 (____90__24877), .Q
       (____00__25558));
  nor2s1 _____0_444259(.DIN1 (________25483), .DIN2 (___0____25287), .Q
       (____99__25557));
  and2s1 _____0_444260(.DIN1 (___9_9__25240), .DIN2 (_____0__23695), .Q
       (____9___25556));
  nnd2s1 _____0_444261(.DIN1 (___0____25282), .DIN2 (__9_____26469), .Q
       (____9___25555));
  nor2s1 _______444262(.DIN1 (___0_____27483), .DIN2 (___0____25293),
       .Q (____9___25554));
  nor2s1 _______444263(.DIN1 (________24567), .DIN2 (___9____25248), .Q
       (____9___25553));
  nor2s1 _______444264(.DIN1 (________24721), .DIN2 (___0____25297), .Q
       (____9___25552));
  xor2s1 _______444265(.DIN1 (______________18870), .DIN2
       (____9___25551), .Q (________25697));
  xnr2s1 _______444266(.DIN1 (_________30341), .DIN2 (_____9__25108),
       .Q (__99_0__27154));
  or2s1 ______444267(.DIN1 (___00____27200), .DIN2 (___9____25222), .Q
       (____9___25550));
  or2s1 _______444268(.DIN1 (__9_____26350), .DIN2 (___00___25272), .Q
       (____90__25549));
  or2s1 ______444269(.DIN1 (___0_0___27561), .DIN2 (___00___25274), .Q
       (_____9__25548));
  nor2s1 ______444270(.DIN1 (________26032), .DIN2 (___00___25278), .Q
       (________25547));
  nor2s1 _______444271(.DIN1 (________22344), .DIN2 (___0____25298), .Q
       (________25546));
  nor2s1 _______444272(.DIN1 (____9___23342), .DIN2 (___9____25256), .Q
       (________25545));
  nnd2s1 _______444273(.DIN1 (___9____25234), .DIN2 (________24497), .Q
       (________25544));
  nnd2s1 _______444274(.DIN1 (___0____25306), .DIN2 (________23686), .Q
       (________25543));
  and2s1 _______444275(.DIN1 (___000__25271), .DIN2 (________25874), .Q
       (________25542));
  nnd2s1 _______444276(.DIN1 (___999__25270), .DIN2 (________24530), .Q
       (________25541));
  nor2s1 _______444277(.DIN1 (________24079), .DIN2 (___99___25269), .Q
       (________25540));
  nnd2s1 _______444278(.DIN1 (___0_9__20742), .DIN2 (___9____25228), .Q
       (_____0__25539));
  nor2s1 _______444279(.DIN1 (___9_0__25251), .DIN2 (___9____25196), .Q
       (_____9__25538));
  nnd2s1 _______444280(.DIN1 (___99___25267), .DIN2 (_____9__24876), .Q
       (________25537));
  nor2s1 _______444281(.DIN1 (________25535), .DIN2 (___0____25292), .Q
       (________25536));
  hi1s1 _____9_444282(.DIN (________25533), .Q (________25534));
  or2s1 _____0_444283(.DIN1 (________25531), .DIN2 (___9____25255), .Q
       (________25532));
  nnd2s1 _____0_444284(.DIN1 (___9_9__25260), .DIN2 (________25004), .Q
       (________25530));
  nnd2s1 _______444285(.DIN1 (___0____25296), .DIN2 (_____9__25528), .Q
       (_____0__25529));
  nnd2s1 ______444286(.DIN1 (___00___25276), .DIN2 (________24571), .Q
       (________25527));
  nor2s1 _______444287(.DIN1 (________25516), .DIN2 (___9____25252), .Q
       (________25526));
  or2s1 _______444288(.DIN1 (________25524), .DIN2 (___00___25275), .Q
       (________25525));
  nor2s1 _______444289(.DIN1 (_____0__24616), .DIN2 (___9_9__25250), .Q
       (________25523));
  and2s1 _______444290(.DIN1 (___99___25266), .DIN2 (_________35046),
       .Q (________25522));
  and2s1 _______444291(.DIN1 (___9____25242), .DIN2 (_____0__25520), .Q
       (________25521));
  nor2s1 _______444292(.DIN1 (___0_____27798), .DIN2 (___0____25285),
       .Q (_____9__25519));
  nor2s1 _______444293(.DIN1 (___9_9__25220), .DIN2 (___9____24287), .Q
       (________25518));
  nor2s1 ______444294(.DIN1 (________25516), .DIN2 (___00___25279), .Q
       (________25517));
  nor2s1 ______444295(.DIN1 (_____9__24181), .DIN2 (___9____25235), .Q
       (________25515));
  nor2s1 _______444296(.DIN1 (________25513), .DIN2 (___9____25232), .Q
       (________25514));
  nnd2s1 _______444297(.DIN1 (___9____25229), .DIN2 (_____0__25790), .Q
       (________25512));
  nnd2s1 _______444298(.DIN1 (___9_9__25230), .DIN2 (_____0__25790), .Q
       (_____0__25511));
  and2s1 _______444299(.DIN1 (___9____25247), .DIN2 (________25509), .Q
       (_____9__25510));
  nor2s1 _____9_444300(.DIN1 (________25507), .DIN2 (________25506), .Q
       (________25508));
  or2s1 _____444301(.DIN1 (________25504), .DIN2 (________25503), .Q
       (________25505));
  xor2s1 _____0_444302(.DIN1 (___0_9__25346), .DIN2 (_________33541),
       .Q (________25502));
  nor2s1 _______444303(.DIN1 (___9____24293), .DIN2 (___9____25238), .Q
       (_____0__25501));
  nor2s1 _______444304(.DIN1 (________25499), .DIN2 (___9____25215), .Q
       (_____9__25500));
  nor2s1 _______444305(.DIN1 (___9____25214), .DIN2 (________22732), .Q
       (________25498));
  nor2s1 _______444306(.DIN1 (________23239), .DIN2 (___9____25219), .Q
       (________25497));
  nnd2s1 _______444307(.DIN1 (________25494), .DIN2 (_____9__23099), .Q
       (________25496));
  nnd2s1 _____9_444308(.DIN1 (________25494), .DIN2 (________24871), .Q
       (________25495));
  and2s1 ____90_444309(.DIN1 (___9____25209), .DIN2 (___0____22601), .Q
       (________25493));
  and2s1 ____99_444310(.DIN1 (___9____25207), .DIN2 (_____9__25928), .Q
       (_____0__25492));
  nor2s1 ____0_444311(.DIN1 (__9_____26472), .DIN2 (___99___25262), .Q
       (_____9__25491));
  nnd2s1 ____0__444312(.DIN1 (___9____25217), .DIN2 (________25643), .Q
       (___00____27233));
  or2s1 _____9_444313(.DIN1 (________25490), .DIN2 (___9_0__25221), .Q
       (________25934));
  nor2s1 _____9_444314(.DIN1 (outData[6]), .DIN2 (________25609), .Q
       (____9___25749));
  xor2s1 _____0_444315(.DIN1 (_____9__25070), .DIN2 (_________28737),
       .Q (________25761));
  nor2s1 _______444316(.DIN1
       (______________________________________0__________0), .DIN2
       (____9___25551), .Q (________25489));
  nnd2s1 _______444317(.DIN1 (_________34802), .DIN2 (________25806),
       .Q (________25488));
  nnd2s1 _______444318(.DIN1 (___90___25182), .DIN2 (________24852), .Q
       (________25487));
  nor2s1 _______444319(.DIN1 (________25985), .DIN2 (___9_0__25194), .Q
       (________25486));
  nor2s1 _____9_444320(.DIN1 (_________35000), .DIN2 (___9_9__25193),
       .Q (________25485));
  nor2s1 _____9_444321(.DIN1 (________25483), .DIN2 (___9____25187), .Q
       (________25484));
  or2s1 _____9_444322(.DIN1 (____9___25551), .DIN2 (___9____24288), .Q
       (_____0__25482));
  nnd2s1 _____444323(.DIN1 (________25143), .DIN2 (________22828), .Q
       (_____9__25481));
  nor2s1 ______444324(.DIN1 (________25401), .DIN2 (___90___25178), .Q
       (________25480));
  nor2s1 _______444325(.DIN1 (________25478), .DIN2 (________25159), .Q
       (________25479));
  and2s1 ______444326(.DIN1 (___900__25174), .DIN2 (________25476), .Q
       (________25477));
  or2s1 _______444327(.DIN1 (________25831), .DIN2 (___90___25175), .Q
       (________25475));
  nor2s1 _______444328(.DIN1 (__9_9___26698), .DIN2 (____99__25173), .Q
       (________25474));
  nor2s1 _______444329(.DIN1 (________23908), .DIN2 (____9___25172), .Q
       (________25473));
  nnd2s1 _______444330(.DIN1 (____9___25171), .DIN2 (________26089), .Q
       (_____0__25472));
  nnd2s1 _______444331(.DIN1 (________25117), .DIN2 (____0___25470), .Q
       (____0___25471));
  nnd2s1 _______444332(.DIN1 (___9_0__25203), .DIN2 (___9____23396), .Q
       (____0___25469));
  nor2s1 _______444333(.DIN1 (________25478), .DIN2 (___9____25204), .Q
       (____0___25468));
  or2s1 _______444334(.DIN1 (________22641), .DIN2 (________25144), .Q
       (____0___25467));
  nnd2s1 _______444335(.DIN1 (________25131), .DIN2 (____0___25465), .Q
       (____0___25466));
  nnd2s1 _______444336(.DIN1 (________25161), .DIN2 (________24812), .Q
       (____00__25464));
  or2s1 ______444337(.DIN1 (________25160), .DIN2 (____9___25462), .Q
       (____99__25463));
  nnd2s1 ______444338(.DIN1 (________25147), .DIN2 (____9___25460), .Q
       (____9___25461));
  nor2s1 _______444339(.DIN1 (____9___25458), .DIN2 (________25157), .Q
       (____9___25459));
  nor2s1 _______444340(.DIN1 (________25442), .DIN2 (___9____25199), .Q
       (____9___25457));
  nor2s1 _______444341(.DIN1 (________24659), .DIN2 (_____9__25155), .Q
       (____9___25456));
  nnd2s1 ______444342(.DIN1 (________20590), .DIN2 (________25120), .Q
       (____90__25455));
  nnd2s1 _______444343(.DIN1 (___9____25192), .DIN2 (________24568), .Q
       (_____9__25454));
  nnd2s1 _______444344(.DIN1 (________25121), .DIN2 (________25452), .Q
       (________25453));
  nor2s1 ______444345(.DIN1 (_____0__24772), .DIN2 (___9____25188), .Q
       (________25450));
  nor2s1 _______444346(.DIN1 (__990___27088), .DIN2 (________25133), .Q
       (________25449));
  nnd2s1 _______444347(.DIN1 (___9____25201), .DIN2 (________25447), .Q
       (________25448));
  nor2s1 _______444348(.DIN1 (________22342), .DIN2 (_____9__25135), .Q
       (_____0__25446));
  and2s1 _______444349(.DIN1 (___9____25185), .DIN2 (________25444), .Q
       (_____9__25445));
  nor2s1 _______444350(.DIN1 (________25442), .DIN2 (________25128), .Q
       (________25443));
  nor2s1 _____444351(.DIN1 (_____0__25694), .DIN2 (________25149), .Q
       (________25441));
  nor2s1 _____9_444352(.DIN1 (_________30104), .DIN2 (____0____30075),
       .Q (________25440));
  nor2s1 _____9_444353(.DIN1 (____99__24517), .DIN2 (___90___25176), .Q
       (________25439));
  or2s1 _____9_444354(.DIN1 (________25437), .DIN2 (_____0__25146), .Q
       (________25438));
  nor2s1 _____444355(.DIN1 (____0___24798), .DIN2 (________25134), .Q
       (_____0__25436));
  nor2s1 _____0_444356(.DIN1 (________25010), .DIN2 (___90___25177), .Q
       (_____9__25435));
  nnd2s1 _____0_444357(.DIN1 (________25138), .DIN2 (___0____25305), .Q
       (________25434));
  and2s1 _____0_444358(.DIN1 (________25141), .DIN2 (________25774), .Q
       (________25433));
  nnd2s1 _____0_444359(.DIN1 (___9____25189), .DIN2 (_____0__23933), .Q
       (________25432));
  nnd2s1 _____444360(.DIN1 (________25140), .DIN2 (__9__0__26494), .Q
       (________25431));
  nor2s1 _______444361(.DIN1 (__9_____26583), .DIN2 (_____0__25136), .Q
       (________25430));
  nor2s1 _______444362(.DIN1 (________25110), .DIN2 (____9___25166), .Q
       (________25429));
  and2s1 _______444363(.DIN1 (_____9__25164), .DIN2 (________25926), .Q
       (________25428));
  nor2s1 ______444364(.DIN1 (________23767), .DIN2 (_________34806), .Q
       (________25427));
  nor2s1 _______444365(.DIN1 (___9_0__25231), .DIN2 (________25130), .Q
       (_____0__25426));
  or2s1 _______444366(.DIN1 (________25424), .DIN2 (___90___25181), .Q
       (_____9__25425));
  xor2s1 _______444367(.DIN1 (________25422), .DIN2 (______9__33856),
       .Q (________25423));
  nor2s1 _______444368(.DIN1 (__9_____26440), .DIN2 (________25151), .Q
       (________25421));
  nnd2s1 _______444369(.DIN1 (___9____25197), .DIN2 (________25419), .Q
       (________25420));
  xor2s1 _______444370(.DIN1 (____0___19308), .DIN2 (________25417), .Q
       (________25418));
  nor2s1 _______444371(.DIN1 (_____9__25415), .DIN2 (_____0__25109), .Q
       (_____0__25416));
  nor2s1 _______444372(.DIN1 (________25413), .DIN2 (________25152), .Q
       (________25414));
  xor2s1 _______444373(.DIN1
       (______________________________________0_____________18890),
       .DIN2 (___________0___18872), .Q (____9_0__29038));
  dffacs1 ___________________444374(.CLRB (reset), .CLK (clk), .DIN
       (____00__25080), .Q (_________34496));
  nor2s1 _______444375(.DIN1 (____0___25083), .DIN2 (_____9__23820), .Q
       (________25412));
  nor2s1 ______444376(.DIN1 (____0___26055), .DIN2 (________25111), .Q
       (________25411));
  nnd2s1 _______444377(.DIN1 (______________18870), .DIN2
       (____9___25551), .Q (________25410));
  nor2s1 _______444378(.DIN1 (_________30104), .DIN2 (____9___25551),
       .Q (________25409));
  nnd2s1 _______444379(.DIN1 (____9___25551), .DIN2 (_________30104),
       .Q (________25408));
  nor2s1 _______444380(.DIN1 (________23123), .DIN2 (___90___25179), .Q
       (________25407));
  nnd2s1 _______444381(.DIN1 (________25153), .DIN2 (________24505), .Q
       (_____0__25406));
  nnd2s1 _______444382(.DIN1 (_________34804), .DIN2 (____9___24515),
       .Q (_____9__25405));
  and2s1 ______444383(.DIN1 (___9____25190), .DIN2 (________25641), .Q
       (________25404));
  or2s1 _______444384(.DIN1 (________25639), .DIN2 (_____0__25119), .Q
       (________25403));
  nor2s1 ______444385(.DIN1 (________25401), .DIN2 (________25114), .Q
       (________25402));
  and2s1 _______444386(.DIN1 (________25122), .DIN2 (________25399), .Q
       (________25400));
  nnd2s1 _______444387(.DIN1 (___0____25301), .DIN2 (____0____30075),
       .Q (________25398));
  nor2s1 _______444388(.DIN1 (________25401), .DIN2 (____9___25169), .Q
       (_____0__25397));
  nor2s1 _______444389(.DIN1 (____9___25551), .DIN2
       (_________________0___18660), .Q (_____9__25396));
  and2s1 ______444390(.DIN1 (________25163), .DIN2 (________25394), .Q
       (________25395));
  and2s1 _____444391(.DIN1 (________25129), .DIN2 (________25392), .Q
       (________25393));
  nor2s1 ____0__444392(.DIN1 (_____0__25967), .DIN2 (________25066), .Q
       (________25391));
  nor2s1 ____0__444393(.DIN1 (________25389), .DIN2 (________25054), .Q
       (________25390));
  nor2s1 ____0__444394(.DIN1 (____9___24605), .DIN2 (________25056), .Q
       (________25388));
  nnd2s1 ____0_444395(.DIN1 (____0___25087), .DIN2 (________25052), .Q
       (_____0__25387));
  nnd2s1 _______444396(.DIN1 (________25057), .DIN2 (____99__21903), .Q
       (_____9__25386));
  or2s1 _______444397(.DIN1 (___9____25198), .DIN2 (________25069), .Q
       (________25385));
  nnd2s1 _______444398(.DIN1 (____0___25088), .DIN2 (inData[0]), .Q
       (________25384));
  nnd2s1 _______444399(.DIN1 (___0____25343), .DIN2 (outData[5]), .Q
       (________25383));
  nor2s1 _______444400(.DIN1 (________24762), .DIN2 (________25059), .Q
       (________25382));
  nnd2s1 _______444401(.DIN1 (________25092), .DIN2 (________25380), .Q
       (________25381));
  nnd2s1 _______444402(.DIN1 (_____0__25051), .DIN2 (________25378), .Q
       (________25379));
  and2s1 ______444403(.DIN1 (________25053), .DIN2 (________21850), .Q
       (_____0__25377));
  nnd2s1 _______444404(.DIN1 (____0___25085), .DIN2 (____0___24705), .Q
       (____09__25376));
  and2s1 _______444405(.DIN1 (____0___25086), .DIN2 (___0_0__24372), .Q
       (____0___25375));
  nor2s1 ______444406(.DIN1 (____0____30075), .DIN2 (_________30374),
       .Q (____0___25374));
  nnd2s1 _______444407(.DIN1 (________25097), .DIN2 (____0___24521), .Q
       (____0___25373));
  nnd2s1 ______444408(.DIN1 (________25096), .DIN2 (___0_09__27665), .Q
       (____0___25372));
  or2s1 _______444409(.DIN1 (____0___25370), .DIN2 (____9___25078), .Q
       (____0___25371));
  nor2s1 _______444410(.DIN1 (____9___25746), .DIN2 (____0___25084), .Q
       (____0___25369));
  nnd2s1 _____9_444411(.DIN1 (______0__34808), .DIN2 (________23929),
       .Q (____0___25368));
  and2s1 _____9_444412(.DIN1 (____9___25076), .DIN2 (___099__25366), .Q
       (____00__25367));
  and2s1 _____9_444413(.DIN1 (____9___25074), .DIN2 (_____0__25127), .Q
       (___09___25365));
  nor2s1 ____9__444414(.DIN1 (________24583), .DIN2 (____9___25072), .Q
       (___09___25364));
  or2s1 ____9__444415(.DIN1 (____9____30867), .DIN2 (_____0__25061), .Q
       (___09___25363));
  and2s1 ____9_444416(.DIN1 (_____9__25099), .DIN2 (___09___25361), .Q
       (___09___25362));
  nnd2s1 ____0__444417(.DIN1 (____09__25089), .DIN2 (________23938), .Q
       (___09___25360));
  and2s1 ____9__444418(.DIN1 (____0___25082), .DIN2 (___09___25358), .Q
       (___09___25359));
  nnd2s1 ____9__444419(.DIN1 (___0_9__25356), .DIN2 (__9__0__27005), .Q
       (___090__25357));
  or2s1 ____9_444420(.DIN1 (___0____25354), .DIN2 (________25062), .Q
       (___0____25355));
  nor2s1 ____9__444421(.DIN1 (________22922), .DIN2 (________25100), .Q
       (___0____25353));
  nor2s1 ____9_444422(.DIN1 (________24968), .DIN2 (____9___25077), .Q
       (___0____25352));
  nnd2s1 ____9__444423(.DIN1 (________25094), .DIN2 (________24531), .Q
       (___0____25351));
  nor2s1 ____9__444424(.DIN1 (__990___27084), .DIN2 (________25063), .Q
       (___0____25350));
  and2s1 ____9_444425(.DIN1 (________25091), .DIN2 (________26068), .Q
       (___0____25349));
  nor2s1 ____9__444426(.DIN1 (___9____22510), .DIN2 (____99__25079), .Q
       (___0____25348));
  nnd2s1 ____9__444427(.DIN1 (___0_9__25346), .DIN2 (________19453), .Q
       (___0_0__25347));
  nor2s1 ____00_444428(.DIN1 (___9____25246), .DIN2 (____0___25081), .Q
       (___0____25345));
  and2s1 ____00_444429(.DIN1 (________25065), .DIN2 (____0___25560), .Q
       (___0____25344));
  nor2s1 _____9_444430(.DIN1 (______18932), .DIN2 (____9___25551), .Q
       (_____9__25615));
  nnd2s1 _____0_444431(.DIN1
       (______________________________________0__________0__18892),
       .DIN2 (____0____30075), .Q (________25613));
  nnd2s1 _____0_444432(.DIN1 (________25150), .DIN2 (____0___24986), .Q
       (________25533));
  nnd2s1 _____9_444433(.DIN1 (____9___25551), .DIN2 (______9__28578),
       .Q (________25610));
  xor2s1 ____0__444434(.DIN1 (________25038), .DIN2 (___000___27171),
       .Q (________25636));
  nnd2s1 ____0__444435(.DIN1 (___0____25343), .DIN2 (____0___24987), .Q
       (_____0___28426));
  dffacs1 ___________________444436(.CLRB (reset), .CLK (clk), .DIN
       (________25093), .QN (_________________18685));
  nor2s1 _______444437(.DIN1 (________24644), .DIN2 (________25023), .Q
       (___0____25342));
  nnd2s1 _______444438(.DIN1 (________25000), .DIN2 (________24830), .Q
       (___0____25341));
  nor2s1 _____9_444439(.DIN1 (___0____22603), .DIN2 (________25030), .Q
       (___0____25340));
  nnd2s1 _______444440(.DIN1 (________24996), .DIN2 (____09__24992), .Q
       (___0____25339));
  nor2s1 _______444441(.DIN1 (___0____25324), .DIN2 (_____9__25021), .Q
       (___0_0__25338));
  or2s1 _______444442(.DIN1 (___0____25336), .DIN2 (________25028), .Q
       (___0_9__25337));
  nnd2s1 _______444443(.DIN1 (________25025), .DIN2 (________23147), .Q
       (___0____25335));
  nnd2s1 _______444444(.DIN1 (________25026), .DIN2 (___0____25333), .Q
       (___0____25334));
  nnd2s1 _______444445(.DIN1 (________25005), .DIN2 (__9_____27021), .Q
       (___0____25332));
  or2s1 ______444446(.DIN1 (_________28775), .DIN2 (________25024), .Q
       (___0____25331));
  and2s1 _______444447(.DIN1 (_____0__25022), .DIN2 (___0____25329), .Q
       (___0____25330));
  nor2s1 ______444448(.DIN1 (__990___27084), .DIN2 (________25009), .Q
       (___0_0__25328));
  nor2s1 _______444449(.DIN1 (________23948), .DIN2 (___0____25323), .Q
       (___0_9__25327));
  and2s1 _______444450(.DIN1 (________25019), .DIN2 (_____0__25520), .Q
       (___0____25326));
  nor2s1 _______444451(.DIN1 (___0____25324), .DIN2 (___0____25323), .Q
       (___0____25325));
  nnd2s1 ______444452(.DIN1 (________25016), .DIN2 (________23236), .Q
       (___0____25322));
  nnd2s1 _______444453(.DIN1 (_____0__25032), .DIN2 (________24220), .Q
       (___0____25321));
  or2s1 _______444454(.DIN1 (_________35060), .DIN2 (________25029), .Q
       (___0____25320));
  nor2s1 ______444455(.DIN1 (___0_9__25318), .DIN2 (________24994), .Q
       (___0_0__25319));
  nnd2s1 _____0_444456(.DIN1 (________24998), .DIN2 (_____0__24120), .Q
       (___0____25317));
  nor2s1 _______444457(.DIN1 (________23050), .DIN2 (_____9__25031), .Q
       (___0____25316));
  nnd2s1 _______444458(.DIN1 (________25048), .DIN2 (________24113), .Q
       (___0____25315));
  nnd2s1 _______444459(.DIN1 (________25018), .DIN2 (________25115), .Q
       (___0____25314));
  nnd2s1 _______444460(.DIN1 (________25003), .DIN2 (______0__34948),
       .Q (___0____25313));
  nnd2s1 _______444461(.DIN1 (_____0__25002), .DIN2 (__9_____26496), .Q
       (___0____25312));
  nor2s1 _______444462(.DIN1 (________24193), .DIN2 (________24999), .Q
       (___0____25311));
  nnd2s1 _______444463(.DIN1 (___________0___18872), .DIN2
       (_________28939), .Q (___0_0__25310));
  nor2s1 _______444464(.DIN1 (_________34974), .DIN2 (________24997),
       .Q (___0_9__25309));
  and2s1 _______444465(.DIN1 (________25008), .DIN2 (___0____25307), .Q
       (___0____25308));
  and2s1 ______444466(.DIN1 (_____9__24925), .DIN2 (___0____25305), .Q
       (___0____25306));
  nor2s1 _______444467(.DIN1 (___0____25303), .DIN2 (_____9__25011), .Q
       (___0____25304));
  nnd2s1 _______444468(.DIN1 (___0____25301), .DIN2
       (_______________18874), .Q (___0____25302));
  nor2s1 _______444469(.DIN1 (________25913), .DIN2 (________24995), .Q
       (___0_0__25300));
  and2s1 _______444470(.DIN1 (________24950), .DIN2 (________24177), .Q
       (___0_9__25299));
  nnd2s1 _______444471(.DIN1 (________24969), .DIN2 (_____9___34922),
       .Q (___0____25298));
  and2s1 _______444472(.DIN1 (________25036), .DIN2 (__9_____26962), .Q
       (___0____25297));
  nor2s1 ______444473(.DIN1 (____0___24990), .DIN2 (________25014), .Q
       (___0____25296));
  xor2s1 _____0_444474(.DIN1 (________22154), .DIN2
       (______________________________________0_____________18886), .Q
       (___0____25295));
  nor2s1 ______444475(.DIN1 (____09__22365), .DIN2 (_________34812), .Q
       (___0____25294));
  nnd2s1 _______444476(.DIN1 (_____9__24955), .DIN2 (________25447), .Q
       (___0____25293));
  nor2s1 _______444477(.DIN1 (___0____25354), .DIN2 (____0___24985), .Q
       (___0____25292));
  nor2s1 _______444478(.DIN1 (___0_0__25290), .DIN2 (____0___24989), .Q
       (___0____25291));
  and2s1 _______444479(.DIN1 (____9___24980), .DIN2 (___0____25288), .Q
       (___0_9__25289));
  nnd2s1 _______444480(.DIN1 (_____9__24935), .DIN2 (________24774), .Q
       (___0____25287));
  nor2s1 _______444481(.DIN1 (________26081), .DIN2 (_____0__24993), .Q
       (___0____25286));
  or2s1 _______444482(.DIN1 (___0____25284), .DIN2 (________24960), .Q
       (___0____25285));
  nor2s1 _______444483(.DIN1 (____09__22998), .DIN2 (____9___24977), .Q
       (___0____25283));
  nnd2s1 _______444484(.DIN1 (____99__24983), .DIN2 (___9____26230), .Q
       (___0____25282));
  and2s1 _______444485(.DIN1 (________24949), .DIN2 (___009__25280), .Q
       (___0_0__25281));
  nnd2s1 _______444486(.DIN1 (________25013), .DIN2 (________24777), .Q
       (___00___25279));
  nnd2s1 _______444487(.DIN1 (________24961), .DIN2 (____00__21904), .Q
       (___00___25278));
  nor2s1 _______444488(.DIN1 (__9_____26713), .DIN2 (________25042), .Q
       (___00___25277));
  xor2s1 _____0_444489(.DIN1 (___________0___18877), .DIN2
       (_______________18879), .Q (__9_____26368));
  nnd2s1 _____444490(.DIN1 (________25034), .DIN2 (________25604), .Q
       (________25573));
  nnd2s1 _____9_444491(.DIN1 (_______________18873), .DIN2
       (___________0___18872), .Q (________25611));
  nnd2s1 _____9_444492(.DIN1 (_______________18874), .DIN2
       (_________29585), .Q (________25612));
  nor2s1 _____9_444493(.DIN1 (___________0___18872), .DIN2
       (______________________________________0__________0), .Q
       (________25614));
  dffacs1 ___________________444494(.CLRB (reset), .CLK (clk), .DIN
       (________24938), .QN (______0__18865));
  nor2s1 ____444495(.DIN1 (___0____24408), .DIN2 (________24948), .Q
       (___00___25276));
  nnd2s1 _______444496(.DIN1 (____0___24991), .DIN2 (________22091), .Q
       (___00___25275));
  or2s1 _____9_444497(.DIN1 (___00___25273), .DIN2 (________24952), .Q
       (___00___25274));
  or2s1 ____90_444498(.DIN1 (_____9__25415), .DIN2 (________24962), .Q
       (___00___25272));
  and2s1 ____90_444499(.DIN1 (________24918), .DIN2 (_____9__24973), .Q
       (___000__25271));
  and2s1 ____444500(.DIN1 (________24972), .DIN2 (__9__0__26394), .Q
       (___999__25270));
  nnd2s1 ____9__444501(.DIN1 (________24971), .DIN2 (___99___25268), .Q
       (___99___25269));
  nor2s1 ____9__444502(.DIN1 (___9____23421), .DIN2 (____0___24988), .Q
       (___99___25267));
  nor2s1 ____9__444503(.DIN1 (________25710), .DIN2 (________25039), .Q
       (___99___25266));
  nnd2s1 ____9__444504(.DIN1 (___99___25264), .DIN2 (___99___25263), .Q
       (___99___25265));
  or2s1 _______444505(.DIN1 (___990__25261), .DIN2 (________25045), .Q
       (___99___25262));
  nor2s1 ____9__444506(.DIN1 (________24170), .DIN2 (___9____25225), .Q
       (___9_9__25260));
  nor2s1 ____9__444507(.DIN1 (________24232), .DIN2 (________25037), .Q
       (___9____25259));
  nnd2s1 ____9_444508(.DIN1 (________24686), .DIN2 (________24942), .Q
       (___9____25258));
  nnd2s1 ____9__444509(.DIN1 (____00__24984), .DIN2 (________22766), .Q
       (___9____25257));
  nnd2s1 ____9__444510(.DIN1 (________24951), .DIN2 (________25068), .Q
       (___9____25256));
  nnd2s1 ____9__444511(.DIN1 (________24963), .DIN2 (____0___24890), .Q
       (___9____25255));
  nor2s1 ____9__444512(.DIN1 (____00__24429), .DIN2 (________24933), .Q
       (___9____25254));
  nor2s1 ____9_444513(.DIN1 (________24958), .DIN2 (________24455), .Q
       (___9____25253));
  nnd2s1 ____9_444514(.DIN1 (________24953), .DIN2 (________24912), .Q
       (___9____25252));
  or2s1 ____9__444515(.DIN1 (__9_____26671), .DIN2 (________24930), .Q
       (___9_0__25251));
  or2s1 ____9__444516(.DIN1 (___9____25249), .DIN2 (_____9__24945), .Q
       (___9_9__25250));
  nnd2s1 ____9__444517(.DIN1 (________24922), .DIN2 (___00___23442), .Q
       (___9____25248));
  nor2s1 ____9__444518(.DIN1 (___9____25246), .DIN2 (________24957), .Q
       (___9____25247));
  nor2s1 ____9__444519(.DIN1
       (______________________________________0_____________18887),
       .DIN2 (________25417), .Q (___9____25245));
  nor2s1 ____444520(.DIN1 (________25101), .DIN2 (________24966), .Q
       (___9____25244));
  nor2s1 ____99_444521(.DIN1 (________24932), .DIN2 (________24444), .Q
       (___9____25243));
  nor2s1 ____99_444522(.DIN1 (___9_0__25241), .DIN2 (________24941), .Q
       (___9____25242));
  nor2s1 ____99_444523(.DIN1 (________25516), .DIN2 (____9___24982), .Q
       (___9_9__25240));
  nor2s1 ____99_444524(.DIN1 (_________31281), .DIN2 (________25417),
       .Q (___9____25239));
  or2s1 _______444525(.DIN1 (___9____25237), .DIN2 (________24934), .Q
       (___9____25238));
  nnd2s1 ____00_444526(.DIN1 (________24927), .DIN2 (___0____21654), .Q
       (___9____25236));
  nnd2s1 ____00_444527(.DIN1 (________24928), .DIN2 (_____9__25118), .Q
       (___9____25235));
  or2s1 ____444528(.DIN1 (____9___19395), .DIN2 (___9____25233), .Q
       (___9____25234));
  or2s1 ____0_444529(.DIN1 (___9_0__25231), .DIN2 (_____0__24926), .Q
       (___9____25232));
  nor2s1 ____0__444530(.DIN1 (___90___26154), .DIN2 (________24920), .Q
       (___9_9__25230));
  nor2s1 ____0__444531(.DIN1 (________25015), .DIN2 (____90__24974), .Q
       (___9____25229));
  or2s1 ____0__444532(.DIN1 (________25417), .DIN2 (____9____31759), .Q
       (___9____25228));
  nnd2s1 ____0__444533(.DIN1 (________24947), .DIN2 (__9_____26875), .Q
       (___9____25227));
  or2s1 ____0_444534(.DIN1 (___0_9___27848), .DIN2 (___9____25225), .Q
       (___9____25226));
  and2s1 ____0_444535(.DIN1 (________24937), .DIN2 (___9____25223), .Q
       (___9____25224));
  nnd2s1 ____0__444536(.DIN1 (________24940), .DIN2 (_________35010),
       .Q (___9____25222));
  and2s1 ____0__444537(.DIN1 (____0____32762), .DIN2 (________25417),
       .Q (___9_0__25221));
  xor2s1 ____0__444538(.DIN1 (___9_9__19754), .DIN2 (_________28661),
       .Q (___9_9__25220));
  nnd2s1 _____9_444539(.DIN1 (________24910), .DIN2 (________23866), .Q
       (___9____25219));
  nnd2s1 ____0__444540(.DIN1 (_____9__26006), .DIN2 (_____00__30456),
       .Q (___9____25218));
  nor2s1 _______444541(.DIN1 (____0___24431), .DIN2 (___9____25216), .Q
       (___9____25217));
  nnd2s1 _______444542(.DIN1 (________24913), .DIN2 (________25058), .Q
       (___9____25215));
  nor2s1 ____09_444543(.DIN1 (________24914), .DIN2 (___9____25213), .Q
       (___9____25214));
  xnr2s1 ____0_444544(.DIN1 (___9_0__25211), .DIN2 (_____0___32851), .Q
       (___9____25212));
  nor2s1 ____0__444545(.DIN1 (________24924), .DIN2 (____9___24789), .Q
       (___9_9__25210));
  and2s1 ____0__444546(.DIN1 (________24917), .DIN2 (___9____25208), .Q
       (___9____25209));
  nor2s1 ____0_444547(.DIN1 (___9____25206), .DIN2 (_____9__24964), .Q
       (___9____25207));
  nnd2s1 _______444548(.DIN1 (________25047), .DIN2 (___0__9__27879),
       .Q (__99____27128));
  nor2s1 _______444549(.DIN1 (__9_____26553), .DIN2 (________24911), .Q
       (________25494));
  nor2s1 ____0__444550(.DIN1 (_________31388), .DIN2 (_____9__26006),
       .Q (________25507));
  nor2s1 ____0__444551(.DIN1 (________25417), .DIN2 (____0____32762),
       .Q (________25490));
  nor2s1 ____0__444552(.DIN1 (_____00__30456), .DIN2 (_____9__26006),
       .Q (________25897));
  nor2s1 ____0__444553(.DIN1
       (______________________________________0_____________18888),
       .DIN2 (_____9__26006), .Q (________25504));
  nnd2s1 ____9__444554(.DIN1 (_____9__25050), .DIN2 (___9____25205), .Q
       (________25609));
  nnd2s1 _____444555(.DIN1 (____0___24800), .DIN2 (___9____23402), .Q
       (___9____25204));
  nor2s1 ____9__444556(.DIN1 (___9_9__25202), .DIN2 (________24807), .Q
       (___9_0__25203));
  nor2s1 ____9__444557(.DIN1 (___9____25200), .DIN2 (_____0__24867), .Q
       (___9____25201));
  or2s1 ____90_444558(.DIN1 (____9___23709), .DIN2 (________24840), .Q
       (___9____25199));
  nor2s1 ____9__444559(.DIN1 (___90___24245), .DIN2 (________24863), .Q
       (___9____25197));
  nnd2s1 _______444560(.DIN1 (________24907), .DIN2 (___9____25195), .Q
       (___9____25196));
  nnd2s1 _______444561(.DIN1 (________24831), .DIN2 (________23040), .Q
       (___9_0__25194));
  nnd2s1 ______444562(.DIN1 (________24834), .DIN2 (____09__22270), .Q
       (___9_9__25193));
  nor2s1 ______444563(.DIN1 (_____0__24541), .DIN2 (____9___24882), .Q
       (___9____25192));
  and2s1 _______444564(.DIN1 (____9___24883), .DIN2 (________25641), .Q
       (___9____25191));
  and2s1 ______444565(.DIN1 (_____9__24771), .DIN2 (________25991), .Q
       (___9____25190));
  nor2s1 _______444566(.DIN1 (_____9___34926), .DIN2 (____9___24879),
       .Q (___9____25189));
  nnd2s1 _______444567(.DIN1 (________24870), .DIN2 (________23922), .Q
       (___9____25188));
  or2s1 ______444568(.DIN1 (___9____25186), .DIN2 (____9___24878), .Q
       (___9____25187));
  nor2s1 _______444569(.DIN1 (___9_0__25184), .DIN2 (________24810), .Q
       (___9____25185));
  nor2s1 ______444570(.DIN1 (__90____26312), .DIN2 (________24849), .Q
       (___909__25183));
  nor2s1 ______444571(.DIN1 (____9___23254), .DIN2 (________24835), .Q
       (___90___25182));
  nnd2s1 _______444572(.DIN1 (________24875), .DIN2 (___90___25180), .Q
       (___90___25181));
  nnd2s1 _______444573(.DIN1 (________24872), .DIN2 (________24115), .Q
       (___90___25179));
  nnd2s1 _______444574(.DIN1 (____0___24799), .DIN2 (____09__22815), .Q
       (___90___25178));
  nnd2s1 _______444575(.DIN1 (________24869), .DIN2 (__9_____26447), .Q
       (___90___25177));
  nnd2s1 _______444576(.DIN1 (________24868), .DIN2 (________26089), .Q
       (___90___25176));
  nnd2s1 _______444577(.DIN1 (____0___24892), .DIN2 (____9___23795), .Q
       (___90___25175));
  nor2s1 _______444578(.DIN1 (___9____22520), .DIN2 (________24826), .Q
       (___900__25174));
  or2s1 _______444579(.DIN1 (__9_9___26505), .DIN2 (_____9__24866), .Q
       (____99__25173));
  nnd2s1 _______444580(.DIN1 (_____9__24857), .DIN2 (________22967), .Q
       (____9___25172));
  nor2s1 _______444581(.DIN1 (_____9__25829), .DIN2 (____9___24885), .Q
       (____9___25171));
  nnd2s1 ______444582(.DIN1 (________24856), .DIN2 (____9___25168), .Q
       (____9___25169));
  and2s1 _____444583(.DIN1 (________24841), .DIN2 (____9___23344), .Q
       (____9___25167));
  or2s1 _____9_444584(.DIN1 (________24002), .DIN2 (____90__25165), .Q
       (____9___25166));
  and2s1 _____9_444585(.DIN1 (________24862), .DIN2 (___0____25305), .Q
       (_____9__25164));
  nor2s1 _____9_444586(.DIN1 (___9____24260), .DIN2 (________24853), .Q
       (________25163));
  nnd2s1 ____444587(.DIN1 (________24873), .DIN2 (_____0__24481), .Q
       (________25162));
  or2s1 ____90_444588(.DIN1 (_____0__25616), .DIN2 (________24846), .Q
       (________25161));
  nnd2s1 ____90_444589(.DIN1 (________24673), .DIN2 (________24844), .Q
       (________25160));
  nnd2s1 ____90_444590(.DIN1 (________24825), .DIN2 (________25158), .Q
       (________25159));
  or2s1 ____90_444591(.DIN1 (_____0__25156), .DIN2 (________24843), .Q
       (________25157));
  or2s1 ____9__444592(.DIN1 (________25710), .DIN2 (_____9__24808), .Q
       (_____9__25155));
  and2s1 ____9__444593(.DIN1 (____9___24881), .DIN2 (________24185), .Q
       (________25154));
  nor2s1 ____9_444594(.DIN1 (_____9__24578), .DIN2 (_________34814), .Q
       (________25153));
  nnd2s1 ____9__444595(.DIN1 (____9___24880), .DIN2 (________25098), .Q
       (________25152));
  nnd2s1 ____9__444596(.DIN1 (________24860), .DIN2 (____0___21911), .Q
       (________25151));
  xor2s1 ____9__444597(.DIN1 (________24586), .DIN2 (_____0__19985), .Q
       (________25150));
  or2s1 ____9__444598(.DIN1 (________25148), .DIN2 (________24823), .Q
       (________25149));
  and2s1 ____9__444599(.DIN1 (________24837), .DIN2 (___9____25208), .Q
       (________25147));
  or2s1 ____9__444600(.DIN1 (_____9__25145), .DIN2 (_____0__24829), .Q
       (_____0__25146));
  nnd2s1 ____9__444601(.DIN1 (________24851), .DIN2 (________22150), .Q
       (________25144));
  nnd2s1 ____9__444602(.DIN1 (________25142), .DIN2
       (_______________18879), .Q (________25143));
  and2s1 ____9__444603(.DIN1 (________24802), .DIN2 (________25447), .Q
       (________25141));
  and2s1 ____9__444604(.DIN1 (_________34816), .DIN2 (________25139),
       .Q (________25140));
  nor2s1 ____9__444605(.DIN1 (________25137), .DIN2 (____0___24891), .Q
       (________25138));
  or2s1 ____9__444606(.DIN1 (__9_9___26414), .DIN2 (____0___24797), .Q
       (_____0__25136));
  nnd2s1 ____9__444607(.DIN1 (____0___24887), .DIN2 (____09__22181), .Q
       (_____9__25135));
  nnd2s1 ____9__444608(.DIN1 (____0___24889), .DIN2 (___0____24403), .Q
       (________25134));
  nnd2s1 ____9__444609(.DIN1 (_____90__34818), .DIN2 (________25132),
       .Q (________25133));
  nor2s1 ____9_444610(.DIN1 (________24207), .DIN2 (________24816), .Q
       (________25131));
  or2s1 ____9__444611(.DIN1 (________25137), .DIN2 (________24813), .Q
       (________25130));
  nor2s1 ____9__444612(.DIN1 (________26072), .DIN2 (________24815), .Q
       (________25129));
  nnd2s1 ____9__444613(.DIN1 (_____0__24848), .DIN2 (________24073), .Q
       (________25128));
  nnd2s1 ____9__444614(.DIN1 (_____0__25127), .DIN2 (________24482), .Q
       (___0_____27539));
  and2s1 _______444615(.DIN1 (___0_____27690), .DIN2 (____9___24509),
       .Q (___099__25366));
  dffacs1 ___________________444616(.CLRB (reset), .CLK (clk), .DIN
       (________24898), .QN
       (______________0______________________18824));
  hi1s1 _____444617(.DIN (_______________18874), .Q (____0____30075));
  hi1s1 ______444618(.DIN (___________0___18872), .Q (____9___25551));
  nnd2s1 ____9__444619(.DIN1 (________24803), .DIN2 (_____0__24560), .Q
       (_____9__25126));
  nor2s1 ____9_444620(.DIN1 (_________31926), .DIN2
       (______________________________________0_____________18886), .Q
       (________25125));
  nor2s1 ____99_444621(.DIN1
       (______________________________________0_____________18886),
       .DIN2
       (______________________________________0_____________18889), .Q
       (________25124));
  nor2s1 ____00_444622(.DIN1 (___9____24314), .DIN2 (________24805), .Q
       (________25122));
  nor2s1 ____00_444623(.DIN1 (___099__22625), .DIN2 (____0___24796), .Q
       (________25121));
  nnd2s1 ____0__444624(.DIN1 (__99____27118), .DIN2
       (_______________18879), .Q (________25120));
  nnd2s1 ____0__444625(.DIN1 (________25116), .DIN2 (_____9__25118), .Q
       (_____0__25119));
  and2s1 ____0__444626(.DIN1 (________25116), .DIN2 (________25115), .Q
       (________25117));
  nnd2s1 ____0__444627(.DIN1 (____09__24801), .DIN2 (________23145), .Q
       (________25114));
  or2s1 ____0__444628(.DIN1 (__90____26312), .DIN2 (________25112), .Q
       (________25113));
  or2s1 ____0__444629(.DIN1 (________24836), .DIN2 (________25110), .Q
       (________25111));
  or2s1 ____0__444630(.DIN1 (___9_0__25231), .DIN2 (________24832), .Q
       (_____0__25109));
  nnd2s1 ____0__444631(.DIN1 (________25107), .DIN2 (_____0__24739), .Q
       (_____9__25108));
  hi1s1 _____0_444632(.DIN (________25105), .Q (________25106));
  nor2s1 ____0_444633(.DIN1 (_____00__30456), .DIN2
       (______________________________________0_____________18886), .Q
       (________25104));
  xor2s1 _____444634(.DIN1 (____9____30860), .DIN2 (_____9___30627), .Q
       (________25103));
  nor2s1 ____0_444635(.DIN1 (________25101), .DIN2 (_____0__24965), .Q
       (________25102));
  nor2s1 _______444636(.DIN1 (____09__22634), .DIN2 (________24897), .Q
       (________25100));
  and2s1 ____0__444637(.DIN1 (____9___24786), .DIN2 (________25098), .Q
       (_____9__25099));
  nor2s1 ____0_444638(.DIN1 (____9___24236), .DIN2 (________24767), .Q
       (________25097));
  nor2s1 ____0__444639(.DIN1 (________25095), .DIN2 (_____0__24906), .Q
       (________25096));
  or2s1 ____0__444640(.DIN1 (______________18868), .DIN2
       (____9___24785), .Q (________25094));
  nnd2s1 ____0__444641(.DIN1 (____9___24787), .DIN2 (________24442), .Q
       (________25093));
  and2s1 ____0__444642(.DIN1 (_____9___34824), .DIN2 (_____0__22128),
       .Q (________25092));
  and2s1 ____0__444643(.DIN1 (________24750), .DIN2 (_____0__25090), .Q
       (________25091));
  nor2s1 ____0__444644(.DIN1 (___9____24250), .DIN2 (________24776), .Q
       (____09__25089));
  nor2s1 ____0__444645(.DIN1 (___9_0__25211), .DIN2 (________22048), .Q
       (____0___25088));
  nor2s1 ____0__444646(.DIN1 (________24909), .DIN2 (________24779), .Q
       (____0___25087));
  nor2s1 ____09_444647(.DIN1 (_____0__24636), .DIN2 (________24770), .Q
       (____0___25086));
  nor2s1 ____09_444648(.DIN1 (________25483), .DIN2 (____09__24895), .Q
       (____0___25085));
  or2s1 ____09_444649(.DIN1 (___9____25198), .DIN2 (_____9__24818), .Q
       (____0___25084));
  nnd2s1 _____444650(.DIN1 (________24900), .DIN2 (_____9__24043), .Q
       (____0___25083));
  and2s1 _____0_444651(.DIN1 (________24768), .DIN2 (___0____25288), .Q
       (____0___25082));
  nnd2s1 _____0_444652(.DIN1 (________24861), .DIN2 (___9____24273), .Q
       (____0___25081));
  nnd2s1 _______444653(.DIN1 (________24766), .DIN2 (_________32156),
       .Q (____00__25080));
  nnd2s1 ______444654(.DIN1 (________24899), .DIN2 (________22770), .Q
       (____99__25079));
  nnd2s1 _______444655(.DIN1 (________24763), .DIN2 (________24122), .Q
       (____9___25078));
  nnd2s1 _______444656(.DIN1 (________24761), .DIN2 (________24760), .Q
       (____9___25077));
  nor2s1 ______444657(.DIN1 (________24759), .DIN2 (____9___25075), .Q
       (____9___25076));
  nor2s1 _______444658(.DIN1 (________24445), .DIN2 (____9___25073), .Q
       (____9___25074));
  or2s1 _______444659(.DIN1 (________22822), .DIN2 (________24758), .Q
       (____9___25072));
  or2s1 ______444660(.DIN1 (outData[4]), .DIN2 (________24769), .Q
       (_____9__25070));
  nnd2s1 _____9_444661(.DIN1 (_____9___34822), .DIN2 (________25068),
       .Q (________25069));
  nor2s1 _____444662(.DIN1 (_____0__24756), .DIN2 (________24734), .Q
       (________25067));
  nnd2s1 ______444663(.DIN1 (________24903), .DIN2 (________25923), .Q
       (________25066));
  nor2s1 _______444664(.DIN1 (________25064), .DIN2 (________24748), .Q
       (________25065));
  nor2s1 _______444665(.DIN1 (____0___24160), .DIN2 (_____0__24764), .Q
       (________25063));
  nnd2s1 _______444666(.DIN1 (________24773), .DIN2 (________24712), .Q
       (________25062));
  nnd2s1 _______444667(.DIN1 (________20579), .DIN2 (_____0__24896), .Q
       (_____0__25061));
  nnd2s1 _______444668(.DIN1 (____9___19200), .DIN2 (_________28661),
       .Q (_____9__25060));
  nnd2s1 ______444669(.DIN1 (____9___24790), .DIN2 (________25058), .Q
       (________25059));
  nor2s1 _______444670(.DIN1 (__9_____26650), .DIN2 (____0___24793), .Q
       (________25057));
  nnd2s1 _______444671(.DIN1 (________24901), .DIN2 (________24452), .Q
       (________25056));
  and2s1 _______444672(.DIN1 (____9___24788), .DIN2 (___9____25223), .Q
       (________25055));
  nnd2s1 _______444673(.DIN1 (________24778), .DIN2 (__9_____26489), .Q
       (________25054));
  and2s1 ______444674(.DIN1 (_____9__24781), .DIN2 (________25052), .Q
       (________25053));
  nor2s1 _______444675(.DIN1 (________24680), .DIN2 (____0___24894), .Q
       (_____0__25051));
  nnd2s1 ____0__444676(.DIN1 (_______________18879), .DIN2
       (_________33835), .Q (________26070));
  hi1s1 ____0__444677(.DIN (_____9__25050), .Q (___0____25343));
  nnd2s1 _____9_444678(.DIN1 (________24747), .DIN2 (____0___21912), .Q
       (___0_9__25356));
  and2s1 _____9_444679(.DIN1 (_____9__24905), .DIN2 (________25049), .Q
       (___0_____27725));
  nnd2s1 _____0_444680(.DIN1 (____90__24782), .DIN2 (___9____24301), .Q
       (___0_9__25346));
  nor2s1 ____0__444681(.DIN1 (_______________18879), .DIN2
       (_____9___30627), .Q (________25503));
  nor2s1 ____0_444682(.DIN1 (_______________18879), .DIN2
       (_______________18880), .Q (________25506));
  nor2s1 ____9__444683(.DIN1 (____90__26137), .DIN2 (________24713), .Q
       (________25048));
  and2s1 _______444684(.DIN1 (________25046), .DIN2 (_____9__24675), .Q
       (________25047));
  nnd2s1 _______444685(.DIN1 (_____0___34832), .DIN2 (________25044),
       .Q (________25045));
  nor2s1 _______444686(.DIN1 (________24574), .DIN2 (_____9__24208), .Q
       (________25043));
  nnd2s1 ______444687(.DIN1 (_____0__25041), .DIN2 (_____9__24198), .Q
       (________25042));
  nor2s1 _______444688(.DIN1 (____0___24610), .DIN2 (_____9__24081), .Q
       (_____9__25040));
  nnd2s1 _______444689(.DIN1 (____9___24606), .DIN2 (____00__24701), .Q
       (________25039));
  nor2s1 _______444690(.DIN1 (_________18852), .DIN2 (_____9___30627),
       .Q (________25038));
  nnd2s1 _______444691(.DIN1 (_____9__24587), .DIN2 (______0__34968),
       .Q (________25037));
  nnd2s1 ______444692(.DIN1 (_____0___34834), .DIN2 (________25035), .Q
       (________25036));
  nor2s1 _______444693(.DIN1 (________25033), .DIN2 (________24663), .Q
       (________25034));
  nor2s1 ______444694(.DIN1 (________24821), .DIN2 (________24670), .Q
       (_____0__25032));
  nnd2s1 _______444695(.DIN1 (_____9__24665), .DIN2 (___9____22506), .Q
       (_____9__25031));
  nnd2s1 _______444696(.DIN1 (________24653), .DIN2 (________24619), .Q
       (________25030));
  nnd2s1 _______444697(.DIN1 (________24667), .DIN2 (_____0__24956), .Q
       (________25029));
  or2s1 _______444698(.DIN1 (________25027), .DIN2 (________24672), .Q
       (________25028));
  nor2s1 _______444699(.DIN1 (________25985), .DIN2 (________24657), .Q
       (________25026));
  nor2s1 ______444700(.DIN1 (___0_0__23481), .DIN2 (____90__24693), .Q
       (________25025));
  nnd2s1 _______444701(.DIN1 (________24641), .DIN2 (_____0__23231), .Q
       (________25024));
  or2s1 _______444702(.DIN1 (________25123), .DIN2 (________24711), .Q
       (________25023));
  and2s1 _______444703(.DIN1 (____9___24696), .DIN2 (___9____23373), .Q
       (_____0__25022));
  or2s1 _______444704(.DIN1 (________23761), .DIN2 (________25020), .Q
       (_____9__25021));
  and2s1 _______444705(.DIN1 (____0___24708), .DIN2 (_____0__24646), .Q
       (________25019));
  nor2s1 ____9_444706(.DIN1 (________24724), .DIN2 (________24714), .Q
       (________25018));
  or2s1 ____9__444707(.DIN1 (__90____26312), .DIN2 (________24715), .Q
       (________25017));
  nor2s1 ____9__444708(.DIN1 (________25015), .DIN2 (____09__24709), .Q
       (________25016));
  or2s1 _____0_444709(.DIN1 (___9____23371), .DIN2 (____0___24609), .Q
       (________25014));
  and2s1 ____09_444710(.DIN1 (____0___24614), .DIN2 (____9___24981), .Q
       (________25013));
  nnd2s1 ____0__444711(.DIN1 (________24658), .DIN2 (______9__32271),
       .Q (_____0__25012));
  or2s1 ____9_444712(.DIN1 (________25010), .DIN2 (____9___24694), .Q
       (_____9__25011));
  nor2s1 ____9__444713(.DIN1 (_____0__24746), .DIN2 (________24647), .Q
       (________25009));
  and2s1 ____9__444714(.DIN1 (________24652), .DIN2 (________25007), .Q
       (________25008));
  nor2s1 _______444715(.DIN1 (_______________18884), .DIN2
       (_____0__24684), .Q (________25006));
  and2s1 ____9__444716(.DIN1 (_____9__24645), .DIN2 (________25004), .Q
       (________25005));
  nor2s1 ____9__444717(.DIN1 (________23749), .DIN2 (________24640), .Q
       (________25003));
  nor2s1 ____9_444718(.DIN1 (_____9__25001), .DIN2 (________24649), .Q
       (_____0__25002));
  nor2s1 ____9__444719(.DIN1 (________22212), .DIN2 (________24654), .Q
       (________25000));
  nnd2s1 ____9__444720(.DIN1 (________24639), .DIN2 (________23234), .Q
       (________24999));
  and2s1 ____99_444721(.DIN1 (________24643), .DIN2 (_________34956),
       .Q (________24998));
  nnd2s1 ____99_444722(.DIN1 (________24648), .DIN2 (________23871), .Q
       (________24997));
  nor2s1 ____0__444723(.DIN1 (________25148), .DIN2 (_____0__24656), .Q
       (________24996));
  or2s1 ____0__444724(.DIN1 (__9__0__26485), .DIN2 (________24650), .Q
       (________24995));
  or2s1 ____0__444725(.DIN1 (____9___26142), .DIN2 (________24671), .Q
       (________24994));
  nnd2s1 ____0_444726(.DIN1 (________24717), .DIN2 (____09__24992), .Q
       (_____0__24993));
  nor2s1 ____0__444727(.DIN1 (____0___24990), .DIN2 (________24617), .Q
       (____0___24991));
  nnd2s1 ____0_444728(.DIN1 (________24633), .DIN2 (______0__34948), .Q
       (____0___24989));
  and2s1 ____0__444729(.DIN1 (________24634), .DIN2 (________24221), .Q
       (____0___24988));
  nnd2s1 ____0__444730(.DIN1 (____0___24986), .DIN2 (outData[4]), .Q
       (____0___24987));
  or2s1 ____0__444731(.DIN1 (__9_____26487), .DIN2 (________24596), .Q
       (____0___24985));
  and2s1 ____0_444732(.DIN1 (________24631), .DIN2 (______0__34968), .Q
       (____00__24984));
  nor2s1 ____0__444733(.DIN1 (________26000), .DIN2 (________24620), .Q
       (____99__24983));
  nnd2s1 ____0__444734(.DIN1 (________24630), .DIN2 (____9___24981), .Q
       (____9___24982));
  and2s1 ____0__444735(.DIN1 (___0____24384), .DIN2 (_________34840),
       .Q (____9___24980));
  nor2s1 _____0_444736(.DIN1 (________24683), .DIN2 (________24692), .Q
       (___0_____27612));
  and2s1 _____0_444737(.DIN1 (________24678), .DIN2 (___09____28113),
       .Q (_________28278));
  nnd2s1 ____9__444738(.DIN1 (____0___24707), .DIN2 (__9__9__27014), .Q
       (___0____25323));
  nnd2s1 ______444739(.DIN1 (____9___24979), .DIN2 (____0___24433), .Q
       (___9____25216));
  hi1s1 ____0__444740(.DIN (_______________18879), .Q (_____9__26006));
  hi1s1 ____0__444741(.DIN
       (______________________________________0_____________18886), .Q
       (________25417));
  dffacs1 _________________444742(.CLRB (reset), .CLK (clk), .DIN
       (________24618), .QN (______________18869));
  dffacs1 _________________444743(.CLRB (reset), .CLK (clk), .DIN
       (________24622), .QN (______________18870));
  dffacs2 ________________0_444744(.CLRB (reset), .CLK (clk), .DIN
       (________24668), .Q (___________0___18872));
  dffacs2 __________________444745(.CLRB (reset), .CLK (clk), .DIN
       (________24664), .Q (_______________18874));
  nor2s1 _______444746(.DIN1
       (______________________________________0_____________18890),
       .DIN2 (_____9___30627), .Q (____9___24978));
  nnd2s1 ______444747(.DIN1 (________24624), .DIN2 (___0____23465), .Q
       (____9___24977));
  or2s1 ______444748(.DIN1 (________24728), .DIN2 (____99__24700), .Q
       (____9___24976));
  or2s1 _______444749(.DIN1 (____9___24699), .DIN2 (________24595), .Q
       (____9___24975));
  nnd2s1 _______444750(.DIN1 (________24573), .DIN2 (____0___23620), .Q
       (____90__24974));
  nor2s1 _______444751(.DIN1 (________24582), .DIN2 (________24730), .Q
       (_____9__24973));
  and2s1 _______444752(.DIN1 (________24590), .DIN2 (________24591), .Q
       (________24972));
  and2s1 _______444753(.DIN1 (_________34840), .DIN2 (________24970),
       .Q (________24971));
  nor2s1 _______444754(.DIN1 (___9____24265), .DIN2 (____9___24599), .Q
       (________24969));
  nnd2s1 _______444755(.DIN1 (________24674), .DIN2 (_____0__23134), .Q
       (________24968));
  nnd2s1 _____0_444756(.DIN1 (________24224), .DIN2 (________24690), .Q
       (________24967));
  hi1s1 ______444757(.DIN (_____0__24965), .Q (________24966));
  or2s1 _____9_444758(.DIN1 (________26125), .DIN2 (____0___24706), .Q
       (_____9__24964));
  and2s1 _______444759(.DIN1 (________25098), .DIN2 (_____0__24579), .Q
       (________24963));
  nnd2s1 ______444760(.DIN1 (________24565), .DIN2 (___0____25305), .Q
       (________24962));
  nor2s1 _____9_444761(.DIN1 (________25015), .DIN2 (________24575), .Q
       (________24961));
  or2s1 _____9_444762(.DIN1 (________24959), .DIN2 (_____0__24626), .Q
       (________24960));
  nor2s1 _____9_444763(.DIN1 (_____0__25616), .DIN2 (______0__34838),
       .Q (________24958));
  nnd2s1 _____444764(.DIN1 (____9___24603), .DIN2 (___090__22617), .Q
       (________24957));
  nor2s1 _____0_444765(.DIN1 (________25010), .DIN2 (________24723), .Q
       (_____9__24955));
  nor2s1 _____0_444766(.DIN1 (________24576), .DIN2 (_____9__24755), .Q
       (________24954));
  nor2s1 _______444767(.DIN1 (________24780), .DIN2 (________24623), .Q
       (________24953));
  nnd2s1 ______444768(.DIN1 (________24731), .DIN2 (________22735), .Q
       (________24952));
  nor2s1 ______444769(.DIN1 (___9____23367), .DIN2 (________24584), .Q
       (________24951));
  nor2s1 _______444770(.DIN1 (_____0__24946), .DIN2 (________24727), .Q
       (________24950));
  nor2s1 _______444771(.DIN1 (________22704), .DIN2 (________24621), .Q
       (________24949));
  nnd2s1 _______444772(.DIN1 (________24594), .DIN2 (________22687), .Q
       (________24948));
  nor2s1 _______444773(.DIN1 (_____0__24946), .DIN2 (________24732), .Q
       (________24947));
  nnd2s1 _______444774(.DIN1 (____09__24615), .DIN2 (________24944), .Q
       (_____9__24945));
  nor2s1 ______444775(.DIN1 (_________34976), .DIN2 (____9___24604), .Q
       (________24943));
  nnd2s1 _______444776(.DIN1 (________23903), .DIN2 (_____0___34836),
       .Q (________24942));
  nnd2s1 _______444777(.DIN1 (________24736), .DIN2 (________25004), .Q
       (________24941));
  and2s1 _______444778(.DIN1 (________24737), .DIN2 (________24939), .Q
       (________24940));
  nnd2s1 _______444779(.DIN1 (_________32156), .DIN2 (____9___24602),
       .Q (________24938));
  nor2s1 ______444780(.DIN1 (_____0__24936), .DIN2 (____0___24612), .Q
       (________24937));
  nor2s1 ______444781(.DIN1 (____0___21990), .DIN2 (________24581), .Q
       (_____9__24935));
  nnd2s1 _______444782(.DIN1 (____00__24608), .DIN2 (________23931), .Q
       (________24934));
  nor2s1 _______444783(.DIN1 (_____0__24720), .DIN2 (________24733), .Q
       (________24933));
  nor2s1 _______444784(.DIN1 (________24589), .DIN2 (________24931), .Q
       (________24932));
  or2s1 ______444785(.DIN1 (________24929), .DIN2 (________24718), .Q
       (________24930));
  and2s1 _______444786(.DIN1 (________24572), .DIN2 (____9___25460), .Q
       (________24928));
  nnd2s1 _______444787(.DIN1 (____0___24613), .DIN2 (__99____27157), .Q
       (________24927));
  nnd2s1 _______444788(.DIN1 (_____0__24570), .DIN2 (_____0__24008), .Q
       (_____0__24926));
  and2s1 _______444789(.DIN1 (_____0__24729), .DIN2 (_____0__25665), .Q
       (_____9__24925));
  nor2s1 _______444790(.DIN1 (_____0___31902), .DIN2 (________24923),
       .Q (________24924));
  nnd2s1 _______444791(.DIN1 (________24921), .DIN2 (_____0__24140), .Q
       (________24922));
  nnd2s1 ______444792(.DIN1 (________24725), .DIN2 (________22139), .Q
       (________24920));
  nnd2s1 _______444793(.DIN1 (________24679), .DIN2 (____9___24697), .Q
       (________24919));
  nor2s1 ______444794(.DIN1 (________24494), .DIN2 (________24685), .Q
       (________24918));
  and2s1 _____0_444795(.DIN1 (_____0__24916), .DIN2 (_____0__23056), .Q
       (________24917));
  xor2s1 _____0_444796(.DIN1 (___9____21609), .DIN2
       (______________________________________0_____________18888), .Q
       (_____9__24915));
  and2s1 _______444797(.DIN1 (_____9___30627), .DIN2 (inData[4]), .Q
       (________24914));
  and2s1 _______444798(.DIN1 (_____00__34828), .DIN2 (________24912),
       .Q (________24913));
  nnd2s1 _____9_444799(.DIN1 (_____0___34830), .DIN2 (__900_), .Q
       (________24911));
  nor2s1 _____444800(.DIN1 (________24909), .DIN2 (________24681), .Q
       (________24910));
  nor2s1 _______444801(.DIN1 (___0____24347), .DIN2 (____0___24702), .Q
       (__9_____26734));
  nor2s1 _____9_444802(.DIN1 (________24908), .DIN2 (________24566), .Q
       (___9____25233));
  or2s1 _______444803(.DIN1 (___9____24268), .DIN2 (__9__0__27035), .Q
       (____9___25462));
  nnd2s1 ______444804(.DIN1 (_____9___30627), .DIN2 (_________18852),
       .Q (________25105));
  nnd2s1 _____9_444805(.DIN1 (________24688), .DIN2 (___0__0__27287),
       .Q (___9____25225));
  hi1s1 _______444806(.DIN (________25107), .Q (________25422));
  nor2s1 _______444807(.DIN1 (___0_____27914), .DIN2
       (______________________________________0___________), .Q
       (__9_0___26805));
  nor2s1 _______444808(.DIN1 (outData[4]), .DIN2 (____0___24986), .Q
       (_____9__25050));
  xor2s1 _____444809(.DIN1 (________24479), .DIN2 (____0____30977), .Q
       (___99___25264));
  nor2s1 _______444810(.DIN1 (________22421), .DIN2 (___0____24394), .Q
       (________24907));
  nnd2s1 ______444811(.DIN1 (___90___26151), .DIN2 (____9___24516), .Q
       (_____0__24906));
  nor2s1 _______444812(.DIN1 (________24904), .DIN2 (________24468), .Q
       (_____9__24905));
  nor2s1 _______444813(.DIN1 (________24902), .DIN2 (____00__24518), .Q
       (________24903));
  nor2s1 _______444814(.DIN1 (____9___23971), .DIN2 (_________34842),
       .Q (________24901));
  nnd2s1 _______444815(.DIN1 (________24441), .DIN2 (____00__19399), .Q
       (________24900));
  nor2s1 _______444816(.DIN1 (_____9__22763), .DIN2 (________24448), .Q
       (________24899));
  nnd2s1 _______444817(.DIN1 (________24457), .DIN2 (_____0__23582), .Q
       (________24898));
  and2s1 ______444818(.DIN1 (______0__34848), .DIN2 (___9____25195), .Q
       (________24897));
  nnd2s1 ______444819(.DIN1 (__99____27118), .DIN2
       (______________________________________0_____________18888), .Q
       (_____0__24896));
  nnd2s1 _______444820(.DIN1 (____0___24893), .DIN2 (________24775), .Q
       (____09__24895));
  nnd2s1 _____444821(.DIN1 (____0___24893), .DIN2 (_____0__22023), .Q
       (____0___24894));
  and2s1 _______444822(.DIN1 (___0_9__24361), .DIN2 (_____0__25520), .Q
       (____0___24892));
  nnd2s1 _______444823(.DIN1 (________24561), .DIN2 (____0___24890), .Q
       (____0___24891));
  nor2s1 _______444824(.DIN1 (____0___24888), .DIN2 (___0_0__24410), .Q
       (____0___24889));
  nor2s1 _______444825(.DIN1 (____00__24886), .DIN2 (___0____24379), .Q
       (____0___24887));
  or2s1 ____0__444826(.DIN1 (____9___24884), .DIN2 (___0____24359), .Q
       (____9___24885));
  and2s1 ____0__444827(.DIN1 (___0____24367), .DIN2 (________25132), .Q
       (____9___24883));
  nnd2s1 ____0__444828(.DIN1 (___00___24335), .DIN2 (________22818), .Q
       (____9___24882));
  nor2s1 ____0__444829(.DIN1 (_____9__23027), .DIN2 (___9____24321), .Q
       (____9___24881));
  nor2s1 ____0__444830(.DIN1 (________24118), .DIN2 (___99___24327), .Q
       (____9___24880));
  or2s1 ____0__444831(.DIN1 (________24528), .DIN2 (___0____24383), .Q
       (____9___24879));
  nnd2s1 ____0__444832(.DIN1 (___0____24348), .DIN2 (____90__24877), .Q
       (____9___24878));
  nor2s1 ____09_444833(.DIN1 (________23758), .DIN2 (___0____24411), .Q
       (_____9__24876));
  and2s1 ____09_444834(.DIN1 (________24554), .DIN2 (________24817), .Q
       (________24875));
  nor2s1 ____444835(.DIN1 (___9____24303), .DIN2 (___0____24373), .Q
       (________24874));
  nnd2s1 _____0_444836(.DIN1 (___0_9__24390), .DIN2 (____99__25750), .Q
       (________24873));
  and2s1 _____0_444837(.DIN1 (________24871), .DIN2 (_____9__23736), .Q
       (________24872));
  nor2s1 _____0_444838(.DIN1 (____00__24886), .DIN2 (___0____24380), .Q
       (________24870));
  and2s1 _______444839(.DIN1 (___0____24366), .DIN2 (_________34964),
       .Q (________24869));
  nor2s1 _______444840(.DIN1 (________24087), .DIN2 (___090__24419), .Q
       (________24868));
  or2s1 _______444841(.DIN1 (________24902), .DIN2 (___0____24363), .Q
       (_____0__24867));
  nnd2s1 _______444842(.DIN1 (___0____24360), .DIN2 (________24865), .Q
       (_____9__24866));
  nor2s1 ______444843(.DIN1 (____9___25945), .DIN2 (___9____24324), .Q
       (________24864));
  nnd2s1 _______444844(.DIN1 (________24556), .DIN2 (________24090), .Q
       (________24863));
  and2s1 _______444845(.DIN1 (___0____24354), .DIN2 (________25132), .Q
       (________24862));
  nor2s1 _______444846(.DIN1 (________23823), .DIN2 (____09__24436), .Q
       (________24861));
  and2s1 _______444847(.DIN1 (___0____24357), .DIN2 (________24859), .Q
       (________24860));
  nnd2s1 _______444848(.DIN1 (___0____24353), .DIN2 (________23539), .Q
       (________24858));
  nor2s1 _______444849(.DIN1 (___99___24329), .DIN2 (___0_9__24381), .Q
       (_____9__24857));
  nor2s1 _______444850(.DIN1 (________24855), .DIN2 (___0____24404), .Q
       (________24856));
  nor2s1 _______444851(.DIN1 (________24135), .DIN2 (________24850), .Q
       (________24854));
  nnd2s1 _______444852(.DIN1 (___0_9__24351), .DIN2 (________24852), .Q
       (________24853));
  nor2s1 _______444853(.DIN1 (________22639), .DIN2 (________24850), .Q
       (________24851));
  nor2s1 _______444854(.DIN1 (________26101), .DIN2 (___0____24413), .Q
       (________24849));
  nor2s1 _______444855(.DIN1 (_____9__24847), .DIN2 (___0____24392), .Q
       (_____0__24848));
  nor2s1 _______444856(.DIN1 (________24845), .DIN2 (________24555), .Q
       (________24846));
  or2s1 _______444857(.DIN1 (___0____24345), .DIN2 (________24931), .Q
       (________24844));
  nnd2s1 _______444858(.DIN1 (___0____24344), .DIN2 (___9____24271), .Q
       (________24843));
  or2s1 _______444859(.DIN1 (________23647), .DIN2 (___0____24385), .Q
       (________24842));
  nnd2s1 ______444860(.DIN1 (___00___24338), .DIN2 (________19520), .Q
       (________24841));
  nnd2s1 ______444861(.DIN1 (___0____24405), .DIN2 (____9___23615), .Q
       (________24840));
  nnd2s1 _______444862(.DIN1 (________24453), .DIN2 (___0____24349), .Q
       (________24839));
  nor2s1 _____0_444863(.DIN1 (______0__35058), .DIN2 (___0_9__24409),
       .Q (________24837));
  nnd2s1 _______444864(.DIN1 (___0____24388), .DIN2 (___09___25358), .Q
       (________24836));
  nnd2s1 _______444865(.DIN1 (___990__24326), .DIN2 (________22741), .Q
       (________24835));
  nor2s1 _______444866(.DIN1 (________24833), .DIN2 (___0____24387), .Q
       (________24834));
  nnd2s1 _____9_444867(.DIN1 (___999__24332), .DIN2 (________23039), .Q
       (________24832));
  and2s1 _____9_444868(.DIN1 (___99___24330), .DIN2 (________24830), .Q
       (________24831));
  or2s1 _____9_444869(.DIN1 (_____9__24828), .DIN2 (___0_9__24371), .Q
       (_____0__24829));
  nnd2s1 _____444870(.DIN1 (___0____24365), .DIN2 (________24470), .Q
       (________24827));
  nnd2s1 _____0_444871(.DIN1 (_____9__24559), .DIN2 (___9____24275), .Q
       (________24826));
  and2s1 _____0_444872(.DIN1 (___0____24356), .DIN2 (________24824), .Q
       (________24825));
  or2s1 _____0_444873(.DIN1 (__9_9___26416), .DIN2 (_____9__24498), .Q
       (________24823));
  nnd2s1 _____0_444874(.DIN1 (_________34846), .DIN2 (______9__28444),
       .Q (_________28671));
  and2s1 _____9_444875(.DIN1 (___09___24421), .DIN2 (________24822), .Q
       (________25112));
  nor2s1 ______444876(.DIN1 (________24821), .DIN2 (___0____24369), .Q
       (________25116));
  nor2s1 _______444877(.DIN1 (_____0__24465), .DIN2 (________24820), .Q
       (___9_0__25211));
  hi1s1 _______444878(.DIN (_____0__24819), .Q (___0_____27690));
  dffacs2 __________________444879(.CLRB (reset), .CLK (clk), .DIN
       (___0____24370), .Q (_______________18879));
  dffacs2 __________________444880(.CLRB (reset), .CLK (clk), .DIN
       (___0____24376), .Q
       (______________________________________0_____________18886));
  nnd2s1 ______444881(.DIN1 (____0___24523), .DIN2 (________24817), .Q
       (_____9__24818));
  nnd2s1 ______444882(.DIN1 (___0____24346), .DIN2 (________25627), .Q
       (________24816));
  or2s1 _______444883(.DIN1 (________24814), .DIN2 (_____0__24437), .Q
       (________24815));
  nnd2s1 _______444884(.DIN1 (___0____24375), .DIN2 (________24830), .Q
       (________24813));
  nnd2s1 ______444885(.DIN1 (____9___24510), .DIN2 (________24558), .Q
       (________24812));
  nnd2s1 _______444886(.DIN1 (___09___24424), .DIN2 (________25098), .Q
       (________24811));
  nnd2s1 _______444887(.DIN1 (___0____24395), .DIN2 (_____0__24809), .Q
       (________24810));
  nnd2s1 _______444888(.DIN1 (_____9__24550), .DIN2 (________24459), .Q
       (_____9__24808));
  or2s1 _______444889(.DIN1 (________24806), .DIN2 (________24544), .Q
       (________24807));
  nnd2s1 _______444890(.DIN1 (___0____24402), .DIN2 (________24804), .Q
       (________24805));
  nor2s1 _______444891(.DIN1 (___99___24331), .DIN2 (___00___24337), .Q
       (________24803));
  nor2s1 _______444892(.DIN1 (__9__0__26346), .DIN2 (________24552), .Q
       (________24802));
  nor2s1 ______444893(.DIN1 (________22410), .DIN2 (________24545), .Q
       (____09__24801));
  nor2s1 ______444894(.DIN1 (________22222), .DIN2 (___09___24426), .Q
       (____0___24800));
  nor2s1 _______444895(.DIN1 (____0___24798), .DIN2 (___000__24333), .Q
       (____0___24799));
  or2s1 _______444896(.DIN1 (__9_____26713), .DIN2 (________24542), .Q
       (____0___24797));
  nnd2s1 _______444897(.DIN1 (________24562), .DIN2 (________22143), .Q
       (____0___24796));
  nor2s1 _______444898(.DIN1
       (______________________________________0_____________18888),
       .DIN2 (_________30104), .Q (____0___24795));
  nor2s1 _____9_444899(.DIN1 (____0___23532), .DIN2 (___09___24422), .Q
       (____0___24794));
  nnd2s1 _______444900(.DIN1 (________24476), .DIN2 (____00__24792), .Q
       (____0___24793));
  or2s1 _______444901(.DIN1 (___0____23448), .DIN2 (________24757), .Q
       (____99__24791));
  and2s1 _______444902(.DIN1 (________24529), .DIN2 (________24912), .Q
       (____9___24790));
  nor2s1 _______444903(.DIN1 (_________31126), .DIN2 (_________33278),
       .Q (____9___24789));
  and2s1 ______444904(.DIN1 (_____0__24456), .DIN2 (___0_____27825), .Q
       (____9___24788));
  nnd2s1 _______444905(.DIN1 (________24535), .DIN2
       (_________________18700), .Q (____9___24787));
  and2s1 _______444906(.DIN1 (________24484), .DIN2 (_____9__22345), .Q
       (____9___24786));
  nnd2s1 _______444907(.DIN1 (____9___24784), .DIN2 (inData[14]), .Q
       (____9___24785));
  and2s1 _______444908(.DIN1 (____9___24784), .DIN2 (inData[2]), .Q
       (____9___24783));
  nor2s1 _______444909(.DIN1 (________24489), .DIN2 (___9____21623), .Q
       (____90__24782));
  nor2s1 _______444910(.DIN1 (________24780), .DIN2 (________24527), .Q
       (_____9__24781));
  or2s1 _______444911(.DIN1 (____9___22348), .DIN2 (_____0__24491), .Q
       (________24779));
  and2s1 _______444912(.DIN1 (____9___24512), .DIN2 (________24777), .Q
       (________24778));
  nnd2s1 _______444913(.DIN1 (________24775), .DIN2 (________24774), .Q
       (________24776));
  nor2s1 ______444914(.DIN1 (_____0__24772), .DIN2 (_____0__24525), .Q
       (________24773));
  nor2s1 _______444915(.DIN1 (___9_0__25231), .DIN2 (___9_9__24325), .Q
       (_____9__24771));
  nor2s1 _______444916(.DIN1 (____0___19116), .DIN2 (________24765), .Q
       (________24770));
  nnd2s1 _______444917(.DIN1 (____0___24435), .DIN2 (___9____25205), .Q
       (________24769));
  and2s1 _______444918(.DIN1 (________24506), .DIN2 (___0____22595), .Q
       (________24768));
  or2s1 _______444919(.DIN1 (________24192), .DIN2 (____0___24519), .Q
       (________24767));
  and2s1 _______444920(.DIN1 (________24765), .DIN2 (________24212), .Q
       (________24766));
  or2s1 _____9_444921(.DIN1 (____9___24695), .DIN2 (________24450), .Q
       (_____0__24764));
  nor2s1 _____0_444922(.DIN1 (________23940), .DIN2 (____9___24514), .Q
       (________24763));
  and2s1 ______444923(.DIN1 (________24487), .DIN2 (____9___24511), .Q
       (________24761));
  nor2s1 _______444924(.DIN1 (_____9__24464), .DIN2 (___9____24270), .Q
       (________24760));
  nnd2s1 _______444925(.DIN1 (________24478), .DIN2 (_____9__24507), .Q
       (________24759));
  nnd2s1 _______444926(.DIN1 (________24757), .DIN2 (________23812), .Q
       (________24758));
  nor2s1 ______444927(.DIN1 (________24504), .DIN2 (_____9__24755), .Q
       (_____0__24756));
  nor2s1 _______444928(.DIN1 (_____0__24499), .DIN2 (________24500), .Q
       (________24754));
  nor2s1 _______444929(.DIN1 (__9_____26953), .DIN2 (________24564), .Q
       (________24753));
  nor2s1 _______444930(.DIN1 (________24496), .DIN2 (________24495), .Q
       (________24752));
  or2s1 _______444931(.DIN1 (________24493), .DIN2 (_____9__24755), .Q
       (________24751));
  nor2s1 _______444932(.DIN1 (________24749), .DIN2 (________24471), .Q
       (________24750));
  nnd2s1 _____0_444933(.DIN1 (________24461), .DIN2 (_____9__25118), .Q
       (________24748));
  nor2s1 _____0_444934(.DIN1 (_____0__24746), .DIN2 (________24460), .Q
       (________24747));
  nnd2s1 _____9_444935(.DIN1 (_____9__24480), .DIN2 (________24221), .Q
       (_____9__24745));
  nor2s1 ______444936(.DIN1 (____90__21438), .DIN2 (________24526), .Q
       (________24744));
  and2s1 _______444937(.DIN1 (________24742), .DIN2 (____0___24432), .Q
       (__9_____27019));
  nor2s1 _______444938(.DIN1 (____9___24238), .DIN2 (________24741), .Q
       (____90__25645));
  nnd2s1 ______444939(.DIN1 (________24740), .DIN2 (________24462), .Q
       (____9___25073));
  or2s1 ______444940(.DIN1 (____90__24508), .DIN2 (___0__0__27994), .Q
       (____9___25075));
  nnd2s1 _____444941(.DIN1 (___0____24417), .DIN2 (________23903), .Q
       (_____0__25127));
  nnd2s1 _____9_444942(.DIN1 (___09___24425), .DIN2 (________24543), .Q
       (____90__25165));
  xor2s1 _____9_444943(.DIN1 (________24176), .DIN2 (____0____31872),
       .Q (_____0__24965));
  and2s1 _____0_444944(.DIN1 (________24548), .DIN2 (_____0__24739), .Q
       (___09____28121));
  xor2s1 _____0_444945(.DIN1 (_________30595), .DIN2 (________24585),
       .Q (________25107));
  hi1s1 _____0_444946(.DIN
       (______________________________________0___________), .Q
       (_________28661));
  nnd2s1 _____9_444947(.DIN1 (________24117), .DIN2 (________24486), .Q
       (_____9__24738));
  nor2s1 ______444948(.DIN1 (___09___24423), .DIN2 (___9____24259), .Q
       (________24737));
  and2s1 _______444949(.DIN1 (________24197), .DIN2 (________24735), .Q
       (________24736));
  nor2s1 ______444950(.DIN1 (________24733), .DIN2 (______0__34868), .Q
       (________24734));
  or2s1 _______444951(.DIN1 (_____0__26127), .DIN2 (___9____24308), .Q
       (________24732));
  nor2s1 _______444952(.DIN1 (____0___23177), .DIN2 (________24214), .Q
       (________24731));
  nor2s1 ______444953(.DIN1 (________24191), .DIN2 (________24931), .Q
       (________24730));
  nor2s1 _______444954(.DIN1 (_________34856), .DIN2 (_____00__34928),
       .Q (_____0__24729));
  nor2s1 _______444955(.DIN1 (___9____24282), .DIN2 (___9____24269), .Q
       (________24728));
  nnd2s1 _______444956(.DIN1 (________24223), .DIN2 (________24726), .Q
       (________24727));
  nor2s1 _______444957(.DIN1 (________24724), .DIN2 (________24184), .Q
       (________24725));
  or2s1 ______444958(.DIN1 (________24722), .DIN2 (____90__24235), .Q
       (________24723));
  nor2s1 _____444959(.DIN1 (__90____26312), .DIN2 (_____9__24234), .Q
       (________24721));
  nor2s1 _____9_444960(.DIN1 (_____9__24719), .DIN2 (________24215), .Q
       (_____0__24720));
  nor2s1 _____9_444961(.DIN1 (____9___19945), .DIN2 (_________34860),
       .Q (________24718));
  nor2s1 _____9_444962(.DIN1 (________25137), .DIN2 (_____0__24199), .Q
       (________24717));
  nor2s1 _____0_444963(.DIN1 (________24221), .DIN2 (________24206), .Q
       (________24716));
  nor2s1 _______444964(.DIN1 (___09___24420), .DIN2 (________24136), .Q
       (________24715));
  or2s1 _______444965(.DIN1 (________23642), .DIN2 (________24133), .Q
       (________24714));
  nnd2s1 _______444966(.DIN1 (_____0__24130), .DIN2 (________24712), .Q
       (________24713));
  or2s1 _______444967(.DIN1 (________23872), .DIN2 (___9____24311), .Q
       (________24711));
  xor2s1 ______444968(.DIN1 (____9____31787), .DIN2 (____00___33677),
       .Q (_____0__24710));
  or2s1 _______444969(.DIN1 (________24821), .DIN2 (________24167), .Q
       (____09__24709));
  nor2s1 ______444970(.DIN1 (________24175), .DIN2 (___0____24358), .Q
       (____0___24708));
  nor2s1 _______444971(.DIN1 (___9____23401), .DIN2 (___0_9__24400), .Q
       (____0___24707));
  nnd2s1 _______444972(.DIN1 (____9___24152), .DIN2 (____0___24705), .Q
       (____0___24706));
  nor2s1 ______444973(.DIN1 (________22840), .DIN2 (____9___24698), .Q
       (____0___24703));
  nor2s1 _______444974(.DIN1 (____00__24701), .DIN2 (____9___24698), .Q
       (____0___24702));
  nor2s1 _______444975(.DIN1 (________23847), .DIN2 (____9___24698), .Q
       (____99__24700));
  nor2s1 _______444976(.DIN1 (________23297), .DIN2 (____9___24698), .Q
       (____9___24699));
  nnd2s1 _______444977(.DIN1 (________24689), .DIN2 (____9___23972), .Q
       (____9___24697));
  nor2s1 _______444978(.DIN1 (____9___24695), .DIN2 (________24638), .Q
       (____9___24696));
  nnd2s1 _______444979(.DIN1 (____9___24148), .DIN2 (________25798), .Q
       (____9___24694));
  or2s1 _______444980(.DIN1 (________24855), .DIN2 (________24134), .Q
       (____90__24693));
  nor2s1 ______444981(.DIN1 (________23561), .DIN2 (____9___24698), .Q
       (________24691));
  nnd2s1 _______444982(.DIN1 (________24689), .DIN2 (___0____23513), .Q
       (________24690));
  nor2s1 _______444983(.DIN1 (________25913), .DIN2 (________24143), .Q
       (________24688));
  nor2s1 _____9_444984(.DIN1 (____9___23076), .DIN2 (________24733), .Q
       (________24687));
  or2s1 _____9_444985(.DIN1 (________23834), .DIN2 (____9___24698), .Q
       (________24686));
  nor2s1 _____444986(.DIN1 (________23210), .DIN2 (____9___24698), .Q
       (________24685));
  nnd2s1 ____90_444987(.DIN1 (________24117), .DIN2 (___0____23497), .Q
       (_____0__24684));
  nor2s1 ____9__444988(.DIN1 (________24682), .DIN2 (____9___24698), .Q
       (________24683));
  or2s1 ____9__444989(.DIN1 (________24680), .DIN2 (_________34862), .Q
       (________24681));
  nnd2s1 ____9_444990(.DIN1 (________24117), .DIN2 (________22841), .Q
       (________24679));
  and2s1 ____9__444991(.DIN1 (_____9__24147), .DIN2 (________25049), .Q
       (________24678));
  nor2s1 ____9__444992(.DIN1 (___9____26163), .DIN2 (____9___24698), .Q
       (________24677));
  nor2s1 ____9__444993(.DIN1 (________22369), .DIN2 (____9___24698), .Q
       (_____0__24676));
  nnd2s1 ____9__444994(.DIN1 (________24689), .DIN2 (________24477), .Q
       (_____9__24675));
  nnd2s1 ____0__444995(.DIN1 (________24117), .DIN2 (________24549), .Q
       (________24674));
  nnd2s1 ____0__444996(.DIN1 (________24117), .DIN2 (___0____23498), .Q
       (________24673));
  nnd2s1 _____444997(.DIN1 (________24125), .DIN2 (________23944), .Q
       (________24672));
  nnd2s1 _____0_444998(.DIN1 (____09__24162), .DIN2 (________24202), .Q
       (________24671));
  nnd2s1 _____0_444999(.DIN1 (________24168), .DIN2 (________24669), .Q
       (________24670));
  nnd2s1 ____09_445000(.DIN1 (_____9__24129), .DIN2 (_____9__23674), .Q
       (________24668));
  and2s1 ____445001(.DIN1 (________24127), .DIN2 (_____0__24666), .Q
       (________24667));
  nor2s1 ____0__445002(.DIN1 (________23198), .DIN2 (________24661), .Q
       (_____9__24665));
  nnd2s1 ____0_445003(.DIN1 (________24128), .DIN2 (_____0__23675), .Q
       (________24664));
  or2s1 ____0_445004(.DIN1 (________24662), .DIN2 (________24661), .Q
       (________24663));
  nnd2s1 _____0_445005(.DIN1 (_____9__24218), .DIN2 (________24660), .Q
       (________24921));
  nor2s1 ____0__445006(.DIN1 (________23097), .DIN2 (________24733), .Q
       (_____0__24819));
  nor2s1 _____0_445007(.DIN1 (________24186), .DIN2 (________24188), .Q
       (________24743));
  nor2s1 _____445008(.DIN1 (___9_9__24305), .DIN2 (______0__28263), .Q
       (_________28298));
  nnd2s1 ____0__445009(.DIN1 (________24117), .DIN2 (________24659), .Q
       (____9___24979));
  or2s1 ____0__445010(.DIN1 (_____9__25674), .DIN2 (____9___24698), .Q
       (________25046));
  nor2s1 _______445011(.DIN1 (________24196), .DIN2 (___0_____27631),
       .Q (___0_____27336));
  nor2s1 _______445012(.DIN1 (____0___22357), .DIN2 (____9___24153), .Q
       (_____0__24916));
  nor2s1 _______445013(.DIN1 (________22031), .DIN2 (____9___24698), .Q
       (__9__0__27035));
  xor2s1 _______445014(.DIN1 (___________0___18883), .DIN2
       (____9____31787), .Q (_____0___31902));
  xor2s1 _______445015(.DIN1 (_____________9___18703), .DIN2
       (_________35111), .Q (_________32226));
  nnd2s1 _______445016(.DIN1 (________24689), .DIN2 (___0____24389), .Q
       (___0__9__27879));
  nnd2s1 ____0_445017(.DIN1 (________24689), .DIN2 (_________34946), .Q
       (___0_____27527));
  nnd2s1 ____0__445018(.DIN1 (____9___24150), .DIN2 (___09____28113),
       .Q (_________28497));
  nnd2s1 ____0__445019(.DIN1 (________24689), .DIN2 (________23300), .Q
       (___0_____27912));
  hi1s1 ______445020(.DIN
       (______________________________________0_____________18888), .Q
       (_____9___30627));
  nor2s1 _____0_445021(.DIN1 (_________________18702), .DIN2
       (____9___24600), .Q (________24658));
  nnd2s1 _______445022(.DIN1 (_____9__24172), .DIN2 (___0____24374), .Q
       (________24657));
  nnd2s1 _______445023(.DIN1 (________24145), .DIN2 (_____9__24655), .Q
       (_____0__24656));
  nnd2s1 _____445024(.DIN1 (________24131), .DIN2 (________24144), .Q
       (________24654));
  nor2s1 _____0_445025(.DIN1 (___0____24378), .DIN2 (________24174), .Q
       (________24653));
  and2s1 _______445026(.DIN1 (___9____24309), .DIN2 (________24651), .Q
       (________24652));
  nnd2s1 _______445027(.DIN1 (________24178), .DIN2 (_________35064),
       .Q (________24650));
  nnd2s1 ______445028(.DIN1 (________24138), .DIN2 (________23022), .Q
       (________24649));
  nor2s1 _______445029(.DIN1 (________24036), .DIN2 (________24137), .Q
       (________24648));
  nnd2s1 _______445030(.DIN1 (____0___24158), .DIN2 (_____0__24646), .Q
       (________24647));
  nor2s1 _______445031(.DIN1 (________24644), .DIN2 (___9____24310), .Q
       (_____9__24645));
  nor2s1 _______445032(.DIN1 (________24642), .DIN2 (___9____24312), .Q
       (________24643));
  nor2s1 _______445033(.DIN1 (________23945), .DIN2 (_________34864),
       .Q (________24641));
  nnd2s1 _______445034(.DIN1 (________24179), .DIN2 (________21790), .Q
       (________24640));
  nor2s1 _______445035(.DIN1 (_________34960), .DIN2 (________24638),
       .Q (________24639));
  and2s1 ______445036(.DIN1 (________24438), .DIN2 (_________34496), .Q
       (________24637));
  and2s1 _______445037(.DIN1 (_____9__24635), .DIN2 (_________34488),
       .Q (_____0__24636));
  nnd2s1 _______445038(.DIN1 (___9_0__24249), .DIN2 (________24440), .Q
       (________24634));
  and2s1 _______445039(.DIN1 (___90___24247), .DIN2 (________24632), .Q
       (________24633));
  and2s1 _______445040(.DIN1 (________24233), .DIN2 (________25068), .Q
       (________24631));
  and2s1 _______445041(.DIN1 (________24629), .DIN2 (________23852), .Q
       (________24630));
  nnd2s1 _______445042(.DIN1 (____9___24239), .DIN2 (________24627), .Q
       (________24628));
  nnd2s1 _______445043(.DIN1 (___9____24294), .DIN2 (_____9__24625), .Q
       (_____0__24626));
  nor2s1 _______445044(.DIN1 (________23831), .DIN2 (___9____24291), .Q
       (________24624));
  nnd2s1 _______445045(.DIN1 (___9____24292), .DIN2 (____9___24151), .Q
       (________24623));
  nnd2s1 _______445046(.DIN1 (________24210), .DIN2 (________23661), .Q
       (________24622));
  nnd2s1 _______445047(.DIN1 (________24580), .DIN2 (_____9__23755), .Q
       (________24621));
  nnd2s1 ______445048(.DIN1 (________24217), .DIN2 (________24619), .Q
       (________24620));
  nnd2s1 ______445049(.DIN1 (___9____24284), .DIN2 (________23658), .Q
       (________24618));
  or2s1 _______445050(.DIN1 (_____0__24616), .DIN2 (___9_9__24256), .Q
       (________24617));
  nor2s1 _______445051(.DIN1 (_____0__22089), .DIN2 (___9_9__24285), .Q
       (____09__24615));
  and2s1 _______445052(.DIN1 (________24629), .DIN2 (________23296), .Q
       (____0___24614));
  and2s1 ______445053(.DIN1 (___9_0__24286), .DIN2 (____9___24981), .Q
       (____0___24613));
  or2s1 _______445054(.DIN1 (____0___24611), .DIN2 (___9____24280), .Q
       (____0___24612));
  or2s1 _______445055(.DIN1 (________22097), .DIN2 (________24213), .Q
       (____0___24610));
  nnd2s1 _______445056(.DIN1 (________24189), .DIN2 (________23071), .Q
       (____0___24609));
  nor2s1 _____9_445057(.DIN1 (________24141), .DIN2 (____0___23891), .Q
       (____00__24608));
  nor2s1 _______445058(.DIN1 (_____0__24190), .DIN2 (________24931), .Q
       (____99__24607));
  nor2s1 _____0_445059(.DIN1 (____9___24605), .DIN2 (___9____24272), .Q
       (____9___24606));
  nnd2s1 _____0_445060(.DIN1 (___9____24251), .DIN2 (___009__23445), .Q
       (____9___24604));
  nor2s1 _______445061(.DIN1 (________23829), .DIN2 (________24225), .Q
       (____9___24603));
  nor2s1 _______445062(.DIN1 (___90___24246), .DIN2 (________24047), .Q
       (____9___24602));
  nor2s1 _______445063(.DIN1 (______9__32271), .DIN2 (____9___24600),
       .Q (____9___24601));
  nnd2s1 ______445064(.DIN1 (________24231), .DIN2 (_____9__22779), .Q
       (____9___24599));
  nor2s1 _______445065(.DIN1 (___9_9__24266), .DIN2 (________24592), .Q
       (____90__24598));
  nor2s1 _______445066(.DIN1 (___9____24264), .DIN2 (________24733), .Q
       (_____9__24597));
  or2s1 _______445067(.DIN1 (________26130), .DIN2 (___9_0__24296), .Q
       (________24596));
  nor2s1 ______445068(.DIN1 (___9____24261), .DIN2 (________24931), .Q
       (________24595));
  nor2s1 ______445069(.DIN1 (___0_9__20770), .DIN2 (________24536), .Q
       (________24594));
  nor2s1 _______445070(.DIN1 (___9____24258), .DIN2 (________24592), .Q
       (________24593));
  nnd2s1 _______445071(.DIN1 (________23904), .DIN2 (___90___24243), .Q
       (________24591));
  nnd2s1 _______445072(.DIN1 (________24689), .DIN2 (___9____24255), .Q
       (________24590));
  and2s1 ______445073(.DIN1 (____9___24240), .DIN2 (_____0__24588), .Q
       (________24589));
  nor2s1 _______445074(.DIN1 (___0____24398), .DIN2 (________24226), .Q
       (_____9__24587));
  and2s1 _______445075(.DIN1 (________24585), .DIN2 (outData[3]), .Q
       (________24586));
  or2s1 _______445076(.DIN1 (________24583), .DIN2 (___9____24252), .Q
       (________24584));
  nor2s1 _______445077(.DIN1 (_________34854), .DIN2 (_____0__25616),
       .Q (________24582));
  nnd2s1 _______445078(.DIN1 (_____9__23571), .DIN2 (________24580), .Q
       (________24581));
  nor2s1 _______445079(.DIN1 (_____9__24578), .DIN2 (_________34852),
       .Q (_____0__24579));
  nnd2s1 _______445080(.DIN1 (________24204), .DIN2 (inData[30]), .Q
       (________24577));
  nor2s1 _____445081(.DIN1 (___9____22458), .DIN2 (________24203), .Q
       (________24576));
  nnd2s1 _____9_445082(.DIN1 (_____0__24182), .DIN2 (________22783), .Q
       (________24575));
  nor2s1 _____9_445083(.DIN1 (___9____24278), .DIN2 (________24733), .Q
       (________24574));
  nor2s1 ______445084(.DIN1 (___9____26179), .DIN2 (________24201), .Q
       (________24573));
  and2s1 _______445085(.DIN1 (___90___24244), .DIN2 (________24571), .Q
       (________24572));
  and2s1 _______445086(.DIN1 (_____9__24569), .DIN2 (________24568), .Q
       (_____0__24570));
  nnd2s1 _______445087(.DIN1 (___0_9__23489), .DIN2 (____9___24237), .Q
       (________24567));
  nnd2s1 _______445088(.DIN1 (______0__34858), .DIN2 (_____9__23311),
       .Q (________24566));
  nor2s1 ______445089(.DIN1 (________24080), .DIN2 (________25110), .Q
       (________24565));
  and2s1 _______445090(.DIN1 (___9____24299), .DIN2 (________25707), .Q
       (_____0__25041));
  nnd2s1 _______445091(.DIN1 (____0___24161), .DIN2 (__9_____26406), .Q
       (________25020));
  or2s1 _______445092(.DIN1 (outData[3]), .DIN2 (________24585), .Q
       (____0___24986));
  dffacs1 _________________445093(.CLRB (reset), .CLK (clk), .DIN
       (___9_9__24295), .Q
       (______________________________________0___________));
  nor2s1 _______445094(.DIN1 (________24563), .DIN2 (________23960), .Q
       (________24564));
  nor2s1 _______445095(.DIN1 (________23635), .DIN2 (_____9__24101), .Q
       (________24562));
  and2s1 _______445096(.DIN1 (________24037), .DIN2 (_____0__24560), .Q
       (________24561));
  nnd2s1 _______445097(.DIN1 (________24085), .DIN2 (________24221), .Q
       (_____9__24559));
  nnd2s1 _______445098(.DIN1 (____0___24066), .DIN2 (________24557), .Q
       (________24558));
  and2s1 _______445099(.DIN1 (___0____24355), .DIN2 (____9___23798), .Q
       (________24556));
  nnd2s1 ______445100(.DIN1 (___0____24416), .DIN2 (________22272), .Q
       (________24555));
  nor2s1 _______445101(.DIN1 (________23131), .DIN2 (________24099), .Q
       (________24554));
  nnd2s1 _______445102(.DIN1 (________24014), .DIN2 (___0____22568), .Q
       (________24553));
  nnd2s1 _______445103(.DIN1 (________24088), .DIN2 (_____0__24551), .Q
       (________24552));
  nor2s1 _______445104(.DIN1 (________24549), .DIN2 (________24021), .Q
       (_____9__24550));
  nnd2s1 _____9_445105(.DIN1 (________24547), .DIN2 (________24546), .Q
       (________24548));
  nnd2s1 _____9_445106(.DIN1 (_____9__24052), .DIN2 (___9____23379), .Q
       (________24545));
  nnd2s1 _____9_445107(.DIN1 (________24543), .DIN2 (________23327), .Q
       (________24544));
  or2s1 _____445108(.DIN1 (_____0__24541), .DIN2 (________24010), .Q
       (________24542));
  xor2s1 _______445109(.DIN1 (_________33530), .DIN2 (_________31290),
       .Q (________24540));
  xor2s1 ______445110(.DIN1 (____0____31818), .DIN2 (_________31290),
       .Q (________24539));
  xor2s1 _______445111(.DIN1 (_________________0___18633), .DIN2
       (_________31290), .Q (________24538));
  xor2s1 _______445112(.DIN1 (_____9___33026), .DIN2 (_________31290),
       .Q (________24537));
  hi1s1 _______445113(.DIN (_________32053), .Q (________24535));
  nnd2s1 ____9__445114(.DIN1 (________23723), .DIN2 (________23935), .Q
       (_____0__24534));
  nnd2s1 _______445115(.DIN1 (_________32344), .DIN2 (inData[3]), .Q
       (_____9__24533));
  nnd2s1 _______445116(.DIN1 (_________32344), .DIN2 (inData[1]), .Q
       (________24532));
  nnd2s1 _______445117(.DIN1 (_________32344), .DIN2 (inData[2]), .Q
       (________24531));
  nnd2s1 _______445118(.DIN1 (________24469), .DIN2 (________23035), .Q
       (________24530));
  nor2s1 _______445119(.DIN1 (________24528), .DIN2 (_____9__23924), .Q
       (________24529));
  nnd2s1 ______445120(.DIN1 (________23985), .DIN2 (___0_0__24382), .Q
       (________24527));
  nor2s1 _______445121(.DIN1 (___00___22540), .DIN2 (_________34874),
       .Q (________24526));
  nnd2s1 ______445122(.DIN1 (____9___23969), .DIN2 (____9___23793), .Q
       (_____0__24525));
  nnd2s1 ______445123(.DIN1 (________23904), .DIN2 (________23249), .Q
       (____09__24524));
  nor2s1 _______445124(.DIN1 (____0___24522), .DIN2 (________23953), .Q
       (____0___24523));
  nor2s1 _______445125(.DIN1 (___0____25324), .DIN2 (____0___24520), .Q
       (____0___24521));
  nnd2s1 _______445126(.DIN1 (________23936), .DIN2 (____9___23966), .Q
       (____0___24519));
  or2s1 _____9_445127(.DIN1 (____99__24517), .DIN2 (_________34876), .Q
       (____00__24518));
  and2s1 _____9_445128(.DIN1 (________23962), .DIN2 (____9___24515), .Q
       (____9___24516));
  nnd2s1 ______445129(.DIN1 (____0___23977), .DIN2 (________23306), .Q
       (____9___24514));
  nor2s1 _______445130(.DIN1 (____9___23967), .DIN2 (____9___23968), .Q
       (____9___24513));
  and2s1 _______445131(.DIN1 (________23939), .DIN2 (________25058), .Q
       (____9___24512));
  nnd2s1 ______445132(.DIN1 (____9___24510), .DIN2 (________22950), .Q
       (____9___24511));
  nnd2s1 _______445133(.DIN1 (____9___24510), .DIN2 (_____9__23608), .Q
       (____9___24509));
  and2s1 _______445134(.DIN1 (____9___24510), .DIN2 (____0___22995), .Q
       (____90__24508));
  nnd2s1 _______445135(.DIN1 (____9___24510), .DIN2 (____0___24065), .Q
       (_____9__24507));
  and2s1 ______445136(.DIN1 (____0___23980), .DIN2 (________24505), .Q
       (________24506));
  nor2s1 _______445137(.DIN1 (________22696), .DIN2 (________24492), .Q
       (________24504));
  or2s1 _______445138(.DIN1 (_____0___31003), .DIN2 (________23995), .Q
       (________24503));
  nnd2s1 _______445139(.DIN1 (____9___24510), .DIN2 (________23846), .Q
       (________24502));
  nor2s1 _______445140(.DIN1 (____9___22801), .DIN2 (_____9__24755), .Q
       (________24501));
  nor2s1 ______445141(.DIN1 (________22761), .DIN2 (_____9__24755), .Q
       (________24500));
  nor2s1 ______445142(.DIN1 (________22662), .DIN2 (________24592), .Q
       (_____0__24499));
  or2s1 _______445143(.DIN1 (_____9__25415), .DIN2 (________24020), .Q
       (_____9__24498));
  or2s1 _______445144(.DIN1 (____09__22634), .DIN2 (_________34884), .Q
       (________24497));
  nor2s1 _______445145(.DIN1 (________22044), .DIN2 (_____9__24755), .Q
       (________24496));
  nor2s1 _______445146(.DIN1 (________22749), .DIN2 (________24458), .Q
       (________24495));
  nor2s1 _______445147(.DIN1 (________23648), .DIN2 (________24592), .Q
       (________24494));
  nor2s1 _______445148(.DIN1 (______0__34938), .DIN2 (________24492),
       .Q (________24493));
  or2s1 _______445149(.DIN1 (_____9__24490), .DIN2 (________23984), .Q
       (_____0__24491));
  and2s1 _______445150(.DIN1 (____0___24434), .DIN2 (________24488), .Q
       (________24489));
  nnd2s1 ______445151(.DIN1 (________23904), .DIN2 (________24486), .Q
       (________24487));
  nor2s1 _______445152(.DIN1 (________23815), .DIN2 (________23955), .Q
       (________24485));
  nor2s1 _______445153(.DIN1 (________24483), .DIN2 (______0__34878),
       .Q (________24484));
  nnd2s1 _____9_445154(.DIN1 (_____0__24481), .DIN2 (___0____23512), .Q
       (________24482));
  or2s1 _____0_445155(.DIN1 (__9_____26773), .DIN2 (_____9__23964), .Q
       (_____9__24480));
  nor2s1 _______445156(.DIN1 (_________32114), .DIN2
       (_______________18884), .Q (________24479));
  nnd2s1 ____9__445157(.DIN1 (_____0__24481), .DIN2 (________24477), .Q
       (________24478));
  nor2s1 ____9__445158(.DIN1 (________24475), .DIN2 (________23930), .Q
       (________24476));
  nnd2s1 ____9__445159(.DIN1 (________23904), .DIN2 (_____9__23240), .Q
       (_____0__24473));
  nor2s1 ____9__445160(.DIN1 (________23557), .DIN2 (_____0__25616), .Q
       (_____9__24472));
  nnd2s1 ____9__445161(.DIN1 (________23963), .DIN2 (________24712), .Q
       (________24471));
  nnd2s1 ____9_445162(.DIN1 (________24469), .DIN2 (___9_9__23412), .Q
       (________24470));
  or2s1 ____9__445163(.DIN1 (_____0___34930), .DIN2 (____9___24149), .Q
       (________24468));
  hi1s1 _______445164(.DIN (________24466), .Q (________24467));
  nor2s1 ______445165(.DIN1 (________23543), .DIN2 (_____0__25616), .Q
       (_____9__24464));
  nnd2s1 _______445166(.DIN1 (_____0__24481), .DIN2 (___0_9__22599), .Q
       (________24463));
  nnd2s1 _______445167(.DIN1 (________23904), .DIN2 (________23192), .Q
       (________24462));
  nor2s1 _______445168(.DIN1 (___0_9__23463), .DIN2 (_____0__23925), .Q
       (________24461));
  nnd2s1 _______445169(.DIN1 (________23949), .DIN2 (___0____25329), .Q
       (________24460));
  or2s1 _______445170(.DIN1 (_______________18884), .DIN2
       (_________32158), .Q (________24457));
  nor2s1 _____445171(.DIN1 (________22968), .DIN2 (________23928), .Q
       (_____0__24456));
  nor2s1 ____90_445172(.DIN1 (________23605), .DIN2 (________24458), .Q
       (________24455));
  nor2s1 ____9__445173(.DIN1 (________23751), .DIN2 (________24592), .Q
       (________24454));
  or2s1 ____9__445174(.DIN1 (________24452), .DIN2 (________24458), .Q
       (________24453));
  or2s1 ____9_445175(.DIN1 (________24001), .DIN2 (________24592), .Q
       (________24451));
  nnd2s1 ____9__445176(.DIN1 (_____9__23957), .DIN2 (____9___24058), .Q
       (________24450));
  nnd2s1 ____9__445177(.DIN1 (________23903), .DIN2 (________23004), .Q
       (________24449));
  or2s1 ____9__445178(.DIN1 (________23121), .DIN2 (_____0__24447), .Q
       (________24448));
  nor2s1 ____9__445179(.DIN1 (________23822), .DIN2 (_____9__24755), .Q
       (_____9__24446));
  nor2s1 ____9__445180(.DIN1 (________22949), .DIN2 (_____9__24755), .Q
       (________24445));
  nor2s1 ____9__445181(.DIN1 (_____0__21876), .DIN2 (________24458), .Q
       (________24444));
  nor2s1 ____9__445182(.DIN1 (_____0__23143), .DIN2 (_____0__25616), .Q
       (________24443));
  nnd2s1 ____9__445183(.DIN1 (___9_9__24315), .DIN2 (____0____31818),
       .Q (________24442));
  nnd2s1 ____9_445184(.DIN1 (________23994), .DIN2 (________24440), .Q
       (________24441));
  nnd2s1 ____9__445185(.DIN1 (_____0__24481), .DIN2 (________23310), .Q
       (________24439));
  or2s1 _____0_445186(.DIN1 (________24546), .DIN2 (________24547), .Q
       (_____0__24739));
  nor2s1 _______445187(.DIN1 (____09__21454), .DIN2 (________24458), .Q
       (___0__9__27520));
  nnd2s1 _______445188(.DIN1 (________23904), .DIN2 (____99__23258), .Q
       (________24740));
  nnd2s1 _______445189(.DIN1 (_______________18884), .DIN2
       (_________32114), .Q (___99___25263));
  nnd2s1 _______445190(.DIN1 (________23947), .DIN2 (__99____27110), .Q
       (____9___25647));
  nor2s1 _______445191(.DIN1 (__9_9___26888), .DIN2 (________23951), .Q
       (________24757));
  nor2s1 _______445192(.DIN1 (____9___23075), .DIN2 (________24458), .Q
       (________24741));
  hi1s1 _______445193(.DIN (________24438), .Q (________24765));
  nnd2s1 _______445194(.DIN1 (_____0__24481), .DIN2 (___9____22483), .Q
       (___0_____27594));
  dffacs1 __________________445195(.CLRB (reset), .CLK (clk), .DIN
       (________23937), .Q
       (______________________________________0_____________18888));
  or2s1 _______445196(.DIN1 (___0____25336), .DIN2 (_____9__24034), .Q
       (_____0__24437));
  nor2s1 ____99_445197(.DIN1 (________19520), .DIN2 (_________34882),
       .Q (____09__24436));
  nor2s1 ____00_445198(.DIN1 (____0___24434), .DIN2 (____00__22718), .Q
       (____0___24435));
  or2s1 ____00_445199(.DIN1 (_____9__25674), .DIN2 (_____9__24755), .Q
       (____0___24433));
  nnd2s1 ____00_445200(.DIN1 (____9___24510), .DIN2 (___90___22452), .Q
       (____0___24432));
  nor2s1 ____00_445201(.DIN1 (________23194), .DIN2 (_____9__24755), .Q
       (____0___24431));
  and2s1 ____0__445202(.DIN1 (_____0__24481), .DIN2 (____9___26142), .Q
       (____0___24430));
  nor2s1 ____99_445203(.DIN1 (____9___23710), .DIN2 (________24592), .Q
       (____00__24429));
  nnd2s1 ______445204(.DIN1 (_____9__24017), .DIN2 (________22936), .Q
       (___099__24428));
  nor2s1 _______445205(.DIN1
       (______________________________________0__________0), .DIN2
       (_____9__24026), .Q (___09___24427));
  nnd2s1 _______445206(.DIN1 (________24013), .DIN2 (________23740), .Q
       (___09___24426));
  nor2s1 _______445207(.DIN1 (____90__24053), .DIN2 (_________34872),
       .Q (___09___24425));
  nor2s1 _______445208(.DIN1 (___09___24423), .DIN2 (________24004), .Q
       (___09___24424));
  nor2s1 _______445209(.DIN1
       (______________________________________0__________0), .DIN2
       (________24023), .Q (___09___24422));
  nor2s1 _______445210(.DIN1 (___09___24420), .DIN2 (________24011), .Q
       (___09___24421));
  or2s1 _______445211(.DIN1 (_________34870), .DIN2 (____0___24520), .Q
       (___090__24419));
  nor2s1 ______445212(.DIN1 (_____0__24018), .DIN2 (________23158), .Q
       (___0_9__24418));
  nnd2s1 _______445213(.DIN1 (___0____24416), .DIN2 (___9____22466), .Q
       (___0____24417));
  nnd2s1 _______445214(.DIN1 (___99___22529), .DIN2 (________24547), .Q
       (___0____24415));
  nor2s1 _____0_445215(.DIN1 (________24039), .DIN2 (___00___23439), .Q
       (___0____24414));
  or2s1 _____0_445216(.DIN1 (___0____24412), .DIN2 (________24028), .Q
       (___0____24413));
  nor2s1 _____0_445217(.DIN1 (____9___19395), .DIN2 (________24025), .Q
       (___0____24411));
  or2s1 _____445218(.DIN1 (________23824), .DIN2 (___9____24317), .Q
       (___0_0__24410));
  or2s1 _____445219(.DIN1 (___0____24408), .DIN2 (________24032), .Q
       (___0_9__24409));
  nor2s1 _____9_445220(.DIN1 (____0___22901), .DIN2 (___0____24406), .Q
       (___0____24407));
  nor2s1 _____9_445221(.DIN1 (________22979), .DIN2 (___0_0__24391), .Q
       (___0____24405));
  nnd2s1 _______445222(.DIN1 (________24084), .DIN2 (___0____24403), .Q
       (___0____24404));
  and2s1 _____9_445223(.DIN1 (___0____24416), .DIN2 (___0____24350), .Q
       (___0____24402));
  nnd2s1 _______445224(.DIN1 (___0____24364), .DIN2 (_________34866),
       .Q (___0____24401));
  nor2s1 _______445225(.DIN1 (___0____24398), .DIN2 (________23990), .Q
       (___0____24399));
  nnd2s1 _____445226(.DIN1 (________24112), .DIN2
       (_________________18702), .Q (___0____24397));
  nnd2s1 _______445227(.DIN1 (________24222), .DIN2 (inData[12]), .Q
       (___0____24396));
  nor2s1 _______445228(.DIN1 (________23670), .DIN2 (________24015), .Q
       (___0____24395));
  nnd2s1 ______445229(.DIN1 (________24046), .DIN2 (___0____24393), .Q
       (___0____24394));
  or2s1 ______445230(.DIN1 (___0_0__24391), .DIN2 (________23848), .Q
       (___0____24392));
  nor2s1 _______445231(.DIN1 (___0____24389), .DIN2 (____0___24067), .Q
       (___0_9__24390));
  and2s1 _______445232(.DIN1 (____9___24056), .DIN2 (___99___25268), .Q
       (___0____24388));
  nnd2s1 _______445233(.DIN1 (_____9__24110), .DIN2 (___0____24386), .Q
       (___0____24387));
  nor2s1 _______445234(.DIN1 (________24221), .DIN2 (________24109), .Q
       (___0____24385));
  nor2s1 ______445235(.DIN1 (________22135), .DIN2 (___00___24341), .Q
       (___0____24384));
  nnd2s1 _______445236(.DIN1 (________24107), .DIN2 (___0_0__24382), .Q
       (___0____24383));
  nnd2s1 _______445237(.DIN1 (____9___24055), .DIN2 (___00___24336), .Q
       (___0_9__24381));
  nnd2s1 ______445238(.DIN1 (________24114), .DIN2 (____0___25661), .Q
       (___0____24380));
  or2s1 ______445239(.DIN1 (___0____24378), .DIN2 (________24106), .Q
       (___0____24379));
  nnd2s1 _______445240(.DIN1 (_____0__24072), .DIN2 (_____0__23942), .Q
       (___0____24377));
  nnd2s1 _______445241(.DIN1 (__9__0__27025), .DIN2 (________24103), .Q
       (___0____24376));
  and2s1 _______445242(.DIN1 (________24050), .DIN2 (___0____24374), .Q
       (___0____24375));
  nor2s1 _______445243(.DIN1 (___0), .DIN2 (___0_0__24372), .Q
       (___0____24373));
  nnd2s1 _______445244(.DIN1 (________24016), .DIN2 (________23321), .Q
       (___0_9__24371));
  nnd2s1 _______445245(.DIN1 (________23987), .DIN2 (___9____23384), .Q
       (___0____24370));
  or2s1 ______445246(.DIN1 (___0____24368), .DIN2 (________24096), .Q
       (___0____24369));
  nor2s1 _______445247(.DIN1 (________25812), .DIN2 (_____0__24092), .Q
       (___0____24367));
  nor2s1 _______445248(.DIN1 (________25027), .DIN2 (________24228), .Q
       (___0____24366));
  nnd2s1 _______445249(.DIN1 (___0____24364), .DIN2 (________24077), .Q
       (___0____24365));
  or2s1 _______445250(.DIN1 (________25010), .DIN2 (___0_0__24362), .Q
       (___0____24363));
  and2s1 ______445251(.DIN1 (____9___24059), .DIN2 (_________34956), .Q
       (___0_9__24361));
  and2s1 _____9_445252(.DIN1 (________24049), .DIN2 (________24726), .Q
       (___0____24360));
  or2s1 _____9_445253(.DIN1 (________24142), .DIN2 (___0____24358), .Q
       (___0____24359));
  nor2s1 _____9_445254(.DIN1 (_____0__25712), .DIN2 (____9___24061), .Q
       (___0____24357));
  and2s1 _____0_445255(.DIN1 (___0____24355), .DIN2 (________25717), .Q
       (___0____24356));
  nor2s1 _____0_445256(.DIN1 (________25413), .DIN2 (_____0__24082), .Q
       (___0____24354));
  nor2s1 _______445257(.DIN1 (___0_0__24352), .DIN2 (________24076), .Q
       (___0____24353));
  and2s1 _______445258(.DIN1 (________23989), .DIN2 (___0____24350), .Q
       (___0_9__24351));
  nnd2s1 _______445259(.DIN1 (________24469), .DIN2 (____0___24070), .Q
       (___0____24349));
  nor2s1 _______445260(.DIN1 (________23853), .DIN2 (________24104), .Q
       (___0____24348));
  nor2s1 _______445261(.DIN1 (____0___24069), .DIN2 (_____0__25616), .Q
       (___0____24347));
  nor2s1 _______445262(.DIN1 (____9___23970), .DIN2 (________24095), .Q
       (___0____24346));
  nor2s1 _______445263(.DIN1 (___0____22609), .DIN2 (________24097), .Q
       (___0____24345));
  nor2s1 _______445264(.DIN1 (___0_0__24343), .DIN2 (_____0__24027), .Q
       (___0____24344));
  nor2s1 _______445265(.DIN1 (___00___24341), .DIN2 (___00___24340), .Q
       (___009__24342));
  nnd2s1 ______445266(.DIN1 (________24469), .DIN2 (____0___24064), .Q
       (___00___24339));
  nnd2s1 _______445267(.DIN1 (___9____24320), .DIN2 (________23005), .Q
       (___00___24338));
  nnd2s1 _______445268(.DIN1 (___00___24336), .DIN2 (_____9__24091), .Q
       (___00___24337));
  nor2s1 _____9_445269(.DIN1 (___00___24334), .DIN2 (____99__24062), .Q
       (___00___24335));
  nnd2s1 _______445270(.DIN1 (________24116), .DIN2 (_____9__25528), .Q
       (___000__24333));
  nor2s1 _______445271(.DIN1 (___99___24331), .DIN2 (________24009), .Q
       (___999__24332));
  nor2s1 _______445272(.DIN1 (___99___24329), .DIN2 (_________34872),
       .Q (___99___24330));
  xor2s1 ______445273(.DIN1 (_________________0___18607), .DIN2
       (________24546), .Q (___99___24328));
  nnd2s1 _______445274(.DIN1 (________24005), .DIN2 (___0____24374), .Q
       (___99___24327));
  nor2s1 _______445275(.DIN1 (________23927), .DIN2 (____0___24068), .Q
       (___990__24326));
  nnd2s1 _______445276(.DIN1 (________24051), .DIN2 (________25139), .Q
       (___9_9__24325));
  nnd2s1 ______445277(.DIN1 (________24086), .DIN2 (___9____24323), .Q
       (___9____24324));
  nnd2s1 _______445278(.DIN1 (________24019), .DIN2 (____9___22889), .Q
       (___9____24322));
  nor2s1 _______445279(.DIN1 (____0___23716), .DIN2 (___9____24320), .Q
       (___9____24321));
  nnd2s1 _______445280(.DIN1 (____0___23712), .DIN2 (________24098), .Q
       (___9____24319));
  nnd2s1 ____0__445281(.DIN1 (____9___24510), .DIN2 (___9____24318), .Q
       (___0_____27709));
  nnd2s1 _______445282(.DIN1 (________24078), .DIN2 (___900__26147), .Q
       (________24850));
  nnd2s1 _______445283(.DIN1 (_____0__24102), .DIN2 (_____9__22022), .Q
       (___0_____27406));
  nor2s1 _______445284(.DIN1 (____0___24990), .DIN2 (___9____24317), .Q
       (________24871));
  nor2s1 ____0__445285(.DIN1 (________25389), .DIN2 (________23923), .Q
       (____0___24893));
  nnd2s1 ____0__445286(.DIN1 (____9___24510), .DIN2 (________22866), .Q
       (________24742));
  and2s1 ____0__445287(.DIN1 (________23934), .DIN2 (____9___25742), .Q
       (________24775));
  nor2s1 ____0__445288(.DIN1 (________22382), .DIN2 (________24458), .Q
       (________24692));
  nor2s1 ____0_445289(.DIN1 (_________31926), .DIN2
       (_______________18884), .Q (________24820));
  nor2s1 ____0__445290(.DIN1 (________25513), .DIN2 (________25989), .Q
       (_____9__24838));
  nor2s1 ____0__445291(.DIN1 (_____9__24119), .DIN2 (_________32344),
       .Q (____9___24784));
  nnd2s1 ____0_445292(.DIN1 (_______________18884), .DIN2
       (_________30612), .Q (_________31126));
  nnd2s1 ____0_445293(.DIN1 (________23904), .DIN2 (___9_9__22516), .Q
       (___0_0___27755));
  nnd2s1 ____0__445294(.DIN1 (________23904), .DIN2 (___99___23434), .Q
       (__9__0__26394));
  nor2s1 ____0_445295(.DIN1 (________24557), .DIN2 (________24458), .Q
       (___0_____27811));
  and2s1 ____0__445296(.DIN1 (____9___24510), .DIN2 (___9_0__24316), .Q
       (___0_____27281));
  nor2s1 ____0__445297(.DIN1 (_____0__24219), .DIN2 (___9_9__24315), .Q
       (_________31949));
  nor2s1 ____0__445298(.DIN1 (________24094), .DIN2 (________24458), .Q
       (___0_____27477));
  nnd2s1 ____0__445299(.DIN1 (________24469), .DIN2 (___9____24314), .Q
       (__9_____26812));
  nnd2s1 ____0_445300(.DIN1 (________23903), .DIN2 (___9____24313), .Q
       (________25874));
  and2s1 ____0__445301(.DIN1 (__90____26306), .DIN2 (________26074), .Q
       (___90___26151));
  nnd2s1 ____0__445302(.DIN1 (________23904), .DIN2 (____9___22800), .Q
       (________25643));
  nor2s1 ____0__445303(.DIN1 (_____0__21103), .DIN2 (_____0__25616), .Q
       (___0_____27698));
  nnd2s1 ______445304(.DIN1 (____0___23895), .DIN2 (___0____22614), .Q
       (___9____24312));
  nnd2s1 _______445305(.DIN1 (________24169), .DIN2 (________23759), .Q
       (___9____24311));
  nnd2s1 _______445306(.DIN1 (________23861), .DIN2 (________24003), .Q
       (___9____24310));
  nor2s1 _______445307(.DIN1 (___0____22606), .DIN2 (________23865), .Q
       (___9____24309));
  or2s1 ____9__445308(.DIN1 (___0_9___27748), .DIN2 (_____9__23774), .Q
       (___9____24308));
  xor2s1 _______445309(.DIN1 (_________________0___18633), .DIN2
       (_________31667), .Q (___9____24307));
  xor2s1 _______445310(.DIN1 (________22320), .DIN2 (_________31667),
       .Q (___9_0__24306));
  nnd2s1 ____9__445311(.DIN1 (____0____28221), .DIN2 (___9____24304),
       .Q (___9_9__24305));
  nor2s1 _______445312(.DIN1 (inData[18]), .DIN2 (___9____24302), .Q
       (___9____24303));
  nnd2s1 ______445313(.DIN1 (____0___23714), .DIN2 (___9____24300), .Q
       (___9____24301));
  and2s1 _______445314(.DIN1 (________23741), .DIN2 (___9____24298), .Q
       (___9____24299));
  nor2s1 _______445315(.DIN1 (_________34474), .DIN2 (___9____24302),
       .Q (___9____24297));
  nnd2s1 _______445316(.DIN1 (_________34896), .DIN2 (________24619),
       .Q (___9_0__24296));
  or2s1 _______445317(.DIN1 (________23568), .DIN2 (_____9__23836), .Q
       (___9_9__24295));
  nor2s1 ______445318(.DIN1 (________23835), .DIN2 (___9____24293), .Q
       (___9____24294));
  nor2s1 ______445319(.DIN1 (____9___22710), .DIN2 (______0__34908), .Q
       (___9____24292));
  or2s1 _______445320(.DIN1 (___9____24290), .DIN2 (_____0__23828), .Q
       (___9____24291));
  nor2s1 _______445321(.DIN1 (_________9_______18811), .DIN2
       (_________31290), .Q (___9____24289));
  or2s1 _______445322(.DIN1 (________23682), .DIN2 (___9____24287), .Q
       (___9____24288));
  and2s1 _______445323(.DIN1 (______0__34888), .DIN2 (____99__23711),
       .Q (___9_0__24286));
  or2s1 _______445324(.DIN1 (___99___23435), .DIN2 (________23825), .Q
       (___9_9__24285));
  or2s1 _______445325(.DIN1 (______________18870), .DIN2
       (___9____24287), .Q (___9____24284));
  nnd2s1 _______445326(.DIN1 (______0__32006), .DIN2 (________19478),
       .Q (___9____24283));
  nor2s1 _______445327(.DIN1 (____9___23252), .DIN2 (________23782), .Q
       (___9____24282));
  or2s1 ______445328(.DIN1 (_____________9___18703), .DIN2
       (_________31290), .Q (___9____24281));
  nnd2s1 _______445329(.DIN1 (________23818), .DIN2 (___9____24279), .Q
       (___9____24280));
  nor2s1 ______445330(.DIN1 (___9____24277), .DIN2 (_________34886), .Q
       (___9____24278));
  nnd2s1 _____9_445331(.DIN1 (_____9__23876), .DIN2 (________19570), .Q
       (___9_0__24276));
  nnd2s1 _____445332(.DIN1 (________23813), .DIN2 (________23757), .Q
       (___9____24275));
  and2s1 _____0_445333(.DIN1 (_________31290), .DIN2
       (_________9_______18811), .Q (___9____24274));
  and2s1 _____0_445334(.DIN1 (________23558), .DIN2 (________23769), .Q
       (___9____24273));
  nnd2s1 _______445335(.DIN1 (____0___23810), .DIN2 (___9____24271), .Q
       (___9____24272));
  nor2s1 _______445336(.DIN1 (________22160), .DIN2 (___9____24269), .Q
       (___9____24270));
  nor2s1 _______445337(.DIN1 (___0____23446), .DIN2 (________24931), .Q
       (___9____24268));
  nor2s1 _______445338(.DIN1 (____9___22982), .DIN2 (________24931), .Q
       (___9_0__24267));
  nor2s1 _______445339(.DIN1 (___9____24265), .DIN2 (___9____23400), .Q
       (___9_9__24266));
  nor2s1 _______445340(.DIN1 (___9____24263), .DIN2 (________23841), .Q
       (___9____24264));
  nnd2s1 _______445341(.DIN1 (___0____24364), .DIN2 (____9___23613), .Q
       (___9____24262));
  nor2s1 _______445342(.DIN1 (___9____24260), .DIN2 (_________34902),
       .Q (___9____24261));
  nnd2s1 _______445343(.DIN1 (____0___23808), .DIN2 (___9____24298), .Q
       (___9____24259));
  nor2s1 _______445344(.DIN1 (__9_____26764), .DIN2 (________23849), .Q
       (___9____24258));
  nor2s1 ______445345(.DIN1 (inData[0]), .DIN2 (_________29386), .Q
       (___9_0__24257));
  or2s1 ______445346(.DIN1 (___0_0__23490), .DIN2 (________23832), .Q
       (___9_9__24256));
  nnd2s1 _______445347(.DIN1 (________23745), .DIN2 (____99__25750), .Q
       (___9____24255));
  nnd2s1 _______445348(.DIN1 (________23838), .DIN2 (inData[0]), .Q
       (___9____24254));
  nnd2s1 _______445349(.DIN1 (________23839), .DIN2 (________23043), .Q
       (___9____24252));
  nor2s1 ______445350(.DIN1 (___9____24250), .DIN2 (________23854), .Q
       (___9____24251));
  and2s1 _______445351(.DIN1 (________23787), .DIN2 (___909__24248), .Q
       (___9_0__24249));
  nor2s1 _______445352(.DIN1 (____9___22986), .DIN2 (________23830), .Q
       (___90___24247));
  nor2s1 _______445353(.DIN1 (___90___19686), .DIN2 (___9____24302), .Q
       (___90___24246));
  nor2s1 _____9_445354(.DIN1 (________23052), .DIN2 (________23730), .Q
       (___90___24244));
  nnd2s1 _____9_445355(.DIN1 (________23874), .DIN2 (___90___24242), .Q
       (___90___24243));
  nor2s1 ____9_445356(.DIN1 (_____9__23325), .DIN2 (________23725), .Q
       (___900__24241));
  nor2s1 ____445357(.DIN1 (_____0___35032), .DIN2 (_________34904), .Q
       (____9___24240));
  nnd2s1 ____90_445358(.DIN1 (________23734), .DIN2 (____0___19400), .Q
       (____9___24239));
  nor2s1 ____90_445359(.DIN1 (____90__23250), .DIN2 (________24931), .Q
       (____9___24238));
  or2s1 ____90_445360(.DIN1 (_________34900), .DIN2 (________23596), .Q
       (____9___24237));
  nnd2s1 ____445361(.DIN1 (________23564), .DIN2 (_________34906), .Q
       (____9___24236));
  nnd2s1 _____9_445362(.DIN1 (________23918), .DIN2 (________23768), .Q
       (____90__24235));
  nor2s1 ______445363(.DIN1 (________21758), .DIN2 (________23722), .Q
       (_____9__24234));
  nor2s1 _______445364(.DIN1 (________23724), .DIN2 (________24232), .Q
       (________24233));
  and2s1 _______445365(.DIN1 (________23739), .DIN2 (________24230), .Q
       (________24231));
  nor2s1 _______445366(.DIN1 (____0___19400), .DIN2 (_____9__23764), .Q
       (_____0__24227));
  nnd2s1 _______445367(.DIN1 (________23743), .DIN2 (________22777), .Q
       (________24226));
  nnd2s1 _______445368(.DIN1 (________23777), .DIN2 (________23069), .Q
       (________24225));
  nnd2s1 ______445369(.DIN1 (___0____24364), .DIN2 (________23542), .Q
       (________24224));
  nor2s1 _______445370(.DIN1 (____0___22813), .DIN2 (_________34892),
       .Q (________24223));
  nnd2s1 _____0_445371(.DIN1 (_____9__23859), .DIN2 (_________35006),
       .Q (________24638));
  nor2s1 _______445372(.DIN1 (_________34488), .DIN2 (___9____24302),
       .Q (________24438));
  hi1s1 ______445373(.DIN (________24222), .Q (____9___24600));
  and2s1 ______445374(.DIN1 (_________34890), .DIN2 (_____90__34918),
       .Q (_____9__24569));
  nnd2s1 _______445375(.DIN1 (________23772), .DIN2 (________24221), .Q
       (___0__0__27890));
  and2s1 _______445376(.DIN1 (_____9__23827), .DIN2 (____9___25742), .Q
       (________24580));
  nor2s1 _______445377(.DIN1 (______9__28588), .DIN2 (________23816),
       .Q (___0_____27705));
  nor2s1 ______445378(.DIN1 (____9___23253), .DIN2 (___9____24269), .Q
       (__999___27167));
  and2s1 _______445379(.DIN1 (____0___23807), .DIN2 (___09____28078),
       .Q (____09___28232));
  nnd2s1 _______445380(.DIN1 (________24220), .DIN2 (________22060), .Q
       (________24536));
  nor2s1 ______445381(.DIN1 (____0__19016), .DIN2 (___9____24302), .Q
       (_____9__24635));
  nnd2s1 ______445382(.DIN1 (______0__32006), .DIN2 (_____0__24219), .Q
       (_________32053));
  nnd2s1 _______445383(.DIN1 (________24546), .DIN2 (___9____24300), .Q
       (________24585));
  nor2s1 ______445384(.DIN1 (________22322), .DIN2 (___9____24269), .Q
       (___0_____27631));
  nor2s1 ____9__445385(.DIN1 (___9_0__26157), .DIN2 (_____9__24139), .Q
       (_____9__24218));
  and2s1 ____9_445386(.DIN1 (_____0__23756), .DIN2 (________24216), .Q
       (________24217));
  or2s1 ____9_445387(.DIN1 (___0_9__25318), .DIN2 (________23748), .Q
       (________24215));
  nor2s1 ____9__445388(.DIN1 (____0___19400), .DIN2 (_____9__23746), .Q
       (________24214));
  nor2s1 ____9__445389(.DIN1 (________19520), .DIN2 (_____9__23784), .Q
       (________24213));
  nnd2s1 ____9__445390(.DIN1 (___9____24302), .DIN2 (_________31926),
       .Q (________24212));
  nor2s1 ____9_445391(.DIN1 (___0____22576), .DIN2 (___9____24269), .Q
       (________24211));
  or2s1 ____9__445392(.DIN1 (___9_0__19755), .DIN2 (___9____24287), .Q
       (________24210));
  nor2s1 ____9__445393(.DIN1 (___09___22624), .DIN2 (___9____24269), .Q
       (_____0__24209));
  and2s1 ____9__445394(.DIN1 (___0____24364), .DIN2 (________24207), .Q
       (_____9__24208));
  nor2s1 ____9_445395(.DIN1 (________24205), .DIN2 (________23993), .Q
       (________24206));
  and2s1 ____9__445396(.DIN1 (_________31261), .DIN2 (___0____19812),
       .Q (________24204));
  nnd2s1 ____9__445397(.DIN1 (________23776), .DIN2 (________24202), .Q
       (________24203));
  or2s1 ____9__445398(.DIN1 (________24200), .DIN2 (________23732), .Q
       (________24201));
  nnd2s1 ____9__445399(.DIN1 (________23766), .DIN2 (_____9__24198), .Q
       (_____0__24199));
  nor2s1 ____9__445400(.DIN1 (____0___23888), .DIN2 (________23873), .Q
       (________24197));
  nor2s1 ____9__445401(.DIN1 (________24195), .DIN2 (___9____24269), .Q
       (________24196));
  nnd2s1 ____9__445402(.DIN1 (_____0__23728), .DIN2 (________24221), .Q
       (________24194));
  or2s1 ____9__445403(.DIN1 (________23779), .DIN2 (________24192), .Q
       (________24193));
  nor2s1 ____9_445404(.DIN1 (________22213), .DIN2 (_________34902), .Q
       (________24191));
  nor2s1 ____9__445405(.DIN1 (_________34904), .DIN2 (___9____23410),
       .Q (_____0__24190));
  nor2s1 ____9__445406(.DIN1 (_____9__21923), .DIN2 (_____0__23737), .Q
       (________24189));
  and2s1 ____9__445407(.DIN1 (___0____24364), .DIN2 (___9____24318), .Q
       (________24188));
  nor2s1 ____99_445408(.DIN1 (_____9__23727), .DIN2 (___9____23409), .Q
       (________24187));
  nor2s1 ____99_445409(.DIN1 (________22963), .DIN2 (________24931), .Q
       (________24186));
  nor2s1 ____445410(.DIN1 (________23128), .DIN2 (_____0__23720), .Q
       (________24185));
  or2s1 ____00_445411(.DIN1 (________24183), .DIN2 (________23750), .Q
       (________24184));
  nor2s1 ____00_445412(.DIN1 (_____9__24181), .DIN2 (____0___23803), .Q
       (_____0__24182));
  nnd2s1 ____00_445413(.DIN1 (______0__32006), .DIN2 (________19651),
       .Q (________24180));
  nor2s1 _______445414(.DIN1 (_________34962), .DIN2 (________23864),
       .Q (________24179));
  and2s1 _______445415(.DIN1 (________23858), .DIN2 (________24177), .Q
       (________24178));
  nnd2s1 ____0__445416(.DIN1 (_____0___35109), .DIN2 (_________31926),
       .Q (________24176));
  or2s1 _______445417(.DIN1 (________23699), .DIN2 (________24124), .Q
       (________24175));
  or2s1 _____445418(.DIN1 (_____0__24173), .DIN2 (________23789), .Q
       (________24174));
  nor2s1 _____9_445419(.DIN1 (________24171), .DIN2 (________24030), .Q
       (_____9__24172));
  nnd2s1 _______445420(.DIN1 (________24169), .DIN2 (____9___23799), .Q
       (________24170));
  nor2s1 _______445421(.DIN1 (___0____24412), .DIN2 (____9___23878), .Q
       (________24168));
  nnd2s1 _______445422(.DIN1 (____99__23886), .DIN2 (________25115), .Q
       (________24167));
  nnd2s1 _______445423(.DIN1 (________24165), .DIN2 (_____0__24163), .Q
       (________24166));
  nor2s1 ______445424(.DIN1 (_____0__24163), .DIN2 (________24165), .Q
       (________24164));
  nor2s1 _______445425(.DIN1 (________24207), .DIN2 (____00__23887), .Q
       (____09__24162));
  nor2s1 _____9_445426(.DIN1 (____0___24160), .DIN2 (____0___24159), .Q
       (____0___24161));
  nor2s1 _____9_445427(.DIN1 (____0___24157), .DIN2 (________23956), .Q
       (____0___24158));
  or2s1 _____445428(.DIN1 (____0___24155), .DIN2 (_____0__23897), .Q
       (____0___24156));
  nnd2s1 ______445429(.DIN1 (____9___23708), .DIN2 (________25864), .Q
       (____9___24153));
  and2s1 _______445430(.DIN1 (_________34910), .DIN2 (____9___24151),
       .Q (____9___24152));
  hi1s1 _______445431(.DIN (____9___24149), .Q (____9___24150));
  and2s1 _______445432(.DIN1 (____0___23892), .DIN2 (___0_____27410),
       .Q (____9___24148));
  and2s1 _______445433(.DIN1 (________24146), .DIN2 (_____0__23915), .Q
       (_____9__24147));
  and2s1 _______445434(.DIN1 (____9___23884), .DIN2 (________24144), .Q
       (________24145));
  or2s1 ____90_445435(.DIN1 (____9___22444), .DIN2 (________24142), .Q
       (________24143));
  and2s1 _____9_445436(.DIN1 (_____0__24140), .DIN2 (_____9__24139), .Q
       (________24141));
  nor2s1 _______445437(.DIN1 (____0___22991), .DIN2 (________24126), .Q
       (________24138));
  nnd2s1 _____0_445438(.DIN1 (________24031), .DIN2 (________23014), .Q
       (________24137));
  or2s1 _______445439(.DIN1 (________24135), .DIN2 (____9___23880), .Q
       (________24136));
  or2s1 _____0_445440(.DIN1 (___0____23488), .DIN2 (____0___23893), .Q
       (________24134));
  or2s1 ______445441(.DIN1 (________24132), .DIN2 (____9___23705), .Q
       (________24133));
  and2s1 _______445442(.DIN1 (____0___23890), .DIN2 (________23235), .Q
       (________24131));
  nor2s1 _______445443(.DIN1 (________23867), .DIN2 (________25033), .Q
       (_____0__24130));
  or2s1 _______445444(.DIN1 (_________29585), .DIN2 (________23901), .Q
       (_____9__24129));
  nnd2s1 _______445445(.DIN1 (____9___23881), .DIN2
       (______________________________________0_____________18890), .Q
       (________24128));
  nor2s1 _______445446(.DIN1 (___9_0__23376), .DIN2 (________24126), .Q
       (________24127));
  nor2s1 ______445447(.DIN1 (________23997), .DIN2 (________24124), .Q
       (________24125));
  nnd2s1 ______445448(.DIN1 (_____0__23276), .DIN2 (________23863), .Q
       (________24123));
  nnd2s1 ______445449(.DIN1 (____9___23706), .DIN2 (________24122), .Q
       (___0__0__27637));
  hi1s1 _______445450(.DIN (________24121), .Q (____0____28219));
  nnd2s1 ____0_445451(.DIN1 (_________31290), .DIN2
       (___________0___18883), .Q (_____9___31088));
  nor2s1 ____0__445452(.DIN1 (_________31926), .DIN2 (_____0___35109),
       .Q (________25101));
  nor2s1 ____0__445453(.DIN1 (____0___23804), .DIN2 (________24546), .Q
       (________24466));
  nnd2s1 _______445454(.DIN1 (____0___23889), .DIN2 (_____0__24120), .Q
       (___0_9__24400));
  nnd2s1 ______445455(.DIN1 (________23790), .DIN2 (___909__22454), .Q
       (________24661));
  nor2s1 ____0__445456(.DIN1
       (______________________________________0_____________18887),
       .DIN2 (_________31290), .Q (_____0__24465));
  nor2s1 ____0__445457(.DIN1 (________21822), .DIN2 (___9____24269), .Q
       (___0__0__27994));
  or2s1 ____0__445458(.DIN1 (____99__25750), .DIN2 (___9____24269), .Q
       (___0_____27536));
  nor2s1 ____0__445459(.DIN1 (________25389), .DIN2 (____90__23877), .Q
       (________24629));
  nnd2s1 ____0__445460(.DIN1 (_________29386), .DIN2 (_____9__24119),
       .Q (_________32356));
  or2s1 ____0__445461(.DIN1 (________24118), .DIN2 (________23786), .Q
       (________25110));
  hi1s1 ____09_445462(.DIN (____9___24510), .Q (________24733));
  hi1s1 ____09_445463(.DIN (________24592), .Q (________24689));
  hi1s1 ____09_445464(.DIN (________24117), .Q (____9___24698));
  and2s1 _____445465(.DIN1 (________24115), .DIN2 (________23149), .Q
       (________24116));
  and2s1 _______445466(.DIN1 (________23657), .DIN2 (________24113), .Q
       (________24114));
  nor2s1 _______445467(.DIN1 (_______18957), .DIN2 (________24111), .Q
       (________24112));
  and2s1 _______445468(.DIN1 (_____9__23563), .DIN2 (________25806), .Q
       (_____9__24110));
  nor2s1 _______445469(.DIN1 (_________34986), .DIN2 (________23538),
       .Q (________24109));
  nnd2s1 ______445470(.DIN1 (________23659), .DIN2 (inData[4]), .Q
       (________24108));
  nor2s1 _______445471(.DIN1 (________23577), .DIN2 (________23851), .Q
       (________24107));
  or2s1 _______445472(.DIN1 (________24105), .DIN2 (________23651), .Q
       (________24106));
  or2s1 _______445473(.DIN1 (________22820), .DIN2 (_____9__23655), .Q
       (________24104));
  nor2s1 _______445474(.DIN1 (________23680), .DIN2 (________23329), .Q
       (________24103));
  nnd2s1 _______445475(.DIN1 (_____0__23999), .DIN2 (________19520), .Q
       (_____0__24102));
  or2s1 _______445476(.DIN1 (________24100), .DIN2 (_____9__23843), .Q
       (_____9__24101));
  nnd2s1 _______445477(.DIN1 (________23649), .DIN2 (_____9__23646), .Q
       (________24099));
  nnd2s1 ______445478(.DIN1 (________23640), .DIN2 (____9___19395), .Q
       (________24098));
  nnd2s1 _______445479(.DIN1 (_____0__23685), .DIN2 (________23698), .Q
       (________24097));
  or2s1 _______445480(.DIN1 (________25582), .DIN2 (________23643), .Q
       (________24096));
  nnd2s1 _______445481(.DIN1 (________24094), .DIN2 (____9___23612), .Q
       (________24095));
  nor2s1 _____445482(.DIN1 (________23287), .DIN2 (________23540), .Q
       (________24093));
  or2s1 _____9_445483(.DIN1 (________25793), .DIN2 (________23671), .Q
       (_____0__24092));
  and2s1 _____9_445484(.DIN1 (________24090), .DIN2 (________24089), .Q
       (_____9__24091));
  nor2s1 _____0_445485(.DIN1 (________24087), .DIN2 (_____0__23545), .Q
       (________24088));
  nor2s1 _____0_445486(.DIN1 (____9___25652), .DIN2 (________23631), .Q
       (________24086));
  nnd2s1 _____0_445487(.DIN1 (________23630), .DIN2 (___9____23394), .Q
       (________24085));
  nor2s1 _______445488(.DIN1 (________24083), .DIN2 (___9____23372), .Q
       (________24084));
  nnd2s1 _______445489(.DIN1 (________23669), .DIN2 (_____9__24198), .Q
       (_____0__24082));
  nnd2s1 _______445490(.DIN1 (____9___23611), .DIN2 (________21960), .Q
       (_____9__24081));
  or2s1 _______445491(.DIN1 (________24079), .DIN2 (________23688), .Q
       (________24080));
  nor2s1 _______445492(.DIN1 (_____0__25997), .DIN2 (____0___23621), .Q
       (________24078));
  nnd2s1 _______445493(.DIN1 (________23653), .DIN2 (___9_0__26177), .Q
       (________24077));
  or2s1 _______445494(.DIN1 (________24075), .DIN2 (________23594), .Q
       (________24076));
  and2s1 _______445495(.DIN1 (____9___23616), .DIN2 (________24073), .Q
       (________24074));
  nnd2s1 _______445496(.DIN1 (____09__24071), .DIN2 (____0___19400), .Q
       (_____0__24072));
  nnd2s1 _______445497(.DIN1 (________23788), .DIN2 (__9_____26354), .Q
       (____0___24070));
  nor2s1 _______445498(.DIN1 (_____9__22233), .DIN2 (________23988), .Q
       (____0___24069));
  nnd2s1 ______445499(.DIN1 (____9___23614), .DIN2 (____0___23809), .Q
       (____0___24068));
  nnd2s1 _______445500(.DIN1 (________23781), .DIN2 (________23216), .Q
       (____0___24067));
  nor2s1 _______445501(.DIN1 (____0___24065), .DIN2 (____90__23609), .Q
       (____0___24066));
  nnd2s1 _______445502(.DIN1 (________23549), .DIN2 (____0___25465), .Q
       (____0___24064));
  nor2s1 ______445503(.DIN1 (____9___24054), .DIN2 (_____0__23765), .Q
       (____00__24063));
  nnd2s1 _______445504(.DIN1 (_____9__23600), .DIN2 (________25717), .Q
       (____99__24062));
  or2s1 _______445505(.DIN1 (____9___24060), .DIN2 (________23599), .Q
       (____9___24061));
  and2s1 _______445506(.DIN1 (____9___24058), .DIN2 (____9___24057), .Q
       (____9___24059));
  nor2s1 _____445507(.DIN1 (____0___21907), .DIN2 (________23844), .Q
       (____9___24056));
  nor2s1 _____9_445508(.DIN1 (____9___24054), .DIN2 (____90__24053), .Q
       (____9___24055));
  nor2s1 _____9_445509(.DIN1 (___0____23452), .DIN2 (________23602), .Q
       (_____9__24052));
  and2s1 _____9_445510(.DIN1 (____0___25566), .DIN2 (_________34916),
       .Q (________24051));
  nor2s1 _____445511(.DIN1 (____0___23979), .DIN2 (________23998), .Q
       (________24050));
  nor2s1 _____0_445512(.DIN1 (___0____25336), .DIN2 (________23584), .Q
       (________24049));
  nnd2s1 _____0_445513(.DIN1 (___0____23456), .DIN2 (________23579), .Q
       (________24048));
  nor2s1 _____0_445514(.DIN1 (_________30612), .DIN2 (_________32122),
       .Q (________24047));
  and2s1 _____0_445515(.DIN1 (________23598), .DIN2 (_____9___35026),
       .Q (________24046));
  nnd2s1 _____9_445516(.DIN1 (_____0__24044), .DIN2 (____0___22266), .Q
       (________24045));
  nnd2s1 _______445517(.DIN1 (____0___23625), .DIN2 (________23814), .Q
       (_____9__24043));
  xnr2s1 ____0__445518(.DIN1 (outData[0]), .DIN2 (____9____30874), .Q
       (________24042));
  xor2s1 ____0_445519(.DIN1 (_________18864), .DIN2 (______9__28560),
       .Q (________24041));
  nor2s1 ____00_445520(.DIN1 (________23588), .DIN2 (___0____23501), .Q
       (________24040));
  and2s1 ____99_445521(.DIN1 (_____0__24140), .DIN2 (________23592), .Q
       (________24039));
  nnd2s1 ____445522(.DIN1 (________23585), .DIN2 (___0____23475), .Q
       (________24038));
  nor2s1 ____9__445523(.DIN1 (________24036), .DIN2 (_____0__24035), .Q
       (________24037));
  nnd2s1 ____9__445524(.DIN1 (_________34914), .DIN2 (__90____26310),
       .Q (_____9__24034));
  nnd2s1 ____9__445525(.DIN1 (________23672), .DIN2 (_________31618),
       .Q (________24033));
  nnd2s1 ____9_445526(.DIN1 (____0___23531), .DIN2 (___9_0__22500), .Q
       (________24032));
  nnd2s1 _______445527(.DIN1 (________23629), .DIN2 (________24221), .Q
       (________24029));
  nnd2s1 _______445528(.DIN1 (________23636), .DIN2 (____9___23879), .Q
       (________24028));
  nnd2s1 _______445529(.DIN1 (____0___23619), .DIN2 (________23697), .Q
       (_____0__24027));
  nnd2s1 _______445530(.DIN1 (________24022), .DIN2 (____90__19196), .Q
       (_____9__24026));
  nor2s1 _______445531(.DIN1 (________22817), .DIN2 (____0___23533), .Q
       (________24025));
  nnd2s1 _______445532(.DIN1 (________24022), .DIN2 (_________28828),
       .Q (________24023));
  or2s1 ______445533(.DIN1 (_____0__25156), .DIN2 (_____0__23555), .Q
       (________24021));
  nnd2s1 _______445534(.DIN1 (________23551), .DIN2 (____0___24890), .Q
       (________24020));
  nor2s1 _______445535(.DIN1 (_____0__23572), .DIN2 (________23334), .Q
       (________24019));
  nnd2s1 _____9_445536(.DIN1 (________23570), .DIN2 (____99__22171), .Q
       (_____0__24018));
  nor2s1 _____9_445537(.DIN1 (___0____23474), .DIN2 (________23546), .Q
       (_____9__24017));
  nor2s1 ____9__445538(.DIN1 (___9____25249), .DIN2 (________23550), .Q
       (________24016));
  nnd2s1 ____9__445539(.DIN1 (_____0__23785), .DIN2 (___9____23403), .Q
       (________24015));
  nnd2s1 ____9__445540(.DIN1 (________23783), .DIN2 (________19520), .Q
       (________24014));
  nor2s1 ____9__445541(.DIN1 (____9___23883), .DIN2 (_____0__23638), .Q
       (________24013));
  nnd2s1 ____9__445542(.DIN1 (________23862), .DIN2 (________23632), .Q
       (________24012));
  nnd2s1 ____9__445543(.DIN1 (________23633), .DIN2 (______0__34948),
       .Q (________24011));
  or2s1 ____9__445544(.DIN1 (____0___26055), .DIN2 (___0____23511), .Q
       (________24010));
  nnd2s1 ____9__445545(.DIN1 (_____0__24008), .DIN2 (_____9__24007), .Q
       (________24009));
  and2s1 ____9_445546(.DIN1 (________23687), .DIN2 (________24505), .Q
       (________24006));
  nor2s1 ____9__445547(.DIN1 (________25978), .DIN2 (________23575), .Q
       (________24005));
  or2s1 ____9__445548(.DIN1 (_________34974), .DIN2 (_________34912),
       .Q (________24004));
  nnd2s1 ____0__445549(.DIN1 (________24003), .DIN2 (________23098), .Q
       (___0_0__24362));
  nnd2s1 _______445550(.DIN1 (_________32122), .DIN2 (____0___19117),
       .Q (___0_0__24372));
  nor2s1 _______445551(.DIN1 (____________0___18686), .DIN2
       (________24111), .Q (________24222));
  or2s1 _______445552(.DIN1 (_____0__24541), .DIN2 (________24002), .Q
       (___00___24340));
  nnd2s1 _______445553(.DIN1 (________23634), .DIN2 (_________28602),
       .Q (___0____24358));
  nnd2s1 _______445554(.DIN1 (________24090), .DIN2 (__9_____26358), .Q
       (___00___24341));
  nnd2s1 _______445555(.DIN1 (____0___23623), .DIN2 (________24001), .Q
       (___0_0__24391));
  nnd2s1 ______445556(.DIN1 (___0____23515), .DIN2 (________24000), .Q
       (__99_0__27144));
  nor2s1 _______445557(.DIN1 (________23132), .DIN2 (_____0__23999), .Q
       (___9____24320));
  and2s1 ____0__445558(.DIN1 (_____9__23590), .DIN2 (_________35010),
       .Q (________24543));
  nnd2s1 ____0_445559(.DIN1 (___090__23518), .DIN2 (____9___21899), .Q
       (___9____24317));
  nor2s1 ____0_445560(.DIN1 (________25772), .DIN2 (________23998), .Q
       (___0____24355));
  nor2s1 ____0__445561(.DIN1 (________23997), .DIN2 (________23565), .Q
       (________24229));
  or2s1 ____0__445562(.DIN1 (__9_____26736), .DIN2 (________23547), .Q
       (___0____24406));
  nnd2s1 ____0__445563(.DIN1 (____0___23534), .DIN2 (_____9__22374), .Q
       (__990___27086));
  or2s1 _______445564(.DIN1 (______9__28588), .DIN2 (________23645), .Q
       (______0__28263));
  nnd2s1 ______445565(.DIN1 (_________32122), .DIN2 (________23996), .Q
       (_________32156));
  or2s1 _______445566(.DIN1 (________________18736), .DIN2
       (______0__32252), .Q (________23995));
  hi1s1 ____0_445567(.DIN (________23993), .Q (________23994));
  nor2s1 _______445568(.DIN1 (________19100), .DIN2 (_____9__23991), .Q
       (_____0__23992));
  or2s1 _____0_445569(.DIN1 (_____0__26057), .DIN2 (___0____23514), .Q
       (________23990));
  nor2s1 _______445570(.DIN1 (________22966), .DIN2 (________23988), .Q
       (________23989));
  or2s1 _______445571(.DIN1 (_________31281), .DIN2 (________25687), .Q
       (________23987));
  nnd2s1 ______445572(.DIN1 (___0_9__23454), .DIN2 (________23034), .Q
       (________23986));
  and2s1 ______445573(.DIN1 (_____9___34924), .DIN2 (________23654), .Q
       (________23985));
  or2s1 _______445574(.DIN1 (____9___21352), .DIN2 (________23912), .Q
       (________23984));
  nnd2s1 _______445575(.DIN1 (________23290), .DIN2 (____0___23981), .Q
       (____0___23982));
  nor2s1 _______445576(.DIN1 (________23753), .DIN2 (____0___23979), .Q
       (____0___23980));
  and2s1 ______445577(.DIN1 (_____9___30454), .DIN2 (____99__20039), .Q
       (____0___23978));
  nor2s1 ______445578(.DIN1 (___0____23451), .DIN2 (____9___22888), .Q
       (____0___23977));
  and2s1 _______445579(.DIN1 (_____9___30454), .DIN2 (_______19023), .Q
       (____0___23976));
  nnd2s1 _______445580(.DIN1 (_____9___30454), .DIN2 (________22239),
       .Q (____0___23975));
  or2s1 _______445581(.DIN1 (_____9__22942), .DIN2 (________23916), .Q
       (____00__23974));
  or2s1 _____445582(.DIN1 (____9___23971), .DIN2 (____9___23970), .Q
       (____9___23972));
  nor2s1 _______445583(.DIN1 (________23139), .DIN2 (___0____23468), .Q
       (____9___23969));
  or2s1 _______445584(.DIN1 (___0____23447), .DIN2 (____9___22891), .Q
       (____9___23968));
  nnd2s1 _______445585(.DIN1 (___0____23467), .DIN2 (_____9__23064), .Q
       (____9___23967));
  nor2s1 ______445586(.DIN1 (____90__23965), .DIN2 (___0____23460), .Q
       (____9___23966));
  or2s1 _______445587(.DIN1 (_________34986), .DIN2 (_____9__23941), .Q
       (_____9__23964));
  nor2s1 _______445588(.DIN1 (____0___21986), .DIN2 (_____9___34920),
       .Q (________23963));
  nor2s1 _______445589(.DIN1 (________23857), .DIN2 (________23961), .Q
       (________23962));
  nnd2s1 _______445590(.DIN1 (___0_0__23464), .DIN2 (____0___25470), .Q
       (________23960));
  or2s1 _______445591(.DIN1 (_____0__23958), .DIN2 (_____0__24044), .Q
       (________23959));
  nor2s1 ______445592(.DIN1 (____0___22993), .DIN2 (________23956), .Q
       (_____9__23957));
  nor2s1 ______445593(.DIN1 (____00__19399), .DIN2 (___0____23457), .Q
       (________23955));
  nor2s1 _______445594(.DIN1 (____9___22987), .DIN2 (___0____23458), .Q
       (________23954));
  or2s1 _____445595(.DIN1 (________24583), .DIN2 (___0____23466), .Q
       (________23953));
  or2s1 _______445596(.DIN1 (________22683), .DIN2 (_____0__23950), .Q
       (________23951));
  nor2s1 _______445597(.DIN1 (____0___23088), .DIN2 (________23948), .Q
       (________23949));
  and2s1 _______445598(.DIN1 (________23946), .DIN2 (_____9__23073), .Q
       (________23947));
  nnd2s1 _____445599(.DIN1 (________23909), .DIN2 (________23944), .Q
       (________23945));
  nnd2s1 _______445600(.DIN1 (___0____23504), .DIN2 (________22420), .Q
       (________23943));
  nnd2s1 _______445601(.DIN1 (_____9__23941), .DIN2 (________24221), .Q
       (_____0__23942));
  nnd2s1 _______445602(.DIN1 (___9____23408), .DIN2 (_____9__23189), .Q
       (________23940));
  and2s1 _______445603(.DIN1 (___00___23440), .DIN2 (________23938), .Q
       (________23939));
  nnd2s1 _______445604(.DIN1 (___0_0__23473), .DIN2 (____0___25758), .Q
       (________23937));
  nor2s1 _______445605(.DIN1 (________22940), .DIN2 (___9_0__25241), .Q
       (________23936));
  nor2s1 _______445606(.DIN1 (___9____23418), .DIN2 (____0___23175), .Q
       (________23935));
  and2s1 _______445607(.DIN1 (___9____23425), .DIN2 (_____0__23933), .Q
       (________23934));
  nor2s1 ______445608(.DIN1 (___99___23433), .DIN2 (___9____23423), .Q
       (________23931));
  nnd2s1 _______445609(.DIN1 (___0____23492), .DIN2 (________23929), .Q
       (________23930));
  nnd2s1 ______445610(.DIN1 (___0____23483), .DIN2 (________22918), .Q
       (________23928));
  or2s1 _______445611(.DIN1 (___9____19762), .DIN2 (______0__32252), .Q
       (________23926));
  nnd2s1 ______445612(.DIN1 (___0____23461), .DIN2 (________22853), .Q
       (_____0__23925));
  nnd2s1 _____9_445613(.DIN1 (___9____23420), .DIN2 (________22276), .Q
       (_____9__23924));
  nnd2s1 _____9_445614(.DIN1 (____0____34553), .DIN2 (________23922),
       .Q (________23923));
  and2s1 _____445615(.DIN1 (___0____23486), .DIN2 (________23920), .Q
       (________23921));
  and2s1 ____0__445616(.DIN1 (________23553), .DIN2 (___09____28074),
       .Q (________26123));
  or2s1 _______445617(.DIN1 (___99___23431), .DIN2 (___09_9__28080), .Q
       (_____0__24936));
  hi1s1 ____0__445618(.DIN (________24546), .Q (____0___24434));
  hi1s1 ____0_445619(.DIN (______0__32006), .Q (___9_9__24315));
  nnd2s1 ____0_445620(.DIN1 (________23918), .DIN2 (____9___23796), .Q
       (________24228));
  nnd2s1 ______445621(.DIN1 (________25049), .DIN2 (___0____23507), .Q
       (________24121));
  nnd2s1 ______445622(.DIN1 (___0____23479), .DIN2 (________23917), .Q
       (_____0__24447));
  nor2s1 _____0_445623(.DIN1 (___0____23505), .DIN2 (________23916), .Q
       (___0_____27902));
  nor2s1 _______445624(.DIN1 (___0____23496), .DIN2 (_____0__23294), .Q
       (___0_____27573));
  nnd2s1 _______445625(.DIN1 (________24474), .DIN2 (_____0__23915), .Q
       (____9___24149));
  nnd2s1 ______445626(.DIN1 (___00___23443), .DIN2 (________22862), .Q
       (___00____27235));
  or2s1 _______445627(.DIN1 (_____9__23914), .DIN2 (___0____23493), .Q
       (___0_____27966));
  nnd2s1 _______445628(.DIN1 (____0____28179), .DIN2 (________23913),
       .Q (________24959));
  and2s1 _______445629(.DIN1 (__9__9__26476), .DIN2 (_____9__22098), .Q
       (_________28381));
  nnd2s1 _______445630(.DIN1 (___0_9__23499), .DIN2 (___9____26223), .Q
       (________24492));
  nor2s1 ____0__445631(.DIN1 (________26008), .DIN2 (________23842), .Q
       (____9___25460));
  and2s1 _______445632(.DIN1 (___0_9__23472), .DIN2 (__9_____26623), .Q
       (________25866));
  nor2s1 ______445633(.DIN1 (_____0__26117), .DIN2 (________23912), .Q
       (____9___24981));
  nor2s1 _______445634(.DIN1 (___0_____27291), .DIN2 (___0____23459),
       .Q (___0_09__27665));
  nnd2s1 ____0__445635(.DIN1 (___0____23516), .DIN2 (__9_____26717), .Q
       (________25516));
  nor2s1 _______445636(.DIN1 (________23911), .DIN2 (___9____23424), .Q
       (__90____26306));
  nor2s1 ____0__445637(.DIN1 (________23910), .DIN2 (________23845), .Q
       (___0____24416));
  nnd2s1 ______445638(.DIN1 (________23909), .DIN2 (________21881), .Q
       (____0___24520));
  nnd2s1 _______445639(.DIN1 (________23902), .DIN2 (________23691), .Q
       (________24117));
  xor2s1 ____0__445640(.DIN1 (outData[2]), .DIN2 (outData[0]), .Q
       (________24547));
  nor2s1 _______445641(.DIN1 (________23908), .DIN2 (____0___23979), .Q
       (________25098));
  nor2s1 _______445642(.DIN1 (________23907), .DIN2 (________23696), .Q
       (_________28537));
  nnd2s1 _____445643(.DIN1 (____0___23981), .DIN2 (________23906), .Q
       (_________32219));
  nor2s1 ______445644(.DIN1 (___0____23494), .DIN2 (________23916), .Q
       (_________28832));
  or2s1 _______445645(.DIN1 (___9_0__26167), .DIN2 (___99___23428), .Q
       (________25989));
  hi1s1 _______445646(.DIN (________23905), .Q (____9____31787));
  hi1s1 ____09_445647(.DIN (________24931), .Q (________24469));
  nnd2s1 _____9_445648(.DIN1 (_____9___30454), .DIN2 (____9____32697),
       .Q (_________31303));
  hi1s1 _____0_445649(.DIN (________23905), .Q (_________35111));
  hi1s1 ____09_445650(.DIN (___9____24269), .Q (_____0__24481));
  hi1s1 ______445651(.DIN (_________29386), .Q (_________32344));
  nor2s1 ______445652(.DIN1 (________23690), .DIN2 (___0____23476), .Q
       (________24592));
  nnd2s1 ____0__445653(.DIN1 (________23641), .DIN2 (___9____20651), .Q
       (____0____31831));
  hi1s1 _____0_445654(.DIN (________23904), .Q (_____9__24755));
  hi1s1 ____09_445655(.DIN (___0____24364), .Q (________24458));
  hi1s1 ____09_445656(.DIN (________23903), .Q (_____0__25616));
  nor2s1 _______445657(.DIN1 (inData[23]), .DIN2 (________23902), .Q
       (____9___24510));
  nnd2s1 _______445658(.DIN1 (________23900), .DIN2 (inData[18]), .Q
       (________23901));
  nnd2s1 _______445659(.DIN1 (___9____23378), .DIN2 (inData[2]), .Q
       (________23899));
  nor2s1 _______445660(.DIN1 (___09___22622), .DIN2 (___9____23369), .Q
       (________23898));
  nnd2s1 _______445661(.DIN1 (___9_0__23356), .DIN2 (____9_0__33597),
       .Q (_____0__23897));
  or2s1 _______445662(.DIN1 (________24722), .DIN2 (_____0__24746), .Q
       (____09__23896));
  nor2s1 _____9_445663(.DIN1 (____0___23894), .DIN2 (___9____23382), .Q
       (____0___23895));
  nnd2s1 _____9_445664(.DIN1 (___9____23380), .DIN2 (________23292), .Q
       (____0___23893));
  nor2s1 _____445665(.DIN1 (____0___24160), .DIN2 (___9____23377), .Q
       (____0___23892));
  nnd2s1 _____0_445666(.DIN1 (____90__22885), .DIN2 (___9_9__23375), .Q
       (____0___23891));
  nor2s1 _____0_445667(.DIN1 (________23593), .DIN2 (____0___23174), .Q
       (____0___23890));
  nor2s1 _____445668(.DIN1 (____0___23888), .DIN2 (___0_____27303), .Q
       (____0___23889));
  or2s1 _______445669(.DIN1 (_____9__23302), .DIN2 (___900__23346), .Q
       (____00__23887));
  and2s1 _______445670(.DIN1 (___9____23360), .DIN2 (____9___23885), .Q
       (____99__23886));
  nor2s1 _______445671(.DIN1 (____9___23883), .DIN2 (________23333), .Q
       (____9___23884));
  and2s1 ______445672(.DIN1 (_________33241), .DIN2 (_________18847),
       .Q (____9___23882));
  and2s1 _____9_445673(.DIN1 (________23900), .DIN2 (inData[24]), .Q
       (____9___23881));
  nnd2s1 _____0_445674(.DIN1 (___9____23363), .DIN2 (____9___23879), .Q
       (____9___23880));
  or2s1 ______445675(.DIN1 (__9_____26440), .DIN2 (___9____23359), .Q
       (____9___23878));
  or2s1 _____9_445676(.DIN1 (___0____24378), .DIN2 (_____0___34936), .Q
       (____90__23877));
  nnd2s1 ______445677(.DIN1 (_____0__23317), .DIN2 (________23875), .Q
       (_____9__23876));
  nor2s1 _______445678(.DIN1 (____9___22799), .DIN2 (_____0__23775), .Q
       (________23874));
  or2s1 _______445679(.DIN1 (________23245), .DIN2 (________23872), .Q
       (________23873));
  xnr2s1 ______445680(.DIN1 (________20546), .DIN2 (____0____31820), .Q
       (________23870));
  nor2s1 _______445681(.DIN1 (____09__22634), .DIN2 (___90___23348), .Q
       (________23869));
  nnd2s1 ____9__445682(.DIN1 (________23866), .DIN2 (_____9__23335), .Q
       (________23867));
  nnd2s1 ____9__445683(.DIN1 (________23866), .DIN2 (________22705), .Q
       (________23865));
  or2s1 ____9_445684(.DIN1 (________23731), .DIN2 (_____9__23703), .Q
       (________23864));
  nnd2s1 ____9_445685(.DIN1 (________23862), .DIN2 (____90__23336), .Q
       (________23863));
  nor2s1 ____9__445686(.DIN1 (________23111), .DIN2 (_____0__23860), .Q
       (________23861));
  and2s1 ____99_445687(.DIN1 (____9___23337), .DIN2 (_____9__25634), .Q
       (_____9__23859));
  nor2s1 ____99_445688(.DIN1 (________23857), .DIN2 (___9____23374), .Q
       (________23858));
  nnd2s1 ____0_445689(.DIN1 (___9____20638), .DIN2 (____9___23340), .Q
       (________23856));
  nnd2s1 ____0__445690(.DIN1 (________23224), .DIN2 (____9_0__33597),
       .Q (________23855));
  or2s1 ______445691(.DIN1 (________23853), .DIN2 (____0___23172), .Q
       (________23854));
  nor2s1 _______445692(.DIN1 (________22228), .DIN2 (________23851), .Q
       (________23852));
  xor2s1 ____0__445693(.DIN1 (____0__19046), .DIN2 (____0____31820), .Q
       (_____0__23850));
  nnd2s1 _______445694(.DIN1 (________23304), .DIN2 (________24195), .Q
       (________23849));
  nnd2s1 _______445695(.DIN1 (___9____23426), .DIN2 (________22405), .Q
       (________23848));
  nor2s1 _______445696(.DIN1 (________23833), .DIN2 (________24549), .Q
       (________23847));
  nnd2s1 _______445697(.DIN1 (_____0__23747), .DIN2 (________23840), .Q
       (________23846));
  nnd2s1 _______445698(.DIN1 (________23205), .DIN2 (___9____24271), .Q
       (________23841));
  nnd2s1 _______445699(.DIN1 (____0___23260), .DIN2 (____09__22634), .Q
       (________23839));
  nor2s1 _______445700(.DIN1 (_________34436), .DIN2 (_____0__23837),
       .Q (________23838));
  nor2s1 _______445701(.DIN1 (inData[4]), .DIN2 (________23693), .Q
       (_____9__23836));
  nnd2s1 _______445702(.DIN1 (____90__23162), .DIN2 (________23272), .Q
       (________23835));
  nor2s1 _______445703(.DIN1 (________23193), .DIN2 (________23833), .Q
       (________23834));
  nnd2s1 _______445704(.DIN1 (________23587), .DIN2 (________23299), .Q
       (________23832));
  nnd2s1 _______445705(.DIN1 (_____0___34932), .DIN2 (_____0__22690),
       .Q (________23830));
  or2s1 _______445706(.DIN1 (________22015), .DIN2 (________23191), .Q
       (________23829));
  or2s1 ______445707(.DIN1 (_____9__22951), .DIN2 (________23742), .Q
       (_____0__23828));
  and2s1 _______445708(.DIN1 (________25007), .DIN2 (____00__22081), .Q
       (_____9__23827));
  or2s1 _______445709(.DIN1 (________23072), .DIN2 (________23150), .Q
       (________23826));
  or2s1 _______445710(.DIN1 (________23824), .DIN2 (____00__23259), .Q
       (________23825));
  nor2s1 _______445711(.DIN1 (____09__22634), .DIN2 (___0____23480), .Q
       (________23823));
  nor2s1 ______445712(.DIN1 (____9___23257), .DIN2 (______0__34938), .Q
       (________23822));
  nnd2s1 _______445713(.DIN1 (________23291), .DIN2 (_________32158),
       .Q (_____0__23821));
  or2s1 _______445714(.DIN1 (________21969), .DIN2 (________23301), .Q
       (_____9__23820));
  nor2s1 _______445715(.DIN1 (________23320), .DIN2 (________23269), .Q
       (________23819));
  nor2s1 _______445716(.DIN1 (________23203), .DIN2 (_____9__23151), .Q
       (________23818));
  or2s1 _____445717(.DIN1 (_____0__23215), .DIN2 (_________31920), .Q
       (________23817));
  nnd2s1 _____445718(.DIN1 (___9____24304), .DIN2 (___09_0__28051), .Q
       (________23816));
  nor2s1 _____445719(.DIN1 (________23814), .DIN2 (_____0__23312), .Q
       (________23815));
  nnd2s1 _____0_445720(.DIN1 (________23812), .DIN2 (_____0__23811), .Q
       (________23813));
  and2s1 _______445721(.DIN1 (____0___23809), .DIN2 (_____0__22291), .Q
       (____0___23810));
  and2s1 _______445722(.DIN1 (___9____23392), .DIN2 (________22691), .Q
       (____0___23808));
  and2s1 _______445723(.DIN1 (____0___23806), .DIN2 (____0___23805), .Q
       (____0___23807));
  and2s1 _______445724(.DIN1 (outData[0]), .DIN2 (outData[1]), .Q
       (____0___23804));
  nnd2s1 _______445725(.DIN1 (________22755), .DIN2 (____9___23797), .Q
       (____0___23803));
  and2s1 _______445726(.DIN1 (___9____23388), .DIN2 (__9__0__26854), .Q
       (_____0__24666));
  or2s1 _____0_445727(.DIN1 (________23278), .DIN2 (____00__23802), .Q
       (___0_____27968));
  nnd2s1 ____0__445728(.DIN1 (____99__23801), .DIN2 (____9___23800), .Q
       (____0___24159));
  nnd2s1 ____0__445729(.DIN1 (___90___23349), .DIN2 (__9_____26496), .Q
       (____0___24157));
  nnd2s1 ____0__445730(.DIN1 (____9___23799), .DIN2 (________25672), .Q
       (________24124));
  nnd2s1 ____0__445731(.DIN1 (____9___23798), .DIN2 (_____9__22336), .Q
       (________24030));
  and2s1 ____0_445732(.DIN1 (________23900), .DIN2 (________19236), .Q
       (___0____25301));
  nor2s1 ____0__445733(.DIN1 (___9_0__25184), .DIN2 (___90___23351), .Q
       (________24031));
  and2s1 _____445734(.DIN1 (____9___23797), .DIN2 (________22378), .Q
       (________24220));
  nor2s1 _______445735(.DIN1 (____0___19400), .DIN2 (___9____23368), .Q
       (______9__28320));
  and2s1 _______445736(.DIN1 (____9___23796), .DIN2 (___0_____27897),
       .Q (________24169));
  nnd2s1 _______445737(.DIN1 (____99__23801), .DIN2 (____9___23795), .Q
       (________24126));
  nnd2s1 _____9_445738(.DIN1 (________22925), .DIN2 (________23146), .Q
       (___0_____27529));
  nnd2s1 _____9_445739(.DIN1 (___9_0__23405), .DIN2 (____9___23794), .Q
       (___9____24265));
  nnd2s1 _____9_445740(.DIN1 (________23283), .DIN2 (_________28294),
       .Q (________23993));
  nnd2s1 _______445741(.DIN1 (____9___23793), .DIN2 (____90__23792), .Q
       (________25033));
  xor2s1 ____0__445742(.DIN1 (_____9__23791), .DIN2 (____0____32807),
       .Q (________24165));
  hi1s1 ____09_445743(.DIN (_________32122), .Q (___9____24302));
  nor2s1 ______445744(.DIN1 (_________34976), .DIN2 (________24528), .Q
       (________23790));
  nnd2s1 _____445745(.DIN1 (___9____23383), .DIN2 (________23007), .Q
       (________23789));
  and2s1 _______445746(.DIN1 (________23771), .DIN2 (____09__23627), .Q
       (________23787));
  hi1s1 ______445747(.DIN (_____0__23785), .Q (________23786));
  hi1s1 _______445748(.DIN (________23783), .Q (_____9__23784));
  hi1s1 _______445749(.DIN (________23781), .Q (________23782));
  nnd2s1 ______445750(.DIN1 (________23763), .DIN2 (____0___19400), .Q
       (________23780));
  or2s1 _______445751(.DIN1 (____9___23973), .DIN2 (____0___24160), .Q
       (________23779));
  or2s1 _______445752(.DIN1 (___9____24300), .DIN2 (outData[0]), .Q
       (________23778));
  nnd2s1 _______445753(.DIN1 (________23289), .DIN2 (____0___19400), .Q
       (________23777));
  nor2s1 ______445754(.DIN1 (________22695), .DIN2 (_____0__23775), .Q
       (________23776));
  nnd2s1 _______445755(.DIN1 (___9____23406), .DIN2 (________23773), .Q
       (_____9__23774));
  nnd2s1 _______445756(.DIN1 (________23771), .DIN2 (________23770), .Q
       (________23772));
  nnd2s1 ______445757(.DIN1 (________23298), .DIN2 (________23154), .Q
       (________23769));
  nor2s1 _____445758(.DIN1 (________23767), .DIN2 (_____9__23214), .Q
       (________23768));
  nor2s1 _____9_445759(.DIN1 (_____0__23765), .DIN2 (________23237), .Q
       (________23766));
  nor2s1 _____9_445760(.DIN1 (________23126), .DIN2 (________23763), .Q
       (_____9__23764));
  nnd2s1 _____9_445761(.DIN1 (________23186), .DIN2 (________23308), .Q
       (________23762));
  nnd2s1 _____9_445762(.DIN1 (________23760), .DIN2 (________23759), .Q
       (________23761));
  nor2s1 _____445763(.DIN1 (________23757), .DIN2 (________23280), .Q
       (________23758));
  and2s1 _____0_445764(.DIN1 (_____9__23755), .DIN2 (________22024), .Q
       (_____0__23756));
  or2s1 _____0_445765(.DIN1 (________24118), .DIN2 (________23753), .Q
       (________23754));
  and2s1 _______445766(.DIN1 (____9___23256), .DIN2 (________24001), .Q
       (________23751));
  or2s1 ______445767(.DIN1 (________23749), .DIN2 (_____0___34934), .Q
       (________23750));
  nnd2s1 ______445768(.DIN1 (_____0__23747), .DIN2 (________22225), .Q
       (________23748));
  nor2s1 _______445769(.DIN1 (___9_9__23422), .DIN2 (________23127), .Q
       (_____9__23746));
  nor2s1 _______445770(.DIN1 (_____0__23303), .DIN2 (________23183), .Q
       (________23745));
  nnd2s1 _______445771(.DIN1 (_____0__23181), .DIN2
       (______________________________________0__________0), .Q
       (________23744));
  nor2s1 ______445772(.DIN1 (________23742), .DIN2 (________23200), .Q
       (________23743));
  and2s1 _______445773(.DIN1 (________23740), .DIN2 (___990__23427), .Q
       (________23741));
  and2s1 _______445774(.DIN1 (____9___23251), .DIN2 (________23738), .Q
       (________23739));
  nnd2s1 ______445775(.DIN1 (____09__22904), .DIN2 (_____9__23736), .Q
       (_____0__23737));
  nnd2s1 ______445776(.DIN1 (________23155), .DIN2 (___0____22569), .Q
       (________23735));
  nnd2s1 _______445777(.DIN1 (____9___23343), .DIN2 (________23733), .Q
       (________23734));
  or2s1 _______445778(.DIN1 (________23731), .DIN2 (_________34944), .Q
       (________23732));
  or2s1 _______445779(.DIN1 (________23729), .DIN2 (_________34942), .Q
       (________23730));
  nnd2s1 ______445780(.DIN1 (________23771), .DIN2 (________21886), .Q
       (_____0__23728));
  nor2s1 _______445781(.DIN1 (________23153), .DIN2 (_____0__23286), .Q
       (_____9__23727));
  nnd2s1 ______445782(.DIN1 (________23135), .DIN2 (____00__23171), .Q
       (________23726));
  nor2s1 _______445783(.DIN1 (___00___22540), .DIN2 (________23118), .Q
       (________23725));
  nnd2s1 _______445784(.DIN1 (__9_____26722), .DIN2 (________23188), .Q
       (________23724));
  nor2s1 ______445785(.DIN1 (____0___22900), .DIN2 (________23117), .Q
       (________23723));
  or2s1 _______445786(.DIN1 (________25064), .DIN2 (________23271), .Q
       (________23722));
  nor2s1 _______445787(.DIN1 (________20289), .DIN2 (_________31241),
       .Q (________23721));
  nor2s1 _______445788(.DIN1 (____9___19945), .DIN2 (________23196), .Q
       (_____0__23720));
  nor2s1 _______445789(.DIN1 (____9___23168), .DIN2 (________23122), .Q
       (____0___23719));
  or2s1 _______445790(.DIN1 (________23309), .DIN2 (_________32604), .Q
       (____0___23718));
  nor2s1 _____9_445791(.DIN1 (____0___23716), .DIN2 (_____9__23133), .Q
       (____0___23717));
  nnd2s1 _____9_445792(.DIN1 (_____9__23124), .DIN2 (________22880), .Q
       (____0___23715));
  nor2s1 _____445793(.DIN1 (outData[0]), .DIN2 (____9___22073), .Q
       (____0___23714));
  nnd2s1 _____0_445794(.DIN1 (________23578), .DIN2 (____9___23165), .Q
       (____0___23713));
  nnd2s1 _____0_445795(.DIN1 (____0___23265), .DIN2 (________23757), .Q
       (____0___23712));
  nor2s1 ___90__445796(.DIN1 (________23217), .DIN2 (____9___23709), .Q
       (____9___23710));
  and2s1 ____9_445797(.DIN1 (_________34940), .DIN2 (____9___23707), .Q
       (____9___23708));
  hi1s1 ____9__445798(.DIN (___09_9__28080), .Q (____9___23706));
  or2s1 ______445799(.DIN1 (____90__23704), .DIN2 (_____9__23703), .Q
       (____9___23705));
  nnd2s1 _______445800(.DIN1 (outData[0]), .DIN2 (___9____24300), .Q
       (________24488));
  and2s1 _______445801(.DIN1 (____0___23806), .DIN2 (________23138), .Q
       (_____9__24625));
  nnd2s1 _______445802(.DIN1 (________23702), .DIN2 (________23129), .Q
       (___9____24293));
  and2s1 ______445803(.DIN1 (_____0__23125), .DIN2 (________23701), .Q
       (________25476));
  nnd2s1 _______445804(.DIN1 (_____0__22635), .DIN2 (_____0__23190), .Q
       (___9____25246));
  or2s1 _______445805(.DIN1 (________23700), .DIN2 (________23699), .Q
       (________24142));
  nnd2s1 _______445806(.DIN1 (________23319), .DIN2 (________19570), .Q
       (________23952));
  nor2s1 ______445807(.DIN1 (____9___22169), .DIN2 (________23141), .Q
       (__9__0__26816));
  nnd2s1 _______445808(.DIN1 (_____9__23285), .DIN2 (________22219), .Q
       (_____9__24139));
  nnd2s1 _______445809(.DIN1 (________23697), .DIN2 (________26084), .Q
       (________24477));
  nor2s1 _______445810(.DIN1 (_____18909), .DIN2 (_____9__23694), .Q
       (________23903));
  hi1s1 _____0_445811(.DIN (_______________18884), .Q (________23905));
  hi1s1 ____9__445812(.DIN (________23696), .Q (________24146));
  nor2s1 _______445813(.DIN1 (________22829), .DIN2 (________23220), .Q
       (__9_9___26987));
  nnd2s1 _____0_445814(.DIN1 (________23322), .DIN2 (________22927), .Q
       (___9____25237));
  nor2s1 _______445815(.DIN1 (inData[23]), .DIN2 (_____9__23694), .Q
       (________23904));
  nor2s1 _______445816(.DIN1 (_________28667), .DIN2 (_____0__23208),
       .Q (____0____28221));
  nor2s1 _______445817(.DIN1 (_____9__22797), .DIN2 (_________32604),
       .Q (_________31261));
  nnd2s1 _______445818(.DIN1 (________23228), .DIN2 (________21232), .Q
       (___09____28113));
  nnd2s1 _______445819(.DIN1 (________23693), .DIN2 (________23692), .Q
       (___9____24287));
  nor2s1 _______445820(.DIN1 (___0_____27696), .DIN2 (________23313),
       .Q (__9_____26389));
  nnd2s1 _____9_445821(.DIN1 (_____9__23293), .DIN2 (___0____22552), .Q
       (_________29386));
  nnd2s1 _______445822(.DIN1 (_____9__23694), .DIN2 (________23691), .Q
       (___0____24364));
  nor2s1 _______445823(.DIN1 (outData[1]), .DIN2 (outData[0]), .Q
       (________24546));
  hi1s1 _______445824(.DIN (_______________18884), .Q (_____0___35109));
  nnd2s1 _______445825(.DIN1 (____0___23263), .DIN2 (________22312), .Q
       (______0__32006));
  ib1s1 _____0_445826(.DIN (_______________18884), .Q (_________31290));
  nnd2s1 _______445827(.DIN1 (________23689), .DIN2 (inData[23]), .Q
       (___9____24269));
  nor2s1 _______445828(.DIN1 (________23690), .DIN2 (________23689), .Q
       (________24931));
  or2s1 _______445829(.DIN1 (___0____23510), .DIN2 (________24483), .Q
       (________23688));
  and2s1 _______445830(.DIN1 (___09___23523), .DIN2 (________23686), .Q
       (________23687));
  nor2s1 _______445831(.DIN1 (________23315), .DIN2 (________23548), .Q
       (_____0__23685));
  and2s1 ______445832(.DIN1 (________23683), .DIN2 (________23682), .Q
       (_____9__23684));
  nor2s1 ______445833(.DIN1 (inData[23]), .DIN2 (________23679), .Q
       (________23681));
  nor2s1 _______445834(.DIN1 (inData[25]), .DIN2 (________23679), .Q
       (________23680));
  nnd2s1 _______445835(.DIN1 (________23676), .DIN2 (inData[15]), .Q
       (________23678));
  nnd2s1 _______445836(.DIN1 (________23676), .DIN2 (inData[12]), .Q
       (________23677));
  nnd2s1 _______445837(.DIN1 (________23676), .DIN2 (inData[13]), .Q
       (_____0__23675));
  nnd2s1 _______445838(.DIN1 (________23676), .DIN2 (inData[10]), .Q
       (_____9__23674));
  nor2s1 ______445839(.DIN1 (_______19051), .DIN2 (________23667), .Q
       (________23673));
  nnd2s1 _______445840(.DIN1 (________22916), .DIN2 (inData[24]), .Q
       (________23672));
  or2s1 _______445841(.DIN1 (________22221), .DIN2 (________23670), .Q
       (________23671));
  nor2s1 _______445842(.DIN1 (________25793), .DIN2 (________23046), .Q
       (________23669));
  nor2s1 ______445843(.DIN1 (____9___23078), .DIN2 (________23667), .Q
       (________23668));
  and2s1 _______445844(.DIN1 (____9_0__33597), .DIN2 (_____9__23665),
       .Q (_____0__23666));
  nnd2s1 _______445845(.DIN1 (________23683), .DIN2 (inData[9]), .Q
       (________23664));
  nor2s1 _______445846(.DIN1 (_____18910), .DIN2 (________23662), .Q
       (________23663));
  nnd2s1 _______445847(.DIN1 (________23683), .DIN2 (inData[6]), .Q
       (________23661));
  and2s1 _______445848(.DIN1 (________23006), .DIN2 (________19520), .Q
       (________23660));
  nor2s1 _______445849(.DIN1 (_________34432), .DIN2 (________23662),
       .Q (________23659));
  nnd2s1 ______445850(.DIN1 (________23683), .DIN2 (inData[5]), .Q
       (________23658));
  and2s1 _______445851(.DIN1 (________23051), .DIN2 (________21380), .Q
       (________23657));
  nor2s1 _______445852(.DIN1 (____0___22084), .DIN2 (________23001), .Q
       (_____0__23656));
  nnd2s1 _______445853(.DIN1 (________23654), .DIN2 (________22661), .Q
       (_____9__23655));
  and2s1 _______445854(.DIN1 (________23652), .DIN2 (________23010), .Q
       (________23653));
  nnd2s1 _______445855(.DIN1 (____0___22996), .DIN2 (________25803), .Q
       (________23651));
  nnd2s1 _______445856(.DIN1 (________23683), .DIN2 (inData[7]), .Q
       (________23650));
  nnd2s1 ______445857(.DIN1 (________23060), .DIN2 (________24221), .Q
       (________23649));
  and2s1 _______445858(.DIN1 (________23020), .DIN2 (________24230), .Q
       (________23648));
  nor2s1 _______445859(.DIN1 (____9___19395), .DIN2 (________23316), .Q
       (________23647));
  or2s1 _______445860(.DIN1 (____0___23716), .DIN2 (________23044), .Q
       (_____9__23646));
  or2s1 _______445861(.DIN1 (________23644), .DIN2 (________24904), .Q
       (________23645));
  or2s1 _______445862(.DIN1 (________23642), .DIN2 (________23053), .Q
       (________23643));
  nor2s1 _______445863(.DIN1 (_____9__22042), .DIN2 (________23068), .Q
       (________23641));
  nnd2s1 _______445864(.DIN1 (_____0__22999), .DIN2 (_____0__23028), .Q
       (________23640));
  and2s1 _____9_445865(.DIN1 (____9_0__33597), .DIN2 (___0____19791),
       .Q (________23639));
  or2s1 _____9_445866(.DIN1 (________23045), .DIN2 (_____9__23637), .Q
       (_____0__23638));
  nor2s1 _____0_445867(.DIN1 (________23036), .DIN2 (________23635), .Q
       (________23636));
  nor2s1 _____0_445868(.DIN1 (_____9__25001), .DIN2 (____9___24695), .Q
       (________23634));
  and2s1 _____0_445869(.DIN1 (_________34954), .DIN2 (________24632),
       .Q (________23633));
  nnd2s1 _____0_445870(.DIN1 (___0_0__23455), .DIN2 (________23059), .Q
       (________23632));
  or2s1 _____0_445871(.DIN1 (____0___23089), .DIN2 (________23583), .Q
       (________23631));
  and2s1 _____0_445872(.DIN1 (_____0__23536), .DIN2 (_____0__23628), .Q
       (________23630));
  nnd2s1 _______445873(.DIN1 (_____0__23628), .DIN2 (____09__23627), .Q
       (________23629));
  nor2s1 _______445874(.DIN1 (________22913), .DIN2 (________23067), .Q
       (____0___23626));
  nnd2s1 _______445875(.DIN1 (___0____24386), .DIN2 (________23580), .Q
       (____0___23625));
  nor2s1 _______445876(.DIN1 (________22937), .DIN2 (____0___22899), .Q
       (____0___23624));
  nor2s1 _______445877(.DIN1 (________22381), .DIN2 (____0___23622), .Q
       (____0___23623));
  nnd2s1 _______445878(.DIN1 (_________34950), .DIN2 (____0___23620),
       .Q (____0___23621));
  nor2s1 _______445879(.DIN1 (____9___23081), .DIN2 (________22823), .Q
       (____0___23619));
  nnd2s1 ______445880(.DIN1 (_____9__22961), .DIN2 (________23016), .Q
       (____00__23618));
  nor2s1 ______445881(.DIN1 (_____09__34430), .DIN2 (_________33180),
       .Q (____99__23617));
  and2s1 _______445882(.DIN1 (_____0__22934), .DIN2 (____9___23615), .Q
       (____9___23616));
  nor2s1 _______445883(.DIN1 (________22293), .DIN2 (________23607), .Q
       (____9___23614));
  or2s1 _______445884(.DIN1 (________23541), .DIN2 (________23604), .Q
       (____9___23613));
  nor2s1 _______445885(.DIN1 (____9___22984), .DIN2 (____0___23622), .Q
       (____9___23612));
  nnd2s1 ______445886(.DIN1 (________23012), .DIN2 (________23757), .Q
       (____9___23611));
  nnd2s1 _______445887(.DIN1 (____9____32719), .DIN2 (_________34437),
       .Q (____9___23610));
  or2s1 _______445888(.DIN1 (_____9__23608), .DIN2 (________23607), .Q
       (____90__23609));
  nnd2s1 ______445889(.DIN1 (________22919), .DIN2 (inData[30]), .Q
       (________23606));
  nor2s1 ______445890(.DIN1 (_____0___35036), .DIN2 (________23604), .Q
       (________23605));
  nnd2s1 _______445891(.DIN1 (_________33177), .DIN2
       (_________________18777), .Q (________23603));
  nnd2s1 _______445892(.DIN1 (________23019), .DIN2 (_____0__23601), .Q
       (________23602));
  nor2s1 _______445893(.DIN1 (________23041), .DIN2 (__990___27088), .Q
       (_____9__23600));
  or2s1 _______445894(.DIN1 (___0____22565), .DIN2 (_____9__23037), .Q
       (________23599));
  nor2s1 _______445895(.DIN1 (________22093), .DIN2 (________22930), .Q
       (________23598));
  or2s1 _______445896(.DIN1 (________22975), .DIN2 (________23596), .Q
       (________23597));
  and2s1 _____0_445897(.DIN1 (____9_0__33597), .DIN2 (___0____19778),
       .Q (________23595));
  or2s1 _______445898(.DIN1 (________23593), .DIN2 (________23670), .Q
       (________23594));
  or2s1 _____0_445899(.DIN1 (_____0__23591), .DIN2 (____0___22896), .Q
       (________23592));
  nor2s1 _____0_445900(.DIN1 (________23589), .DIN2 (___99___24329), .Q
       (_____9__23590));
  nor2s1 _____445901(.DIN1 (________23587), .DIN2 (___0____23495), .Q
       (________23588));
  nnd2s1 _____9_445902(.DIN1 (____00__22895), .DIN2 (____9___19395), .Q
       (________23586));
  nnd2s1 _______445903(.DIN1 (________23862), .DIN2 (________23093), .Q
       (________23585));
  or2s1 _______445904(.DIN1 (________22970), .DIN2 (________23583), .Q
       (________23584));
  nnd2s1 _______445905(.DIN1 (_________32158), .DIN2 (___09___22619),
       .Q (_____0__23582));
  nor2s1 _______445906(.DIN1 (____9___19395), .DIN2 (________23580), .Q
       (_____9__23581));
  nnd2s1 _______445907(.DIN1 (________23578), .DIN2 (_________34952),
       .Q (________23579));
  nnd2s1 _______445908(.DIN1 (________23061), .DIN2 (___0_9__21675), .Q
       (________23577));
  nnd2s1 _______445909(.DIN1 (________23862), .DIN2 (________22973), .Q
       (________23576));
  nnd2s1 _______445910(.DIN1 (________23740), .DIN2 (_____0__24560), .Q
       (________23575));
  nor2s1 ______445911(.DIN1 (________19521), .DIN2 (________23667), .Q
       (________23574));
  nor2s1 ______445912(.DIN1 (________24221), .DIN2 (________23537), .Q
       (________23573));
  nor2s1 _______445913(.DIN1 (____09__22634), .DIN2 (_____0__23223), .Q
       (_____0__23572));
  nor2s1 _______445914(.DIN1 (________22325), .DIN2 (_____9__22923), .Q
       (_____9__23571));
  or2s1 _______445915(.DIN1 (____0___23716), .DIN2 (___09___23524), .Q
       (________23570));
  nnd2s1 _______445916(.DIN1 (_________33177), .DIN2 (_______18995), .Q
       (________23569));
  nor2s1 _______445917(.DIN1 (____0___22633), .DIN2 (________23683), .Q
       (________23568));
  hi1s1 _______445918(.DIN (________23566), .Q (________23567));
  hi1s1 _______445919(.DIN (________23564), .Q (________23565));
  nor2s1 _______445920(.DIN1 (________23562), .DIN2 (________23032), .Q
       (_____9__23563));
  nor2s1 _______445921(.DIN1 (________23209), .DIN2 (________24486), .Q
       (________23561));
  nor2s1 _______445922(.DIN1 (________20102), .DIN2 (________23667), .Q
       (________23560));
  nor2s1 _______445923(.DIN1 (____0___22990), .DIN2 (____9___22985), .Q
       (________23559));
  nnd2s1 _______445924(.DIN1 (________23029), .DIN2 (____9___19395), .Q
       (________23558));
  nor2s1 ______445925(.DIN1 (________23556), .DIN2 (____9___22983), .Q
       (________23557));
  or2s1 _______445926(.DIN1 (___00___21635), .DIN2 (_____9__23554), .Q
       (_____0__23555));
  nor2s1 _______445927(.DIN1 (________23552), .DIN2 (________22877), .Q
       (________23553));
  nor2s1 _______445928(.DIN1 (________22282), .DIN2 (___9_9__25202), .Q
       (________23551));
  nnd2s1 _______445929(.DIN1 (________23042), .DIN2 (_____0__23601), .Q
       (________23550));
  nor2s1 _______445930(.DIN1 (___9____23411), .DIN2 (________23548), .Q
       (________23549));
  or2s1 _____9_445931(.DIN1 (____0___22359), .DIN2 (________23767), .Q
       (________23547));
  nor2s1 _____9_445932(.DIN1 (_____0__23065), .DIN2 (________23227), .Q
       (________23546));
  nnd2s1 _____9_445933(.DIN1 (________23023), .DIN2 (_____9__23544), .Q
       (_____0__23545));
  nor2s1 _____0_445934(.DIN1 (________22343), .DIN2 (________22932), .Q
       (________23543));
  or2s1 _____0_445935(.DIN1 (________23541), .DIN2 (________23011), .Q
       (________23542));
  nor2s1 _____0_445936(.DIN1 (____0___23086), .DIN2 (________23202), .Q
       (________23540));
  nnd2s1 _______445937(.DIN1 (________23537), .DIN2 (_____0__23536), .Q
       (________23538));
  nor2s1 _______445938(.DIN1 (____0___23716), .DIN2 (________22850), .Q
       (____09__23535));
  nnd2s1 _______445939(.DIN1 (________22939), .DIN2 (____0___23716), .Q
       (____0___23534));
  nnd2s1 _______445940(.DIN1 (___999__26246), .DIN2 (________22944), .Q
       (____0___23533));
  nor2s1 ______445941(.DIN1 (______18932), .DIN2 (________22921), .Q
       (____0___23532));
  nor2s1 _______445942(.DIN1 (_____9__22854), .DIN2 (_________34962),
       .Q (____0___23531));
  and2s1 _______445943(.DIN1 (____0____31820), .DIN2 (_________30807),
       .Q (____0___23530));
  nnd2s1 _______445944(.DIN1 (_____0__23018), .DIN2 (_________35046),
       .Q (________23988));
  nnd2s1 _____9_445945(.DIN1 (________23048), .DIN2 (____0___23529), .Q
       (___0__9__27819));
  or2s1 _____9_445946(.DIN1 (____00__23528), .DIN2 (___099__23527), .Q
       (____09__24071));
  nnd2s1 _____445947(.DIN1 (____9___23079), .DIN2 (___09___23526), .Q
       (________24662));
  nnd2s1 _____0_445948(.DIN1 (___09___23525), .DIN2 (_____9__23017), .Q
       (________23845));
  nnd2s1 _____0_445949(.DIN1 (___09___23524), .DIN2 (________22781), .Q
       (_____0__23999));
  nnd2s1 _____0_445950(.DIN1 (________22977), .DIN2 (______0__28974),
       .Q (________23844));
  nnd2s1 _____0_445951(.DIN1 (___09___23523), .DIN2 (__9_____26555), .Q
       (________24002));
  nor2s1 _____445952(.DIN1 (___9____24260), .DIN2 (____0___22897), .Q
       (________23788));
  nnd2s1 _______445953(.DIN1 (________22868), .DIN2 (___09___23522), .Q
       (________23842));
  nor2s1 _______445954(.DIN1 (____0___23087), .DIN2 (___09___23521), .Q
       (__99____27100));
  nnd2s1 _______445955(.DIN1 (________23013), .DIN2 (___900__26147), .Q
       (_____9__23843));
  nor2s1 _______445956(.DIN1 (___09___23520), .DIN2 (________22978), .Q
       (_____0__24809));
  and2s1 _______445957(.DIN1 (___09___23519), .DIN2 (___0____25333), .Q
       (________24090));
  nnd2s1 _______445958(.DIN1 (_____9__23230), .DIN2 (________23679), .Q
       (________25687));
  xnr2s1 ____0__445959(.DIN1 (__9__0__26618), .DIN2 (____000__32751),
       .Q (_____0__24044));
  and2s1 ______445960(.DIN1 (_____0__25665), .DIN2 (___09___23519), .Q
       (________25717));
  nor2s1 _______445961(.DIN1 (____9___21808), .DIN2 (_____0__23038), .Q
       (____0____31863));
  dffacs2 __________________445962(.CLRB (reset), .CLK (clk), .DIN
       (________23054), .Q (_______________18884));
  nnd2s1 ______445963(.DIN1 (________23002), .DIN2 (________22249), .Q
       (_________32122));
  nnd2s1 _______445964(.DIN1 (________23049), .DIN2 (_____9__22679), .Q
       (_________31667));
  and2s1 _____0_445965(.DIN1 (________22881), .DIN2 (________24660), .Q
       (___090__23518));
  nnd2s1 _____0_445966(.DIN1 (___0____23506), .DIN2 (_____0__22905), .Q
       (___0_9__23517));
  nor2s1 ______445967(.DIN1 (_____0__24173), .DIN2 (_____9__23008), .Q
       (___0____23516));
  nnd2s1 _______445968(.DIN1 (________22908), .DIN2 (____09__22634), .Q
       (___0____23515));
  or2s1 _______445969(.DIN1 (________23562), .DIN2 (________23094), .Q
       (___0____23514));
  or2s1 _____9_445970(.DIN1 (___0____23512), .DIN2 (____9___22988), .Q
       (___0____23513));
  or2s1 _______445971(.DIN1 (___0____23510), .DIN2 (___9_9__25202), .Q
       (___0____23511));
  nor2s1 _______445972(.DIN1 (_______18954), .DIN2 (_________33180), .Q
       (___0_0__23509));
  nnd2s1 ___9___445973(.DIN1 (___0____23506), .DIN2 (________22388), .Q
       (___0____23507));
  and2s1 ___9___445974(.DIN1 (___0____23506), .DIN2 (__90____26258), .Q
       (___0____23505));
  nnd2s1 ___9___445975(.DIN1 (________22860), .DIN2 (____9___19945), .Q
       (___0____23504));
  nor2s1 ___9___445976(.DIN1 (___0____23502), .DIN2 (___0____23450), .Q
       (___0____23503));
  nor2s1 ___9___445977(.DIN1 (___0_0__23500), .DIN2 (___000__23437), .Q
       (___0____23501));
  nor2s1 ___9___445978(.DIN1 (___0____23498), .DIN2 (___0____23497), .Q
       (___0_9__23499));
  nor2s1 ___9__445979(.DIN1 (___0_0__22608), .DIN2 (___0____23495), .Q
       (___0____23496));
  nor2s1 ___9__445980(.DIN1 (________21760), .DIN2 (____0___22810), .Q
       (___0____23494));
  and2s1 ___9___445981(.DIN1 (___0____23482), .DIN2 (____0___24798), .Q
       (___0____23493));
  nor2s1 ___9___445982(.DIN1 (___9____22469), .DIN2 (_____0__22848), .Q
       (___0____23492));
  and2s1 ___9_445983(.DIN1 (___0____23453), .DIN2 (___0_0__23490), .Q
       (___0____23491));
  nnd2s1 ___9_0_445984(.DIN1 (___0____23506), .DIN2 (___0____23488), .Q
       (___0_9__23489));
  nor2s1 ___9_0_445985(.DIN1 (________22329), .DIN2 (____0___22810), .Q
       (___0____23487));
  nnd2s1 ___445986(.DIN1 (___0____23506), .DIN2 (_____9__25145), .Q
       (___0____23486));
  nor2s1 ___909_445987(.DIN1 (___0____23484), .DIN2 (___0____23495), .Q
       (___0____23485));
  nnd2s1 ___909_445988(.DIN1 (___0____23482), .DIN2 (___0_0__23481), .Q
       (___0____23483));
  nor2s1 ___90_445989(.DIN1 (___9_0__23413), .DIN2 (________22839), .Q
       (___0____23479));
  nnd2s1 ___90__445990(.DIN1 (___0____23477), .DIN2 (_______18992), .Q
       (___0____23478));
  hi1s1 _______445991(.DIN (_____9__23694), .Q (___0____23476));
  or2s1 ___90__445992(.DIN1 (___0____22578), .DIN2 (___0____23495), .Q
       (___0____23475));
  nor2s1 _______445993(.DIN1 (_____9__22070), .DIN2 (___0____23495), .Q
       (___0____23474));
  nor2s1 _______445994(.DIN1 (_____9__22825), .DIN2 (________22738), .Q
       (___0_0__23473));
  nor2s1 _______445995(.DIN1 (___0____23471), .DIN2 (________22846), .Q
       (___0_9__23472));
  nnd2s1 _______445996(.DIN1 (______0__33058), .DIN2 (______18919), .Q
       (___0____23470));
  nnd2s1 _______445997(.DIN1 (________23114), .DIN2 (________23274), .Q
       (___0____23468));
  nnd2s1 _______445998(.DIN1 (___0____23506), .DIN2 (________23305), .Q
       (___0____23467));
  nnd2s1 _______445999(.DIN1 (________23031), .DIN2 (___0____23465), .Q
       (___0____23466));
  nor2s1 ______446000(.DIN1 (________22640), .DIN2 (___0_9__23463), .Q
       (___0_0__23464));
  nnd2s1 ___90__446001(.DIN1 (_____0__24140), .DIN2 (___0____22577), .Q
       (___0____23462));
  nor2s1 _____0_446002(.DIN1 (________23182), .DIN2 (________23113), .Q
       (___0____23461));
  nnd2s1 _____0_446003(.DIN1 (___0_____27410), .DIN2 (_____0__24120),
       .Q (___0____23460));
  nnd2s1 _______446004(.DIN1 (_____0__24120), .DIN2 (________22773), .Q
       (___0____23459));
  and2s1 _______446005(.DIN1 (___0____23506), .DIN2 (___990), .Q
       (___0____23458));
  and2s1 _______446006(.DIN1 (________22844), .DIN2 (________24440), .Q
       (___0____23457));
  or2s1 _______446007(.DIN1 (___0_0__23455), .DIN2 (___00___23441), .Q
       (___0____23456));
  nnd2s1 _______446008(.DIN1 (___0____23453), .DIN2 (___0____23452), .Q
       (___0_9__23454));
  nor2s1 _______446009(.DIN1 (___9____22493), .DIN2 (___0____23450), .Q
       (___0____23451));
  nnd2s1 _______446010(.DIN1 (________25424), .DIN2 (___0____23448), .Q
       (___0____23449));
  nor2s1 _______446011(.DIN1 (___9_0__22465), .DIN2 (____0___22810), .Q
       (___0____23447));
  nor2s1 _______446012(.DIN1 (___9____24260), .DIN2 (_____0__22875), .Q
       (___0____23446));
  nor2s1 ___90__446013(.DIN1 (________22390), .DIN2 (_____9__22864), .Q
       (___00___23443));
  or2s1 ___9_0_446014(.DIN1 (___00___23438), .DIN2 (___00___23441), .Q
       (___00___23442));
  nor2s1 ___90_446015(.DIN1 (_____0__22855), .DIN2 (________22863), .Q
       (___00___23440));
  nor2s1 ___90__446016(.DIN1 (___00___23438), .DIN2 (___000__23437), .Q
       (___00___23439));
  nnd2s1 ___90__446017(.DIN1 (___0____23453), .DIN2 (___99___23435), .Q
       (___999__23436));
  or2s1 ___90__446018(.DIN1 (________23247), .DIN2 (___0____23497), .Q
       (___99___23434));
  and2s1 ___90__446019(.DIN1 (___0____23453), .DIN2 (___99___23432), .Q
       (___99___23433));
  nor2s1 ___90__446020(.DIN1 (___9____26159), .DIN2 (____0___22810), .Q
       (___99___23431));
  nor2s1 ___90__446021(.DIN1 (___99___23429), .DIN2 (___000__23437), .Q
       (___99___23430));
  hi1s1 ____9__446022(.DIN (___990__23427), .Q (___99___23428));
  and2s1 ___90__446023(.DIN1 (________22856), .DIN2 (________24651), .Q
       (___9____23425));
  nnd2s1 ____9__446024(.DIN1 (__9_____26447), .DIN2 (__9_____26875), .Q
       (___9____23424));
  nor2s1 ____9__446025(.DIN1 (________23057), .DIN2 (___000__23437), .Q
       (___9____23423));
  nor2s1 ____9__446026(.DIN1 (________24221), .DIN2 (_____9__22874), .Q
       (___9____23421));
  and2s1 ____9__446027(.DIN1 (____9___22803), .DIN2 (______0__34958),
       .Q (___9____23420));
  nor2s1 ____9__446028(.DIN1 (________22415), .DIN2 (___0____23450), .Q
       (___9____23419));
  nor2s1 ____9__446029(.DIN1 (___9____22475), .DIN2 (___0____23495), .Q
       (___9____23418));
  nor2s1 ___90_446030(.DIN1 (___9____23416), .DIN2 (___00___23441), .Q
       (___9____23417));
  nor2s1 ____9_446031(.DIN1 (__9_____26828), .DIN2 (___00___23441), .Q
       (___9____23415));
  nnd2s1 ___900_446032(.DIN1 (___0____23453), .DIN2 (___9_0__23413), .Q
       (___9____23414));
  or2s1 ___900_446033(.DIN1 (___9____23411), .DIN2 (___9____23410), .Q
       (___9_9__23412));
  and2s1 ___90_446034(.DIN1 (___0____23482), .DIN2 (________25524), .Q
       (___9____23409));
  nnd2s1 ___90_446035(.DIN1 (_____0__24140), .DIN2 (____0___21723), .Q
       (___9____23408));
  and2s1 _______446036(.DIN1 (____0___22902), .DIN2 (__9__0__26854), .Q
       (____9___24058));
  dffacs1 __________________446037(.CLRB (reset), .CLK (clk), .DIN
       (________23024), .QN (_______________18882));
  nor2s1 _______446038(.DIN1 (___9____23407), .DIN2 (________22974), .Q
       (_____0__23785));
  xnr2s1 ____0__446039(.DIN1 (_________33385), .DIN2 (______18945), .Q
       (_____9__23991));
  nnd2s1 _______446040(.DIN1 (________23314), .DIN2 (_________34994),
       .Q (_____0__24035));
  nnd2s1 ______446041(.DIN1 (_____0__24956), .DIN2 (_________34964), .Q
       (________24192));
  nnd2s1 _______446042(.DIN1 (____90__22981), .DIN2 (________19570), .Q
       (___0__0__27792));
  or2s1 ______446043(.DIN1 (____9___22439), .DIN2 (________25424), .Q
       (_____0__23950));
  nnd2s1 _______446044(.DIN1 (______0__34958), .DIN2 (________22275),
       .Q (________23912));
  nnd2s1 _______446045(.DIN1 (________22830), .DIN2 (________23773), .Q
       (________23956));
  nnd2s1 _______446046(.DIN1 (________22883), .DIN2 (____0___22903), .Q
       (___0_9___27557));
  hi1s1 _______446047(.DIN (________23689), .Q (________23902));
  hi1s1 _______446048(.DIN (___9____23406), .Q (________23961));
  hi1s1 _____0_446049(.DIN (___9_0__23405), .Q (____9___23970));
  nor2s1 ___9___446050(.DIN1 (____99__21074), .DIN2 (____0___22810), .Q
       (________23696));
  nor2s1 ___9_9_446051(.DIN1 (________23058), .DIN2 (___000__23437), .Q
       (___0_____27549));
  or2s1 ___9_9_446052(.DIN1 (__9_____26828), .DIN2 (___000__23437), .Q
       (________23913));
  nor2s1 ______446053(.DIN1 (________21883), .DIN2 (___9_9__23404), .Q
       (_____0__25625));
  nnd2s1 _______446054(.DIN1 (___9____23403), .DIN2 (___9____23402), .Q
       (____9___24054));
  nor2s1 _______446055(.DIN1 (___9____23401), .DIN2 (________22851), .Q
       (________24003));
  nor2s1 ______446056(.DIN1 (___0_____27291), .DIN2 (________22935), .Q
       (________23918));
  nor2s1 _______446057(.DIN1 (_____0__22216), .DIN2 (___9____23400), .Q
       (________23781));
  nor2s1 _______446058(.DIN1 (___9____23399), .DIN2 (________22928), .Q
       (_____0__24008));
  xor2s1 _______446059(.DIN1 (_______________18873), .DIN2
       (_____99__31353), .Q (________24022));
  and2s1 _______446060(.DIN1 (_____9__23047), .DIN2 (____9___26043), .Q
       (________24115));
  nnd2s1 _______446061(.DIN1 (___9____23398), .DIN2 (__9_____26862), .Q
       (________23998));
  nnd2s1 ______446062(.DIN1 (____9___23080), .DIN2 (___9____23397), .Q
       (________23783));
  nnd2s1 _______446063(.DIN1 (________23211), .DIN2 (___9____23396), .Q
       (____90__24053));
  nor2s1 ___9___446064(.DIN1 (____09__22088), .DIN2 (___000__23437), .Q
       (___0____25284));
  nor2s1 ___9__446065(.DIN1 (___9____26182), .DIN2 (________23583), .Q
       (________23909));
  or2s1 ___9___446066(.DIN1 (________23917), .DIN2 (___000__23437), .Q
       (________24122));
  or2s1 ___9___446067(.DIN1 (__9_____26548), .DIN2 (_________34960), .Q
       (________23948));
  nnd2s1 ___9___446068(.DIN1 (___0____23453), .DIN2 (___9_9__23395), .Q
       (________23946));
  or2s1 ___9___446069(.DIN1 (_________35054), .DIN2 (____0___22810), .Q
       (_____0__23915));
  nnd2s1 ___9___446070(.DIN1 (_____9__22832), .DIN2 (___9____23394), .Q
       (_____9__23941));
  nnd2s1 ___9__446071(.DIN1 (___0____23482), .DIN2 (________21087), .Q
       (________24474));
  or2s1 _______446072(.DIN1 (___0_0__23455), .DIN2 (___000__23437), .Q
       (___09____28105));
  or2s1 ___9___446073(.DIN1 (________23917), .DIN2 (___00___23441), .Q
       (____0____28179));
  or2s1 ___9___446074(.DIN1 (__9_____26597), .DIN2 (________22861), .Q
       (___9_0__25241));
  or2s1 ___9__446075(.DIN1 (___00____27182), .DIN2 (____0___22810), .Q
       (___0_____27873));
  or2s1 ___9__446076(.DIN1 (__9__0__26749), .DIN2 (__9_____26831), .Q
       (____0___23979));
  nnd2s1 ___9___446077(.DIN1 (________22842), .DIN2 (________23757), .Q
       (__9__9__26476));
  nor2s1 ______446078(.DIN1 (___9____21594), .DIN2 (___0____23495), .Q
       (________23916));
  nor2s1 _______446079(.DIN1 (________22769), .DIN2 (___0____23450), .Q
       (___0_9___27940));
  and2s1 _______446080(.DIN1 (______0__33058), .DIN2 (________23100),
       .Q (_____0___33034));
  nnd2s1 _______446081(.DIN1 (________22837), .DIN2 (___00___23438), .Q
       (________24083));
  hi1s1 _______446082(.DIN (_____0___32294), .Q (____0___23981));
  nnd2s1 _______446083(.DIN1 (_________32158), .DIN2 (___09___22620),
       .Q (________24111));
  nnd2s1 ______446084(.DIN1 (____9_0__33597), .DIN2 (___909__23355), .Q
       (____9____33613));
  nor2s1 ___9___446085(.DIN1 (____00__21719), .DIN2 (____0___22810), .Q
       (___09_9__28080));
  or2s1 ___9___446086(.DIN1 (__900_), .DIN2 (___0____23495), .Q
       (____0____28153));
  or2s1 ___9___446087(.DIN1 (___9____23416), .DIN2 (___000__23437), .Q
       (_________28478));
  or2s1 ___9___446088(.DIN1 (___0____21652), .DIN2 (____0___22810), .Q
       (________25049));
  nor2s1 ___9___446089(.DIN1 (________21107), .DIN2 (___00___23441), .Q
       (_________28461));
  or2s1 ____9__446090(.DIN1 (___9____23393), .DIN2 (_________34966), .Q
       (______0__32252));
  hi1s1 ____9__446091(.DIN (_________31241), .Q (_____9___30454));
  nor2s1 _______446092(.DIN1 (___9____23391), .DIN2 (_____0__22833), .Q
       (___9____23392));
  xor2s1 ____0__446093(.DIN1 (___0____22548), .DIN2 (___9____23389), .Q
       (___9____23390));
  nor2s1 _______446094(.DIN1 (___9____23387), .DIN2 (________25963), .Q
       (___9____23388));
  and2s1 _______446095(.DIN1 (______0__33918), .DIN2 (______18946), .Q
       (___9_0__23386));
  or2s1 _______446096(.DIN1 (inData[11]), .DIN2 (__9_____27027), .Q
       (___9_9__23385));
  nnd2s1 _______446097(.DIN1 (__9_____26675), .DIN2 (inData[22]), .Q
       (___9____23384));
  nor2s1 ______446098(.DIN1 (________22958), .DIN2 (________22656), .Q
       (___9____23383));
  or2s1 _____9_446099(.DIN1 (___00___22543), .DIN2 (___9____23381), .Q
       (___9____23382));
  and2s1 _____9_446100(.DIN1 (_____9__22771), .DIN2 (___9____23379), .Q
       (___9____23380));
  and2s1 _____9_446101(.DIN1 (______0__33336), .DIN2 (________22759),
       .Q (___9____23378));
  or2s1 _____9_446102(.DIN1 (____0___22811), .DIN2 (___9_0__23376), .Q
       (___9____23377));
  nnd2s1 _____0_446103(.DIN1 (________23862), .DIN2 (___0____22557), .Q
       (___9_9__23375));
  nnd2s1 ______446104(.DIN1 (_____9__22971), .DIN2 (___9____23373), .Q
       (___9____23374));
  or2s1 _______446105(.DIN1 (___9____23371), .DIN2 (_____0__22764), .Q
       (___9____23372));
  and2s1 _______446106(.DIN1 (__9_____26675), .DIN2 (_____09__31192),
       .Q (___9____23370));
  nor2s1 _______446107(.DIN1 (________19520), .DIN2 (________22778), .Q
       (___9____23369));
  nor2s1 ______446108(.DIN1 (________22767), .DIN2 (___9____23367), .Q
       (___9____23368));
  nnd2s1 _______446109(.DIN1 (__9_____26675), .DIN2 (inData[24]), .Q
       (___9_0__23366));
  nnd2s1 _______446110(.DIN1 (______0__33918), .DIN2 (___9____22509),
       .Q (___9_9__23365));
  nnd2s1 _______446111(.DIN1 (________22757), .DIN2 (____0_9__32819),
       .Q (___9____23364));
  nor2s1 _______446112(.DIN1 (___9____23362), .DIN2 (________22756), .Q
       (___9____23363));
  or2s1 _______446113(.DIN1 (inData[14]), .DIN2 (__9_____27027), .Q
       (___9____23361));
  nor2s1 ______446114(.DIN1 (_____0__22754), .DIN2 (________23749), .Q
       (___9____23360));
  or2s1 _______446115(.DIN1 (____9___24060), .DIN2 (________22867), .Q
       (___9____23359));
  nnd2s1 _______446116(.DIN1 (__9_____26675), .DIN2 (inData[27]), .Q
       (___9____23358));
  nnd2s1 _______446117(.DIN1 (______0__33336), .DIN2 (___0_0__19793),
       .Q (___9____23357));
  nor2s1 _____9_446118(.DIN1 (________19172), .DIN2 (___909__23355), .Q
       (___9_0__23356));
  or2s1 _______446119(.DIN1 (___90___23353), .DIN2 (___90___23352), .Q
       (___90___23354));
  nnd2s1 _______446120(.DIN1 (________22703), .DIN2 (___90___23350), .Q
       (___90___23351));
  nor2s1 _______446121(.DIN1 (___9____25200), .DIN2 (________25831), .Q
       (___90___23349));
  nor2s1 ______446122(.DIN1 (___90___23347), .DIN2 (________25881), .Q
       (___90___23348));
  nnd2s1 _______446123(.DIN1 (____99__23345), .DIN2 (________21975), .Q
       (___900__23346));
  nnd2s1 _______446124(.DIN1 (________25881), .DIN2 (____09__22634), .Q
       (____9___23344));
  nor2s1 ___446125(.DIN1 (_____9___35022), .DIN2 (____9___23342), .Q
       (____9___23343));
  xor2s1 _____0_446126(.DIN1 (_________9_), .DIN2 (_________32624), .Q
       (____9___23341));
  xor2s1 _______446127(.DIN1 (______0__34491), .DIN2
       (______________0______________________18826), .Q
       (____9___23340));
  xor2s1 _______446128(.DIN1 (_______19038), .DIN2 (_________33444), .Q
       (____9___23339));
  nnd2s1 _______446129(.DIN1 (_____9__23275), .DIN2 (________22785), .Q
       (____9___23338));
  nor2s1 _______446130(.DIN1 (________23144), .DIN2 (____9___25945), .Q
       (____9___23337));
  nnd2s1 _______446131(.DIN1 (________22972), .DIN2 (___00___23438), .Q
       (____90__23336));
  and2s1 ______446132(.DIN1 (________23229), .DIN2 (____99__23711), .Q
       (_____9__23335));
  nor2s1 _______446133(.DIN1 (________19520), .DIN2 (_____9__22708), .Q
       (________23334));
  nnd2s1 _____446134(.DIN1 (________23332), .DIN2 (________23871), .Q
       (________23333));
  and2s1 _____9_446135(.DIN1 (________23330), .DIN2 (________23757), .Q
       (________23331));
  nor2s1 _____9_446136(.DIN1 (_______19021), .DIN2 (__9_____26675), .Q
       (________23329));
  nnd2s1 _____9_446137(.DIN1 (________23327), .DIN2 (_____0__23326), .Q
       (________23328));
  nor2s1 _____0_446138(.DIN1 (____09__22634), .DIN2 (________22707), .Q
       (_____9__23325));
  xnr2s1 _______446139(.DIN1 (________19922), .DIN2 (____0_9__30961),
       .Q (________23324));
  xor2s1 _______446140(.DIN1 (_________34442), .DIN2 (_________32624),
       .Q (________23323));
  or2s1 _____446141(.DIN1 (________23321), .DIN2 (_____0__23241), .Q
       (________23322));
  and2s1 _____9_446142(.DIN1 (________22731), .DIN2 (___00___22540), .Q
       (________23320));
  or2s1 _____9_446143(.DIN1 (________23318), .DIN2 (_____0__22790), .Q
       (________23319));
  nor2s1 _____446144(.DIN1 (___9____22522), .DIN2 (________23279), .Q
       (_____0__23317));
  hi1s1 _____0_446145(.DIN (___09___23523), .Q (________23313));
  and2s1 _______446146(.DIN1 (________22747), .DIN2 (_____9__23311), .Q
       (_____0__23312));
  nnd2s1 _______446147(.DIN1 (________22660), .DIN2 (________22693), .Q
       (________23310));
  nor2s1 _______446148(.DIN1 (________20288), .DIN2 (____90__22798), .Q
       (________23309));
  or2s1 ______446149(.DIN1 (_____0__23199), .DIN2 (________23307), .Q
       (________23308));
  nnd2s1 _______446150(.DIN1 (________23578), .DIN2 (________23305), .Q
       (________23306));
  nor2s1 _______446151(.DIN1 (_____0__23303), .DIN2 (_____9__23302), .Q
       (________23304));
  and2s1 _______446152(.DIN1 (____9___25746), .DIN2 (___00___22540), .Q
       (________23301));
  nnd2s1 _______446153(.DIN1 (________24230), .DIN2 (_____9__21947), .Q
       (________23300));
  nor2s1 ______446154(.DIN1 (___9____22470), .DIN2 (____0___22808), .Q
       (________23299));
  nnd2s1 _______446155(.DIN1 (________23307), .DIN2 (___0_____27862),
       .Q (________23298));
  nor2s1 _______446156(.DIN1 (_____9__22743), .DIN2 (____0___22809), .Q
       (________23297));
  and2s1 _______446157(.DIN1 (____0___25754), .DIN2 (________23295), .Q
       (________23296));
  nor2s1 _______446158(.DIN1 (____9___25168), .DIN2 (____0___23266), .Q
       (_____0__23294));
  nor2s1 ______446159(.DIN1 (_____9__19917), .DIN2 (____0___23262), .Q
       (_____9__23293));
  nnd2s1 _______446160(.DIN1 (___09___22621), .DIN2 (inData[26]), .Q
       (________23291));
  nnd2s1 _______446161(.DIN1 (____09__22724), .DIN2 (inData[16]), .Q
       (________23290));
  or2s1 _____446162(.DIN1 (___0____22567), .DIN2 (________23288), .Q
       (________23289));
  nor2s1 _____9_446163(.DIN1 (________22100), .DIN2 (_____0__23286), .Q
       (________23287));
  nor2s1 _____446164(.DIN1 (________23284), .DIN2 (_____0__23152), .Q
       (_____9__23285));
  and2s1 _____0_446165(.DIN1 (________23277), .DIN2 (________23770), .Q
       (________23283));
  nnd2s1 ______446166(.DIN1 (____0___23178), .DIN2 (_____9__22290), .Q
       (________23282));
  nor2s1 _______446167(.DIN1 (____09__23267), .DIN2 (________23062), .Q
       (________23281));
  nor2s1 _______446168(.DIN1 (_____0__22670), .DIN2 (________23279), .Q
       (________23280));
  nor2s1 _______446169(.DIN1 (________24221), .DIN2 (________23277), .Q
       (________23278));
  nnd2s1 _______446170(.DIN1 (_____9__23275), .DIN2 (________22286), .Q
       (_____0__23276));
  nnd2s1 ______446171(.DIN1 (________23137), .DIN2 (____0___21815), .Q
       (________23272));
  nnd2s1 _______446172(.DIN1 (________23270), .DIN2 (___9____21557), .Q
       (________23271));
  nor2s1 _______446173(.DIN1 (________23757), .DIN2 (___90___25180), .Q
       (________23269));
  nor2s1 _______446174(.DIN1 (____09__23267), .DIN2 (____0___23266), .Q
       (_____0__23268));
  nnd2s1 _______446175(.DIN1 (___90___25180), .DIN2 (________23030), .Q
       (____0___23265));
  nnd2s1 _______446176(.DIN1 (___0____22580), .DIN2 (________22728), .Q
       (____0___23264));
  nor2s1 _______446177(.DIN1 (________19317), .DIN2 (____0___23262), .Q
       (____0___23263));
  and2s1 _______446178(.DIN1 (________23578), .DIN2 (________22740), .Q
       (____0___23261));
  or2s1 _______446179(.DIN1 (________23919), .DIN2 (___9____25198), .Q
       (____0___23260));
  nnd2s1 _______446180(.DIN1 (________23102), .DIN2 (_________34980),
       .Q (____00__23259));
  or2s1 _______446181(.DIN1 (____9___23257), .DIN2 (________22760), .Q
       (____99__23258));
  nor2s1 _______446182(.DIN1 (____9___23255), .DIN2 (____9___23254), .Q
       (____9___23256));
  nor2s1 _______446183(.DIN1 (__9_____26764), .DIN2 (____9___23252), .Q
       (____9___23253));
  and2s1 _______446184(.DIN1 (___9____22512), .DIN2 (____90__23250), .Q
       (____9___23251));
  or2s1 _______446185(.DIN1 (________23248), .DIN2 (________23247), .Q
       (________23249));
  nor2s1 ______446186(.DIN1 (_________18845), .DIN2 (____0_0__32780),
       .Q (________23246));
  nnd2s1 _______446187(.DIN1 (________23244), .DIN2 (________23243), .Q
       (________23245));
  nnd2s1 ______446188(.DIN1 (___90___23352), .DIN2 (___90___23353), .Q
       (________23242));
  nor2s1 _____0_446189(.DIN1 (inData[23]), .DIN2 (___00____27202), .Q
       (________23690));
  nor2s1 ______446190(.DIN1 (___90___23347), .DIN2 (_____0__22734), .Q
       (___0____23480));
  nor2s1 _______446191(.DIN1 (____0___24065), .DIN2 (_____0__22780), .Q
       (_____0__23747));
  nor2s1 ______446192(.DIN1 (________22186), .DIN2 (_____0__23241), .Q
       (____0___25370));
  or2s1 _______446193(.DIN1 (_____9__23240), .DIN2 (________23248), .Q
       (________23833));
  nor2s1 ___9_9_446194(.DIN1 (________23103), .DIN2 (____9___26142), .Q
       (___9____23426));
  nor2s1 _______446195(.DIN1 (____0___23716), .DIN2 (________22782), .Q
       (________24929));
  nor2s1 ______446196(.DIN1 (________23239), .DIN2 (________22762), .Q
       (____9___23793));
  nor2s1 ______446197(.DIN1 (________23238), .DIN2 (________24118), .Q
       (____9___23798));
  hi1s1 _____0_446198(.DIN (________23237), .Q (___00___24336));
  nnd2s1 _______446199(.DIN1 (________22702), .DIN2 (________23236), .Q
       (_____9__23703));
  hi1s1 _____446200(.DIN (________23235), .Q (________23753));
  hi1s1 _______446201(.DIN (________23683), .Q (________23693));
  nnd2s1 _______446202(.DIN1 (________23234), .DIN2 (_____0__22366), .Q
       (_____0__23860));
  or2s1 _______446203(.DIN1 (__9_____26472), .DIN2 (________22784), .Q
       (________24135));
  xnr2s1 _______446204(.DIN1 (_____9___32930), .DIN2 (________19084),
       .Q (________23566));
  nor2s1 ______446205(.DIN1 (_____0__22700), .DIN2 (________25963), .Q
       (____9___23796));
  nor2s1 _______446206(.DIN1 (________23233), .DIN2 (_________28775),
       .Q (____9___23799));
  nor2s1 _______446207(.DIN1 (__9090), .DIN2 (____9___22711), .Q
       (____9___24057));
  nor2s1 ______446208(.DIN1 (___0____22589), .DIN2 (________22791), .Q
       (________23812));
  nor2s1 _______446209(.DIN1 (__9_____26548), .DIN2 (____90__22709), .Q
       (________23564));
  nnd2s1 _______446210(.DIN1 (________22774), .DIN2 (__9__0__26854), .Q
       (_____0__24746));
  hi1s1 ______446211(.DIN (_________31060), .Q (______9__28560));
  and2s1 ______446212(.DIN1 (______0__33336), .DIN2 (________23232), .Q
       (_________33241));
  nnd2s1 _______446213(.DIN1 (________23234), .DIN2 (_____0__23231), .Q
       (___0_____27303));
  nor2s1 _______446214(.DIN1 (________24105), .DIN2 (____0___23090), .Q
       (________23866));
  nor2s1 _______446215(.DIN1 (________22122), .DIN2 (________26072), .Q
       (____99__23801));
  nnd2s1 _______446216(.DIN1 (____9___22714), .DIN2 (__9__0__26739), .Q
       (___09___24423));
  nor2s1 ___9___446217(.DIN1 (_________34970), .DIN2 (_________33442),
       .Q (____9____33647));
  or2s1 _______446218(.DIN1 (__9_____26675), .DIN2 (_____9__23230), .Q
       (__9__0__27025));
  nnd2s1 _______446219(.DIN1 (________23229), .DIN2 (___9____22505), .Q
       (________24528));
  nnd2s1 _______446220(.DIN1 (______0__33918), .DIN2 (_________34996),
       .Q (_________33916));
  nor2s1 _______446221(.DIN1 (___9____26194), .DIN2 (________22821), .Q
       (___0____24374));
  hi1s1 _______446222(.DIN (_________32442), .Q (____0____30977));
  and2s1 _____9_446223(.DIN1 (__9_____26677), .DIN2 (__9_____27027), .Q
       (________23900));
  nnd2s1 _______446224(.DIN1 (______0__33336), .DIN2 (________22758),
       .Q (_________33379));
  nor2s1 ___90__446225(.DIN1 (____0___20142), .DIN2 (________23227), .Q
       (________23228));
  nor2s1 _______446226(.DIN1 (____9___19395), .DIN2 (________22786), .Q
       (________23225));
  nor2s1 ______446227(.DIN1 (________20108), .DIN2 (___909__23355), .Q
       (________23224));
  nor2s1 ___9__446228(.DIN1 (___0____21654), .DIN2 (___0__9__27771), .Q
       (________23221));
  nor2s1 ___9_0_446229(.DIN1 (________23219), .DIN2 (__9_____26621), .Q
       (________23220));
  hi1s1 ___9___446230(.DIN (________23216), .Q (________23217));
  nor2s1 ___9___446231(.DIN1 (________19088), .DIN2 (________23212), .Q
       (_____0__23215));
  or2s1 ___9__446232(.DIN1 (___09___21712), .DIN2 (________23857), .Q
       (_____9__23214));
  or2s1 ___9___446233(.DIN1 (_________________18731), .DIN2
       (________23212), .Q (________23213));
  hi1s1 ____9__446234(.DIN (________23209), .Q (________23210));
  hi1s1 ____9__446235(.DIN (___09_0__28051), .Q (_____0__23208));
  nor2s1 ____9__446236(.DIN1 (____09__22634), .DIN2 (________22654), .Q
       (________23206));
  nor2s1 ____9__446237(.DIN1 (___9____22459), .DIN2 (________23204), .Q
       (________23205));
  nor2s1 ____9__446238(.DIN1 (________22065), .DIN2 (________23202), .Q
       (________23203));
  and2s1 ___90__446239(.DIN1 (________23200), .DIN2 (_____0__23199), .Q
       (________23201));
  nnd2s1 ____9_446240(.DIN1 (________23195), .DIN2 (____09__22634), .Q
       (________23197));
  nor2s1 ____9__446241(.DIN1 (________22906), .DIN2 (________23195), .Q
       (________23196));
  nor2s1 ____9__446242(.DIN1 (________23193), .DIN2 (________23192), .Q
       (________23194));
  nor2s1 ____9__446243(.DIN1 (________24221), .DIN2 (____0___23176), .Q
       (________23191));
  or2s1 ____99_446244(.DIN1 (________23814), .DIN2 (___999__26246), .Q
       (_____0__23190));
  nnd2s1 ____99_446245(.DIN1 (____99__23170), .DIN2 (________22123), .Q
       (_____9__23189));
  or2s1 ____99_446246(.DIN1 (____9___19395), .DIN2 (___999__26246), .Q
       (________23188));
  nor2s1 ___446247(.DIN1 (____90__22071), .DIN2 (________23156), .Q
       (________23187));
  or2s1 ___900_446248(.DIN1 (________19520), .DIN2 (____99__25654), .Q
       (________23186));
  nor2s1 ___900_446249(.DIN1 (____9___23164), .DIN2 (________23202), .Q
       (________23185));
  nnd2s1 ___446250(.DIN1 (________22645), .DIN2 (____0___22175), .Q
       (________23184));
  or2s1 ___90__446251(.DIN1 (_____9__22933), .DIN2 (____9___23709), .Q
       (________23183));
  nor2s1 ___90_446252(.DIN1 (________22920), .DIN2 (_____99__31353), .Q
       (_____0__23181));
  or2s1 ___90__446253(.DIN1 (________24660), .DIN2 (_____0__23286), .Q
       (____09__23180));
  and2s1 ___90__446254(.DIN1 (____0___23178), .DIN2 (________25401), .Q
       (____0___23179));
  nor2s1 ___90__446255(.DIN1 (____00__19399), .DIN2 (____0___23176), .Q
       (____0___23177));
  nor2s1 ___90__446256(.DIN1 (________22642), .DIN2 (________22941), .Q
       (____0___23175));
  nnd2s1 ______446257(.DIN1 (____0___23173), .DIN2 (____0___21909), .Q
       (____0___23174));
  nnd2s1 ___90__446258(.DIN1 (________22852), .DIN2 (___00___22538), .Q
       (____0___23172));
  nnd2s1 ___90__446259(.DIN1 (____99__23170), .DIN2 (____9___23169), .Q
       (____00__23171));
  nor2s1 ___90__446260(.DIN1 (__9_____26639), .DIN2 (____0___23266), .Q
       (____9___23168));
  or2s1 ___90__446261(.DIN1 (___99___26242), .DIN2 (____0___23266), .Q
       (____9___23167));
  nor2s1 ___90__446262(.DIN1 (________24944), .DIN2 (________23202), .Q
       (____9___23166));
  nnd2s1 ___90_446263(.DIN1 (____9___23164), .DIN2 (________21950), .Q
       (____9___23165));
  nnd2s1 ___90__446264(.DIN1 (____99__22806), .DIN2 (_____9__23161), .Q
       (____90__23162));
  or2s1 ___90__446265(.DIN1 (____0___19400), .DIN2 (___0__0__27609), .Q
       (________23160));
  nnd2s1 ___90__446266(.DIN1 (_____9__23275), .DIN2 (___99___23432), .Q
       (________23159));
  and2s1 ___90_446267(.DIN1 (__9__0__26637), .DIN2 (____0___23716), .Q
       (________23158));
  nor2s1 ___90_446268(.DIN1 (__9_____26937), .DIN2 (________23156), .Q
       (________23157));
  nnd2s1 ___90__446269(.DIN1 (________23200), .DIN2 (________23154), .Q
       (________23155));
  nor2s1 ___90__446270(.DIN1 (________22069), .DIN2 (_____0__23152), .Q
       (________23153));
  nor2s1 ___90__446271(.DIN1 (____0___22265), .DIN2 (_____0__23241), .Q
       (_____9__23151));
  nor2s1 ___90__446272(.DIN1 (________23149), .DIN2 (________23202), .Q
       (________23150));
  or2s1 ___90_446273(.DIN1 (________23147), .DIN2 (_____0__23241), .Q
       (________23148));
  or2s1 ___90__446274(.DIN1 (________23145), .DIN2 (____0___23266), .Q
       (________23146));
  and2s1 ___90__446275(.DIN1 (________24804), .DIN2 (_____9__23142), .Q
       (_____0__23143));
  nor2s1 ___90__446276(.DIN1 (________23140), .DIN2 (_____0__23241), .Q
       (________23141));
  nnd2s1 ___90__446277(.DIN1 (________23137), .DIN2 (________23136), .Q
       (________23138));
  nnd2s1 ___9___446278(.DIN1 (_____9__23275), .DIN2 (___9_9__23395), .Q
       (________23135));
  nnd2s1 ___909_446279(.DIN1 (________22673), .DIN2 (___9____24314), .Q
       (_____0__23134));
  nor2s1 ___909_446280(.DIN1 (___0_____27804), .DIN2 (________23132),
       .Q (_____9__23133));
  nnd2s1 ___9_0_446281(.DIN1 (________22423), .DIN2 (________23130), .Q
       (________23131));
  nnd2s1 ___9___446282(.DIN1 (________23862), .DIN2 (____99__22355), .Q
       (________23129));
  and2s1 ___9___446283(.DIN1 (____9___23342), .DIN2 (___00___22540), .Q
       (________23128));
  or2s1 ___9___446284(.DIN1 (____9___23342), .DIN2 (________23126), .Q
       (________23127));
  nnd2s1 ___9___446285(.DIN1 (________23288), .DIN2 (___00___22540), .Q
       (_____0__23125));
  nnd2s1 ___9___446286(.DIN1 (_____9__23275), .DIN2 (________23123), .Q
       (_____9__23124));
  and2s1 ___9___446287(.DIN1 (________23862), .DIN2 (________23121), .Q
       (________23122));
  nor2s1 ___9___446288(.DIN1 (________23119), .DIN2 (_____0__23286), .Q
       (________23120));
  and2s1 ___9__446289(.DIN1 (___0__0__27609), .DIN2 (___0_0___27563),
       .Q (________23118));
  nor2s1 ___9___446290(.DIN1 (___0____23484), .DIN2 (_____0__23286), .Q
       (________23117));
  nnd2s1 ___9___446291(.DIN1 (________23095), .DIN2 (_____0__23115), .Q
       (________23116));
  nnd2s1 ____446292(.DIN1 (________23137), .DIN2 (_____9__22107), .Q
       (________23112));
  or2s1 _______446293(.DIN1 (___0____23498), .DIN2 (_____0__22744), .Q
       (_____0__23775));
  nor2s1 _______446294(.DIN1 (________23111), .DIN2 (____9___25652), .Q
       (________23760));
  nnd2s1 _______446295(.DIN1 (____0___22628), .DIN2 (_____0__22200), .Q
       (________25814));
  or2s1 ______446296(.DIN1 (__9_9___26511), .DIN2 (________22834), .Q
       (________23699));
  nnd2s1 _______446297(.DIN1 (________22646), .DIN2 (________23110), .Q
       (______9__28301));
  nor2s1 _____9_446298(.DIN1 (____90__23965), .DIN2 (____0___23894), .Q
       (___9____23406));
  nnd2s1 _______446299(.DIN1 (________24777), .DIN2 (________22318), .Q
       (________23851));
  and2s1 _______446300(.DIN1 (___09___22618), .DIN2 (________23109), .Q
       (__9_____27041));
  nor2s1 _______446301(.DIN1 (________23729), .DIN2 (_____9__22789), .Q
       (____9___23797));
  nor2s1 ___9___446302(.DIN1 (________22742), .DIN2 (___09___22623), .Q
       (________23697));
  nor2s1 ___9___446303(.DIN1 (____0___22264), .DIN2 (________23227), .Q
       (___0_____27284));
  nor2s1 ___9___446304(.DIN1 (___0_0__23481), .DIN2 (____0___22629), .Q
       (_____9__23736));
  hi1s1 ____9__446305(.DIN (_________33177), .Q (_____0__23837));
  nor2s1 ___9___446306(.DIN1 (________21758), .DIN2 (_____9__22652), .Q
       (________23929));
  nor2s1 ___9__446307(.DIN1 (________23757), .DIN2 (_____0__23108), .Q
       (___0_9___27459));
  nnd2s1 ___9___446308(.DIN1 (_____9__23107), .DIN2 (________22678), .Q
       (________23742));
  nor2s1 ___9___446309(.DIN1 (_____0__21401), .DIN2 (____0___23266), .Q
       (________23907));
  nnd2s1 ___9___446310(.DIN1 (________23578), .DIN2 (__9__9__26921), .Q
       (________23920));
  nor2s1 ___9__446311(.DIN1 (________23106), .DIN2 (________23105), .Q
       (___0_9___27357));
  nnd2s1 ___9__446312(.DIN1 (________22658), .DIN2 (___9____23396), .Q
       (_____0__23765));
  nnd2s1 ___9___446313(.DIN1 (________22668), .DIN2 (________25524), .Q
       (___9____24279));
  nnd2s1 ___9___446314(.DIN1 (_____9__23275), .DIN2 (________22220), .Q
       (________23702));
  nor2s1 ___9___446315(.DIN1 (________23104), .DIN2 (____9___22804), .Q
       (_____9__23755));
  nor2s1 ___9_9_446316(.DIN1 (___0_0__22600), .DIN2 (_________34974),
       .Q (___990__23427));
  or2s1 _______446317(.DIN1 (________22730), .DIN2 (________23288), .Q
       (________23763));
  nnd2s1 _______446318(.DIN1 (________22673), .DIN2 (inData[23]), .Q
       (________23691));
  nor2s1 _______446319(.DIN1 (___9____24277), .DIN2 (_____0__22725), .Q
       (____0___23809));
  nor2s1 _______446320(.DIN1 (________23103), .DIN2 (_____9__23302), .Q
       (___9_0__23405));
  nor2s1 ___9___446321(.DIN1 (___0____22607), .DIN2 (________23156), .Q
       (___0_____27711));
  nnd2s1 ___9___446322(.DIN1 (_____9__23275), .DIN2 (________21845), .Q
       (___0_____27780));
  nor2s1 ___9___446323(.DIN1 (________21928), .DIN2 (_____0__23241), .Q
       (___0_____27877));
  and2s1 ___9___446324(.DIN1 (________23578), .DIN2 (____0___23085), .Q
       (___0_____27730));
  nor2s1 ___9___446325(.DIN1 (_________34986), .DIN2 (________22831),
       .Q (________23771));
  nnd2s1 ___9___446326(.DIN1 (____9___22805), .DIN2 (__9_____26784), .Q
       (___0_90__27938));
  or2s1 ___9___446327(.DIN1 (________23102), .DIN2 (________23070), .Q
       (___0_____27825));
  and2s1 ___9___446328(.DIN1 (____0___23178), .DIN2 (_____0__24616), .Q
       (_________28483));
  nnd2s1 ___9__446329(.DIN1 (________22666), .DIN2 (_________34982), .Q
       (_____9__25829));
  nor2s1 ___9___446330(.DIN1 (________26018), .DIN2 (________23156), .Q
       (___0_9___28034));
  nnd2s1 ___9_446331(.DIN1 (________23137), .DIN2 (________23101), .Q
       (____0___23806));
  or2s1 _______446332(.DIN1 (________23757), .DIN2 (________22671), .Q
       (__99____27150));
  nnd2s1 _______446333(.DIN1 (________23578), .DIN2 (________21951), .Q
       (____0_9__28185));
  nnd2s1 ___9_0_446334(.DIN1 (_____9__23275), .DIN2 (___9____20678), .Q
       (___9____24304));
  nor2s1 ___9_0_446335(.DIN1 (___90___23347), .DIN2 (________22858), .Q
       (________25509));
  nor2s1 ___9_0_446336(.DIN1 (____0___23716), .DIN2 (____99__25654), .Q
       (__9_____26671));
  nnd2s1 ___9_0_446337(.DIN1 (_________33236), .DIN2 (_________34970),
       .Q (_________33350));
  nor2s1 ___9_0_446338(.DIN1 (________24001), .DIN2 (___00____27202),
       .Q (___0_____27505));
  nor2s1 _____446339(.DIN1 (________23100), .DIN2 (_________34972), .Q
       (_____0___33037));
  nor2s1 _____9_446340(.DIN1 (________22947), .DIN2 (_________32925),
       .Q (______9__30207));
  and2s1 _____9_446341(.DIN1 (________22736), .DIN2 (_________35062),
       .Q (________25007));
  nor2s1 ____90_446342(.DIN1 (inData[1]), .DIN2 (___00____27202), .Q
       (________23689));
  nor2s1 ___9___446343(.DIN1 (________22655), .DIN2 (________24075), .Q
       (___09___25358));
  or2s1 _____9_446344(.DIN1 (_____9__23099), .DIN2 (________23227), .Q
       (__99____27110));
  and2s1 ___9_446345(.DIN1 (________23578), .DIN2 (_____9__21782), .Q
       (_____00__28331));
  nnd2s1 ____90_446346(.DIN1 (________23098), .DIN2 (____9___23795), .Q
       (____0___24160));
  nor2s1 ___9___446347(.DIN1 (________21457), .DIN2 (________23156), .Q
       (_________28667));
  nnd2s1 _____446348(.DIN1 (________22673), .DIN2 (inData[1]), .Q
       (_____9__23694));
  nor2s1 ___9___446349(.DIN1 (____0____29098), .DIN2 (________22664),
       .Q (_________31241));
  or2s1 ___99__446350(.DIN1 (_________28837), .DIN2 (__9_____26621), .Q
       (___0_____27485));
  nnd2s1 ____9__446351(.DIN1 (____0___22722), .DIN2 (________23097), .Q
       (_________28942));
  nnd2s1 ___9___446352(.DIN1 (________23578), .DIN2 (___9____21602), .Q
       (______9__28444));
  nnd2s1 ____9_446353(.DIN1 (________22750), .DIN2 (___9____22524), .Q
       (_____0___32294));
  nor2s1 ___9___446354(.DIN1 (________21893), .DIN2 (_____9__22733), .Q
       (_________31920));
  nor2s1 ___9___446355(.DIN1 (________22341), .DIN2 (____0___22627), .Q
       (_________32604));
  dffacs1 _____________0_(.CLRB (reset), .CLK (clk), .DIN
       (________22729), .QN (outData[0]));
  hi1s1 ___9__446356(.DIN (________23095), .Q (________23096));
  nnd2s1 _______446357(.DIN1 (___0____22558), .DIN2 (___90___22448), .Q
       (________23094));
  nnd2s1 ____9__446358(.DIN1 (___9____22471), .DIN2 (__9_____26828), .Q
       (________23093));
  xor2s1 _______446359(.DIN1 (_________34437), .DIN2 (____9____31746),
       .Q (_____0__23092));
  or2s1 ____9__446360(.DIN1 (___00____27182), .DIN2 (________23596), .Q
       (____09__23091));
  or2s1 ____9_446361(.DIN1 (__9_____26535), .DIN2 (____0___23088), .Q
       (____0___23089));
  nor2s1 ____9__446362(.DIN1 (___0_____27696), .DIN2 (___00___22539),
       .Q (____0___23087));
  nor2s1 ____9_446363(.DIN1 (____0___23085), .DIN2 (________22430), .Q
       (____0___23086));
  nnd2s1 _______446364(.DIN1 (_____0__22400), .DIN2 (inData[6]), .Q
       (____00__23084));
  or2s1 _______446365(.DIN1 (_________________18741), .DIN2
       (_________32492), .Q (____99__23083));
  or2s1 _______446366(.DIN1 (_________________18744), .DIN2
       (_________32492), .Q (____9___23082));
  nnd2s1 _______446367(.DIN1 (___999__22535), .DIN2 (_____0__21455), .Q
       (____9___23081));
  nor2s1 _______446368(.DIN1 (_____9__22223), .DIN2 (________22957), .Q
       (____9___23080));
  nor2s1 _______446369(.DIN1 (____00__24886), .DIN2 (___9____22486), .Q
       (____9___23079));
  nnd2s1 ______446370(.DIN1 (___9_0__22508), .DIN2 (inData[16]), .Q
       (____9___23078));
  nnd2s1 ______446371(.DIN1 (____0____31829), .DIN2 (_____9__19389), .Q
       (____9___23077));
  and2s1 _______446372(.DIN1 (____9___23075), .DIN2 (___9_0__26177), .Q
       (____9___23076));
  nor2s1 _______446373(.DIN1 (____09__21820), .DIN2 (_____9__23055), .Q
       (____90__23074));
  nnd2s1 _______446374(.DIN1 (________23033), .DIN2 (________23101), .Q
       (_____9__23073));
  nor2s1 ______446375(.DIN1 (________23071), .DIN2 (________23070), .Q
       (________23072));
  nor2s1 _______446376(.DIN1 (____0___22086), .DIN2 (________22418), .Q
       (________23069));
  nnd2s1 _______446377(.DIN1 (___9____22514), .DIN2 (___90___20612), .Q
       (________23068));
  and2s1 _______446378(.DIN1 (________23066), .DIN2 (____00__19399), .Q
       (________23067));
  nor2s1 _______446379(.DIN1 (________23101), .DIN2 (___9____22511), .Q
       (_____0__23065));
  or2s1 ______446380(.DIN1 (________23063), .DIN2 (________23062), .Q
       (_____9__23064));
  nor2s1 ______446381(.DIN1 (____0___21987), .DIN2 (_____0__22772), .Q
       (________23061));
  or2s1 _______446382(.DIN1 (________22194), .DIN2 (________23066), .Q
       (________23060));
  and2s1 _______446383(.DIN1 (________23058), .DIN2 (________23057), .Q
       (________23059));
  nor2s1 _______446384(.DIN1 (________20996), .DIN2 (_____9__23055), .Q
       (_____0__23056));
  nnd2s1 _______446385(.DIN1 (___00___22537), .DIN2 (___9____21563), .Q
       (________23054));
  or2s1 _______446386(.DIN1 (________23052), .DIN2 (___9____22474), .Q
       (________23053));
  nor2s1 ______446387(.DIN1 (___9____22504), .DIN2 (________23050), .Q
       (________23051));
  nor2s1 _______446388(.DIN1 (___999__21632), .DIN2 (________22402), .Q
       (________23049));
  nnd2s1 _______446389(.DIN1 (________25728), .DIN2 (___00___22540), .Q
       (________23048));
  and2s1 _______446390(.DIN1 (________22917), .DIN2 (____9___25168), .Q
       (_____9__23047));
  or2s1 _______446391(.DIN1 (___90___24245), .DIN2 (________23045), .Q
       (________23046));
  and2s1 _______446392(.DIN1 (________22849), .DIN2 (________23043), .Q
       (________23044));
  nor2s1 _______446393(.DIN1 (________23123), .DIN2 (________22230), .Q
       (________23042));
  nnd2s1 _______446394(.DIN1 (________23040), .DIN2 (________23039), .Q
       (________23041));
  nnd2s1 _______446395(.DIN1 (___9____22502), .DIN2 (_____9__21522), .Q
       (_____0__23038));
  or2s1 ______446396(.DIN1 (____0___21817), .DIN2 (________23036), .Q
       (_____9__23037));
  nnd2s1 _____9_446397(.DIN1 (________24852), .DIN2 (________22158), .Q
       (________23035));
  nnd2s1 _____9_446398(.DIN1 (________23033), .DIN2 (________22106), .Q
       (________23034));
  nnd2s1 _____9_446399(.DIN1 (________23031), .DIN2 (________23030), .Q
       (________23032));
  nnd2s1 _____9_446400(.DIN1 (________23026), .DIN2 (_____0__23028), .Q
       (________23029));
  nor2s1 _____9_446401(.DIN1 (________23814), .DIN2 (________23026), .Q
       (_____9__23027));
  nor2s1 _____0_446402(.DIN1 (________23015), .DIN2 (________23070), .Q
       (________23025));
  nnd2s1 _____0_446403(.DIN1 (___000__22536), .DIN2 (___9____21581), .Q
       (________23024));
  and2s1 _____0_446404(.DIN1 (________23022), .DIN2 (________23021), .Q
       (________23023));
  and2s1 _____446405(.DIN1 (___0____22615), .DIN2 (____9___23794), .Q
       (________23020));
  nor2s1 _______446406(.DIN1 (________22387), .DIN2 (___9____23371), .Q
       (________23019));
  and2s1 _______446407(.DIN1 (_____9__23017), .DIN2 (____9___22354), .Q
       (_____0__23018));
  nnd2s1 ______446408(.DIN1 (________23015), .DIN2 (__9_____26937), .Q
       (________23016));
  and2s1 _______446409(.DIN1 (_____9__22399), .DIN2 (____0___23620), .Q
       (________23013));
  nnd2s1 _______446410(.DIN1 (_____9__22980), .DIN2 (________22876), .Q
       (________23012));
  nnd2s1 _______446411(.DIN1 (________23010), .DIN2 (________22748), .Q
       (________23011));
  nnd2s1 _______446412(.DIN1 (____0____31829), .DIN2 (________19089),
       .Q (_____0__23009));
  nnd2s1 ______446413(.DIN1 (____0___24704), .DIN2 (________23007), .Q
       (_____9__23008));
  nnd2s1 _______446414(.DIN1 (__9_00), .DIN2 (________23005), .Q
       (________23006));
  nnd2s1 ____9_446415(.DIN1 (________23003), .DIN2 (_____9__22689), .Q
       (________23004));
  nor2s1 _______446416(.DIN1 (________20005), .DIN2 (___0____22556), .Q
       (________23002));
  and2s1 _______446417(.DIN1 (________23000), .DIN2 (____09__22634), .Q
       (________23001));
  nor2s1 ______446418(.DIN1 (________22943), .DIN2 (____09__22998), .Q
       (_____0__22999));
  nnd2s1 ______446419(.DIN1 (________22909), .DIN2 (_____9__22251), .Q
       (____0___22997));
  nor2s1 _______446420(.DIN1 (____0___22362), .DIN2 (___9_9__22507), .Q
       (____0___22996));
  nnd2s1 ______446421(.DIN1 (____9___23075), .DIN2 (________21921), .Q
       (____0___22995));
  nnd2s1 ______446422(.DIN1 (_________32049), .DIN2 (___0_____27914),
       .Q (____0___22994));
  or2s1 _______446423(.DIN1 (____0___22992), .DIN2 (____0___22991), .Q
       (____0___22993));
  and2s1 _______446424(.DIN1 (__9_____26469), .DIN2 (___9_0__22481), .Q
       (____0___22990));
  nnd2s1 _______446425(.DIN1 (________22403), .DIN2 (____9___19945), .Q
       (____00__22989));
  or2s1 _______446426(.DIN1 (________22142), .DIN2 (________22659), .Q
       (____9___22988));
  nor2s1 _______446427(.DIN1 (________21761), .DIN2 (________23596), .Q
       (____9___22987));
  nor2s1 _______446428(.DIN1 (___0____22562), .DIN2 (________25535), .Q
       (____9___22985));
  nnd2s1 _______446429(.DIN1 (________22768), .DIN2 (________22315), .Q
       (____9___22984));
  nnd2s1 _______446430(.DIN1 (________25394), .DIN2 (____9___22982), .Q
       (____9___22983));
  nnd2s1 _______446431(.DIN1 (_____9__22980), .DIN2 (_____0__22327), .Q
       (____90__22981));
  nnd2s1 _______446432(.DIN1 (___9____22484), .DIN2 (____9___22254), .Q
       (________22979));
  nnd2s1 _____9_446433(.DIN1 (___9____22485), .DIN2 (________22217), .Q
       (________22978));
  and2s1 _____9_446434(.DIN1 (________22964), .DIN2 (________24824), .Q
       (________22977));
  nnd2s1 _____9_446435(.DIN1 (____0____31829), .DIN2 (________20586),
       .Q (________22976));
  nor2s1 _____446436(.DIN1 (___0_0__23481), .DIN2 (________22775), .Q
       (________22975));
  hi1s1 ____9__446437(.DIN (________23327), .Q (________22974));
  hi1s1 ____9_446438(.DIN (________22972), .Q (________22973));
  nnd2s1 ___9_0_446439(.DIN1 (_____0__22680), .DIN2 (________22969), .Q
       (________22970));
  nor2s1 ___9___446440(.DIN1 (________25973), .DIN2 (________23596), .Q
       (________22968));
  nor2s1 _____446441(.DIN1 (___9_0__26207), .DIN2 (________23066), .Q
       (________23537));
  and2s1 _______446442(.DIN1 (___09___25361), .DIN2 (________22967), .Q
       (________24568));
  nor2s1 _______446443(.DIN1 (___9____21573), .DIN2 (________22966), .Q
       (___09___23525));
  nor2s1 _______446444(.DIN1 (________22965), .DIN2 (________22959), .Q
       (____09__23627));
  or2s1 _______446445(.DIN1 (___99___22528), .DIN2 (__90____26275), .Q
       (___9____24290));
  nnd2s1 _______446446(.DIN1 (___09___25361), .DIN2 (__9_____26917), .Q
       (_____9__23637));
  and2s1 ______446447(.DIN1 (________23040), .DIN2 (________22964), .Q
       (___9____23398));
  nor2s1 _______446448(.DIN1 (___9____21597), .DIN2 (____9___22890), .Q
       (________23644));
  nnd2s1 _______446449(.DIN1 (________23003), .DIN2 (________22963), .Q
       (________23548));
  nor2s1 _______446450(.DIN1 (____00__19399), .DIN2 (________22380), .Q
       (___00___25273));
  nnd2s1 _______446451(.DIN1 (________24852), .DIN2 (_________35046),
       .Q (________23315));
  nor2s1 _______446452(.DIN1 (_____0__22962), .DIN2 (________23000), .Q
       (_____0__23223));
  nnd2s1 _______446453(.DIN1 (________24202), .DIN2 (___9____22461), .Q
       (_____9__23554));
  nnd2s1 _______446454(.DIN1 (_____9__22961), .DIN2 (________22373), .Q
       (___0_____27524));
  nnd2s1 ______446455(.DIN1 (________22301), .DIN2 (________22960), .Q
       (___0__0__27714));
  nor2s1 ______446456(.DIN1 (________25478), .DIN2 (___9____22521), .Q
       (________23314));
  nor2s1 _______446457(.DIN1 (________22959), .DIN2 (____0___24522), .Q
       (_____0__23536));
  nor2s1 _______446458(.DIN1 (________22958), .DIN2 (___9____22513), .Q
       (________23654));
  nnd2s1 _______446459(.DIN1 (___9_9__22480), .DIN2 (________23814), .Q
       (___0_____27473));
  nnd2s1 _______446460(.DIN1 (________23039), .DIN2 (________22948), .Q
       (________23237));
  nnd2s1 ___9__446461(.DIN1 (________23010), .DIN2 (________21280), .Q
       (________23607));
  nor2s1 _______446462(.DIN1 (________22144), .DIN2 (___9____26209), .Q
       (________23235));
  nor2s1 _______446463(.DIN1 (__9_9___26511), .DIN2 (________24722), .Q
       (________23226));
  nnd2s1 ___9__446464(.DIN1 (___9____22518), .DIN2 (___9____26163), .Q
       (________23209));
  nor2s1 _____0_446465(.DIN1 (________22311), .DIN2 (________22957), .Q
       (___09___23524));
  nnd2s1 _______446466(.DIN1 (___9____22501), .DIN2 (___90___22451), .Q
       (________23604));
  hi1s1 ____9__446467(.DIN (________22956), .Q (_____0__24163));
  nor2s1 _____0_446468(.DIN1 (_____0__20474), .DIN2 (___9____22525), .Q
       (________23996));
  nor2s1 _____0_446469(.DIN1 (___0_0__22573), .DIN2 (___9____22488), .Q
       (________23316));
  or2s1 ______446470(.DIN1 (____09__23983), .DIN2 (________25728), .Q
       (___099__23527));
  nor2s1 _______446471(.DIN1 (___9____26213), .DIN2 (___00___22542), .Q
       (___09___23523));
  nnd2s1 _______446472(.DIN1 (________22406), .DIN2 (___99___22527), .Q
       (___0_____27816));
  nnd2s1 ______446473(.DIN1 (____90__25840), .DIN2 (________24824), .Q
       (________23670));
  nor2s1 _______446474(.DIN1 (________22954), .DIN2 (________23062), .Q
       (___0_____28002));
  nnd2s1 ______446475(.DIN1 (________22953), .DIN2 (_____0__22952), .Q
       (____9___24695));
  nor2s1 _______446476(.DIN1 (_____9__22951), .DIN2 (________23932), .Q
       (________24817));
  and2s1 _______446477(.DIN1 (___9____22498), .DIN2 (________22960), .Q
       (__9_____26722));
  nor2s1 _____9_446478(.DIN1 (___9____24263), .DIN2 (________22950), .Q
       (________23652));
  nor2s1 _____9_446479(.DIN1 (________23757), .DIN2 (___9____22523), .Q
       (___0_____27783));
  nor2s1 _____9_446480(.DIN1 (_____0__25156), .DIN2 (___9____24318), .Q
       (________24094));
  nor2s1 _____9_446481(.DIN1 (________23292), .DIN2 (________23596), .Q
       (___09____28066));
  hi1s1 ___9___446482(.DIN (________22949), .Q (___0____23497));
  nnd2s1 _______446483(.DIN1 (________22953), .DIN2 (________26099), .Q
       (___0____25324));
  hi1s1 _______446484(.DIN (__9_____26675), .Q (________23679));
  nnd2s1 _______446485(.DIN1 (________24202), .DIN2 (____9___23794), .Q
       (____0___23622));
  or2s1 _______446486(.DIN1 (__9_____26597), .DIN2 (___9____23401), .Q
       (________23767));
  nnd2s1 ______446487(.DIN1 (________22953), .DIN2 (________22095), .Q
       (________25027));
  nnd2s1 ______446488(.DIN1 (___9____23402), .DIN2 (________22948), .Q
       (________23593));
  nnd2s1 _______446489(.DIN1 (____0____31829), .DIN2 (________22947),
       .Q (________23662));
  nnd2s1 _______446490(.DIN1 (____00__25948), .DIN2 (____90__25840), .Q
       (________24483));
  nor2s1 _______446491(.DIN1 (____9___22170), .DIN2 (___99___22534), .Q
       (________25068));
  hi1s1 ______446492(.DIN (______0__33918), .Q (________23667));
  nnd2s1 ____90_446493(.DIN1 (____00__25948), .DIN2 (________22946), .Q
       (________25812));
  nnd2s1 ____9__446494(.DIN1 (___9____22515), .DIN2 (____9___22438), .Q
       (_________32442));
  hi1s1 ____9__446495(.DIN (__9_____27027), .Q (________23676));
  nnd2s1 ____9__446496(.DIN1 (___9____23402), .DIN2 (________22945), .Q
       (________25793));
  nor2s1 ____9__446497(.DIN1 (__9_____26754), .DIN2 (___9____26209), .Q
       (________25991));
  nnd2s1 ____90_446498(.DIN1 (___9____23373), .DIN2 (_____0__22952), .Q
       (________26092));
  nor2s1 ____9__446499(.DIN1 (________22332), .DIN2 (___9____22489), .Q
       (_________31060));
  or2s1 ____9_446500(.DIN1 (________23097), .DIN2 (___0_0___27659), .Q
       (____9____29042));
  hi1s1 _______446501(.DIN (_________29736), .Q (____0____32807));
  hi1s1 ___9__446502(.DIN (________23862), .Q (___00___23441));
  nor2s1 ____9__446503(.DIN1 (_____0__19918), .DIN2 (___0____22561), .Q
       (____0____32777));
  nor2s1 ____9__446504(.DIN1 (________21127), .DIN2 (___9____22519), .Q
       (____0____31820));
  nor2s1 ____9__446505(.DIN1 (____0___21813), .DIN2 (___9____22494), .Q
       (________23683));
  nnd2s1 ____9__446506(.DIN1 (___9_9__22499), .DIN2 (________22672), .Q
       (____9_0__33597));
  nor2s1 ____9__446507(.DIN1 (____9___22352), .DIN2 (________22943), .Q
       (________22944));
  nor2s1 ____9__446508(.DIN1 (________21949), .DIN2 (________22941), .Q
       (_____9__22942));
  nnd2s1 ____99_446509(.DIN1 (__9_00), .DIN2 (________22938), .Q
       (________22939));
  nor2s1 ____99_446510(.DIN1 (_____9__21933), .DIN2 (________23062), .Q
       (________22937));
  nnd2s1 ____99_446511(.DIN1 (_____9__22961), .DIN2 (________22392), .Q
       (________22936));
  nnd2s1 ___900_446512(.DIN1 (___0____22545), .DIN2 (________25672), .Q
       (________22935));
  nor2s1 ___900_446513(.DIN1 (_____9__22933), .DIN2 (________22407), .Q
       (_____0__22934));
  nnd2s1 ___900_446514(.DIN1 (________22931), .DIN2 (___9____22456), .Q
       (________22932));
  nnd2s1 ___900_446515(.DIN1 (________23031), .DIN2 (___0____22613), .Q
       (________22930));
  nor2s1 ___90_446516(.DIN1 (________24221), .DIN2 (________22414), .Q
       (________22929));
  nnd2s1 ___90__446517(.DIN1 (________25861), .DIN2 (____0___21910), .Q
       (________22928));
  nnd2s1 ___90__446518(.DIN1 (________23033), .DIN2 (___9____22492), .Q
       (________22927));
  nnd2s1 ___90__446519(.DIN1 (________23033), .DIN2 (_____9__24828), .Q
       (________22926));
  nnd2s1 ___90__446520(.DIN1 (_____9__22961), .DIN2 (_____0__22924), .Q
       (________22925));
  nnd2s1 ___90__446521(.DIN1 (_____0__22816), .DIN2 (________22765), .Q
       (_____9__22923));
  nor2s1 ___90__446522(.DIN1 (_____0__23199), .DIN2 (___9____22497), .Q
       (________22922));
  nnd2s1 ___90__446523(.DIN1 (_________33444), .DIN2 (________22920),
       .Q (________22921));
  nor2s1 ___90__446524(.DIN1 (_____9__21344), .DIN2 (___99___22531), .Q
       (________22919));
  or2s1 ___90__446525(.DIN1 (________22917), .DIN2 (________23070), .Q
       (________22918));
  nor2s1 ___90_446526(.DIN1 (________19222), .DIN2 (________22915), .Q
       (________22916));
  nor2s1 ___90__446527(.DIN1 (____9___19395), .DIN2 (_____9__22426), .Q
       (_____0__22914));
  and2s1 ___90__446528(.DIN1 (________22957), .DIN2 (________19520), .Q
       (________22913));
  or2s1 ___90__446529(.DIN1 (____0___22085), .DIN2 (________23596), .Q
       (________22912));
  nor2s1 ___90__446530(.DIN1 (___9____26159), .DIN2 (________23596), .Q
       (________22911));
  nnd2s1 ___90__446531(.DIN1 (________22909), .DIN2 (_____0__21934), .Q
       (________22910));
  or2s1 ___90__446532(.DIN1 (________22907), .DIN2 (________22906), .Q
       (________22908));
  nnd2s1 ___90__446533(.DIN1 (____09__22904), .DIN2 (________23149), .Q
       (_____0__22905));
  or2s1 ___90__446534(.DIN1 (________22103), .DIN2 (________23062), .Q
       (____0___22903));
  nor2s1 ___90__446535(.DIN1 (___9____23387), .DIN2 (____0___22901), .Q
       (____0___22902));
  nor2s1 ___909_446536(.DIN1 (____0___21993), .DIN2 (________23596), .Q
       (____0___22900));
  nor2s1 ___909_446537(.DIN1 (_____0__22148), .DIN2 (________22941), .Q
       (____0___22899));
  or2s1 ___909_446538(.DIN1 (__9_____26639), .DIN2 (________23062), .Q
       (____0___22898));
  nnd2s1 ___9_0_446539(.DIN1 (____0___22721), .DIN2 (____9___22353), .Q
       (____0___22897));
  nnd2s1 ___9_0_446540(.DIN1 (________22411), .DIN2 (________23119), .Q
       (____0___22896));
  or2s1 ___9_0_446541(.DIN1 (____99__22894), .DIN2 (________22419), .Q
       (____00__22895));
  nnd2s1 ___9___446542(.DIN1 (________22422), .DIN2 (________23814), .Q
       (____9___22893));
  nor2s1 ___9___446543(.DIN1 (____0___22179), .DIN2 (________23070), .Q
       (____9___22892));
  nor2s1 ___9___446544(.DIN1 (________23147), .DIN2 (____9___22890), .Q
       (____9___22891));
  nor2s1 ___9___446545(.DIN1 (___0_9__22572), .DIN2 (_____0__22271), .Q
       (____9___22889));
  nor2s1 ___9___446546(.DIN1 (____0___22262), .DIN2 (____9___22890), .Q
       (____9___22888));
  nor2s1 ___9__446547(.DIN1 (____9___22886), .DIN2 (________23596), .Q
       (____9___22887));
  or2s1 ___9__446548(.DIN1 (_____9__22884), .DIN2 (____9___22890), .Q
       (____90__22885));
  or2s1 ___9___446549(.DIN1 (________22882), .DIN2 (____9___22890), .Q
       (________22883));
  and2s1 ___9___446550(.DIN1 (___0____22555), .DIN2 (________23119), .Q
       (________22881));
  nnd2s1 ___9__446551(.DIN1 (_____9__22961), .DIN2 (_____9__23161), .Q
       (________22880));
  and2s1 ___9___446552(.DIN1 (________25139), .DIN2 (____0___24890), .Q
       (________22879));
  and2s1 ___9___446553(.DIN1 (_____9__22961), .DIN2 (________22146), .Q
       (________22878));
  nor2s1 ___9___446554(.DIN1 (________19570), .DIN2 (________22876), .Q
       (________22877));
  hi1s1 ___9___446555(.DIN (________24804), .Q (_____0__22875));
  nor2s1 ___9_446556(.DIN1 (________22685), .DIN2 (__9_____26773), .Q
       (_____9__22874));
  nnd2s1 _____9_446557(.DIN1 (________22787), .DIN2 (________22872), .Q
       (________22873));
  nnd2s1 ______446558(.DIN1 (________22870), .DIN2 (________22869), .Q
       (________22871));
  hi1s1 _____9_446559(.DIN (________22867), .Q (________22868));
  or2s1 _____9_446560(.DIN1 (___0_0__22564), .DIN2 (________23541), .Q
       (________22866));
  nnd2s1 _______446561(.DIN1 (________22404), .DIN2 (inData[30]), .Q
       (_____0__22865));
  nor2s1 ___9___446562(.DIN1 (_____0__21995), .DIN2 (__90____26312), .Q
       (_____9__22864));
  nnd2s1 ___9___446563(.DIN1 (________22845), .DIN2 (________21935), .Q
       (________22863));
  nnd2s1 ___9__446564(.DIN1 (__9_____26962), .DIN2 (________24183), .Q
       (________22862));
  nnd2s1 ___9___446565(.DIN1 (________26121), .DIN2 (___0____21662), .Q
       (________22861));
  or2s1 ___9___446566(.DIN1 (________22859), .DIN2 (________22858), .Q
       (________22860));
  nor2s1 ___9_9_446567(.DIN1 (___0____19799), .DIN2 (________22835), .Q
       (________22857));
  nor2s1 ___9___446568(.DIN1 (_____0__22855), .DIN2 (________22819), .Q
       (________22856));
  nnd2s1 ___9___446569(.DIN1 (_____9__22847), .DIN2 (________22853), .Q
       (_____9__22854));
  or2s1 ____9__446570(.DIN1 (__9__0__26346), .DIN2 (___9____22468), .Q
       (________22851));
  and2s1 ____9__446571(.DIN1 (________22849), .DIN2 (_____0__22138), .Q
       (________22850));
  nnd2s1 ___9___446572(.DIN1 (_____9__22847), .DIN2 (________22151), .Q
       (_____0__22848));
  nnd2s1 ___9___446573(.DIN1 (________22845), .DIN2 (____90__24877), .Q
       (________22846));
  nor2s1 ___9___446574(.DIN1 (________22196), .DIN2 (__9_____26773), .Q
       (________22844));
  nor2s1 ___9___446575(.DIN1 (________19239), .DIN2 (____0____32793),
       .Q (________22843));
  nnd2s1 ___9_0_446576(.DIN1 (________22372), .DIN2 (_____0__23811), .Q
       (________22842));
  nnd2s1 ___9_9_446577(.DIN1 (_____0__22384), .DIN2 (________22840), .Q
       (________22841));
  nnd2s1 ___9_9_446578(.DIN1 (____00__22807), .DIN2 (_________34980),
       .Q (________22839));
  nnd2s1 ___9_9_446579(.DIN1 (___9____25213), .DIN2 (inData[20]), .Q
       (_____9__22838));
  and2s1 ___9___446580(.DIN1 (________22377), .DIN2 (___9____23416), .Q
       (________22837));
  nor2s1 ___9___446581(.DIN1 (______18939), .DIN2 (________22835), .Q
       (________22836));
  hi1s1 ___9___446582(.DIN (________22831), .Q (_____9__22832));
  hi1s1 ___9_9_446583(.DIN (________24024), .Q (________22830));
  nor2s1 ___9___446584(.DIN1 (____09__21994), .DIN2 (__90____26312), .Q
       (________22829));
  nnd2s1 ___9__446585(.DIN1 (___9____25213), .DIN2 (inData[21]), .Q
       (________22828));
  nnd2s1 ___9__446586(.DIN1 (___9____25213), .DIN2 (inData[16]), .Q
       (________22827));
  nnd2s1 ___9___446587(.DIN1 (________22395), .DIN2 (inData[0]), .Q
       (_____0__22826));
  nor2s1 ___9___446588(.DIN1
       (______________________________________0_____________18891),
       .DIN2 (___9____25213), .Q (_____9__22825));
  nnd2s1 ___9___446589(.DIN1 (________22396), .DIN2 (inData[28]), .Q
       (________22824));
  or2s1 ___9___446590(.DIN1 (________22152), .DIN2 (________22823), .Q
       (___9____23400));
  hi1s1 ___9___446591(.DIN (________22822), .Q (___0____23465));
  and2s1 ___9___446592(.DIN1 (___9____22477), .DIN2 (____0___25560), .Q
       (____9___23879));
  hi1s1 ______446593(.DIN (________22821), .Q (___09___23519));
  nor2s1 ___9__446594(.DIN1 (________22285), .DIN2 (________23070), .Q
       (____0___24611));
  nor2s1 ___9___446595(.DIN1 (_____0__24541), .DIN2 (____90__25939), .Q
       (___9____23403));
  nor2s1 ___9___446596(.DIN1 (________25715), .DIN2 (________25413), .Q
       (________23211));
  nnd2s1 ___9___446597(.DIN1 (______0__34978), .DIN2 (__9_____26370),
       .Q (________23113));
  nor2s1 ___9___446598(.DIN1 (________22820), .DIN2 (________22819), .Q
       (________23114));
  nnd2s1 ___9___446599(.DIN1 (________23003), .DIN2 (________25394), .Q
       (___9____23410));
  nnd2s1 ___9_9_446600(.DIN1 (________22379), .DIN2 (___09___23522), .Q
       (__9_0___26427));
  nor2s1 ___9___446601(.DIN1 (___0____22590), .DIN2 (________22835), .Q
       (___0____23477));
  nnd2s1 ___9_446602(.DIN1 (__9_____26469), .DIN2 (____0___22176), .Q
       (__9__9__26691));
  nnd2s1 ___9_9_446603(.DIN1 (________22385), .DIN2 (________22818), .Q
       (________24171));
  nor2s1 ___9___446604(.DIN1 (_____0__22427), .DIN2 (___0____22570), .Q
       (_____0___28337));
  nnd2s1 ___9_9_446605(.DIN1 (________24669), .DIN2 (________21736), .Q
       (___0_9__23463));
  nor2s1 ___9___446606(.DIN1 (________22394), .DIN2 (________21758), .Q
       (__9_____26959));
  nor2s1 ___9___446607(.DIN1 (___90___22453), .DIN2 (_____0__23303), .Q
       (________23216));
  nor2s1 ___9__446608(.DIN1 (________22817), .DIN2 (________22413), .Q
       (________23580));
  and2s1 ___9___446609(.DIN1 (________23033), .DIN2 (__9_____26553), .Q
       (_____9__23914));
  nnd2s1 ___9___446610(.DIN1 (___9____22473), .DIN2 (________23236), .Q
       (________23635));
  nor2s1 ___9___446611(.DIN1 (_____0__22816), .DIN2 (________25535), .Q
       (___09___23521));
  nnd2s1 ___9_9_446612(.DIN1 (________22909), .DIN2 (__9_____26784), .Q
       (____0___23805));
  nnd2s1 ___9___446613(.DIN1 (___00___22541), .DIN2 (____0___23529), .Q
       (___9_9__23404));
  nnd2s1 ___9___446614(.DIN1 (________22389), .DIN2 (____09__22815), .Q
       (____0___24990));
  nnd2s1 ___9_0_446615(.DIN1 (_____9__22961), .DIN2 (____0___22363), .Q
       (___0_____27915));
  nnd2s1 ___9___446616(.DIN1 (________22429), .DIN2 (________24440), .Q
       (________24232));
  nor2s1 ___9_0_446617(.DIN1 (________23145), .DIN2 (________23062), .Q
       (___0_____27921));
  and2s1 ___9___446618(.DIN1 (_____0__22417), .DIN2 (________22946), .Q
       (____0___25566));
  nor2s1 ___9___446619(.DIN1 (____00__21446), .DIN2 (____9___22890), .Q
       (________24904));
  nor2s1 ___9___446620(.DIN1 (___0____22602), .DIN2 (___9____25213), .Q
       (________25142));
  nor2s1 ___9_446621(.DIN1 (________23140), .DIN2 (____9___22890), .Q
       (___0_____27798));
  nnd2s1 ___9___446622(.DIN1 (_____9__25596), .DIN2 (____9___21805), .Q
       (________23583));
  and2s1 ___9__446623(.DIN1 (________25861), .DIN2 (_________35056), .Q
       (________23740));
  or2s1 ___9__446624(.DIN1 (________22029), .DIN2 (________23070), .Q
       (___9____25223));
  or2s1 ___9___446625(.DIN1 (_____0__25694), .DIN2 (___9____22467), .Q
       (___99___24329));
  and2s1 ___9___446626(.DIN1 (___0____22560), .DIN2 (_________28602),
       .Q (________25004));
  or2s1 ___9___446627(.DIN1 (____0___22814), .DIN2 (________23070), .Q
       (___0__9__27839));
  nor2s1 ___9___446628(.DIN1 (_________33103), .DIN2 (________22915),
       .Q (____9____32719));
  nnd2s1 ___9___446629(.DIN1 (_____9__22961), .DIN2 (___9____21605), .Q
       (___09_0__28051));
  and2s1 ___9___446630(.DIN1 (_____9__24655), .DIN2 (___0____25333), .Q
       (_____0__25665));
  nor2s1 ___9__446631(.DIN1 (____0___22813), .DIN2 (________22386), .Q
       (_____0__24120));
  nnd2s1 ___9___446632(.DIN1 (________22909), .DIN2 (___0____21700), .Q
       (___09____28078));
  nor2s1 ___9___446633(.DIN1 (__9_____26937), .DIN2 (________23070), .Q
       (___0__0__28004));
  nor2s1 ___9__446634(.DIN1 (___99___21631), .DIN2 (____9___22890), .Q
       (______9__28588));
  hi1s1 ___9___446635(.DIN (____0___22810), .Q (___0____23482));
  or2s1 ___990_446636(.DIN1 (____0___22812), .DIN2 (________22383), .Q
       (________25424));
  nor2s1 ___99_446637(.DIN1 (___9____21559), .DIN2 (_____9__22391), .Q
       (__9_____26447));
  hi1s1 ___9_0_446638(.DIN (________23137), .Q (___0____23450));
  hi1s1 _______446639(.DIN (______0__33336), .Q (_________33180));
  nor2s1 ___99_446640(.DIN1 (____0___22811), .DIN2 (________22940), .Q
       (_____0__25520));
  nnd2s1 ___9___446641(.DIN1 (_____9__24007), .DIN2 (________22340), .Q
       (___9_9__25202));
  nor2s1 ___99__446642(.DIN1 (_____9__22215), .DIN2 (________22397), .Q
       (__9_____26831));
  nor2s1 ___9__446643(.DIN1 (________21422), .DIN2 (_________33153), .Q
       (_________33177));
  hi1s1 ___9___446644(.DIN (_____0__23286), .Q (_____0__24140));
  dffacs1 __________________446645(.CLRB (reset), .CLK (clk), .DIN
       (________22428), .Q (______________0___________________0));
  hi1s1 ___9_446646(.DIN (_____0__23241), .Q (___0____23453));
  hi1s1 ____9__446647(.DIN (_________33325), .Q (______9__32620));
  hi1s1 ___9__446648(.DIN (________23202), .Q (___0____23506));
  hi1s1 ___9___446649(.DIN (____99__23170), .Q (___0____23495));
  nnd2s1 ___9___446650(.DIN1 (___0_9__22553), .DIN2 (________22000), .Q
       (_________32158));
  hi1s1 ___9___446651(.DIN (____0___23178), .Q (___000__23437));
  hi1s1 ___9___446652(.DIN (_________34972), .Q (______0__33058));
  nnd2s1 ___9___446653(.DIN1 (___9_0__22517), .DIN2 (___0____22587), .Q
       (____0___22809));
  nnd2s1 ___9___446654(.DIN1 (____00__22807), .DIN2 (___0_0__22554), .Q
       (____0___22808));
  hi1s1 ___9___446655(.DIN (________23070), .Q (____99__22806));
  hi1s1 ___9___446656(.DIN (________23062), .Q (____9___22805));
  hi1s1 ___9__446657(.DIN (____9___22803), .Q (____9___22804));
  nnd2s1 ___9___446658(.DIN1 (____0___22174), .DIN2 (inData[8]), .Q
       (____9___22802));
  nor2s1 ___9___446659(.DIN1 (________24659), .DIN2 (________22697), .Q
       (____9___22801));
  or2s1 ___9___446660(.DIN1 (____9___22799), .DIN2 (_____9__22241), .Q
       (____9___22800));
  or2s1 ___9___446661(.DIN1 (____________9___18758), .DIN2
       (_____9__22797), .Q (____90__22798));
  nor2s1 ___9___446662(.DIN1 (________24221), .DIN2 (________22195), .Q
       (________22796));
  nor2s1 ___9__446663(.DIN1 (inData[19]), .DIN2 (________22737), .Q
       (________22795));
  and2s1 ___9___446664(.DIN1 (_____0___32572), .DIN2 (___0___18984), .Q
       (________22794));
  xor2s1 _______446665(.DIN1 (____9___22072), .DIN2 (___90___23353), .Q
       (________22793));
  xor2s1 _______446666(.DIN1 (_________34448), .DIN2 (_________33333),
       .Q (________22792));
  hi1s1 ___9___446667(.DIN (________23030), .Q (________22791));
  hi1s1 ___9_446668(.DIN (_____9__22980), .Q (_____0__22790));
  nnd2s1 ___9___446669(.DIN1 (________22288), .DIN2 (________23219), .Q
       (_____9__22789));
  hi1s1 _____9_446670(.DIN (________22787), .Q (________22788));
  nor2s1 ______446671(.DIN1 (________22817), .DIN2 (________23831), .Q
       (________22786));
  or2s1 _______446672(.DIN1 (___9_9__23395), .DIN2 (___0____23452), .Q
       (________22785));
  nnd2s1 _______446673(.DIN1 (_____9__22753), .DIN2 (________22783), .Q
       (________22784));
  and2s1 _______446674(.DIN1 (________22781), .DIN2 (________22776), .Q
       (________22782));
  hi1s1 ___9__446675(.DIN (_____9__22779), .Q (_____0__22780));
  and2s1 _______446676(.DIN1 (________22777), .DIN2 (________22776), .Q
       (________22778));
  and2s1 _____0_446677(.DIN1 (___0_____27897), .DIN2 (________22773),
       .Q (________22774));
  and2s1 _______446678(.DIN1 (________22770), .DIN2 (________22769), .Q
       (_____9__22771));
  nnd2s1 _______446679(.DIN1 (________22283), .DIN2 (________22766), .Q
       (________22767));
  or2s1 _______446680(.DIN1 (________23824), .DIN2 (_____9__22763), .Q
       (_____0__22764));
  or2s1 _______446681(.DIN1 (________22958), .DIN2 (_____9__22299), .Q
       (________22762));
  nor2s1 ___9___446682(.DIN1 (___0____21679), .DIN2 (________22760), .Q
       (________22761));
  nor2s1 ______446683(.DIN1 (___0___18987), .DIN2 (________22758), .Q
       (________22759));
  nor2s1 ______446684(.DIN1 (_____0___29362), .DIN2 (________22676), .Q
       (________22757));
  nnd2s1 _____9_446685(.DIN1 (________22755), .DIN2 (____9___22351), .Q
       (________22756));
  nnd2s1 _____9_446686(.DIN1 (_____9__22753), .DIN2 (____0___21814), .Q
       (_____0__22754));
  nnd2s1 ___9___446687(.DIN1 (____0_9__32819), .DIN2 (________19319),
       .Q (________22752));
  and2s1 ___9___446688(.DIN1 (_________31464), .DIN2 (______9__30169),
       .Q (________22751));
  nor2s1 ___9__446689(.DIN1 (________22183), .DIN2 (_____9__22199), .Q
       (________22750));
  and2s1 ___9_0_446690(.DIN1 (________22748), .DIN2 (________22237), .Q
       (________22749));
  and2s1 ___9_0_446691(.DIN1 (___0____24386), .DIN2 (_____0__22014), .Q
       (________22747));
  nnd2s1 ___9_0_446692(.DIN1 (________22692), .DIN2 (________22745), .Q
       (________22746));
  or2s1 ___9_9_446693(.DIN1 (____0___22178), .DIN2 (_____9__22743), .Q
       (_____0__22744));
  nnd2s1 ___9_446694(.DIN1 (________22741), .DIN2 (___0____22585), .Q
       (________22742));
  nnd2s1 ___9__446695(.DIN1 (________22739), .DIN2 (___0____22611), .Q
       (________22740));
  nor2s1 ___9___446696(.DIN1 (inData[18]), .DIN2 (________22737), .Q
       (________22738));
  nor2s1 ___9___446697(.DIN1 (________24749), .DIN2 (_____0__22182), .Q
       (________22736));
  nnd2s1 ___9___446698(.DIN1 (_____0__22734), .DIN2 (____09__22634), .Q
       (________22735));
  nnd2s1 ___9___446699(.DIN1 (____9___22168), .DIN2 (________22663), .Q
       (_____9__22733));
  nor2s1 ___9___446700(.DIN1 (inData[17]), .DIN2 (________22737), .Q
       (________22732));
  or2s1 ___9___446701(.DIN1 (________22730), .DIN2 (___9_9__23422), .Q
       (________22731));
  or2s1 ___9___446702(.DIN1 (_____9__22062), .DIN2 (________22245), .Q
       (________22729));
  nnd2s1 ___9___446703(.DIN1 (________22727), .DIN2 (________23757), .Q
       (________22728));
  nnd2s1 ___9___446704(.DIN1 (____0_9__32819), .DIN2 (_________29646),
       .Q (________22726));
  and2s1 ___9___446705(.DIN1 (________22190), .DIN2
       (______________________18672), .Q (_____0__22725));
  and2s1 ___9___446706(.DIN1 (________23906), .DIN2 (_________34486),
       .Q (____09__22724));
  hi1s1 ___9_9_446707(.DIN
       (______________0______________________18826), .Q
       (____0___22723));
  hi1s1 ___9_9_446708(.DIN (___0_0___27659), .Q (____0___22722));
  xnr2s1 ___9_446709(.DIN1 (_________________18774), .DIN2
       (_________35012), .Q (____0___22720));
  xor2s1 ___9___446710(.DIN1 (_________34445), .DIN2 (_________35012),
       .Q (____0___22719));
  xor2s1 ____9__446711(.DIN1 (________19237), .DIN2 (_________35002),
       .Q (____00__22718));
  xor2s1 ____9__446712(.DIN1 (________20580), .DIN2 (_________35002),
       .Q (____99__22717));
  xor2s1 ____9__446713(.DIN1 (________20583), .DIN2 (_________35002),
       .Q (____9___22716));
  nnd2s1 ____99_446714(.DIN1 (________22273), .DIN2 (________22274), .Q
       (____9___22715));
  and2s1 ____446715(.DIN1 (________25451), .DIN2 (_________35056), .Q
       (____9___22714));
  nor2s1 ___90__446716(.DIN1 (____0___22267), .DIN2 (____9___22712), .Q
       (____9___22713));
  nnd2s1 ___90_446717(.DIN1 (_____9__25634), .DIN2 (_____90__35018), .Q
       (____9___22711));
  nnd2s1 ___90_446718(.DIN1 (___009__22544), .DIN2 (________21799), .Q
       (____9___22710));
  nnd2s1 ___90__446719(.DIN1 (_____9__25634), .DIN2 (________22665), .Q
       (____90__22709));
  nor2s1 ___90__446720(.DIN1 (_________35000), .DIN2 (____9___22442),
       .Q (_____9__22708));
  and2s1 ___90_446721(.DIN1 (___9____25195), .DIN2 (________22706), .Q
       (________22707));
  nor2s1 ___90_446722(.DIN1 (________22704), .DIN2 (________23050), .Q
       (________22705));
  nor2s1 ___90__446723(.DIN1 (________22218), .DIN2 (___9____23407), .Q
       (________22703));
  nor2s1 ___909_446724(.DIN1 (__9_____26632), .DIN2 (________22284), .Q
       (________22702));
  nor2s1 ___90__446725(.DIN1 (____00__19399), .DIN2 (________22317), .Q
       (________22701));
  nnd2s1 ___9___446726(.DIN1 (____00__22261), .DIN2 (________23875), .Q
       (________23330));
  nnd2s1 ___9___446727(.DIN1 (_____9__22408), .DIN2 (_________35006),
       .Q (___9____23381));
  nor2s1 ___9___446728(.DIN1 (________23284), .DIN2 (_____9__22763), .Q
       (________23587));
  nor2s1 ___9__446729(.DIN1 (_____0__22700), .DIN2 (_____9__22699), .Q
       (_____9__22971));
  nnd2s1 ___9___446730(.DIN1 (________22188), .DIN2 (________22674), .Q
       (____0___23262));
  nnd2s1 ___9_0_446731(.DIN1 (________22367), .DIN2 (________25926), .Q
       (_____0__22833));
  nnd2s1 ___9_9_446732(.DIN1 (___0____22616), .DIN2 (________22698), .Q
       (________22834));
  or2s1 ___9_9_446733(.DIN1 (________22697), .DIN2 (________22696), .Q
       (____9___23257));
  or2s1 ___9___446734(.DIN1 (________22696), .DIN2 (________22695), .Q
       (________23247));
  and2s1 ___9___446735(.DIN1 (________22694), .DIN2 (____09__21728), .Q
       (____0____28183));
  nor2s1 ___9___446736(.DIN1 (___900__22446), .DIN2 (_____9__22669), .Q
       (_____0__23108));
  xor2s1 ___9__446737(.DIN1 (____9___19112), .DIN2 (_____0___32570), .Q
       (________22956));
  nnd2s1 ___9___446738(.DIN1 (____9___22350), .DIN2 (________22693), .Q
       (____9___23252));
  nnd2s1 ___9___446739(.DIN1 (________22692), .DIN2 (________22247), .Q
       (____9_0__32685));
  hi1s1 ___9___446740(.DIN (________22691), .Q (___0____23510));
  hi1s1 ___9___446741(.DIN (________22876), .Q (________23279));
  nnd2s1 ___9___446742(.DIN1 (____0___25752), .DIN2 (_____0__22690), .Q
       (________24100));
  and2s1 ___9___446743(.DIN1 (___0____21706), .DIN2 (________23063), .Q
       (____09__23267));
  hi1s1 ___9___446744(.DIN (_____9__22689), .Q (________23910));
  nor2s1 ___9_9_446745(.DIN1 (________22688), .DIN2 (________25401), .Q
       (________22972));
  hi1s1 ___9_446746(.DIN (__9_____26354), .Q (________23556));
  and2s1 ___9___446747(.DIN1 (________23738), .DIN2 (____0___21448), .Q
       (____99__23345));
  nnd2s1 _____0_446748(.DIN1 (________22303), .DIN2 (________22687), .Q
       (________22867));
  or2s1 _______446749(.DIN1 (________22686), .DIN2 (________24087), .Q
       (___9_0__23376));
  nor2s1 _______446750(.DIN1 (________22685), .DIN2 (________22305), .Q
       (_____0__23628));
  nnd2s1 _______446751(.DIN1 (_____9__22326), .DIN2 (_____0__23695), .Q
       (____0___23090));
  and2s1 _______446752(.DIN1 (____9___22443), .DIN2 (________25704), .Q
       (____0___23173));
  nor2s1 _______446753(.DIN1 (_____0__22300), .DIN2 (________26094), .Q
       (________23229));
  nor2s1 _______446754(.DIN1 (________22094), .DIN2 (____9___22166), .Q
       (____0___25656));
  nor2s1 ______446755(.DIN1 (________21889), .DIN2 (________22314), .Q
       (________22821));
  xor2s1 _______446756(.DIN1 (________22684), .DIN2 (_________33333),
       .Q (___90___23352));
  nor2s1 ___9_0_446757(.DIN1 (_____0__25694), .DIN2 (____9___22441), .Q
       (________24970));
  nor2s1 ___9___446758(.DIN1 (________21997), .DIN2 (________26081), .Q
       (________23327));
  nor2s1 ___9___446759(.DIN1 (_____0__24541), .DIN2 (________22338), .Q
       (________23332));
  nor2s1 ___9___446760(.DIN1 (________23757), .DIN2 (________22328), .Q
       (___0_9___27648));
  and2s1 _______446761(.DIN1 (_________34982), .DIN2 (________22682),
       .Q (________23234));
  nnd2s1 _______446762(.DIN1 (__9__0__26854), .DIN2 (_____0__22952), .Q
       (________23872));
  nnd2s1 ___9__446763(.DIN1 (________25451), .DIN2 (________22681), .Q
       (________25978));
  hi1s1 ___9___446764(.DIN (_____0__22680), .Q (____90__23965));
  nnd2s1 ____9__446765(.DIN1 (_____9__22309), .DIN2 (_____9__22679), .Q
       (_________29736));
  or2s1 ___9___446766(.DIN1 (________25478), .DIN2 (________24806), .Q
       (________24118));
  nnd2s1 ____90_446767(.DIN1 (__9__9__27014), .DIN2 (__9_____27021), .Q
       (________25963));
  or2s1 ____90_446768(.DIN1 (________21952), .DIN2 (__9_____26535), .Q
       (_________28775));
  nnd2s1 ___9___446769(.DIN1 (________22307), .DIN2 (_________35084),
       .Q (_________33325));
  nnd2s1 ____90_446770(.DIN1 (___9____25195), .DIN2 (________22678), .Q
       (________25881));
  or2s1 ___9___446771(.DIN1 (________22279), .DIN2 (___0_9___27848), .Q
       (__9_9___26698));
  or2s1 ____446772(.DIN1 (________22675), .DIN2 (__9_____27037), .Q
       (________25831));
  nnd2s1 ____446773(.DIN1 (_____0__22281), .DIN2 (________22677), .Q
       (__9_____26647));
  or2s1 ___9___446774(.DIN1 (___0____22591), .DIN2 (________23045), .Q
       (__990___27088));
  hi1s1 ___9___446775(.DIN (_________33444), .Q (_____99__31353));
  nnd2s1 ____9__446776(.DIN1 (_____0__23231), .DIN2 (__9_____26406), .Q
       (____9___25945));
  nnd2s1 ___9__446777(.DIN1 (____0_9__32819), .DIN2 (________22676), .Q
       (_________32874));
  nnd2s1 ____9__446778(.DIN1 (________25798), .DIN2 (________25447), .Q
       (________26072));
  or2s1 ____9__446779(.DIN1 (________25722), .DIN2 (________22675), .Q
       (__9__0__26485));
  hi1s1 ___9_0_446780(.DIN (____0____31829), .Q (_________32925));
  nnd2s1 ___9___446781(.DIN1 (________22313), .DIN2 (________21733), .Q
       (__9_____27027));
  nnd2s1 ____9__446782(.DIN1 (________22298), .DIN2 (_____0__20079), .Q
       (_________33385));
  nnd2s1 ____9__446783(.DIN1 (________22308), .DIN2 (________22333), .Q
       (____000__32751));
  hi1s1 ___9___446784(.DIN (____9___22890), .Q (_____9__23275));
  nnd2s1 ____9_446785(.DIN1 (________22306), .DIN2 (________20390), .Q
       (____9_9__31781));
  nnd2s1 ____9__446786(.DIN1 (________22184), .DIN2 (________22674), .Q
       (__9_____26675));
  hi1s1 ___9___446787(.DIN (________22673), .Q (___00____27202));
  nnd2s1 ____9__446788(.DIN1 (_____0__22157), .DIN2 (________22672), .Q
       (______0__33918));
  nnd2s1 ____9__446789(.DIN1 (________22155), .DIN2 (________22672), .Q
       (______0__33336));
  nor2s1 ___9___446790(.DIN1 (_____0__22670), .DIN2 (_____9__22669), .Q
       (________22671));
  hi1s1 ___9_0_446791(.DIN (________23596), .Q (________22668));
  nnd2s1 ___9__446792(.DIN1 (____0_9__32819), .DIN2 (____0___20228), .Q
       (________22667));
  and2s1 ___9___446793(.DIN1 (________22665), .DIN2 (_____0__24551), .Q
       (________22666));
  nnd2s1 ___9___446794(.DIN1 (____9___22256), .DIN2 (________22663), .Q
       (________22664));
  nor2s1 ___9_0_446795(.DIN1 (___0____23512), .DIN2 (__9_____26764), .Q
       (________22662));
  hi1s1 ___9___446796(.DIN (________22659), .Q (________22660));
  hi1s1 ___9___446797(.DIN (________22657), .Q (________22658));
  nnd2s1 _____446798(.DIN1 (___0_0__24382), .DIN2 (____0___22269), .Q
       (________22656));
  hi1s1 ___99__446799(.DIN (_____9__24655), .Q (________22655));
  and2s1 ___9___446800(.DIN1 (___00___23444), .DIN2 (_____0__22653), .Q
       (________22654));
  or2s1 ___9__446801(.DIN1 (___09___24420), .DIN2 (________22638), .Q
       (_____9__22652));
  and2s1 ___9___446802(.DIN1 (_____0___32572), .DIN2 (________19080),
       .Q (________22651));
  nor2s1 ___9___446803(.DIN1 (______9__28887), .DIN2 (________22648),
       .Q (________22650));
  nor2s1 ___9___446804(.DIN1 (_________30710), .DIN2 (________22648),
       .Q (________22649));
  or2s1 ___9_9_446805(.DIN1 (________23757), .DIN2 (________26020), .Q
       (________22647));
  nnd2s1 ___9_9_446806(.DIN1 (_________34986), .DIN2 (________24221),
       .Q (________22646));
  or2s1 ___9_446807(.DIN1 (________19570), .DIN2 (________26020), .Q
       (________22645));
  nor2s1 ___9_0_446808(.DIN1 (___0____23448), .DIN2 (___0____22593), .Q
       (_____0__22644));
  nnd2s1 ___9___446809(.DIN1 (____00__23528), .DIN2 (____0___19400), .Q
       (_____9__22643));
  nor2s1 ___9___446810(.DIN1 (________25437), .DIN2 (________22202), .Q
       (________22642));
  or2s1 ___9___446811(.DIN1 (________22639), .DIN2 (________22638), .Q
       (________22640));
  nor2s1 ___9___446812(.DIN1 (_________35062), .DIN2 (__99_9__27116),
       .Q (________22637));
  nnd2s1 ___9___446813(.DIN1 (________22193), .DIN2 (______9__32927),
       .Q (________22636));
  or2s1 ___9___446814(.DIN1 (____09__22634), .DIN2 (___00___23444), .Q
       (_____0__22635));
  and2s1 ___9___446815(.DIN1 (________23692), .DIN2 (____0___19500), .Q
       (____0___22633));
  nor2s1 ___9___446816(.DIN1 (________22686), .DIN2 (___0____22612), .Q
       (____0___22632));
  nor2s1 ___9___446817(.DIN1 (________19074), .DIN2 (_____9__22797), .Q
       (____0___22631));
  nnd2s1 ___9__446818(.DIN1 (____0___22177), .DIN2 (____9___22886), .Q
       (____0___22629));
  or2s1 ___9___446819(.DIN1 (____9___19395), .DIN2 (__9__9__27043), .Q
       (____0___22628));
  or2s1 ___9___446820(.DIN1 (____0____29098), .DIN2 (________22692), .Q
       (____0___22627));
  or2s1 ___9___446821(.DIN1 (___099__22625), .DIN2 (________22641), .Q
       (____00__22626));
  nor2s1 ___9__446822(.DIN1 (__9_____26764), .DIN2 (___09___22623), .Q
       (___09___22624));
  nor2s1 ___9___446823(.DIN1 (____9___19945), .DIN2 (___00___23444), .Q
       (___09___22622));
  and2s1 ___9___446824(.DIN1 (___09___22620), .DIN2 (________19126), .Q
       (___09___22621));
  nnd2s1 ___9___446825(.DIN1 (___09___22620), .DIN2 (_____0__19331), .Q
       (___09___22619));
  or2s1 ___9___446826(.DIN1 (________23814), .DIN2 (___090__22617), .Q
       (___09___22618));
  nnd2s1 ___9___446827(.DIN1 (___0_____27862), .DIN2 (_____0__23811),
       .Q (________22822));
  nnd2s1 ___0___446828(.DIN1 (__9_____26445), .DIN2 (___0____22616), .Q
       (________23111));
  hi1s1 ___9_9_446829(.DIN (___0____22615), .Q (____9___23254));
  nnd2s1 ___9___446830(.DIN1 (__9_____26372), .DIN2 (________25392), .Q
       (________23997));
  hi1s1 ___9__446831(.DIN (________22959), .Q (________23277));
  nnd2s1 ___9___446832(.DIN1 (________22197), .DIN2 (________22316), .Q
       (________22831));
  nnd2s1 ___0___446833(.DIN1 (________22161), .DIN2 (inData[10]), .Q
       (________23212));
  nnd2s1 ___9___446834(.DIN1 (___0_0__22582), .DIN2 (________22433), .Q
       (____0___22810));
  hi1s1 ___9___446835(.DIN (___0____22614), .Q (____0___23888));
  hi1s1 ___9___446836(.DIN (___0____22613), .Q (________23126));
  hi1s1 ___9___446837(.DIN (__9_____26736), .Q (________23098));
  nor2s1 ___9___446838(.DIN1 (_____9___35024), .DIN2 (___0____22612),
       .Q (________23944));
  and2s1 ___9___446839(.DIN1 (___0____22611), .DIN2 (________25726), .Q
       (____9___23164));
  nor2s1 ___9__446840(.DIN1 (________22153), .DIN2 (__9_____26953), .Q
       (____0___23176));
  nnd2s1 ___9___446841(.DIN1 (___00____27220), .DIN2 (___0____22610),
       .Q (________23752));
  nor2s1 ___9___446842(.DIN1 (________23154), .DIN2 (___0_____27862),
       .Q (________23105));
  and2s1 ___9___446843(.DIN1 (________21735), .DIN2 (____0___25752), .Q
       (________23270));
  nor2s1 ___9___446844(.DIN1 (___0____22609), .DIN2 (___9____24313), .Q
       (____90__23250));
  nnd2s1 ___9_9_446845(.DIN1 (________22938), .DIN2 (________22776), .Q
       (________23132));
  nnd2s1 ___9_9_446846(.DIN1 (___0____22604), .DIN2 (________22226), .Q
       (________23204));
  xnr2s1 ___9_446847(.DIN1 (______0__35008), .DIN2 (_____9__19095), .Q
       (________23095));
  nor2s1 ___9_0_446848(.DIN1 (_____9__21513), .DIN2 (____9___22252), .Q
       (________23192));
  nnd2s1 ___9_0_446849(.DIN1 (___0____23484), .DIN2 (___0_0__22608), .Q
       (_____0__23152));
  or2s1 ___9___446850(.DIN1 (__9_____26472), .DIN2 (____9___22255), .Q
       (________24200));
  nor2s1 ___9___446851(.DIN1 (________25913), .DIN2 (____00__22172), .Q
       (________23244));
  and2s1 ___9___446852(.DIN1 (____9___21899), .DIN2 (___0____22607), .Q
       (________23102));
  nor2s1 ___9__446853(.DIN1 (________23104), .DIN2 (___0____22606), .Q
       (________22852));
  nnd2s1 ___9___446854(.DIN1 (___0____22605), .DIN2 (________23154), .Q
       (________23130));
  and2s1 ___9__446855(.DIN1 (__9_____26877), .DIN2 (_____0__25770), .Q
       (___0____23469));
  nnd2s1 ___9_0_446856(.DIN1 (___00___23444), .DIN2 (___0____21672), .Q
       (________23195));
  or2s1 ___9___446857(.DIN1 (____9___25458), .DIN2 (____9___22164), .Q
       (________23927));
  nnd2s1 ___9___446858(.DIN1 (___0____22605), .DIN2 (_____0__23199), .Q
       (_____9__23107));
  and2s1 ___9___446859(.DIN1 (___0____22604), .DIN2 (______0__34998),
       .Q (____9___23615));
  nnd2s1 ___99__446860(.DIN1 (________22198), .DIN2 (________22131), .Q
       (________22949));
  nor2s1 _______446861(.DIN1 (___0____22603), .DIN2 (________22277), .Q
       (____9___24154));
  nnd2s1 ___9___446862(.DIN1 (________22737), .DIN2 (___0____22602), .Q
       (____0___25758));
  nnd2s1 ___9__446863(.DIN1 (________22323), .DIN2 (___0____22601), .Q
       (_____0__25712));
  or2s1 ___9___446864(.DIN1 (_____0__25967), .DIN2 (___0____22612), .Q
       (_____0__26127));
  or2s1 ___9___446865(.DIN1 (________23908), .DIN2 (___0_0__22600), .Q
       (________25772));
  nnd2s1 ___9___446866(.DIN1 (________22250), .DIN2 (________22110), .Q
       (__9_____26677));
  or2s1 ___9___446867(.DIN1 (____9___23255), .DIN2 (___0_9__22599), .Q
       (____9___23709));
  nnd2s1 ___9_446868(.DIN1 (__9_____26406), .DIN2 (________22238), .Q
       (________24644));
  nnd2s1 ___9_9_446869(.DIN1 (__9_____27045), .DIN2 (________25980), .Q
       (___0_0___27272));
  nnd2s1 ___9_9_446870(.DIN1 (_____0___32572), .DIN2 (_________32487),
       .Q (_____0___32574));
  xor2s1 ___990_446871(.DIN1 (___00), .DIN2 (______0__35008), .Q
       (_____9___31345));
  nnd2s1 ___9___446872(.DIN1 (________23097), .DIN2 (________22235), .Q
       (___9_0__24316));
  nor2s1 ___9___446873(.DIN1 (________23193), .DIN2 (________22287), .Q
       (________25627));
  nor2s1 _______446874(.DIN1 (________22227), .DIN2 (________22304), .Q
       (___909__23355));
  and2s1 ___9___446875(.DIN1 (__9__9__26540), .DIN2 (___0____22598), .Q
       (____0___25754));
  and2s1 ___9___446876(.DIN1 (____9___24605), .DIN2
       (_____________________18664), .Q (_____9__23302));
  nnd2s1 ___9___446877(.DIN1 (___0_____27862), .DIN2 (___9____22496),
       .Q (________23200));
  nor2s1 ___9___446878(.DIN1 (___0____22597), .DIN2 (________22371), .Q
       (________24712));
  nor2s1 ___9___446879(.DIN1 (___0____22605), .DIN2 (___0____22596), .Q
       (________23307));
  and2s1 ___9__446880(.DIN1 (___0____22595), .DIN2 (__9_____26358), .Q
       (___99___25268));
  nnd2s1 ___9___446881(.DIN1 (____0_9__32819), .DIN2 (___0____22594),
       .Q (____0_0__32780));
  nnd2s1 ___9__446882(.DIN1 (_________35006), .DIN2 (____9___22258), .Q
       (________24024));
  nor2s1 ___9___446883(.DIN1 (____9___21981), .DIN2 (___0____22606), .Q
       (________24777));
  nnd2s1 ___0___446884(.DIN1 (___0____22616), .DIN2 (__9_____26496), .Q
       (________23857));
  nnd2s1 ___9__446885(.DIN1 (___0____22593), .DIN2 (___99___22532), .Q
       (________23562));
  nor2s1 ___9___446886(.DIN1 (__9_____26905), .DIN2 (________24079), .Q
       (___0____25288));
  or2s1 ___9___446887(.DIN1 (________23814), .DIN2 (__9__9__27043), .Q
       (___0_____27998));
  nor2s1 ___99_446888(.DIN1 (________22334), .DIN2 (___0____22584), .Q
       (____99__23170));
  or2s1 ___99__446889(.DIN1 (___0____22592), .DIN2 (___0____22591), .Q
       (___9_0__25231));
  nor2s1 ___99__446890(.DIN1 (_____0___35034), .DIN2 (___0_9__22599),
       .Q (________24230));
  nor2s1 ___99__446891(.DIN1 (________25531), .DIN2 (________22115), .Q
       (_____9__24198));
  hi1s1 ___00__446892(.DIN (__90____26312), .Q (__9_____26576));
  nnd2s1 ___99__446893(.DIN1 (___0____22588), .DIN2 (________22938), .Q
       (__9__0__26637));
  or2s1 ___99__446894(.DIN1 (________23238), .DIN2 (____9___25943), .Q
       (____0___26055));
  or2s1 ___99__446895(.DIN1 (_____9___35022), .DIN2 (___9_9__23422), .Q
       (________23288));
  nor2s1 ___99_446896(.DIN1 (_____0___35032), .DIN2 (________22324), .Q
       (________24804));
  and2s1 ___99__446897(.DIN1 (__9_9___26604), .DIN2 (________25419), .Q
       (________24830));
  nnd2s1 ___9__446898(.DIN1 (____90__22436), .DIN2 (___0____22583), .Q
       (____0___23178));
  hi1s1 ___9_0_446899(.DIN (________23033), .Q (________23227));
  nnd2s1 ___99__446900(.DIN1 (__9_____27045), .DIN2 (____00__21075), .Q
       (_____9___28517));
  nnd2s1 ___99__446901(.DIN1 (_________31464), .DIN2 (___0____22590),
       .Q (_____9___31443));
  nnd2s1 ___99__446902(.DIN1 (___0_0___27563), .DIN2 (___0____22586),
       .Q (____9___25746));
  nor2s1 ___9___446903(.DIN1 (___0____22589), .DIN2 (________22727), .Q
       (___90___25180));
  and2s1 ___9__446904(.DIN1 (___0____22588), .DIN2 (________23005), .Q
       (____99__25654));
  nnd2s1 ___9___446905(.DIN1 (________22368), .DIN2 (___0_____27600),
       .Q (__9_9___26505));
  nnd2s1 ___9___446906(.DIN1 (___0____22587), .DIN2 (____00__24701), .Q
       (________23248));
  nnd2s1 ___99_446907(.DIN1 (_____0__22653), .DIN2 (________22706), .Q
       (___9____25198));
  nnd2s1 ___9___446908(.DIN1 (___0____22586), .DIN2 (________22766), .Q
       (____9___23342));
  nnd2s1 ___99__446909(.DIN1 (________24195), .DIN2 (___0____22585), .Q
       (____9___26142));
  nor2s1 ___99__446910(.DIN1 (____0________________18591), .DIN2
       (_________34984), .Q (___90___23347));
  nnd2s1 ___9_0_446911(.DIN1 (___0____22584), .DIN2 (___0____22583), .Q
       (________23137));
  hi1s1 ___9___446912(.DIN (___09___23520), .Q (__99____27091));
  hi1s1 ___9___446913(.DIN (_____9__22961), .Q (________23156));
  hi1s1 ___00__446914(.DIN (___0_9__22581), .Q (___00____27211));
  nor2s1 ___9_9_446915(.DIN1 (________22112), .DIN2 (________22236), .Q
       (___999__26246));
  nor2s1 ___99__446916(.DIN1 (________22331), .DIN2 (___0_0__22582), .Q
       (_____0__23286));
  nor2s1 ___9_0_446917(.DIN1 (____00__23528), .DIN2 (________24833), .Q
       (___0__0__27609));
  hi1s1 ___9___446918(.DIN (________22909), .Q (____0___23266));
  nor2s1 ___99__446919(.DIN1 (________22330), .DIN2 (___0_0__22582), .Q
       (________23202));
  nor2s1 ___9___446920(.DIN1 (________22432), .DIN2 (___0_0__22582), .Q
       (_____0__23241));
  nnd2s1 ___99__446921(.DIN1 (_____9__22191), .DIN2 (____9___19940), .Q
       (_____9___33026));
  hi1s1 ___00__446922(.DIN (__9_____26962), .Q (__9_____26621));
  nnd2s1 ___99__446923(.DIN1 (_____9__22797), .DIN2 (________21871), .Q
       (____9____32723));
  hi1s1 ___00_446924(.DIN (__9__0__27005), .Q (__990___27084));
  nor2s1 ___9__446925(.DIN1 (____9___22437), .DIN2 (___0____22584), .Q
       (________23862));
  hi1s1 ___00_446926(.DIN (__9_____27061), .Q (___0__9__27771));
  hi1s1 ___9__446927(.DIN (________22941), .Q (________23578));
  hi1s1 ___00__446928(.DIN (___0_____27386), .Q (_____0___28805));
  nnd2s1 ___9___446929(.DIN1 (___0____22579), .DIN2 (____0___19400), .Q
       (___0____22580));
  nor2s1 ___9___446930(.DIN1 (_____0__22099), .DIN2 (___0____22577), .Q
       (___0____22578));
  and2s1 ___9___446931(.DIN1 (___9____22482), .DIN2 (________24001), .Q
       (___0____22576));
  nnd2s1 ___9___446932(.DIN1 (____9___22076), .DIN2 (____9___19945), .Q
       (___0____22575));
  and2s1 ___9__446933(.DIN1 (___0_0__22573), .DIN2 (________23814), .Q
       (___0____22574));
  and2s1 ___9___446934(.DIN1 (___0____22571), .DIN2 (________23757), .Q
       (___0_9__22572));
  nor2s1 ___9_0_446935(.DIN1 (____00__19399), .DIN2 (____9___22079), .Q
       (___0____22570));
  nnd2s1 ___9_0_446936(.DIN1 (___0____22579), .DIN2 (___00___22540), .Q
       (___0____22569));
  nnd2s1 ___9_0_446937(.DIN1 (___0____22567), .DIN2 (___00___22540), .Q
       (___0____22568));
  nor2s1 ___9___446938(.DIN1 (___0____22565), .DIN2 (___0_0__25290), .Q
       (___0____22566));
  or2s1 ___9_0_446939(.DIN1 (___0_9__22563), .DIN2 (____0___24065), .Q
       (___0_0__22564));
  nor2s1 ___9___446940(.DIN1 (________22058), .DIN2 (________21966), .Q
       (___0____22562));
  nnd2s1 ___9__446941(.DIN1 (________22040), .DIN2 (________19376), .Q
       (___0____22561));
  nor2s1 ___9__446942(.DIN1 (____0___22813), .DIN2 (___0____22559), .Q
       (___0____22560));
  or2s1 ______446943(.DIN1 (____0___23716), .DIN2 (________22777), .Q
       (___0____22558));
  nnd2s1 ______446944(.DIN1 (________22092), .DIN2 (___0_0__23500), .Q
       (___0____22557));
  nnd2s1 ___9___446945(.DIN1 (________22104), .DIN2 (________20272), .Q
       (___0____22556));
  and2s1 ___9_0_446946(.DIN1 (___0_0__22554), .DIN2 (___9____22460), .Q
       (___0____22555));
  and2s1 ___9_446947(.DIN1 (________22101), .DIN2 (___0____22552), .Q
       (___0_9__22553));
  and2s1 ____9__446948(.DIN1 (________21943), .DIN2 (_________29873),
       .Q (___0____22551));
  xnr2s1 ___9___446949(.DIN1 (___0____22549), .DIN2 (______0__31325),
       .Q (___0____22550));
  xor2s1 ___9___446950(.DIN1 (___0____22547), .DIN2 (___0____22546), .Q
       (___0____22548));
  nor2s1 ___9_9_446951(.DIN1 (________25872), .DIN2 (____0___22811), .Q
       (___0____22545));
  hi1s1 ___9_9_446952(.DIN (__9_____26840), .Q (___00___22542));
  nnd2s1 ___9__446953(.DIN1 (___9____23367), .DIN2 (___00___22540), .Q
       (___00___22541));
  and2s1 ___9___446954(.DIN1 (___00___22538), .DIN2 (_________35072),
       .Q (___00___22539));
  nnd2s1 ___9___446955(.DIN1 (________22049), .DIN2 (inData[10]), .Q
       (___00___22537));
  nnd2s1 ___9___446956(.DIN1 (________22007), .DIN2 (inData[4]), .Q
       (___000__22536));
  nor2s1 ___9___446957(.DIN1 (___0____21647), .DIN2 (________22064), .Q
       (___999__22535));
  nnd2s1 ___9___446958(.DIN1 (___99___22533), .DIN2 (___99___22532), .Q
       (___99___22534));
  nor2s1 ___9___446959(.DIN1 (_____0__19187), .DIN2 (________21964), .Q
       (___99___22531));
  nnd2s1 ___9__446960(.DIN1 (___99___22529), .DIN2 (___99___19768), .Q
       (___99___22530));
  and2s1 ___9__446961(.DIN1 (________22683), .DIN2 (___99___22527), .Q
       (___99___22528));
  nnd2s1 ___9___446962(.DIN1 (___9____22457), .DIN2 (____9___19395), .Q
       (___990__22526));
  nnd2s1 ___9___446963(.DIN1 (________22057), .DIN2 (___9____22524), .Q
       (___9____22525));
  nor2s1 ___9___446964(.DIN1 (________23318), .DIN2 (___9____22522), .Q
       (___9____22523));
  nnd2s1 ___9___446965(.DIN1 (___9____23396), .DIN2 (________22948), .Q
       (___9____22521));
  nor2s1 ___9___446966(.DIN1 (____9___19945), .DIN2 (___90___22449), .Q
       (___9____22520));
  nnd2s1 ___9___446967(.DIN1 (________21953), .DIN2 (________21847), .Q
       (___9____22519));
  and2s1 ___9__446968(.DIN1 (___9_0__22517), .DIN2 (______0__34998), .Q
       (___9____22518));
  nnd2s1 ___9__446969(.DIN1 (______0__34998), .DIN2 (________22145), .Q
       (___9_9__22516));
  nor2s1 ___9___446970(.DIN1 (________22434), .DIN2 (_____0__22005), .Q
       (___9____22515));
  nor2s1 ___9___446971(.DIN1 (____09__19861), .DIN2 (_____9__22013), .Q
       (___9____22514));
  nnd2s1 ___9__446972(.DIN1 (___9____22503), .DIN2 (________21791), .Q
       (___9____22513));
  and2s1 ___9___446973(.DIN1 (____9___22077), .DIN2 (_____9__21139), .Q
       (___9____22512));
  or2s1 ___9__446974(.DIN1 (___9____22510), .DIN2 (___9_0__22491), .Q
       (___9____22511));
  nor2s1 ___9__446975(.DIN1 (_____0__19225), .DIN2 (_________34996), .Q
       (___9____22509));
  nor2s1 ___9___446976(.DIN1 (_____9__19379), .DIN2 (_________34996),
       .Q (___9_0__22508));
  nnd2s1 ___9___446977(.DIN1 (___9____22506), .DIN2 (___9____22505), .Q
       (___9_9__22507));
  nnd2s1 ___9___446978(.DIN1 (________24774), .DIN2 (___9____22503), .Q
       (___9____22504));
  and2s1 ___9___446979(.DIN1 (________22046), .DIN2 (_________35084),
       .Q (___9____22502));
  nor2s1 ___9_9_446980(.DIN1 (___9____24277), .DIN2 (___9____24263), .Q
       (___9____22501));
  nor2s1 ___9_0_446981(.DIN1 (________21306), .DIN2 (_____9__22032), .Q
       (___9_9__22499));
  or2s1 ___9___446982(.DIN1 (____9___19395), .DIN2 (___9____22487), .Q
       (___9____22498));
  and2s1 ___9___446983(.DIN1 (___9____22496), .DIN2 (___9____22495), .Q
       (___9____22497));
  nnd2s1 ___9___446984(.DIN1 (________22003), .DIN2 (________22187), .Q
       (___9____22494));
  nor2s1 ___9___446985(.DIN1 (___9____22492), .DIN2 (___9_0__22491), .Q
       (___9____22493));
  nor2s1 ___9___446986(.DIN1 (____________0___18786), .DIN2
       (_________33442), .Q (___9_9__22490));
  nnd2s1 ___9___446987(.DIN1 (________21945), .DIN2 (___0____20763), .Q
       (___9____22489));
  nnd2s1 ___9___446988(.DIN1 (___9____22487), .DIN2 (___9_9__22464), .Q
       (___9____22488));
  nnd2s1 ___9___446989(.DIN1 (________24113), .DIN2 (_____0__23695), .Q
       (___9____22486));
  nor2s1 ___9___446990(.DIN1 (_____9__25684), .DIN2 (________22162), .Q
       (___9____22485));
  or2s1 ___9___446991(.DIN1 (_________34393), .DIN2 (________22009), .Q
       (___9____22484));
  nnd2s1 ___9___446992(.DIN1 (___9____22482), .DIN2 (________22693), .Q
       (___9____22483));
  nnd2s1 ___9__446993(.DIN1 (_____9___28891), .DIN2 (________21827), .Q
       (___9_0__22481));
  nnd2s1 ___9___446994(.DIN1 (___9____22487), .DIN2 (________22370), .Q
       (___9_9__22480));
  and2s1 ___9___446995(.DIN1 (___9____22478), .DIN2 (_________29330),
       .Q (___9____22479));
  nor2s1 ___9___446996(.DIN1 (______0__35058), .DIN2 (________22204),
       .Q (___9____22477));
  nor2s1 ___9___446997(.DIN1 (_________29330), .DIN2 (___9____22478),
       .Q (___9____22476));
  nor2s1 ___9__446998(.DIN1 (___9_0__26157), .DIN2 (___0____22577), .Q
       (___9____22475));
  nnd2s1 ___9___446999(.DIN1 (________22321), .DIN2 (________21390), .Q
       (___9____22474));
  nor2s1 ___9___447000(.DIN1 (___9_0__22472), .DIN2 (________22205), .Q
       (___9____22473));
  nor2s1 ___9___447001(.DIN1 (________22688), .DIN2 (___9____22470), .Q
       (___9____22471));
  or2s1 ___9___447002(.DIN1 (_____0__25967), .DIN2 (________22020), .Q
       (___9____22468));
  or2s1 ___9___447003(.DIN1 (_____9__25684), .DIN2 (______0__28551), .Q
       (___9____22467));
  nnd2s1 _______447004(.DIN1 (___9_0__22455), .DIN2 (___9____24300), .Q
       (________22870));
  nnd2s1 ___9___447005(.DIN1 (___9_0__22465), .DIN2 (____9___22886), .Q
       (________22775));
  nnd2s1 ___9___447006(.DIN1 (____0___22083), .DIN2 (________21461), .Q
       (________22964));
  nnd2s1 ___9___447007(.DIN1 (_____0__22053), .DIN2 (___9____19711), .Q
       (_____9__23230));
  and2s1 ___9_9_447008(.DIN1 (________22010), .DIN2 (__9_____26717), .Q
       (___009__25280));
  nnd2s1 ___9_9_447009(.DIN1 (________22055), .DIN2 (____9___23707), .Q
       (________23036));
  nnd2s1 ___9_447010(.DIN1 (___9_9__22464), .DIN2 (___9____22463), .Q
       (_____9__22951));
  nnd2s1 ___9_447011(.DIN1 (___9____22462), .DIN2 (___9____22461), .Q
       (________22659));
  and2s1 ___9_0_447012(.DIN1 (________22698), .DIN2 (__9_0___26517), .Q
       (________23243));
  and2s1 ___9_0_447013(.DIN1 (___9_0__26177), .DIN2 (________24459), .Q
       (________23840));
  and2s1 ___9_0_447014(.DIN1 (________22739), .DIN2 (___9____22460), .Q
       (____09__22904));
  nnd2s1 ___9_447015(.DIN1 (________22683), .DIN2 (___0____23448), .Q
       (________24627));
  nnd2s1 ___9__447016(.DIN1 (____99__22445), .DIN2 (________22292), .Q
       (____0___22721));
  nor2s1 ___9___447017(.DIN1 (___9____22459), .DIN2 (________25442), .Q
       (_____9__22779));
  nor2s1 ___9___447018(.DIN1 (___9____22458), .DIN2 (________24549), .Q
       (_____9__25606));
  nor2s1 ___9___447019(.DIN1 (____99__22894), .DIN2 (___9____22457), .Q
       (________23026));
  hi1s1 ___9___447020(.DIN (___9____22456), .Q (___9____23411));
  nnd2s1 _____0_447021(.DIN1 (___9_0__22455), .DIN2 (__________), .Q
       (________22787));
  nnd2s1 _____0_447022(.DIN1 (________22096), .DIN2 (________22061), .Q
       (________23552));
  nnd2s1 ___9___447023(.DIN1 (________22105), .DIN2
       (__________________0___18670), .Q (_____9__22689));
  nor2s1 ___9___447024(.DIN1 (____00__22356), .DIN2 (________24814), .Q
       (________23021));
  nor2s1 ___9__447025(.DIN1 (____9___25458), .DIN2 (_____0__22234), .Q
       (________22768));
  nnd2s1 ___9___447026(.DIN1 (________22019), .DIN2
       (_____________________18665), .Q (_____9__23017));
  nor2s1 ___9___447027(.DIN1 (________23239), .DIN2 (___9____24250), .Q
       (________22765));
  nnd2s1 ___9___447028(.DIN1 (________22027), .DIN2 (___909__22454), .Q
       (_____0__22772));
  nor2s1 ___9__447029(.DIN1 (____9___21440), .DIN2 (_________35000), .Q
       (________22849));
  nnd2s1 ___9___447030(.DIN1 (_____0__22033), .DIN2 (_____0__20382), .Q
       (________22673));
  nor2s1 ___9___447031(.DIN1 (___0____23512), .DIN2 (___90___22453), .Q
       (___0____22615));
  nor2s1 ___9___447032(.DIN1 (_____0__22670), .DIN2 (___9____22522), .Q
       (_____9__22980));
  nor2s1 ___9___447033(.DIN1 (__9_____26452), .DIN2 (___0____22559), .Q
       (_____0__24956));
  nor2s1 ___9__447034(.DIN1 (____9___21982), .DIN2 (___90___22452), .Q
       (____9___23075));
  nnd2s1 ___9___447035(.DIN1 (________24113), .DIN2 (________25380), .Q
       (___9____25186));
  nnd2s1 ___9___447036(.DIN1 (________24452), .DIN2 (___90___22451), .Q
       (________22950));
  nnd2s1 ___9___447037(.DIN1 (________22840), .DIN2 (___0_9__21685), .Q
       (________24486));
  nnd2s1 ___9___447038(.DIN1 (________24833), .DIN2 (___00___22540), .Q
       (___09____28103));
  nnd2s1 ___9___447039(.DIN1 (____09__21913), .DIN2 (________25707), .Q
       (___90___24245));
  nor2s1 ___9___447040(.DIN1 (____0___25853), .DIN2 (___90___22450), .Q
       (___9____23373));
  and2s1 ___9___447041(.DIN1 (__9_____26591), .DIN2 (________21779), .Q
       (________23039));
  nnd2s1 ___9___447042(.DIN1 (________22012), .DIN2 (___0_____27720),
       .Q (___0_0___27561));
  nnd2s1 ___9___447043(.DIN1 (___90___22449), .DIN2 (___90___22448), .Q
       (________23000));
  nnd2s1 ___9___447044(.DIN1 (___90___22447), .DIN2 (____0___19400), .Q
       (_________28353));
  dffacs1 ___________________447045(.CLRB (reset), .CLK (clk), .DIN
       (________22068), .QN
       (______________0______________________18826));
  and2s1 ___9___447046(.DIN1 (__9__0__26739), .DIN2 (________25704), .Q
       (_____9__24007));
  nnd2s1 ___9__447047(.DIN1 (___9____26200), .DIN2 (____09__24992), .Q
       (_____9__24578));
  nor2s1 ___9___447048(.DIN1 (___9____25206), .DIN2 (________22025), .Q
       (____0___24704));
  nnd2s1 ___9___447049(.DIN1 (_____9__22004), .DIN2 (____0___21453), .Q
       (___9____24271));
  nnd2s1 ___9___447050(.DIN1 (________24619), .DIN2 (__9_____26489), .Q
       (________24762));
  nor2s1 ___9___447051(.DIN1 (___0____22571), .DIN2 (___900__22446), .Q
       (________23030));
  nnd2s1 ___9__447052(.DIN1 (____99__22445), .DIN2 (_____9__22147), .Q
       (____9___22982));
  nnd2s1 ___9___447053(.DIN1 (________21972), .DIN2 (____9___21803), .Q
       (____00__25948));
  nnd2s1 ___9___447054(.DIN1 (__9_____26572), .DIN2
       (_____________________18663), .Q (________24852));
  hi1s1 ___9__447055(.DIN (____9___22444), .Q (________25923));
  hi1s1 ___9___447056(.DIN (____9___22443), .Q (__9_____26713));
  nnd2s1 ___9___447057(.DIN1 (_________34990), .DIN2
       (__________________0___18670), .Q (________24202));
  nor2s1 ___9___447058(.DIN1 (____9___22347), .DIN2 (____9___23973), .Q
       (__90____26310));
  nnd2s1 ___9___447059(.DIN1 (________22038), .DIN2 (___0____21698), .Q
       (____90__25840));
  nnd2s1 ____90_447060(.DIN1 (_____9__23544), .DIN2 (__9_____26401), .Q
       (________25010));
  and2s1 ____9_447061(.DIN1 (________24177), .DIN2 (___9____24323), .Q
       (________26089));
  hi1s1 ___9___447062(.DIN (____9___22442), .Q (__9_00));
  hi1s1 ___9__447063(.DIN (__9_9___26507), .Q (___9____23387));
  nnd2s1 ___9___447064(.DIN1 (________24177), .DIN2 (____90__21895), .Q
       (________24722));
  nnd2s1 ___9_447065(.DIN1 (________22748), .DIN2 (____90__22346), .Q
       (________24207));
  nor2s1 ___9___447066(.DIN1 (________25593), .DIN2 (____9___22441), .Q
       (___09___25361));
  nnd2s1 ___9___447067(.DIN1 (________22036), .DIN2 (________21208), .Q
       (___9____26218));
  nor2s1 ___9___447068(.DIN1 (________22113), .DIN2 (________22045), .Q
       (___9____26209));
  nnd2s1 ___9__447069(.DIN1 (________22028), .DIN2 (___0____21684), .Q
       (___9____23402));
  nor2s1 ___9___447070(.DIN1 (____9___22257), .DIN2 (________24814), .Q
       (___0_____27410));
  nnd2s1 ___9___447071(.DIN1 (_________28636), .DIN2 (_____9___28891),
       .Q (___0_0___27659));
  or2s1 ___9___447072(.DIN1 (________22730), .DIN2 (____9___22440), .Q
       (________25728));
  nnd2s1 ___9__447073(.DIN1 (____99__22445), .DIN2 (________22141), .Q
       (____0___25465));
  and2s1 ___9___447074(.DIN1 (____9___22439), .DIN2 (___99___22527), .Q
       (______9__28464));
  nnd2s1 ___9_447075(.DIN1 (__9_____26572), .DIN2 (____9___22253), .Q
       (__9_____26354));
  nnd2s1 ___9___447076(.DIN1 (________22047), .DIN2 (____9___22438), .Q
       (____0_9__30961));
  nor2s1 ___9_0_447077(.DIN1 (____9___22437), .DIN2 (____90__22436), .Q
       (________23033));
  nor2s1 ___9___447078(.DIN1 (________21458), .DIN2 (_____0__22043), .Q
       (_____00__30545));
  nnd2s1 ___9__447079(.DIN1 (_____9__22052), .DIN2 (_____9__22435), .Q
       (____0____31829));
  and2s1 ___9_0_447080(.DIN1 (________22021), .DIN2 (_____0__21831), .Q
       (_________33153));
  nor2s1 ___9___447081(.DIN1 (________22039), .DIN2 (________22034), .Q
       (_____9___32930));
  nor2s1 ___9___447082(.DIN1 (________22434), .DIN2 (________22018), .Q
       (_________32049));
  nor2s1 ___9___447083(.DIN1 (_____9__20303), .DIN2 (________22051), .Q
       (_________33444));
  nnd2s1 ___9___447084(.DIN1 (________22431), .DIN2 (________22433), .Q
       (____9___22890));
  nor2s1 ___9_447085(.DIN1 (________22432), .DIN2 (________22431), .Q
       (________23596));
  nnd2s1 ___9___447086(.DIN1 (________22201), .DIN2 (________22149), .Q
       (________22430));
  nor2s1 ___9___447087(.DIN1 (__9_9___26888), .DIN2 (________22111), .Q
       (________22429));
  nnd2s1 ___9___447088(.DIN1 (________21944), .DIN2 (_____9___30173),
       .Q (________22428));
  and2s1 ___9___447089(.DIN1 (__9_9___26888), .DIN2 (___99___22527), .Q
       (_____0__22427));
  nor2s1 ___9___447090(.DIN1 (________22425), .DIN2 (________22424), .Q
       (_____9__22426));
  nnd2s1 ___9___447091(.DIN1 (________22424), .DIN2 (____9___19395), .Q
       (________22423));
  or2s1 ___9___447092(.DIN1 (________22421), .DIN2 (___0_0__22573), .Q
       (________22422));
  nnd2s1 ___9___447093(.DIN1 (_________35000), .DIN2 (____0___23716),
       .Q (________22420));
  nnd2s1 ___9___447094(.DIN1 (___0____24393), .DIN2 (___9____26220), .Q
       (________22419));
  nor2s1 ___9___447095(.DIN1 (____0___19400), .DIN2 (________23733), .Q
       (________22418));
  and2s1 ___9___447096(.DIN1 (_____9__22416), .DIN2 (_____0__23326), .Q
       (_____0__22417));
  nor2s1 ___9___447097(.DIN1 (____0___22263), .DIN2 (___9____22510), .Q
       (________22415));
  nor2s1 ___9___447098(.DIN1 (__9_____26953), .DIN2 (________24205), .Q
       (________22414));
  or2s1 ___9___447099(.DIN1 (________22412), .DIN2 (___0_0__22573), .Q
       (________22413));
  nor2s1 ___9___447100(.DIN1 (________22410), .DIN2 (____9___23169), .Q
       (________22411));
  nor2s1 ___9___447101(.DIN1 (________20256), .DIN2 (_________33442),
       .Q (________22409));
  nor2s1 ___9_9_447102(.DIN1 (_____0__22063), .DIN2 (____0___22360), .Q
       (________22407));
  or2s1 ___9___447103(.DIN1 (____0___22812), .DIN2 (____9___22439), .Q
       (________22406));
  nnd2s1 ___9___447104(.DIN1 (_____9__21956), .DIN2 (___0____20730), .Q
       (________22405));
  and2s1 ___9___447105(.DIN1 (___99___22529), .DIN2 (_______18998), .Q
       (________22404));
  nnd2s1 ___9___447106(.DIN1 (____9___22165), .DIN2 (___90___22449), .Q
       (________22403));
  nnd2s1 ___9__447107(.DIN1 (________22011), .DIN2 (________20859), .Q
       (________22402));
  and2s1 ___9___447108(.DIN1 (____09__22998), .DIN2 (____9___19395), .Q
       (________22401));
  and2s1 ___9___447109(.DIN1 (___99___22529), .DIN2
       (_________9_______18812), .Q (_____0__22400));
  nor2s1 ___9___447110(.DIN1 (___0_0__25290), .DIN2 (________22398), .Q
       (_____9__22399));
  nnd2s1 ___0___447111(.DIN1 (________22335), .DIN2 (________21369), .Q
       (________22397));
  nor2s1 ___0___447112(.DIN1 (________19190), .DIN2 (_________35004),
       .Q (________22396));
  nor2s1 ___0___447113(.DIN1 (____9___19679), .DIN2 (_________35004),
       .Q (________22395));
  nor2s1 ___0__447114(.DIN1 (________22393), .DIN2 (________22392), .Q
       (________22394));
  and2s1 ___0___447115(.DIN1 (_____0__21940), .DIN2 (________22339), .Q
       (_____9__22391));
  nor2s1 ___0___447116(.DIN1 (________21405), .DIN2 (__9_____26953), .Q
       (________22390));
  nor2s1 ___0___447117(.DIN1 (________22388), .DIN2 (________22387), .Q
       (________22389));
  hi1s1 ___0___447118(.DIN (_____0__24551), .Q (________22386));
  hi1s1 ___0___447119(.DIN (________25531), .Q (________22385));
  hi1s1 ___0___447120(.DIN (___0_0__24343), .Q (_____0__22384));
  hi1s1 ___0___447121(.DIN (___0____22593), .Q (________22383));
  nor2s1 ___0___447122(.DIN1 (_____9__24719), .DIN2 (________22381), .Q
       (________22382));
  nor2s1 ___9__447123(.DIN1 (________22965), .DIN2 (________24205), .Q
       (________22380));
  and2s1 ___0___447124(.DIN1 (________21932), .DIN2 (________22378), .Q
       (________22379));
  and2s1 ___0__447125(.DIN1 (________21929), .DIN2 (___9____26159), .Q
       (________22377));
  nnd2s1 ___0___447126(.DIN1 (________21927), .DIN2 (inData[30]), .Q
       (________22376));
  or2s1 ___0_0_447127(.DIN1 (_________________18728), .DIN2
       (_________35004), .Q (_____0__22375));
  nnd2s1 ___9___447128(.DIN1 (________22424), .DIN2 (________23814), .Q
       (_____9__22374));
  nnd2s1 ___0_0_447129(.DIN1 (____9___21899), .DIN2 (____09__22815), .Q
       (________22373));
  hi1s1 ___99__447130(.DIN (_____9__22669), .Q (________22372));
  nnd2s1 ___9__447131(.DIN1 (________21954), .DIN2 (________22370), .Q
       (________22943));
  hi1s1 ___00__447132(.DIN (______0__34988), .Q (___0_____27896));
  or2s1 ___9_0_447133(.DIN1 (__90_9), .DIN2 (___90___22450), .Q
       (____0___22991));
  and2s1 ___9___447134(.DIN1 (_____0__24588), .DIN2 (________22369), .Q
       (________24073));
  hi1s1 ___99__447135(.DIN (________22368), .Q (________25095));
  nor2s1 ___99__447136(.DIN1 (________24642), .DIN2 (_____9__23868), .Q
       (_____0__22680));
  hi1s1 ___0__447137(.DIN (________22367), .Q (________24036));
  and2s1 ___9__447138(.DIN1 (___0____25307), .DIN2 (________23938), .Q
       (_____0__22816));
  nnd2s1 ___9_9_447139(.DIN1 (_____0__21948), .DIN2 (_____0__22366), .Q
       (________23144));
  or2s1 ___9_9_447140(.DIN1 (____09__22365), .DIN2 (___9____26182), .Q
       (____0___22992));
  and2s1 ___9_0_447141(.DIN1 (________23071), .DIN2 (________21496), .Q
       (________22917));
  nnd2s1 ___9_447142(.DIN1 (___9____22506), .DIN2 (____0___22364), .Q
       (________23139));
  nnd2s1 ___9__447143(.DIN1 (___0_____27894), .DIN2 (_____0__23199), .Q
       (________23701));
  nor2s1 ___9_447144(.DIN1 (____0___22363), .DIN2 (________22030), .Q
       (________23015));
  nor2s1 ___9__447145(.DIN1 (____09__23983), .DIN2 (____9___22440), .Q
       (___0____22613));
  and2s1 ___9___447146(.DIN1 (____0___22087), .DIN2 (__9_____26828), .Q
       (________23057));
  nor2s1 ___9___447147(.DIN1 (____0___22362), .DIN2 (________25499), .Q
       (____9___22803));
  nor2s1 ___9___447148(.DIN1 (__9__9__27073), .DIN2 (__9__0__26449), .Q
       (________22691));
  nnd2s1 ___0__447149(.DIN1 (____9___21899), .DIN2 (inData[11]), .Q
       (___0_9__22581));
  nor2s1 ___0___447150(.DIN1 (________21178), .DIN2 (___0090__27257),
       .Q (________23022));
  and2s1 ___9___447151(.DIN1 (_____0__24588), .DIN2 (_____9__23142), .Q
       (___0____24350));
  nnd2s1 ___9___447152(.DIN1 (________24144), .DIN2 (_________35010),
       .Q (________22657));
  hi1s1 ___9_0_447153(.DIN (___9____25195), .Q (________22906));
  hi1s1 ___0___447154(.DIN (____0___22361), .Q (____0___23088));
  nor2s1 ___9___447155(.DIN1 (_____9__21979), .DIN2 (____0___22360), .Q
       (________22966));
  nnd2s1 ___9___447156(.DIN1 (__9_9___26888), .DIN2 (___0____23448), .Q
       (___0__9__27324));
  nor2s1 ___9___447157(.DIN1 (____0___22359), .DIN2 (__9_____26838), .Q
       (___0____22614));
  hi1s1 ___0__447158(.DIN (_____0__22653), .Q (________22858));
  or2s1 ___0___447159(.DIN1 (___0____22559), .DIN2 (___0090__27257), .Q
       (____0___22901));
  or2s1 ___0___447160(.DIN1 (____0___22362), .DIN2 (__9_____26487), .Q
       (________22819));
  nor2s1 ___0___447161(.DIN1 (____0___22358), .DIN2 (________25389), .Q
       (________22661));
  nor2s1 ___0___447162(.DIN1 (____0___22357), .DIN2 (_____9__21939), .Q
       (_____9__22847));
  nor2s1 ___0_0_447163(.DIN1 (__9__0__26749), .DIN2 (___9____23399), .Q
       (________24089));
  nor2s1 ___0_447164(.DIN1 (__9_____26597), .DIN2 (____00__22356), .Q
       (__9_____26362));
  nnd2s1 ___9__447165(.DIN1 (___90___22447), .DIN2 (___00___22540), .Q
       (________23110));
  nor2s1 ___9___447166(.DIN1 (__9_____26655), .DIN2 (____99__22355), .Q
       (________23058));
  nor2s1 ___9___447167(.DIN1 (________22136), .DIN2 (____0___22360), .Q
       (________22823));
  nnd2s1 ___9___447168(.DIN1 (___9_0__22500), .DIN2 (________22203), .Q
       (_____9__23055));
  and2s1 ___9___447169(.DIN1 (____9___22354), .DIN2 (____9___22353), .Q
       (________22931));
  or2s1 ___9___447170(.DIN1 (________22859), .DIN2 (________25983), .Q
       (________22907));
  nnd2s1 ___9__447171(.DIN1 (________23207), .DIN2 (____9___21809), .Q
       (________23749));
  nnd2s1 ___9___447172(.DIN1 (________21958), .DIN2 (________23140), .Q
       (________23123));
  nnd2s1 ___9___447173(.DIN1 (____9___22352), .DIN2 (________23814), .Q
       (________22960));
  nnd2s1 ___9___447174(.DIN1 (________22066), .DIN2 (____9___21073), .Q
       (________22957));
  hi1s1 ___0_0_447175(.DIN (_________31464), .Q (________22835));
  nor2s1 ___9___447176(.DIN1 (________22102), .DIN2 (_____9__21884), .Q
       (____99__23711));
  or2s1 ___0__447177(.DIN1 (____99__24517), .DIN2 (__9_____26935), .Q
       (________22940));
  hi1s1 ___0_9_447178(.DIN (__9_9___26604), .Q (____90__25939));
  nnd2s1 ___9___447179(.DIN1 (________22090), .DIN2 (___99___26242), .Q
       (___9____23371));
  nnd2s1 ___0___447180(.DIN1 (_____9___28891), .DIN2 (________25913),
       .Q (____90___28999));
  and2s1 ___0___447181(.DIN1 (____9___22351), .DIN2 (___9____21583), .Q
       (________24669));
  and2s1 ___0_0_447182(.DIN1 (_____9___28891), .DIN2 (____0___22364),
       .Q (____9___24151));
  nor2s1 ___9__447183(.DIN1 (__9_9___26695), .DIN2 (___90___22450), .Q
       (________24735));
  hi1s1 ___0___447184(.DIN (____9___22350), .Q (_____0__23303));
  nor2s1 ___9__447185(.DIN1 (____0___22812), .DIN2 (________22207), .Q
       (________23031));
  nor2s1 ___9___447186(.DIN1 (________21283), .DIN2 (____99__22080), .Q
       (________22915));
  or2s1 ___9___447187(.DIN1 (____9___22349), .DIN2 (___0_____27483), .Q
       (____9___24884));
  hi1s1 ___0___447188(.DIN (___0____22609), .Q (________25399));
  hi1s1 ___9_9_447189(.DIN (__9_____26372), .Q (___9____23401));
  nor2s1 ___0___447190(.DIN1 (________21938), .DIN2 (____9___22348), .Q
       (________22845));
  or2s1 ___0___447191(.DIN1 (________23911), .DIN2 (____9___22347), .Q
       (___0_9___27748));
  nor2s1 ___9_9_447192(.DIN1 (__9_____27023), .DIN2 (___0_____27483),
       .Q (_____0__24646));
  dffacs1 ___________________447193(.CLRB (reset), .CLK (clk), .DIN
       (________22006), .Q (_________________18682));
  nnd2s1 ___9_9_447194(.DIN1 (________22121), .DIN2 (_________35064),
       .Q (________25123));
  and2s1 ___9_9_447195(.DIN1 (________24459), .DIN2 (____90__22346), .Q
       (________23010));
  nor2s1 ___99_447196(.DIN1 (___0____22571), .DIN2 (________22124), .Q
       (________22876));
  nor2s1 ___99__447197(.DIN1 (____0________________18592), .DIN2
       (________21968), .Q (________22959));
  nnd2s1 ___99__447198(.DIN1 (_____9__22345), .DIN2 (_________34994),
       .Q (___09___23520));
  nor2s1 ___9___447199(.DIN1 (____9___25943), .DIN2 (__9_0___26338), .Q
       (________23014));
  nnd2s1 ___990_447200(.DIN1 (________21965), .DIN2 (________22818), .Q
       (________25137));
  nor2s1 ___0___447201(.DIN1 (________22344), .DIN2 (________22343), .Q
       (________23003));
  nor2s1 ___0___447202(.DIN1 (________22342), .DIN2 (________21936), .Q
       (__9_0___26424));
  and2s1 ___99__447203(.DIN1 (___9____24253), .DIN2 (________23539), .Q
       (________25861));
  and2s1 ___0___447204(.DIN1 (________21941), .DIN2 (________22341), .Q
       (__9_9___26511));
  and2s1 ___99__447205(.DIN1 (__9_____26686), .DIN2 (__9__0__26494), .Q
       (____0___24890));
  nnd2s1 ___99__447206(.DIN1 (________22431), .DIN2 (________21917), .Q
       (________22941));
  and2s1 ___990_447207(.DIN1 (__9_____26591), .DIN2 (__9_____26387), .Q
       (________25641));
  or2s1 ___99_447208(.DIN1 (________25910), .DIN2 (___0____22592), .Q
       (________25413));
  and2s1 ___990_447209(.DIN1 (___00____27220), .DIN2 (________22340),
       .Q (________25139));
  or2s1 ___99__447210(.DIN1 (________22685), .DIN2 (________24205), .Q
       (________23066));
  and2s1 ___0__447211(.DIN1 (_____9___28891), .DIN2 (___9____26235), .Q
       (________26079));
  nnd2s1 ___0___447212(.DIN1 (________21931), .DIN2 (________22339), .Q
       (_____9__25596));
  nor2s1 ___9___447213(.DIN1 (________22338), .DIN2 (________25593), .Q
       (___0____25305));
  hi1s1 ___9_447214(.DIN (_____9__22699), .Q (________22953));
  nor2s1 ___9___447215(.DIN1 (____09__23983), .DIN2 (___90___22447), .Q
       (________25806));
  nnd2s1 ___99__447216(.DIN1 (_____0__22337), .DIN2 (_____9__22336), .Q
       (_____9__25415));
  nnd2s1 ___99__447217(.DIN1 (_____9__22416), .DIN2 (________25836), .Q
       (__9_9___26416));
  nor2s1 ___99__447218(.DIN1 (____9___21898), .DIN2 (____0___22360), .Q
       (___9____24318));
  hi1s1 ___00__447219(.DIN (__9_____27045), .Q (________25535));
  nor2s1 ___99__447220(.DIN1 (________21505), .DIN2 (_____0__21962), .Q
       (__9_____26736));
  hi1s1 ___9_0_447221(.DIN (____0____30965), .Q (_________30131));
  nnd2s1 ___0___447222(.DIN1 (________22335), .DIN2 (_____0__20254), .Q
       (_____9__24655));
  nor2s1 ___0___447223(.DIN1 (inData[24]), .DIN2 (_____9__21884), .Q
       (___0_____27386));
  dffacs1 ___________________447224(.CLRB (reset), .CLK (clk), .DIN
       (________22008), .Q
       (______________0___________________9__18827));
  dffacs1 ___________________447225(.CLRB (reset), .CLK (clk), .DIN
       (________21946), .Q (_________________18683));
  nor2s1 ___99__447226(.DIN1 (________22334), .DIN2 (____90__22436), .Q
       (________22909));
  and2s1 ___0__447227(.DIN1 (________22969), .DIN2 (________21873), .Q
       (________26121));
  nnd2s1 ___0___447228(.DIN1 (________21886), .DIN2 (_________28294),
       .Q (__9_____26773));
  or2s1 ___99__447229(.DIN1 (____9____32697), .DIN2 (_________32440),
       .Q (_________32492));
  hi1s1 ___00__447230(.DIN (__99_9__27116), .Q (__9_____26469));
  nnd2s1 ___9___447231(.DIN1 (________21963), .DIN2 (________22333), .Q
       (_________30166));
  nor2s1 ___0___447232(.DIN1 (inData[13]), .DIN2 (__9_____26953), .Q
       (__9_____26962));
  nor2s1 ___0___447233(.DIN1 (inData[11]), .DIN2 (________22146), .Q
       (__9_____27061));
  hi1s1 ___0_0_447234(.DIN (________22737), .Q (___9____25213));
  nor2s1 ___99_447235(.DIN1 (________22332), .DIN2 (________22016), .Q
       (_________32624));
  nor2s1 ___0___447236(.DIN1 (____0___24155), .DIN2 (_____9__21884), .Q
       (__9__0__27005));
  nor2s1 ___99_447237(.DIN1 (________22331), .DIN2 (________22431), .Q
       (________23062));
  hi1s1 ___00__447238(.DIN (________22692), .Q (____0____32793));
  nor2s1 ___99_447239(.DIN1 (____0___19211), .DIN2 (____90__22436), .Q
       (_____9__22961));
  nnd2s1 ___0___447240(.DIN1 (________21886), .DIN2 (inData[13]), .Q
       (__90____26312));
  nor2s1 ___99__447241(.DIN1 (________22330), .DIN2 (________22431), .Q
       (________23070));
  and2s1 ___9___447242(.DIN1 (___099__21718), .DIN2 (____9___22886), .Q
       (________22329));
  and2s1 ___9__447243(.DIN1 (_____0__22327), .DIN2 (___9____22463), .Q
       (________22328));
  nor2s1 ___9__447244(.DIN1 (________21780), .DIN2 (________22325), .Q
       (_____9__22326));
  hi1s1 ___0___447245(.DIN (____9___22353), .Q (________22324));
  hi1s1 ___0___447246(.DIN (________22398), .Q (________22323));
  nor2s1 ___9_0_447247(.DIN1 (________22159), .DIN2 (________21764), .Q
       (________22322));
  nnd2s1 ___9_9_447248(.DIN1 (_____0__22319), .DIN2 (________20094), .Q
       (________22320));
  nor2s1 ___9___447249(.DIN1 (________22114), .DIN2 (________22820), .Q
       (________22318));
  and2s1 ___9___447250(.DIN1 (___909__24248), .DIN2 (________22316), .Q
       (________22317));
  nor2s1 ___9___447251(.DIN1 (____9___22163), .DIN2 (________21731), .Q
       (________22315));
  nnd2s1 ___9__447252(.DIN1 (________21837), .DIN2 (_____0__21885), .Q
       (________22314));
  and2s1 ___9___447253(.DIN1 (_____0__21849), .DIN2 (________22312), .Q
       (________22313));
  nnd2s1 ___9_9_447254(.DIN1 (_____0__22224), .DIN2 (____00__21985), .Q
       (________22311));
  and2s1 ___9_9_447255(.DIN1 (________21737), .DIN2 (____0___21722), .Q
       (_____0__22310));
  nor2s1 ___9_447256(.DIN1 (____9___20978), .DIN2 (________21833), .Q
       (_____9__22309));
  nor2s1 ___9_447257(.DIN1 (_____0__22206), .DIN2 (_____9__21830), .Q
       (________22308));
  nor2s1 ___9___447258(.DIN1 (_____9__21102), .DIN2 (____0___21727), .Q
       (________22307));
  and2s1 ___9___447259(.DIN1 (________21828), .DIN2 (________22333), .Q
       (________22306));
  nnd2s1 ___9___447260(.DIN1 (________22316), .DIN2 (________21915), .Q
       (________22305));
  nnd2s1 ___9___447261(.DIN1 (________21835), .DIN2 (____90__20217), .Q
       (________22304));
  nor2s1 ___9___447262(.DIN1 (________21823), .DIN2 (________22302), .Q
       (________22303));
  and2s1 ___9___447263(.DIN1 (____0___21726), .DIN2 (________23109), .Q
       (________22301));
  or2s1 ___9___447264(.DIN1 (__9_____26660), .DIN2 (________21851), .Q
       (_____0__22300));
  or2s1 ___9__447265(.DIN1 (________23853), .DIN2 (____0___22268), .Q
       (_____9__22299));
  nor2s1 ___9___447266(.DIN1 (________20359), .DIN2 (________21856), .Q
       (________22298));
  nor2s1 ___9__447267(.DIN1 (________19247), .DIN2 (________22296), .Q
       (________22297));
  nnd2s1 ___0___447268(.DIN1 (________21878), .DIN2 (inData[26]), .Q
       (________22295));
  nnd2s1 ___0___447269(.DIN1 (________21745), .DIN2 (inData[4]), .Q
       (________22294));
  and2s1 ___0___447270(.DIN1 (________22189), .DIN2 (________22292), .Q
       (________22293));
  nnd2s1 ___0___447271(.DIN1 (___0____21710), .DIN2 (________22292), .Q
       (_____0__22291));
  nnd2s1 ___0___447272(.DIN1 (___0_0__23500), .DIN2 (________22289), .Q
       (_____9__22290));
  nor2s1 ___0___447273(.DIN1 (________21926), .DIN2 (_____0__21757), .Q
       (________22288));
  nnd2s1 ___0_0_447274(.DIN1 (___9____22461), .DIN2 (________21863), .Q
       (________22287));
  nnd2s1 ___0_447275(.DIN1 (________23140), .DIN2 (________23321), .Q
       (________22286));
  and2s1 ___9___447276(.DIN1 (___0____22607), .DIN2 (________26018), .Q
       (________22285));
  nnd2s1 ___9__447277(.DIN1 (________24859), .DIN2 (_____0__21220), .Q
       (________22284));
  nor2s1 ___9___447278(.DIN1 (_____9___35022), .DIN2 (________21959),
       .Q (________22283));
  nnd2s1 ___9___447279(.DIN1 (_____9__22345), .DIN2 (________21916), .Q
       (________22282));
  nor2s1 ___9_447280(.DIN1 (_____9__22280), .DIN2 (___0____24398), .Q
       (_____0__22281));
  nnd2s1 ___9_9_447281(.DIN1 (_____9___35020), .DIN2 (________26074),
       .Q (________22279));
  nor2s1 ___9_9_447282(.DIN1 (________23757), .DIN2 (_____9___35026),
       .Q (________22278));
  nnd2s1 ___9___447283(.DIN1 (________22276), .DIN2 (________22275), .Q
       (________22277));
  nnd2s1 ___9_0_447284(.DIN1 (____99__22894), .DIN2 (____9___19395), .Q
       (________22274));
  nnd2s1 ___9___447285(.DIN1 (___0____22596), .DIN2 (________23154), .Q
       (________22273));
  nor2s1 ___9__447286(.DIN1 (________22231), .DIN2 (________22343), .Q
       (________22272));
  nor2s1 ___9___447287(.DIN1 (___00___22540), .DIN2 (____09__22270), .Q
       (_____0__22271));
  nor2s1 ___9___447288(.DIN1 (___0____21703), .DIN2 (____0___22268), .Q
       (____0___22269));
  nor2s1 ___9___447289(.DIN1 (________19520), .DIN2 (___0____23508), .Q
       (____0___22267));
  or2s1 ___9__447290(.DIN1 (_________________0___18607), .DIN2
       (_____0__23958), .Q (____0___22266));
  nor2s1 ___9__447291(.DIN1 (________22185), .DIN2 (___9_9__23395), .Q
       (____0___22265));
  nor2s1 ___9__447292(.DIN1 (____0___22263), .DIN2 (________23101), .Q
       (____0___22264));
  nor2s1 ___9___447293(.DIN1 (________21957), .DIN2 (___9_0__23413), .Q
       (____0___22262));
  and2s1 ___9___447294(.DIN1 (_____9___35026), .DIN2 (___9____22463),
       .Q (____00__22261));
  xor2s1 ___9___447295(.DIN1 (_____09__34430), .DIN2 (_________31486),
       .Q (____99__22260));
  xor2s1 ___9__447296(.DIN1 (____9__18996), .DIN2 (______0__30591), .Q
       (____9___22259));
  nor2s1 ___009_447297(.DIN1 (____9___22257), .DIN2 (________25722), .Q
       (____9___22258));
  nor2s1 ___00__447298(.DIN1 (________21175), .DIN2 (____9___22167), .Q
       (____9___22256));
  nnd2s1 ___00__447299(.DIN1 (_____9__22137), .DIN2 (________22783), .Q
       (____9___22255));
  nnd2s1 ___00__447300(.DIN1 (_____0__21763), .DIN2 (____9___22253), .Q
       (____9___22254));
  or2s1 ___00__447301(.DIN1 (__________________0___18670), .DIN2
       (________21842), .Q (____9___22252));
  nnd2s1 ___00__447302(.DIN1 (___99___26242), .DIN2 (________22954), .Q
       (_____9__22251));
  and2s1 ___00_447303(.DIN1 (________22249), .DIN2 (________22134), .Q
       (________22250));
  nnd2s1 ___00__447304(.DIN1 (________22244), .DIN2 (________20924), .Q
       (________22248));
  nnd2s1 ___00__447305(.DIN1 (________22246), .DIN2 (inData[6]), .Q
       (________22247));
  nor2s1 ___00__447306(.DIN1 (__________0__0_), .DIN2 (________22244),
       .Q (________22245));
  nnd2s1 ___00__447307(.DIN1 (_____0__22242), .DIN2
       (__________0___0___18823), .Q (________22243));
  nor2s1 ___00__447308(.DIN1 (_____________________18666), .DIN2
       (___0____21707), .Q (_____9__22241));
  and2s1 ___00__447309(.DIN1 (_____0__22192), .DIN2 (_________18856),
       .Q (________22240));
  nor2s1 ___00__447310(.DIN1 (______9__34470), .DIN2 (____9____32697),
       .Q (________22239));
  hi1s1 ___447311(.DIN (__9_____26838), .Q (________22238));
  hi1s1 ___999_447312(.DIN (___9____24277), .Q (________22237));
  hi1s1 ___99__447313(.DIN (___9_9__22464), .Q (________22236));
  hi1s1 ___99__447314(.DIN (_____0__22234), .Q (________22235));
  nor2s1 ___9__447315(.DIN1 (_____9__22233), .DIN2 (________21798), .Q
       (___9____22466));
  or2s1 ___9___447316(.DIN1 (___9____26215), .DIN2 (________22232), .Q
       (________23731));
  and2s1 ___9_0_447317(.DIN1 (________21834), .DIN2
       (_____________________18664), .Q (_____9__24119));
  nor2s1 ___0__447318(.DIN1 (____0___23085), .DIN2 (___9____25249), .Q
       (____00__22807));
  nor2s1 ___9___447319(.DIN1 (________22231), .DIN2 (___9____24314), .Q
       (________22963));
  hi1s1 ___9___447320(.DIN (________22230), .Q (________22770));
  nor2s1 ___9___447321(.DIN1 (_____0__23199), .DIN2 (________22229), .Q
       (____9___22712));
  hi1s1 ___0__447322(.DIN (________24939), .Q (___0____22591));
  nor2s1 ___9___447323(.DIN1 (___9_0__22491), .DIN2 (_____9__24828), .Q
       (________22769));
  or2s1 ___0__447324(.DIN1 (________23919), .DIN2 (________22859), .Q
       (_____0__22734));
  nor2s1 ___9___447325(.DIN1 (__9_____26660), .DIN2 (________22228), .Q
       (___009__22544));
  nor2s1 ___9___447326(.DIN1 (________22227), .DIN2 (________21826), .Q
       (________22676));
  nor2s1 ___9__447327(.DIN1 (________20338), .DIN2 (________21829), .Q
       (________22758));
  nnd2s1 ___9_9_447328(.DIN1 (________24865), .DIN2 (____9___23800), .Q
       (___00___22543));
  nnd2s1 ___9_9_447329(.DIN1 (___09___21713), .DIN2 (___0_____27905),
       .Q (________22675));
  nnd2s1 ___9_0_447330(.DIN1 (________22226), .DIN2 (________22225), .Q
       (_____9__23608));
  and2s1 ___9_0_447331(.DIN1 (_____0__22224), .DIN2 (___09___21716), .Q
       (________23043));
  nor2s1 ___9_0_447332(.DIN1 (_____9__22223), .DIN2 (___09___21717), .Q
       (________22781));
  nnd2s1 ___9___447333(.DIN1 (________22739), .DIN2 (____0___21358), .Q
       (________23305));
  nor2s1 ___9___447334(.DIN1 (____9___23163), .DIN2 (________24845), .Q
       (___9____22456));
  nor2s1 ___0___447335(.DIN1 (____9___22253), .DIN2 (_____9__21839), .Q
       (________22760));
  nnd2s1 ___0___447336(.DIN1 (________22246), .DIN2 (____90___29904),
       .Q (________22745));
  hi1s1 ___00__447337(.DIN (_________35002), .Q (________22648));
  hi1s1 ___000_447338(.DIN (________22948), .Q (________23589));
  nnd2s1 ___0___447339(.DIN1 (_____0__23933), .DIN2 (___0____22598), .Q
       (________22371));
  nor2s1 ___9___447340(.DIN1 (____09__22365), .DIN2 (_____9___35024),
       .Q (________23759));
  or2s1 ___0___447341(.DIN1 (___99___23432), .DIN2 (________21846), .Q
       (___0_0__23490));
  nor2s1 ___9_9_447342(.DIN1 (_____0__24946), .DIN2 (__9_____27037), .Q
       (_____9__22408));
  hi1s1 ___99__447343(.DIN (____9___22352), .Q (_____9__23311));
  nor2s1 ___99_447344(.DIN1 (________22222), .DIN2 (____0____34554), .Q
       (____9___22443));
  nnd2s1 ___99__447345(.DIN1 (_____0__26077), .DIN2 (________21786), .Q
       (____9___22444));
  nnd2s1 ___0__447346(.DIN1 (________21469), .DIN2 (____9___22437), .Q
       (___0____22583));
  nor2s1 ___0___447347(.DIN1 (________22221), .DIN2 (___00___24334), .Q
       (________23686));
  nnd2s1 ___9___447348(.DIN1 (________22276), .DIN2 (___0____21702), .Q
       (________23050));
  nnd2s1 ___99__447349(.DIN1 (_____9__21961), .DIN2 (________22211), .Q
       (__9_9___26507));
  or2s1 ___9__447350(.DIN1 (________22387), .DIN2 (_____9__24828), .Q
       (________23824));
  nnd2s1 ___9___447351(.DIN1 (________22773), .DIN2 (________22214), .Q
       (________24087));
  nor2s1 ___9_9_447352(.DIN1 (_____0___32299), .DIN2 (________21762),
       .Q (_____9__22699));
  nor2s1 ___9___447353(.DIN1 (___9_0__23413), .DIN2 (________22220), .Q
       (________23147));
  or2s1 ___9___447354(.DIN1 (________25513), .DIN2 (__9_____26583), .Q
       (________23045));
  hi1s1 ___000_447355(.DIN (__9_0___26422), .Q (___9____26230));
  nor2s1 ___9___447356(.DIN1 (________23757), .DIN2 (_____0__22327), .Q
       (___0_____27446));
  nor2s1 ___9___447357(.DIN1 (_____9__21756), .DIN2 (________26032), .Q
       (___9____25208));
  hi1s1 ___00__447358(.DIN (_________33442), .Q (_________33236));
  nor2s1 ___9___447359(.DIN1 (___0____21671), .DIN2 (________22209), .Q
       (________24806));
  nnd2s1 ___9__447360(.DIN1 (________22219), .DIN2 (________24660), .Q
       (_____9__22763));
  nor2s1 ___9___447361(.DIN1 (________22218), .DIN2 (__90_0__26318), .Q
       (___9____24298));
  or2s1 ___990_447362(.DIN1 (________25715), .DIN2 (____0____34554), .Q
       (___99___24331));
  and2s1 ___990_447363(.DIN1 (____99__22894), .DIN2 (________23814), .Q
       (____0____28172));
  nnd2s1 ___447364(.DIN1 (________22217), .DIN2 (________22946), .Q
       (____9___23883));
  nor2s1 ___9_9_447365(.DIN1 (_____0__22216), .DIN2 (________22231), .Q
       (________23738));
  nnd2s1 ___9_9_447366(.DIN1 (________21888), .DIN2 (________25419), .Q
       (___9____23407));
  nor2s1 ___9_9_447367(.DIN1 (____0___21720), .DIN2 (____0___24798), .Q
       (________23292));
  nnd2s1 ___9___447368(.DIN1 (________25672), .DIN2 (__9_____26401), .Q
       (____9___25652));
  nnd2s1 ___99__447369(.DIN1 (________21882), .DIN2 (________21797), .Q
       (________25451));
  hi1s1 ___00_447370(.DIN (____00___31812), .Q (_____0___31005));
  nnd2s1 ___9___447371(.DIN1 (________21860), .DIN2 (_____9__22679), .Q
       (____0____30965));
  nor2s1 ___99_447372(.DIN1 (_____9__22215), .DIN2 (________21825), .Q
       (________26081));
  and2s1 ___9___447373(.DIN1 (________22214), .DIN2 (________24865), .Q
       (___0_____27897));
  hi1s1 ___447374(.DIN (________22213), .Q (________25394));
  nnd2s1 ___9_9_447375(.DIN1 (________22210), .DIN2 (________22119), .Q
       (__9_____26372));
  nor2s1 ___447376(.DIN1 (________22212), .DIN2 (____9___21896), .Q
       (________25132));
  nor2s1 ___99__447377(.DIN1 (___0____25303), .DIN2 (_____9___35024),
       .Q (_____9__25634));
  or2s1 ___99__447378(.DIN1 (________19570), .DIN2 (_____9___35026), .Q
       (___09____28074));
  nnd2s1 ___99__447379(.DIN1 (_____0__21924), .DIN2 (________22289), .Q
       (________25401));
  nnd2s1 ___9_9_447380(.DIN1 (____0___21725), .DIN2 (_____0__22118), .Q
       (__9_____26840));
  nnd2s1 ___9_9_447381(.DIN1 (________22208), .DIN2 (________22211), .Q
       (_________28602));
  nnd2s1 ___9_9_447382(.DIN1 (________22210), .DIN2 (________22339), .Q
       (________25447));
  nor2s1 ___9_9_447383(.DIN1 (________21014), .DIN2 (________22209), .Q
       (_____0__25694));
  nor2s1 ___99_447384(.DIN1 (________21788), .DIN2 (________22209), .Q
       (_____0__24541));
  nnd2s1 ___9_0_447385(.DIN1 (_____9__21858), .DIN2 (________22050), .Q
       (___9____25195));
  nnd2s1 ___9_447386(.DIN1 (________22208), .DIN2 (________22109), .Q
       (__9__9__27014));
  hi1s1 ___00__447387(.DIN (________22207), .Q (___00___23444));
  nnd2s1 ___99__447388(.DIN1 (________22120), .DIN2 (________21774), .Q
       (__9__0__26854));
  nor2s1 ___9___447389(.DIN1 (_____0__22206), .DIN2 (_____0__21859), .Q
       (____9____31746));
  hi1s1 ___0___447390(.DIN (________22201), .Q (________22202));
  nnd2s1 ___9___447391(.DIN1 (________23318), .DIN2 (________19570), .Q
       (_____0__22200));
  nnd2s1 ___00__447392(.DIN1 (________21861), .DIN2 (___9____20620), .Q
       (_____9__22199));
  hi1s1 ___0__447393(.DIN (____0___22360), .Q (________22198));
  hi1s1 ___99__447394(.DIN (________22196), .Q (________22197));
  nnd2s1 ___00__447395(.DIN1 (________22194), .DIN2 (__________0__0_),
       .Q (________22195));
  nnd2s1 ___0___447396(.DIN1 (_____0__22192), .DIN2 (________19082), .Q
       (________22193));
  nor2s1 ___0___447397(.DIN1 (___0_9__20715), .DIN2 (________21848), .Q
       (_____9__22191));
  and2s1 ___0__447398(.DIN1 (________22189), .DIN2 (____0___19599), .Q
       (________22190));
  and2s1 ___0___447399(.DIN1 (________21874), .DIN2 (________22187), .Q
       (________22188));
  nor2s1 ___0__447400(.DIN1 (________22185), .DIN2 (___99___23432), .Q
       (________22186));
  nor2s1 ___9___447401(.DIN1 (________22183), .DIN2 (________21769), .Q
       (________22184));
  nnd2s1 ___0__447402(.DIN1 (____09__22181), .DIN2 (____0___22180), .Q
       (_____0__22182));
  and2s1 ___0___447403(.DIN1 (________26018), .DIN2 (___0____24403), .Q
       (____0___22179));
  nnd2s1 ___0___447404(.DIN1 (________21937), .DIN2 (________24682), .Q
       (____0___22178));
  and2s1 ___0__447405(.DIN1 (____0___22814), .DIN2 (___9____23379), .Q
       (____0___22177));
  nnd2s1 ___0___447406(.DIN1 (___0_0__21705), .DIN2 (_________35062),
       .Q (____0___22176));
  nnd2s1 ___0___447407(.DIN1 (________22421), .DIN2 (____9___19395), .Q
       (____0___22175));
  and2s1 ___0___447408(.DIN1 (________22246), .DIN2 (________19240), .Q
       (____0___22174));
  nnd2s1 ___0___447409(.DIN1 (________22246), .DIN2 (________19637), .Q
       (____0___22173));
  or2s1 ___0___447410(.DIN1 (_____0__22242), .DIN2 (___0_____27291), .Q
       (____00__22172));
  nnd2s1 ___0___447411(.DIN1 (____9___22170), .DIN2 (____09__22634), .Q
       (____99__22171));
  nor2s1 ___0__447412(.DIN1 (_____9__22884), .DIN2 (________21758), .Q
       (____9___22169));
  nor2s1 ___00__447413(.DIN1 (________21922), .DIN2 (____9___22167), .Q
       (____9___22168));
  nor2s1 ___9___447414(.DIN1 (____09__22634), .DIN2 (____9___22165), .Q
       (____9___22166));
  or2s1 ___0___447415(.DIN1 (_____0__22216), .DIN2 (____9___22163), .Q
       (____9___22164));
  hi1s1 ___0___447416(.DIN (_________35004), .Q (________22161));
  nor2s1 ___9___447417(.DIN1 (________22159), .DIN2 (____9___23255), .Q
       (________22160));
  hi1s1 ______447418(.DIN (________22344), .Q (________22158));
  nor2s1 ___9___447419(.DIN1 (_____9__22156), .DIN2 (________21843), .Q
       (_____0__22157));
  nor2s1 ___9___447420(.DIN1 (________21890), .DIN2 (________21832), .Q
       (________22155));
  xor2s1 ___9__447421(.DIN1 (_____9___30624), .DIN2 (_________31281),
       .Q (________22154));
  nnd2s1 ___0___447422(.DIN1 (________24440), .DIN2 (___9____23394), .Q
       (________22153));
  nor2s1 ___0___447423(.DIN1 (_________35016), .DIN2 (___9____21558),
       .Q (________22368));
  hi1s1 ___0___447424(.DIN (________23541), .Q (___0____22604));
  hi1s1 ___0___447425(.DIN (________25910), .Q (___0____22610));
  hi1s1 ___0___447426(.DIN (__9__9__27073), .Q (________22945));
  hi1s1 ___0__447427(.DIN (___0____22567), .Q (___0____22586));
  or2s1 ___0___447428(.DIN1 (_____0___35034), .DIN2 (________22152), .Q
       (____9___23971));
  nnd2s1 ___0___447429(.DIN1 (________22151), .DIN2 (___0____22601), .Q
       (________23182));
  hi1s1 ___0_447430(.DIN (________22424), .Q (__9_____26846));
  or2s1 ___0___447431(.DIN1 (________24221), .DIN2 (_________28294), .Q
       (________22694));
  nor2s1 ___0_447432(.DIN1 (________22037), .DIN2 (________21768), .Q
       (___0_0__22600));
  nnd2s1 ___0__447433(.DIN1 (________22150), .DIN2 (________22130), .Q
       (________22638));
  and2s1 ___0___447434(.DIN1 (________22149), .DIN2 (_____0__22148), .Q
       (___0____22611));
  nnd2s1 ___0___447435(.DIN1 (________22189), .DIN2 (_____9__22147), .Q
       (___0____22587));
  nnd2s1 ___0___447436(.DIN1 (___99___23429), .DIN2 (___0_0__23500), .Q
       (________23121));
  nnd2s1 ___0___447437(.DIN1 (________22145), .DIN2 (___09___21715), .Q
       (________22697));
  nnd2s1 ___0___447438(.DIN1 (________22133), .DIN2 (__9_____26623), .Q
       (_____9__24490));
  nor2s1 ___0_9_447439(.DIN1 (________22144), .DIN2 (___00___24334), .Q
       (________22367));
  nor2s1 ___0__447440(.DIN1 (________22126), .DIN2 (________22425), .Q
       (___090__22617));
  nor2s1 ___0___447441(.DIN1 (_________35060), .DIN2 (____9___22349),
       .Q (____0___22361));
  hi1s1 ___0___447442(.DIN (___9____22462), .Q (___09___22623));
  and2s1 ___9__447443(.DIN1 (________22143), .DIN2 (________21225), .Q
       (________22755));
  hi1s1 ___99_447444(.DIN (________22142), .Q (___0____22585));
  nnd2s1 ___0___447445(.DIN1 (________22189), .DIN2 (________22141), .Q
       (____9___22350));
  and2s1 ___9___447446(.DIN1 (________22140), .DIN2 (________22139), .Q
       (_____9__22753));
  hi1s1 ___447447(.DIN (_________35000), .Q (___0____22588));
  nnd2s1 ___99__447448(.DIN1 (_____0__22138), .DIN2 (___09___21714), .Q
       (____9___22442));
  hi1s1 ___00_447449(.DIN (_________33894), .Q (_________29762));
  nnd2s1 ___0__447450(.DIN1 (________22249), .DIN2 (____9___20602), .Q
       (________23692));
  nor2s1 ___0___447451(.DIN1 (_____9__21772), .DIN2 (________22125), .Q
       (________22727));
  nnd2s1 ___0___447452(.DIN1 (______0__35038), .DIN2 (_____0__21914),
       .Q (___0____22612));
  and2s1 ___0___447453(.DIN1 (_____9__22137), .DIN2 (____0___25470), .Q
       (_____9__25118));
  nnd2s1 ___0___447454(.DIN1 (________22249), .DIN2 (___0_0), .Q
       (________23906));
  nor2s1 ___0___447455(.DIN1 (________22136), .DIN2 (________21753), .Q
       (___0____22609));
  or2s1 ___9___447456(.DIN1 (___99___23432), .DIN2 (________22220), .Q
       (___0____23452));
  hi1s1 ___0_0_447457(.DIN (________25983), .Q (________22706));
  and2s1 ___0___447458(.DIN1 (________21469), .DIN2 (________23136), .Q
       (___0_____27767));
  dffacs1 ______________0_447459(.CLRB (reset), .CLK (clk), .DIN
       (________21844), .QN (_________0___18904));
  or2s1 ___9___447460(.DIN1 (____0___23716), .DIN2 (___0____23508), .Q
       (___0_____27800));
  nor2s1 ___0___447461(.DIN1 (__________________0___18670), .DIN2
       (_________35014), .Q (____9___24605));
  nor2s1 ___0___447462(.DIN1 (________22212), .DIN2 (___0_____27696),
       .Q (_____0__24560));
  nnd2s1 ___0__447463(.DIN1 (_____9__25928), .DIN2 (___0____21704), .Q
       (___0____22606));
  nor2s1 ___0__447464(.DIN1 (________22135), .DIN2 (___0_0__24352), .Q
       (___0____22595));
  or2s1 ___0___447465(.DIN1 (__9_9___26414), .DIN2 (__9_____26499), .Q
       (________24075));
  nnd2s1 ___0__447466(.DIN1 (________22134), .DIN2 (________20436), .Q
       (___09___22620));
  and2s1 ___0___447467(.DIN1 (________22133), .DIN2 (________26068), .Q
       (________24912));
  or2s1 ___0_9_447468(.DIN1 (_____9__22127), .DIN2 (____9___26144), .Q
       (________24079));
  nor2s1 ___0_9_447469(.DIN1 (____0___21991), .DIN2 (________21751), .Q
       (________22696));
  hi1s1 _____0_447470(.DIN (________25739), .Q (___0____22616));
  hi1s1 _______447471(.DIN (__9_____26935), .Q (__9_____26445));
  or2s1 _______447472(.DIN1 (________22132), .DIN2 (___990__25261), .Q
       (________22641));
  and2s1 ___0_9_447473(.DIN1 (_____0__21749), .DIN2 (________22131), .Q
       (___0_9__22599));
  nnd2s1 ___0_447474(.DIN1 (________21865), .DIN2 (____90__21801), .Q
       (___0____22593));
  nnd2s1 ___0_0_447475(.DIN1 (________22130), .DIN2 (________23222), .Q
       (____9___24060));
  nnd2s1 ___9___447476(.DIN1 (________21754), .DIN2 (________22129), .Q
       (_____0__23231));
  nnd2s1 ___0_0_447477(.DIN1 (________22369), .DIN2 (___90___24242), .Q
       (___0_0__24343));
  hi1s1 ___0_9_447478(.DIN (__9_____26917), .Q (________23238));
  and2s1 ___0_447479(.DIN1 (__9_0___26707), .DIN2 (_____0__22128), .Q
       (___0_0__24382));
  and2s1 ___0_9_447480(.DIN1 (________22954), .DIN2 (__9_____26639), .Q
       (________23063));
  nnd2s1 ___9___447481(.DIN1 (___0_____27973), .DIN2 (___0_____27289),
       .Q (____0___23894));
  nor2s1 ___9___447482(.DIN1 (_____9__22127), .DIN2 (________22222), .Q
       (________23871));
  hi1s1 ___00__447483(.DIN (________22431), .Q (___0____22584));
  hi1s1 ___00_447484(.DIN (________23932), .Q (________22776));
  or2s1 ___9_447485(.DIN1 (_____9__22280), .DIN2 (________22126), .Q
       (________23831));
  hi1s1 ___9___447486(.DIN (_________33333), .Q (____9____31752));
  nor2s1 ___0_0_447487(.DIN1 (__90_9__26308), .DIN2 (____00__22356), .Q
       (___0____25329));
  nor2s1 ___9___447488(.DIN1 (____9___19945), .DIN2 (____9___22165), .Q
       (___09____28117));
  nor2s1 ___0_0_447489(.DIN1 (____9___21804), .DIN2 (________22125), .Q
       (_____9__22669));
  hi1s1 ___0___447490(.DIN (________22124), .Q (________26020));
  hi1s1 ___00__447491(.DIN (____90__22436), .Q (___0_0__22582));
  hi1s1 ___0_0_447492(.DIN (_________35006), .Q (__9090));
  nor2s1 ___0__447493(.DIN1 (________22410), .DIN2 (________22123), .Q
       (___0____23484));
  nor2s1 ___0___447494(.DIN1 (____0___22359), .DIN2 (________22122), .Q
       (________24726));
  hi1s1 ___00__447495(.DIN (_________32081), .Q (_________30595));
  hi1s1 ___0___447496(.DIN (________22121), .Q (__9__0__26346));
  nnd2s1 ___0___447497(.DIN1 (________21880), .DIN2 (________22116), .Q
       (________22938));
  hi1s1 ___0_0_447498(.DIN (________23733), .Q (____00__23528));
  and2s1 ___99__447499(.DIN1 (________22120), .DIN2 (________22119), .Q
       (__9_____26535));
  nnd2s1 ___0_0_447500(.DIN1 (_____0___35030), .DIN2 (_____0__22118),
       .Q (__9_9___26604));
  hi1s1 ___0___447501(.DIN (_____9__22117), .Q (___0____22605));
  nnd2s1 ___0_9_447502(.DIN1 (________21744), .DIN2 (________22116), .Q
       (_____0__22653));
  hi1s1 ___0_0_447503(.DIN (___0____22579), .Q (___0_0___27563));
  nnd2s1 ___0___447504(.DIN1 (_________32487), .DIN2 (_____9__21875),
       .Q (________22692));
  nnd2s1 ___99__447505(.DIN1 (________22120), .DIN2 (________22339), .Q
       (________25798));
  nnd2s1 ___0___447506(.DIN1 (________21732), .DIN2 (________22129), .Q
       (_____0__24551));
  hi1s1 ___0___447507(.DIN (________22115), .Q (_____0__25770));
  nor2s1 ___0__447508(.DIN1 (____0____29098), .DIN2 (_____9__21867), .Q
       (_____9__22797));
  nor2s1 ___0___447509(.DIN1 (________22114), .DIN2 (_____0__24772), .Q
       (__9__9__26540));
  nor2s1 ___0___447510(.DIN1 (________21766), .DIN2 (___0____24408), .Q
       (____0___25752));
  nnd2s1 ___0___447511(.DIN1 (________21740), .DIN2 (____0___21988), .Q
       (________24195));
  nor2s1 ___0___447512(.DIN1 (________22113), .DIN2 (_____9__21748), .Q
       (________25531));
  nor2s1 ___0___447513(.DIN1 (________22221), .DIN2 (________25148), .Q
       (________25926));
  hi1s1 ___0_0_447514(.DIN (______9__34123), .Q (_____0___31184));
  nor2s1 ___0___447515(.DIN1 (________22112), .DIN2 (________22126), .Q
       (___0____24386));
  nor2s1 ___0___447516(.DIN1 (________21862), .DIN2 (________21841), .Q
       (___9_9__23422));
  hi1s1 ___447517(.DIN (________22111), .Q (__9__9__27043));
  nnd2s1 ___0___447518(.DIN1 (________21734), .DIN2 (________22110), .Q
       (________22737));
  nnd2s1 ___0___447519(.DIN1 (________21743), .DIN2 (________22109), .Q
       (__9_____26406));
  nnd2s1 ___99__447520(.DIN1 (___00____27196), .DIN2 (_____0__22108),
       .Q (___0_9___27848));
  nnd2s1 ___0___447521(.DIN1 (________21864), .DIN2 (_____0__21504), .Q
       (__9_____27021));
  and2s1 ___0_0_447522(.DIN1 (________22189), .DIN2 (________21188), .Q
       (__9_____26764));
  nnd2s1 ___0___447523(.DIN1 (________21747), .DIN2 (________21499), .Q
       (___0_____27862));
  nnd2s1 ___0___447524(.DIN1 (___0____21654), .DIN2 (inData[21]), .Q
       (__99_9__27116));
  dffacs1 ________________9_447525(.CLRB (reset), .CLK (clk), .DIN
       (________21854), .QN
       (______________________________________0_____________18887));
  and2s1 ___0___447526(.DIN1 (____9____32697), .DIN2 (________21248),
       .Q (_____0___32572));
  nnd2s1 ___0__447527(.DIN1 (________21872), .DIN2 (____9____32697), .Q
       (_________31464));
  hi1s1 ___00__447528(.DIN (____00___32758), .Q (____0_9__32819));
  nor2s1 ___0__447529(.DIN1 (inData[21]), .DIN2 (___0_____27696), .Q
       (__9_____27045));
  or2s1 ___0___447530(.DIN1 (________22106), .DIN2 (__9_____26553), .Q
       (_____9__22107));
  nor2s1 ___0___447531(.DIN1 (________22017), .DIN2 (________21515), .Q
       (________22105));
  nnd2s1 ___0_9_447532(.DIN1 (________21394), .DIN2 (___0_9__20732), .Q
       (________22104));
  and2s1 ___0_447533(.DIN1 (___99___26242), .DIN2 (________23145), .Q
       (________22103));
  or2s1 ___0__447534(.DIN1 (________21415), .DIN2 (___0____24378), .Q
       (________22102));
  nor2s1 ___0___447535(.DIN1 (________22056), .DIN2 (___0____21642), .Q
       (________22101));
  nor2s1 ___9___447536(.DIN1 (________22123), .DIN2 (_____0__22099), .Q
       (________22100));
  or2s1 ___9___447537(.DIN1 (____0___23716), .DIN2 (________22677), .Q
       (_____9__22098));
  nor2s1 ___9___447538(.DIN1 (_____0__23199), .DIN2 (___9____22495), .Q
       (________22097));
  or2s1 ___9_447539(.DIN1 (________19570), .DIN2 (___0____21688), .Q
       (________22096));
  nor2s1 ___9__447540(.DIN1 (____9___22347), .DIN2 (____0___25853), .Q
       (________22095));
  and2s1 ___9___447541(.DIN1 (________22093), .DIN2 (________23154), .Q
       (________22094));
  and2s1 ___9___447542(.DIN1 (________22091), .DIN2 (___9____23416), .Q
       (________22092));
  nor2s1 ___0___447543(.DIN1 (_____0__22089), .DIN2 (_____0__23591), .Q
       (________22090));
  nor2s1 ___0___447544(.DIN1 (________22688), .DIN2 (__9_____26655), .Q
       (____09__22088));
  and2s1 ___0___447545(.DIN1 (___00___23438), .DIN2 (________23917), .Q
       (____0___22087));
  nor2s1 ___0___447546(.DIN1 (____9___19395), .DIN2 (______0__35048),
       .Q (____0___22086));
  nor2s1 ___0__447547(.DIN1 (___0_0__23481), .DIN2 (___0____21670), .Q
       (____0___22085));
  nor2s1 ___9__447548(.DIN1 (________23154), .DIN2 (___99___22533), .Q
       (____0___22084));
  nor2s1 ___009_447549(.DIN1 (___0_0__21696), .DIN2 (________22035), .Q
       (____0___22083));
  xnr2s1 ___9_447550(.DIN1 (_________31395), .DIN2 (____99___31805), .Q
       (____0___22082));
  nor2s1 ___00__447551(.DIN1 (________25622), .DIN2 (____0___21989), .Q
       (____00__22081));
  nnd2s1 ___0___447552(.DIN1 (___9____21603), .DIN2 (___09___20783), .Q
       (____99__22080));
  nor2s1 ___0___447553(.DIN1 (________22965), .DIN2 (____9___22078), .Q
       (____9___22079));
  or2s1 ___0___447554(.DIN1 (________21730), .DIN2 (________21996), .Q
       (____9___22077));
  nnd2s1 ___0___447555(.DIN1 (________22678), .DIN2 (__9_9___26791), .Q
       (____9___22076));
  xor2s1 ___9___447556(.DIN1 (____9___22074), .DIN2 (____9___22073), .Q
       (____9___22075));
  xnr2s1 ___9___447557(.DIN1 (_________30496), .DIN2 (_________28737),
       .Q (____9___22072));
  nor2s1 ___0___447558(.DIN1 (_____0__22924), .DIN2 (_____9__23161), .Q
       (____90__22071));
  nor2s1 ___0___447559(.DIN1 (________22069), .DIN2 (________22123), .Q
       (_____9__22070));
  nnd2s1 ___0___447560(.DIN1 (____9___21540), .DIN2 (________22067), .Q
       (________22068));
  or2s1 ___0___447561(.DIN1 (____9___21980), .DIN2 (___99___21630), .Q
       (________22066));
  nor2s1 ___0___447562(.DIN1 (____0___23085), .DIN2 (__9__9__26921), .Q
       (________22065));
  nor2s1 ___0__447563(.DIN1 (_____0__22063), .DIN2 (___00___21636), .Q
       (________22064));
  nor2s1 ___0___447564(.DIN1 (___99___20692), .DIN2 (_________34159),
       .Q (_____9__22062));
  nnd2s1 ___0___447565(.DIN1 (___0_____27804), .DIN2 (____0___23716),
       .Q (________22061));
  hi1s1 ___0_9_447566(.DIN (________26032), .Q (________22060));
  nnd2s1 ___0___447567(.DIN1 (________21315), .DIN2 (___90___21548), .Q
       (________22059));
  and2s1 ___00__447568(.DIN1 (___9____25206), .DIN2 (_____18908), .Q
       (________22058));
  nor2s1 ___00_447569(.DIN1 (___00___21640), .DIN2 (________22056), .Q
       (________22057));
  and2s1 ___00__447570(.DIN1 (________22054), .DIN2 (________22783), .Q
       (________22055));
  nor2s1 ___00__447571(.DIN1 (____9___21253), .DIN2 (___0_0__21686), .Q
       (_____0__22053));
  nor2s1 ___00__447572(.DIN1 (___00___20705), .DIN2 (___9____21586), .Q
       (_____9__22052));
  nor2s1 ___00__447573(.DIN1 (________22050), .DIN2 (________21516), .Q
       (________22051));
  nor2s1 ___00_447574(.DIN1 (___999), .DIN2 (________22048), .Q
       (________22049));
  nor2s1 ___00__447575(.DIN1 (________19911), .DIN2 (___000__21633), .Q
       (________22047));
  nor2s1 ___00__447576(.DIN1 (________21331), .DIN2 (___9____21585), .Q
       (________22046));
  nnd2s1 ___00_447577(.DIN1 (___0____21645), .DIN2 (________21824), .Q
       (________22045));
  nor2s1 ___00_447578(.DIN1 (________21919), .DIN2 (___9____22458), .Q
       (________22044));
  or2s1 ___00__447579(.DIN1 (_____9__22042), .DIN2 (___00___21637), .Q
       (_____0__22043));
  nnd2s1 ___00__447580(.DIN1 (________22112), .DIN2 (____9___19395), .Q
       (________22041));
  nor2s1 ___00_447581(.DIN1 (________22039), .DIN2 (_____0__21410), .Q
       (________22040));
  nor2s1 ___00__447582(.DIN1 (________22037), .DIN2 (_____9__21970), .Q
       (________22038));
  nor2s1 ___00__447583(.DIN1 (_____0__21971), .DIN2 (________22035), .Q
       (________22036));
  nnd2s1 ___009_447584(.DIN1 (___0____21646), .DIN2 (________21528), .Q
       (________22034));
  nor2s1 ___009_447585(.DIN1 (_____9__20180), .DIN2 (____9___21902), .Q
       (_____0__22033));
  nnd2s1 ___009_447586(.DIN1 (___9____21613), .DIN2 (_____9__20575), .Q
       (_____9__22032));
  nor2s1 ___009_447587(.DIN1 (_____0__21783), .DIN2 (_____9__22743), .Q
       (________22031));
  nnd2s1 ___0_0_447588(.DIN1 (____09__22815), .DIN2 (________22029), .Q
       (________22030));
  nor2s1 ___0_0_447589(.DIN1 (___9____20617), .DIN2 (________22035), .Q
       (________22028));
  and2s1 ___0_0_447590(.DIN1 (________21998), .DIN2 (________22026), .Q
       (________22027));
  nnd2s1 ___0_447591(.DIN1 (________22024), .DIN2 (_____0__22023), .Q
       (________22025));
  nnd2s1 ___0__447592(.DIN1 (________22112), .DIN2 (________23814), .Q
       (_____9__22022));
  nor2s1 ___0___447593(.DIN1 (________21379), .DIN2 (___0____21653), .Q
       (________22021));
  nnd2s1 ___0___447594(.DIN1 (___9____24323), .DIN2 (____9___21901), .Q
       (________22020));
  and2s1 ___0__447595(.DIN1 (________21436), .DIN2 (________22131), .Q
       (________22019));
  nnd2s1 ___0__447596(.DIN1 (___9_0__21553), .DIN2 (____90__21533), .Q
       (________22018));
  nnd2s1 ___0___447597(.DIN1 (___9_0__21571), .DIN2 (________21855), .Q
       (________22016));
  nor2s1 ___0___447598(.DIN1 (________23814), .DIN2 (_____0__22014), .Q
       (________22015));
  and2s1 ___0___447599(.DIN1 (___90___21551), .DIN2
       (__________________0___18628), .Q (_____9__22013));
  nnd2s1 ___0__447600(.DIN1 (___9_0__26207), .DIN2 (________24221), .Q
       (________22012));
  nor2s1 ___0__447601(.DIN1 (________20092), .DIN2 (___9____21604), .Q
       (________22011));
  and2s1 ___0___447602(.DIN1 (________22026), .DIN2 (________23007), .Q
       (________22010));
  nnd2s1 ___0__447603(.DIN1 (____0___21906), .DIN2 (________21976), .Q
       (________22009));
  nnd2s1 ___0___447604(.DIN1 (___9_9__21560), .DIN2 (________22067), .Q
       (________22008));
  nor2s1 ___0___447605(.DIN1 (___9___19031), .DIN2 (________22048), .Q
       (________22007));
  nnd2s1 ___0___447606(.DIN1 (________21521), .DIN2 (________19629), .Q
       (________22006));
  nnd2s1 ___0___447607(.DIN1 (___9_9__21579), .DIN2 (____0___20892), .Q
       (_____0__22005));
  nor2s1 ___0___447608(.DIN1 (_____0__21429), .DIN2 (________22002), .Q
       (_____9__22004));
  nor2s1 ___0___447609(.DIN1 (___0____20718), .DIN2 (___0_0__21649), .Q
       (________22003));
  nor2s1 ___0_0_447610(.DIN1 (________21974), .DIN2 (____9___21983), .Q
       (________22111));
  nor2s1 ___0___447611(.DIN1 (____9___21900), .DIN2 (________21526), .Q
       (________22196));
  nor2s1 ___0___447612(.DIN1 (________21471), .DIN2 (________22002), .Q
       (_____0__22234));
  nor2s1 ___0___447613(.DIN1 (____99__21542), .DIN2 (________21973), .Q
       (___9____23393));
  nor2s1 ___0___447614(.DIN1 (________22001), .DIN2 (___0____22603), .Q
       (________23274));
  nor2s1 ___0___447615(.DIN1 (___9____21600), .DIN2 (____9___22348), .Q
       (___9____22503));
  and2s1 ___0___447616(.DIN1 (___9____21572), .DIN2 (________22000), .Q
       (___0____22602));
  nnd2s1 ___0___447617(.DIN1 (___090__21711), .DIN2 (___9____21596), .Q
       (________22947));
  and2s1 ___0_447618(.DIN1 (________21838), .DIN2 (________22131), .Q
       (________22695));
  nnd2s1 ___0_9_447619(.DIN1 (________21999), .DIN2 (_____0__22014), .Q
       (___9____22457));
  nnd2s1 ___0_9_447620(.DIN1 (________21998), .DIN2 (________25817), .Q
       (________22704));
  or2s1 ___0_9_447621(.DIN1 (________21997), .DIN2 (___9____26213), .Q
       (___9____23391));
  and2s1 ___0__447622(.DIN1 (__9_____26358), .DIN2 (__9_00__26798), .Q
       (________25444));
  nor2s1 ___0_0_447623(.DIN1 (___9____21584), .DIN2 (___9____26215), .Q
       (________22321));
  nor2s1 ___0_0_447624(.DIN1 (________19613), .DIN2 (________21996), .Q
       (___90___22452));
  nor2s1 ___0_9_447625(.DIN1 (___99___21628), .DIN2 (____0___21908), .Q
       (___00___22538));
  nnd2s1 ___0_9_447626(.DIN1 (________22289), .DIN2 (___00___23438), .Q
       (___9____22470));
  nnd2s1 ___0_9_447627(.DIN1 (________21765), .DIN2 (________22139), .Q
       (________22639));
  nnd2s1 ___0_9_447628(.DIN1 (________22818), .DIN2 (__9_____26779), .Q
       (________22162));
  nnd2s1 ___0_9_447629(.DIN1 (_____0__21995), .DIN2 (____09__21994), .Q
       (________22205));
  nnd2s1 ___9__447630(.DIN1 (________22091), .DIN2 (____0___21993), .Q
       (________22230));
  nor2s1 ___0__447631(.DIN1 (________22433), .DIN2 (________21758), .Q
       (________22432));
  xor2s1 ___9_0_447632(.DIN1 (outData[4]), .DIN2 (_________32606), .Q
       (___9_0__22455));
  nor2s1 ___9___447633(.DIN1 (_____0__23199), .DIN2 (___99___22533), .Q
       (____00__23802));
  nor2s1 ___9___447634(.DIN1 (____0___23716), .DIN2 (___9____23397), .Q
       (________23106));
  nor2s1 ___0___447635(.DIN1 (_____________________18665), .DIN2
       (________21431), .Q (________22142));
  hi1s1 ___0___447636(.DIN (__9_0___26707), .Q (___0____23471));
  hi1s1 ___999_447637(.DIN (___0____22596), .Q (___9____22496));
  nor2s1 ___0__447638(.DIN1 (________20561), .DIN2 (________21520), .Q
       (________22207));
  nor2s1 ___0__447639(.DIN1 (____0___21992), .DIN2 (________25524), .Q
       (___9_0__22465));
  nor2s1 ___0_447640(.DIN1 (___90___21544), .DIN2 (________21977), .Q
       (________22213));
  nnd2s1 ___0_9_447641(.DIN1 (___9____21593), .DIN2 (____0___21991), .Q
       (________22693));
  nor2s1 ___0___447642(.DIN1 (______18933), .DIN2 (___9____21588), .Q
       (____9___22352));
  nnd2s1 ___0_447643(.DIN1 (________21998), .DIN2 (________24216), .Q
       (___9____24250));
  nor2s1 ___0_0_447644(.DIN1 (____0___20888), .DIN2 (________21524), .Q
       (___9____22522));
  nnd2s1 ___0_0_447645(.DIN1 (___9____21555), .DIN2 (____0___21816), .Q
       (________22698));
  nor2s1 ___0___447646(.DIN1 (____0___21990), .DIN2 (____0___21989), .Q
       (________24651));
  nnd2s1 ___0___447647(.DIN1 (___9____21554), .DIN2 (____0___21988), .Q
       (________22741));
  nor2s1 ___0___447648(.DIN1 (___0____22603), .DIN2 (________25887), .Q
       (____90__24877));
  or2s1 ___0___447649(.DIN1 (____0___21987), .DIN2 (____0___21986), .Q
       (________22958));
  or2s1 ___0__447650(.DIN1 (________21131), .DIN2 (____9___21442), .Q
       (________22682));
  nor2s1 ___0__447651(.DIN1 (____0___23716), .DIN2 (____00__21985), .Q
       (_____0__26057));
  and2s1 ___9__447652(.DIN1 (________22091), .DIN2 (_____9__21209), .Q
       (___0_0__23455));
  nnd2s1 ___0___447653(.DIN1 (_____0__21523), .DIN2 (________21776), .Q
       (___9____22487));
  nnd2s1 ___9___447654(.DIN1 (________22093), .DIN2 (_____0__23199), .Q
       (___00____27213));
  and2s1 ___9___447655(.DIN1 (_____0__22138), .DIN2 (________22677), .Q
       (________22777));
  nor2s1 ___9__447656(.DIN1 (________23154), .DIN2 (___9____22495), .Q
       (__90____26275));
  nnd2s1 ___0___447657(.DIN1 (_____0__22014), .DIN2 (______0__35048),
       .Q (____09__22998));
  nor2s1 ___0___447658(.DIN1 (____9___22253), .DIN2 (___0____21709), .Q
       (____99__22445));
  nor2s1 ___0__447659(.DIN1 (________24659), .DIN2 (___9____22458), .Q
       (________22840));
  nnd2s1 ___0_0_447660(.DIN1 (________22026), .DIN2 (_________35072),
       .Q (__9_0___26422));
  nor2s1 ___9__447661(.DIN1 (________23233), .DIN2 (___0_0___27370), .Q
       (_____9__23544));
  nor2s1 ___0___447662(.DIN1 (____9___21984), .DIN2 (____9___21983), .Q
       (___9____23367));
  hi1s1 ___99__447663(.DIN (____9___21982), .Q (________22748));
  nnd2s1 ___0___447664(.DIN1 (________21967), .DIN2 (____0___20983), .Q
       (___90___22449));
  nor2s1 ___0__447665(.DIN1 (____9___21981), .DIN2 (____0___26053), .Q
       (_____0__25090));
  hi1s1 ___0___447666(.DIN (________22338), .Q (__9_00__26419));
  hi1s1 ___0___447667(.DIN (_____9___35020), .Q (________25872));
  nor2s1 ___0___447668(.DIN1 (____9___21980), .DIN2 (________21467), .Q
       (________22683));
  nor2s1 ___0___447669(.DIN1 (____9___21444), .DIN2 (________20252), .Q
       (_________32081));
  nor2s1 ___0___447670(.DIN1 (_____0__21298), .DIN2 (___9_9__21598), .Q
       (________25593));
  nor2s1 ___0___447671(.DIN1 (________19613), .DIN2 (_____9__21428), .Q
       (____0___24065));
  nor2s1 ___0___447672(.DIN1 (________22001), .DIN2 (________21403), .Q
       (________24619));
  or2s1 ___99__447673(.DIN1 (________19520), .DIN2 (___9____23397), .Q
       (___0__0__27802));
  hi1s1 ___000_447674(.DIN (________22217), .Q (__9_____26743));
  nor2s1 ___0__447675(.DIN1 (________21978), .DIN2 (________22002), .Q
       (___0____23512));
  nor2s1 ___0___447676(.DIN1 (____0____________0_), .DIN2
       (_____9__21437), .Q (________23932));
  nor2s1 ___0__447677(.DIN1 (________21857), .DIN2 (____9___21443), .Q
       (________24833));
  nnd2s1 ___99__447678(.DIN1 (________25734), .DIN2 (___9____26174), .Q
       (________25985));
  nnd2s1 ___0___447679(.DIN1 (________21918), .DIN2
       (____0____________0_), .Q (________23733));
  nnd2s1 ___990_447680(.DIN1 (___9____21611), .DIN2 (____9___19587), .Q
       (________24177));
  nnd2s1 ___0___447681(.DIN1 (________21432), .DIN2 (____9___21897), .Q
       (________25707));
  or2s1 ___0__447682(.DIN1 (_____9__25001), .DIN2 (_________35060), .Q
       (____9___23973));
  nor2s1 ___0___447683(.DIN1 (_____9__21894), .DIN2 (________21423), .Q
       (__9_____26452));
  nnd2s1 ___0___447684(.DIN1 (________21426), .DIN2
       (__________________0___18628), .Q (________22948));
  nor2s1 ___0__447685(.DIN1 (________24909), .DIN2 (________21433), .Q
       (________24113));
  nor2s1 ___0___447686(.DIN1 (_____9__21979), .DIN2 (________21925), .Q
       (_____0__25156));
  nor2s1 ___0___447687(.DIN1 (_____0__20923), .DIN2 (_________34159),
       .Q (___99___22529));
  nor2s1 ___0___447688(.DIN1 (______18933), .DIN2 (___9____21574), .Q
       (___90___22447));
  nor2s1 ___0_9_447689(.DIN1 (_____________________18664), .DIN2
       (___909__21552), .Q (__9_____26572));
  nor2s1 ___0_9_447690(.DIN1 (________21978), .DIN2 (________21977), .Q
       (___9____24263));
  and2s1 ___0_9_447691(.DIN1 (___9_9__21570), .DIN2
       (__________________0___18628), .Q (______0__28551));
  nor2s1 ___0_447692(.DIN1 (________21976), .DIN2 (________21975), .Q
       (___9____24277));
  nnd2s1 ___0___447693(.DIN1 (________21469), .DIN2 (inData[17]), .Q
       (____90__22436));
  nor2s1 ___0_9_447694(.DIN1 (________21974), .DIN2 (___90___21550), .Q
       (________24205));
  nor2s1 ___0_0_447695(.DIN1 (____0____________0_), .DIN2
       (___9____21562), .Q (____09__23983));
  nor2s1 ___99__447696(.DIN1 (___9_0__21561), .DIN2 (___9____21612), .Q
       (_________33333));
  nor2s1 ___0___447697(.DIN1 (inData[17]), .DIN2 (________21758), .Q
       (________22431));
  nnd2s1 ___0___447698(.DIN1 (___9____21576), .DIN2 (________21241), .Q
       (__9__0__26739));
  nor2s1 ___0__447699(.DIN1 (________20205), .DIN2 (___00___21638), .Q
       (_____0___32570));
  nor2s1 ___0__447700(.DIN1 (___9_9__20623), .DIN2 (________21529), .Q
       (_________33894));
  nor2s1 ___0___447701(.DIN1 (_____9__20464), .DIN2 (____9___21539), .Q
       (____00___31812));
  nor2s1 ___0___447702(.DIN1 (________20395), .DIN2 (________21434), .Q
       (____0____31872));
  nor2s1 ___0___447703(.DIN1 (________22434), .DIN2 (____9___21534), .Q
       (______0__30283));
  nor2s1 ___0___447704(.DIN1 (________20911), .DIN2 (________21973), .Q
       (_________32440));
  nor2s1 ___0___447705(.DIN1 (________21328), .DIN2 (________21836), .Q
       (_________33442));
  hi1s1 ___0___447706(.DIN (____9___21899), .Q (________22146));
  nor2s1 ___00__447707(.DIN1 (_____0__21971), .DIN2 (_____9__21970), .Q
       (________21972));
  nor2s1 ___00__447708(.DIN1 (________19520), .DIN2 (________23005), .Q
       (________21969));
  nnd2s1 ___0__447709(.DIN1 (________21967), .DIN2 (____00__20226), .Q
       (________21968));
  and2s1 ___00__447710(.DIN1 (________23273), .DIN2 (_________34447),
       .Q (________21966));
  hi1s1 ___999_447711(.DIN (__90_0__26318), .Q (________21965));
  and2s1 ___00_447712(.DIN1 (_________29668), .DIN2 (_____9__19186), .Q
       (________21964));
  nor2s1 ___00__447713(.DIN1 (________20441), .DIN2 (___9____21565), .Q
       (________21963));
  hi1s1 ___0___447714(.DIN (_____9__21961), .Q (_____0__21962));
  nnd2s1 ___0___447715(.DIN1 (________21959), .DIN2 (____0___19400), .Q
       (________21960));
  nor2s1 ___0___447716(.DIN1 (________22185), .DIN2 (________21957), .Q
       (________21958));
  nor2s1 ___0___447717(.DIN1 (___9____19712), .DIN2 (________21977), .Q
       (_____9__21956));
  hi1s1 ___0_0_447718(.DIN (____99__22894), .Q (________21954));
  nor2s1 ___0___447719(.DIN1 (________21036), .DIN2 (_____9__21532), .Q
       (________21953));
  hi1s1 ___999_447720(.DIN (________25774), .Q (________21952));
  nnd2s1 ___0___447721(.DIN1 (________21950), .DIN2 (________21949), .Q
       (________21951));
  and2s1 ___0___447722(.DIN1 (____9___25170), .DIN2 (________26099), .Q
       (_____0__21948));
  hi1s1 ___99_447723(.DIN (____9___23255), .Q (_____9__21947));
  nnd2s1 ___00_447724(.DIN1 (_________35052), .DIN2 (________19650), .Q
       (________21946));
  nor2s1 ___0___447725(.DIN1 (___9____21577), .DIN2 (___0____20775), .Q
       (________21945));
  nor2s1 ___00__447726(.DIN1 (________21427), .DIN2 (___9____21578), .Q
       (________21944));
  xor2s1 ___9___447727(.DIN1 (___0_____27735), .DIN2 (________21942),
       .Q (________21943));
  nor2s1 ______447728(.DIN1 (________21887), .DIN2 (___9_0__21617), .Q
       (________21941));
  nor2s1 ______447729(.DIN1 (________20353), .DIN2 (________21930), .Q
       (_____0__21940));
  nnd2s1 _______447730(.DIN1 (____9___21806), .DIN2 (________23222), .Q
       (_____9__21939));
  hi1s1 ___0___447731(.DIN (_____0__22128), .Q (________21938));
  hi1s1 _______447732(.DIN (________21935), .Q (________21936));
  hi1s1 _______447733(.DIN (_____9__21933), .Q (_____0__21934));
  nor2s1 ___0___447734(.DIN1 (________21755), .DIN2 (________21398), .Q
       (________21932));
  nor2s1 ___0___447735(.DIN1 (____0___21263), .DIN2 (________21930), .Q
       (________21931));
  and2s1 ___09__447736(.DIN1 (________23321), .DIN2 (________21928), .Q
       (________21929));
  or2s1 ___09__447737(.DIN1 (________20466), .DIN2 (_____0__21393), .Q
       (________21927));
  or2s1 ___0__447738(.DIN1 (________21796), .DIN2 (_____0__24173), .Q
       (________23218));
  nor2s1 ___0__447739(.DIN1 (________21926), .DIN2 (________21418), .Q
       (________22203));
  hi1s1 ___000_447740(.DIN (____9___22165), .Q (_____0__22962));
  hi1s1 ___000_447741(.DIN (__9_____26754), .Q (________22681));
  nor2s1 ___0___447742(.DIN1 (______18933), .DIN2 (___0____21643), .Q
       (________22124));
  nnd2s1 ___0___447743(.DIN1 (____0___21452), .DIN2 (__9_0), .Q
       (________22121));
  nnd2s1 ___0___447744(.DIN1 (___9_0__21599), .DIN2 (________21397), .Q
       (________22687));
  hi1s1 ___999_447745(.DIN (________22773), .Q (__90_0));
  nor2s1 ___0___447746(.DIN1 (________25901), .DIN2 (___0____23488), .Q
       (________22201));
  hi1s1 _______447747(.DIN (__9_____26381), .Q (________22340));
  nor2s1 ___0___447748(.DIN1 (___9____21575), .DIN2 (________21462), .Q
       (________22115));
  hi1s1 ___0___447749(.DIN (___9____26194), .Q (_____0__22337));
  hi1s1 _____9_447750(.DIN (_____0__22148), .Q (________22388));
  hi1s1 _____447751(.DIN (_____9__22336), .Q (__9__0__26356));
  xor2s1 ___9___447752(.DIN1 (____9___22073), .DIN2 (____0___19310), .Q
       (_________28628));
  nor2s1 _______447753(.DIN1 (________21391), .DIN2 (________25639), .Q
       (____9___22351));
  or2s1 ___0___447754(.DIN1 (________22136), .DIN2 (________21925), .Q
       (____9___22354));
  hi1s1 ___0___447755(.DIN (_____0__21924), .Q (____99__22355));
  and2s1 ___0___447756(.DIN1 (________21469), .DIN2 (________22334), .Q
       (________22331));
  nor2s1 ___0_0_447757(.DIN1 (_____0__22089), .DIN2 (_____9__21923), .Q
       (___0_0__22554));
  nor2s1 ___0___447758(.DIN1 (________23642), .DIN2 (________21143), .Q
       (________22853));
  hi1s1 _____447759(.DIN (_____0___35036), .Q (____90__22346));
  nor2s1 ___0___447760(.DIN1 (________21922), .DIN2 (________21973), .Q
       (___0____22590));
  hi1s1 _______447761(.DIN (________21921), .Q (___0_9__22563));
  nnd2s1 ___0___447762(.DIN1 (________25035), .DIN2 (__9_____26871), .Q
       (________22204));
  nnd2s1 ___0___447763(.DIN1 (________21920), .DIN2 (____9___21802), .Q
       (___9____22469));
  hi1s1 ___0___447764(.DIN (________25437), .Q (___9____22460));
  nor2s1 ___0__447765(.DIN1 (________21919), .DIN2 (___0____21678), .Q
       (___9_0__22517));
  hi1s1 ___0___447766(.DIN (________22369), .Q (_____9__23240));
  nnd2s1 ___0__447767(.DIN1 (_____0__21840), .DIN2 (________22116), .Q
       (___99___22532));
  hi1s1 ___0__447768(.DIN (___0_0__23500), .Q (________22393));
  nnd2s1 ___0___447769(.DIN1 (________21469), .DIN2 (___0____22601), .Q
       (___9____23362));
  nor2s1 ___099_447770(.DIN1 (___0____20722), .DIN2 (________21892), .Q
       (________22335));
  and2s1 ___0___447771(.DIN1 (____9___23707), .DIN2 (__9_____26631), .Q
       (____0___22630));
  or2s1 ___0___447772(.DIN1 (____0___22263), .DIN2 (__9_____26553), .Q
       (___9____22492));
  nnd2s1 ___0__447773(.DIN1 (________21918), .DIN2 (______18933), .Q
       (_____9__22117));
  nor2s1 ___0___447774(.DIN1 (________21917), .DIN2 (________21758), .Q
       (________22330));
  and2s1 ___0___447775(.DIN1 (__9_____26779), .DIN2 (________21916), .Q
       (________24505));
  or2s1 ___0___447776(.DIN1 (____00__19399), .DIN2 (________21915), .Q
       (___0_____27720));
  nor2s1 ___0___447777(.DIN1 (_____0__22924), .DIN2 (___0____21683), .Q
       (________23071));
  hi1s1 ___0___447778(.DIN (__99____27141), .Q (________23911));
  nnd2s1 ___0___447779(.DIN1 (________21959), .DIN2 (___00___22540), .Q
       (____0___23529));
  and2s1 ___9___447780(.DIN1 (__9_____26877), .DIN2 (________21916), .Q
       (________23040));
  hi1s1 _____0_447781(.DIN (_____0__21914), .Q (___9____25200));
  hi1s1 _______447782(.DIN (__9__0__26664), .Q (________23908));
  hi1s1 _______447783(.DIN (________24557), .Q (_____9__24719));
  nor2s1 ___0___447784(.DIN1 (________21476), .DIN2 (_________35040),
       .Q (____0___22813));
  nor2s1 ___0___447785(.DIN1 (_____9__24181), .DIN2 (_____9__25918), .Q
       (___9_0__22500));
  hi1s1 ___0__447786(.DIN (____09__21913), .Q (__9_0___26338));
  hi1s1 ___999_447787(.DIN (____09__22270), .Q (____9___22440));
  nnd2s1 ___0___447788(.DIN1 (____0___21912), .DIN2 (_________35064),
       .Q (________22686));
  or2s1 ___0__447789(.DIN1 (________24902), .DIN2 (____09__22365), .Q
       (____0___22811));
  nnd2s1 ___0___447790(.DIN1 (________25035), .DIN2 (____0___21911), .Q
       (___099__22625));
  nnd2s1 ___9___447791(.DIN1 (________23770), .DIN2 (___0____21708), .Q
       (____0___24522));
  nor2s1 ___0___447792(.DIN1 (__9_0___26897), .DIN2 (________21413), .Q
       (________24144));
  nor2s1 ______447793(.DIN1 (________21134), .DIN2 (________21396), .Q
       (________22344));
  or2s1 _______447794(.DIN1 (____00__20136), .DIN2 (________21930), .Q
       (________22969));
  nnd2s1 _____9_447795(.DIN1 (________21412), .DIN2 (________21794), .Q
       (____0___22364));
  nor2s1 ___0__447796(.DIN1 (__90_9__26308), .DIN2 (___0_____27430), .Q
       (____9___24515));
  and2s1 ___0_447797(.DIN1 (____0___21910), .DIN2 (____0___21909), .Q
       (_____9__22416));
  nor2s1 ___0___447798(.DIN1 (________20237), .DIN2 (___9____21621), .Q
       (____9___22439));
  or2s1 ___0___447799(.DIN1 (________22106), .DIN2 (________23136), .Q
       (___9____22510));
  or2s1 ___0_9_447800(.DIN1 (____0___21908), .DIN2 (________24680), .Q
       (________25499));
  nor2s1 ___0_9_447801(.DIN1 (____0___21907), .DIN2 (__9_____26350), .Q
       (_____0__23326));
  nor2s1 ___0_9_447802(.DIN1 (________23104), .DIN2 (_____0__26117), .Q
       (___9____22506));
  hi1s1 ___000_447803(.DIN (________22229), .Q (___0_____27894));
  nor2s1 _______447804(.DIN1 (________20345), .DIN2 (________21930), .Q
       (________25739));
  nnd2s1 ___0_9_447805(.DIN1 (________21767), .DIN2 (________22332), .Q
       (___9____24253));
  and2s1 ___0_0_447806(.DIN1 (________22150), .DIN2 (________24822), .Q
       (________23207));
  or2s1 ___0___447807(.DIN1 (________23284), .DIN2 (___9_0__26157), .Q
       (____9___23169));
  dffacs1 _________________0_447808(.CLRB (reset), .CLK (clk), .DIN
       (___9____21564), .QN (_____________0___18684));
  nor2s1 ___0___447809(.DIN1 (___0____25303), .DIN2 (________23233), .Q
       (________23773));
  nnd2s1 ___0___447810(.DIN1 (____0___21906), .DIN2 (____0___21905), .Q
       (________24452));
  nor2s1 ___0___447811(.DIN1 (________21508), .DIN2 (___0____21650), .Q
       (_____9__23868));
  hi1s1 ___0_9_447812(.DIN (________22817), .Q (___9____26220));
  nnd2s1 ___0_0_447813(.DIN1 (___00___21639), .DIN2
       (____0____________0_), .Q (___9_9__22464));
  nnd2s1 ___0___447814(.DIN1 (___9____21569), .DIN2 (____0___21905), .Q
       (____9___22353));
  nor2s1 ___0___447815(.DIN1 (________24105), .DIN2 (____0___26053), .Q
       (________24774));
  hi1s1 ___0_447816(.DIN (__9__0__26449), .Q (__9_____26686));
  nor2s1 ___0__447817(.DIN1 (_____9__21923), .DIN2 (________25901), .Q
       (________23149));
  nnd2s1 ___0___447818(.DIN1 (____9___21536), .DIN2 (___0____21664), .Q
       (___9____22462));
  nnd2s1 ___0___447819(.DIN1 (___909__22454), .DIN2 (___99___21629), .Q
       (____90__26137));
  nnd2s1 ___0___447820(.DIN1 (____00__21904), .DIN2 (____99__21903), .Q
       (________22398));
  nnd2s1 ___0___447821(.DIN1 (________23119), .DIN2 (__900_), .Q
       (___0____22577));
  nor2s1 ___0_0_447822(.DIN1 (________21096), .DIN2 (_____0__22855), .Q
       (___0____25307));
  xor2s1 ___0___447823(.DIN1 (________19087), .DIN2 (_________31295),
       .Q (___9____22478));
  nor2s1 ___0__447824(.DIN1 (____0____________0_), .DIN2
       (_____0__21465), .Q (___0____22567));
  nnd2s1 ___0___447825(.DIN1 (________21416), .DIN2 (_________35074),
       .Q (________24780));
  nor2s1 ___0___447826(.DIN1 (___9____21592), .DIN2 (________22002), .Q
       (________25442));
  or2s1 ___0___447827(.DIN1 (______0__35058), .DIN2 (________24132), .Q
       (___0_0__25290));
  nnd2s1 ___0___447828(.DIN1 (________21466), .DIN2 (________22131), .Q
       (_____0__24588));
  hi1s1 ___999_447829(.DIN (_____90__35018), .Q (___90___22450));
  nor2s1 ___0__447830(.DIN1 (________21407), .DIN2 (____9___21902), .Q
       (________24814));
  nor2s1 ___0___447831(.DIN1 (________20901), .DIN2 (___0_0__21641), .Q
       (________25910));
  nor2s1 ___0___447832(.DIN1 (____0____________0_), .DIN2
       (___9____21601), .Q (___0____22571));
  nor2s1 ___0___447833(.DIN1 (___0____21659), .DIN2 (________21996), .Q
       (________24549));
  nor2s1 ___0___447834(.DIN1 (____0___21362), .DIN2 (___9____21615), .Q
       (________26008));
  nnd2s1 ___0___447835(.DIN1 (________21430), .DIN2 (________21375), .Q
       (________23097));
  nnd2s1 ___0___447836(.DIN1 (__9_____26496), .DIN2 (____9___21901), .Q
       (___0____25336));
  nor2s1 ___0__447837(.DIN1 (________22113), .DIN2 (________21459), .Q
       (__9__9__27073));
  nor2s1 ___0___447838(.DIN1 (____9___21900), .DIN2 (_____9__21464), .Q
       (___0_0__22573));
  nnd2s1 ___0__447839(.DIN1 (____9___21538), .DIN2 (_____0__21821), .Q
       (________24459));
  nnd2s1 ___0___447840(.DIN1 (___9_9__21616), .DIN2 (___0____21677), .Q
       (__9_____26591));
  and2s1 ___0___447841(.DIN1 (___0_0__21667), .DIN2 (________22149), .Q
       (________24944));
  nor2s1 ___0__447842(.DIN1 (____9___21898), .DIN2 (________21925), .Q
       (___9____24313));
  nnd2s1 ___0___447843(.DIN1 (___9____21619), .DIN2 (_____0__22118), .Q
       (________24939));
  nor2s1 ___0___447844(.DIN1 (________19613), .DIN2 (________21517), .Q
       (________23541));
  nnd2s1 ___0_9_447845(.DIN1 (________21460), .DIN2 (____9___21897), .Q
       (__9_____26917));
  hi1s1 ___0___447846(.DIN (____9___21896), .Q (___9____26200));
  nor2s1 _____0_447847(.DIN1 (________19910), .DIN2 (________21930), .Q
       (__9_____26935));
  nor2s1 _______447848(.DIN1 (__9_____26650), .DIN2 (___0____24412), .Q
       (____9___23885));
  nor2s1 ___0_447849(.DIN1 (________21388), .DIN2 (___9____21606), .Q
       (________25983));
  nor2s1 ___0___447850(.DIN1 (____0___21167), .DIN2 (________21531), .Q
       (___0____22579));
  nnd2s1 ___0___447851(.DIN1 (_____0__21514), .DIN2 (___0____20727), .Q
       (______9__34123));
  hi1s1 ___0___447852(.DIN (____90__21895), .Q (__9_____27023));
  nnd2s1 ___0_0_447853(.DIN1 (___0____24393), .DIN2 (________22370), .Q
       (________22424));
  nor2s1 ___0___447854(.DIN1 (_____9__21894), .DIN2 (___9____21567), .Q
       (___9____26182));
  nor2s1 _______447855(.DIN1 (________20307), .DIN2 (___99___21626), .Q
       (__9_____26487));
  nnd2s1 ___0___447856(.DIN1 (___90___21547), .DIN2 (____0___21988), .Q
       (________24001));
  nnd2s1 ___0___447857(.DIN1 (___90___21545), .DIN2
       (_____________________18665), .Q (____0___22360));
  nor2s1 _____0_447858(.DIN1 (________21144), .DIN2 (________21892), .Q
       (__9__0__26749));
  hi1s1 ___0___447859(.DIN (________21891), .Q (________25389));
  nor2s1 ___0___447860(.DIN1 (________21890), .DIN2 (_____0__21419), .Q
       (____00___32758));
  nor2s1 ___0___447861(.DIN1 (____9___21071), .DIN2 (________21408), .Q
       (_____0__25967));
  nor2s1 _____447862(.DIN1 (________21421), .DIN2 (________21339), .Q
       (__9_____26597));
  nor2s1 ___0_447863(.DIN1 (________21889), .DIN2 (________21404), .Q
       (__9_____26905));
  hi1s1 ___0_9_447864(.DIN (________21888), .Q (___00____27200));
  nor2s1 ___0_0_447865(.DIN1 (________21887), .DIN2 (___00___21634), .Q
       (__9_____26838));
  hi1s1 ___0___447866(.DIN (________21886), .Q (__9_____26953));
  nor2s1 _______447867(.DIN1 (____9___20131), .DIN2 (________21930), .Q
       (___0090__27257));
  nor2s1 ___0_447868(.DIN1 (________20868), .DIN2 (____9___21902), .Q
       (___0_____27483));
  nor2s1 ___0_0_447869(.DIN1 (_____0__21475), .DIN2 (___9_0__21590), .Q
       (__9_9___26888));
  nnd2s1 ___0_0_447870(.DIN1 (________21414), .DIN2 (____9___21897), .Q
       (__9_____26862));
  nor2s1 ___0___447871(.DIN1 (________21337), .DIN2 (___9_9__21625), .Q
       (_________31951));
  hi1s1 _______447872(.DIN (_____9__21884), .Q (_____9___28891));
  nor2s1 ___0___447873(.DIN1 (________19570), .DIN2 (________23875), .Q
       (________21883));
  nor2s1 ___0___447874(.DIN1 (_____9__22215), .DIN2 (________21151), .Q
       (________21882));
  hi1s1 _______447875(.DIN (___0_____27430), .Q (________21881));
  nor2s1 ___09__447876(.DIN1 (________21879), .DIN2 (________21746), .Q
       (________21880));
  nnd2s1 ___09__447877(.DIN1 (_____0__21183), .DIN2 (_____0__20107), .Q
       (________21878));
  nor2s1 ___09_447878(.DIN1 (outData[18]), .DIN2 (_________34116), .Q
       (________21877));
  hi1s1 _______447879(.DIN (________22381), .Q (_____0__21876));
  and2s1 ___09__447880(.DIN1 (________21866), .DIN2 (________20910), .Q
       (_____9__21875));
  nor2s1 ___09__447881(.DIN1 (________20430), .DIN2 (________21185), .Q
       (________21874));
  hi1s1 _______447882(.DIN (______0__28751), .Q (________21873));
  and2s1 ___09__447883(.DIN1 (________21871), .DIN2 (___0_9__21657), .Q
       (________21872));
  nnd2s1 ___090_447884(.DIN1 (____00__21811), .DIN2 (_________34448),
       .Q (________21870));
  nor2s1 ___0_9_447885(.DIN1 (________20370), .DIN2 (_________34116),
       .Q (________21869));
  nnd2s1 ___0___447886(.DIN1 (_____9__21249), .DIN2 (inData[26]), .Q
       (________21868));
  nnd2s1 ___0___447887(.DIN1 (________21866), .DIN2 (________22663), .Q
       (_____9__21867));
  nor2s1 ___0___447888(.DIN1 (_____0__21230), .DIN2 (___0____21691), .Q
       (________21865));
  nor2s1 ___0___447889(.DIN1 (_____9__21229), .DIN2 (________21741), .Q
       (________21864));
  nnd2s1 ___0___447890(.DIN1 (_________35070), .DIN2 (________21233),
       .Q (________21863));
  nor2s1 ___0___447891(.DIN1 (___00___19771), .DIN2 (________21116), .Q
       (________21861));
  nor2s1 ___0___447892(.DIN1 (_____9__19350), .DIN2 (________21152), .Q
       (________21860));
  nnd2s1 ___0_0_447893(.DIN1 (________21244), .DIN2 (________21016), .Q
       (_____0__21859));
  nor2s1 ___00__447894(.DIN1 (________21857), .DIN2 (________21296), .Q
       (_____9__21858));
  nnd2s1 ___00__447895(.DIN1 (________21304), .DIN2 (________21855), .Q
       (________21856));
  nnd2s1 ___00__447896(.DIN1 (_____0__21270), .DIN2 (____9___21159), .Q
       (________21854));
  xor2s1 ___9_9_447897(.DIN1 (_________18850), .DIN2 (_________29500),
       .Q (________21853));
  xor2s1 ___9_0_447898(.DIN1 (_________29688), .DIN2 (_________31326),
       .Q (________21852));
  nnd2s1 ___00__447899(.DIN1 (________21850), .DIN2 (___0____21674), .Q
       (________21851));
  and2s1 ___00__447900(.DIN1 (____9___21254), .DIN2 (________20271), .Q
       (_____0__21849));
  nnd2s1 ___0___447901(.DIN1 (_____9__21297), .DIN2 (________21847), .Q
       (________21848));
  or2s1 ___0___447902(.DIN1 (________21845), .DIN2 (___0____21668), .Q
       (________21846));
  nnd2s1 ___0___447903(.DIN1 (________21329), .DIN2 (_____9__19871), .Q
       (________21844));
  or2s1 ___00__447904(.DIN1 (________21123), .DIN2 (_____9__21239), .Q
       (________21843));
  nnd2s1 ___0_0_447905(.DIN1 (_____0__21739), .DIN2 (________20204), .Q
       (________21842));
  hi1s1 ___0___447906(.DIN (_____0__21840), .Q (________21841));
  hi1s1 ___0___447907(.DIN (________21838), .Q (_____9__21839));
  nor2s1 ___00_447908(.DIN1 (________22113), .DIN2 (________21242), .Q
       (________21837));
  nor2s1 ___00_447909(.DIN1 (________21245), .DIN2 (________21284), .Q
       (________21835));
  and2s1 ___00__447910(.DIN1 (____9___21251), .DIN2 (________22110), .Q
       (________21834));
  nnd2s1 ___00_447911(.DIN1 (________21097), .DIN2 (________19997), .Q
       (________21833));
  nnd2s1 ___447912(.DIN1 (_____0__21831), .DIN2 (____9___21255), .Q
       (________21832));
  nnd2s1 ___0_0_447913(.DIN1 (________21289), .DIN2 (________19619), .Q
       (_____9__21830));
  nnd2s1 ___0___447914(.DIN1 (_____9__21307), .DIN2 (________21237), .Q
       (________21829));
  and2s1 ___0___447915(.DIN1 (________21128), .DIN2 (________20211), .Q
       (________21828));
  nnd2s1 ___0___447916(.DIN1 (____0___21261), .DIN2 (___0____21694), .Q
       (________21827));
  or2s1 ___0__447917(.DIN1 (________21890), .DIN2 (________21246), .Q
       (________21826));
  nnd2s1 ___0___447918(.DIN1 (____9___21160), .DIN2 (________21824), .Q
       (________21825));
  nnd2s1 ___0___447919(.DIN1 (________21417), .DIN2 (____0___21819), .Q
       (________21823));
  nnd2s1 ___0___447920(.DIN1 (____90__21250), .DIN2 (_____0__21821), .Q
       (________21822));
  nnd2s1 ___0___447921(.DIN1 (_____0__21147), .DIN2 (____0___21819), .Q
       (____09__21820));
  xor2s1 ___0___447922(.DIN1 (_____________18900), .DIN2
       (_________35086), .Q (____0___21818));
  xor2s1 ___9___447923(.DIN1 (____0___19120), .DIN2 (_________31134),
       .Q (_____0__22319));
  nnd2s1 _______447924(.DIN1 (________21286), .DIN2 (________21784), .Q
       (________21891));
  hi1s1 ___0___447925(.DIN (_____0__22099), .Q (________22219));
  hi1s1 _____0_447926(.DIN (___909__22454), .Q (___9____26171));
  nor2s1 ___0__447927(.DIN1 (________21742), .DIN2 (____9___21807), .Q
       (________22208));
  nnd2s1 ___0___447928(.DIN1 (________21850), .DIN2 (________21435), .Q
       (________22228));
  nnd2s1 ___0_9_447929(.DIN1 (_____9__21190), .DIN2 (____0___21812), .Q
       (________22226));
  nor2s1 ___0_0_447930(.DIN1 (________21978), .DIN2 (________21106), .Q
       (_____9__22233));
  nor2s1 ___0_0_447931(.DIN1 (________20278), .DIN2 (___0____21701), .Q
       (_____9__21961));
  or2s1 ___0___447932(.DIN1 (________25582), .DIN2 (____0___21817), .Q
       (________22232));
  xor2s1 ___0___447933(.DIN1 (___0___18986), .DIN2 (_________33278), .Q
       (________22296));
  nnd2s1 ___0___447934(.DIN1 (________21795), .DIN2 (___9____21624), .Q
       (_____0__21924));
  nnd2s1 ___0__447935(.DIN1 (________21275), .DIN2 (________21785), .Q
       (____09__21913));
  nnd2s1 ___0___447936(.DIN1 (___9____22505), .DIN2 (___00___20702), .Q
       (________22325));
  nor2s1 ___0___447937(.DIN1 (___0____21699), .DIN2 (________21285), .Q
       (____9___21982));
  nor2s1 ___0___447938(.DIN1 (___9____19718), .DIN2 (________21091), .Q
       (_____9__24847));
  nnd2s1 ___0_9_447939(.DIN1 (___0____21673), .DIN2 (________21530), .Q
       (_____0__22224));
  nnd2s1 ___0___447940(.DIN1 (_____9__21792), .DIN2 (________21778), .Q
       (________22214));
  nnd2s1 _______447941(.DIN1 (________21187), .DIN2 (________19257), .Q
       (_____0__21914));
  nor2s1 ___0___447942(.DIN1 (____0___21815), .DIN2 (________22106), .Q
       (_____9__23099));
  hi1s1 ___0___447943(.DIN (_________31956), .Q (___0____22546));
  hi1s1 ___0__447944(.DIN (___0____21656), .Q (________21955));
  and2s1 ___09__447945(.DIN1 (____0___21814), .DIN2 (________21789), .Q
       (________22151));
  or2s1 ___09__447946(.DIN1 (________20860), .DIN2 (___0____24368), .Q
       (__90____26265));
  and2s1 ___09__447947(.DIN1 (________21386), .DIN2 (____0___21911), .Q
       (_____9__22137));
  or2s1 ___447948(.DIN1 (________21142), .DIN2 (____0___21813), .Q
       (_____0__24219));
  nnd2s1 ___099_447949(.DIN1 (________21111), .DIN2 (____0___21812), .Q
       (________22145));
  and2s1 ____447950(.DIN1 (____00__21811), .DIN2 (____99__21810), .Q
       (_____0__22192));
  nnd2s1 ____00_447951(.DIN1 (________25817), .DIN2 (________21149), .Q
       (________23198));
  nnd2s1 ____0__447952(.DIN1 (________21179), .DIN2 (________21777), .Q
       (________22225));
  nnd2s1 ___0___447953(.DIN1 (____0___21168), .DIN2 (______18933), .Q
       (_____0__22327));
  nnd2s1 ___0___447954(.DIN1 (____00__24792), .DIN2 (____9___21809), .Q
       (___9____26179));
  hi1s1 ______447955(.DIN (____0___22363), .Q (____9___26043));
  nnd2s1 ___0_9_447956(.DIN1 (________21090), .DIN2 (____9___21808), .Q
       (____09__22270));
  nor2s1 ___0___447957(.DIN1 (________20311), .DIN2 (____9___21807), .Q
       (________22120));
  nor2s1 ___0___447958(.DIN1 (____0___21724), .DIN2 (____9___21157), .Q
       (________22338));
  nnd2s1 ____447959(.DIN1 (________21420), .DIN2 (________21385), .Q
       (__99____27141));
  hi1s1 ____0__447960(.DIN (____9___21806), .Q (___990__25261));
  hi1s1 ___0__447961(.DIN (____9___21805), .Q (_____0__24946));
  hi1s1 ___0___447962(.DIN (______0__35048), .Q (________22421));
  hi1s1 ___0___447963(.DIN (___9____26223), .Q (________23193));
  hi1s1 ___0___447964(.DIN (______9__33828), .Q (_________33264));
  hi1s1 ___000_447965(.DIN (___90___22451), .Q (___0_9__25318));
  hi1s1 ___0___447966(.DIN (________22122), .Q (__9_____26525));
  hi1s1 ___0__447967(.DIN (________23698), .Q (____9___23163));
  nor2s1 ___0___447968(.DIN1 (____9___21804), .DIN2 (________21125), .Q
       (_____9__22280));
  nnd2s1 _______447969(.DIN1 (___0____21693), .DIN2 (________21050), .Q
       (_____9__22336));
  hi1s1 ____0__447970(.DIN (________23922), .Q (__9_____26435));
  nnd2s1 ___0___447971(.DIN1 (____0___21264), .DIN2 (________19257), .Q
       (___0_____27973));
  nnd2s1 ___0___447972(.DIN1 (____0___21266), .DIN2 (____9___21803), .Q
       (________22217));
  nnd2s1 ___0_0_447973(.DIN1 (__9_____26871), .DIN2 (____9___21802), .Q
       (___0____22565));
  nnd2s1 ___0___447974(.DIN1 (___09___23526), .DIN2 (____90__23792), .Q
       (________22820));
  and2s1 ___0_447975(.DIN1 (________26059), .DIN2 (________23770), .Q
       (___909__24248));
  nnd2s1 ___0__447976(.DIN1 (________21787), .DIN2 (____90__21801), .Q
       (________22229));
  nnd2s1 ___0_0_447977(.DIN1 (_____9__21800), .DIN2 (________21799), .Q
       (____0___22268));
  nor2s1 ___0___447978(.DIN1 (________21793), .DIN2 (____0___24888), .Q
       (_____0__23601));
  nnd2s1 ___0___447979(.DIN1 (____9___21348), .DIN2 (________23875), .Q
       (________24583));
  hi1s1 _______447980(.DIN (________21798), .Q (_____9__23142));
  nnd2s1 ___0___447981(.DIN1 (________21299), .DIN2 (________21797), .Q
       (________22209));
  nor2s1 ___0_9_447982(.DIN1 (________26000), .DIN2 (________21796), .Q
       (________25378));
  nnd2s1 ___0___447983(.DIN1 (________21795), .DIN2 (________21480), .Q
       (___0____22607));
  nor2s1 ___0___447984(.DIN1 (____0___21082), .DIN2 (___09___24420), .Q
       (________25452));
  nor2s1 ___0_0_447985(.DIN1 (________21976), .DIN2 (____09__21269), .Q
       (________22231));
  nnd2s1 ___0_0_447986(.DIN1 (____0___21081), .DIN2 (________21509), .Q
       (___0_____27905));
  nnd2s1 ___0_447987(.DIN1 (________21181), .DIN2 (________21373), .Q
       (_____9__22345));
  nnd2s1 ____0__447988(.DIN1 (_____0__21317), .DIN2 (________21794), .Q
       (_____0__22128));
  nnd2s1 ____0__447989(.DIN1 (_____0__21374), .DIN2 (____0___23620), .Q
       (____90__23704));
  nor2s1 ____0__447990(.DIN1 (________21793), .DIN2 (____0___21815), .Q
       (_____9__25528));
  nnd2s1 ____0__447991(.DIN1 (________21871), .DIN2 (____9___20877), .Q
       (____9___22167));
  nnd2s1 ____0__447992(.DIN1 (___0____21697), .DIN2 (________21218), .Q
       (___0____22598));
  or2s1 ___0___447993(.DIN1 (________24221), .DIN2 (________26059), .Q
       (_________28626));
  nnd2s1 ___0___447994(.DIN1 (________21775), .DIN2 (________22339), .Q
       (____9___23795));
  nnd2s1 ___0___447995(.DIN1 (____9___21072), .DIN2 (____9___19587), .Q
       (__9_____26401));
  nor2s1 ___0_9_447996(.DIN1 (____0____________0_), .DIN2
       (________21121), .Q (___0____22596));
  nor2s1 ___0___447997(.DIN1 (____0____________0_), .DIN2
       (____0___21268), .Q (________23318));
  nor2s1 ___0___447998(.DIN1 (________21750), .DIN2 (________21154), .Q
       (_____9__25684));
  nnd2s1 ___0___447999(.DIN1 (________21247), .DIN2
       (____0____________0_), .Q (___0____23508));
  nor2s1 ___0__448000(.DIN1 (________19613), .DIN2 (_____0__21729), .Q
       (________24845));
  nnd2s1 ___0_9_448001(.DIN1 (_____9__21792), .DIN2 (________21486), .Q
       (________22773));
  nnd2s1 ___0___448002(.DIN1 (________25803), .DIN2 (________21791), .Q
       (________26094));
  nnd2s1 ____0__448003(.DIN1 (________21790), .DIN2 (________21789), .Q
       (_____0__25997));
  nor2s1 ___0___448004(.DIN1 (________24475), .DIN2 (____9___22986), .Q
       (________24859));
  nor2s1 ___0_0_448005(.DIN1 (________21788), .DIN2 (________21781), .Q
       (__9_____26754));
  nor2s1 ___0__448006(.DIN1 (________21788), .DIN2 (___0_9__21695), .Q
       (___9____26194));
  nnd2s1 ___0_0_448007(.DIN1 (________21787), .DIN2 (_____0__21365), .Q
       (____9___22165));
  hi1s1 _______448008(.DIN (________21786), .Q (__90_9));
  nor2s1 ___0_9_448009(.DIN1 (____9___21804), .DIN2 (________21771), .Q
       (________22817));
  nor2s1 ___0___448010(.DIN1 (_____________________18666), .DIN2
       (________21325), .Q (________25710));
  nnd2s1 ___0___448011(.DIN1 (________21301), .DIN2 (________21785), .Q
       (___9____23396));
  nnd2s1 ____0_448012(.DIN1 (_____0__21773), .DIN2 (________21193), .Q
       (________22954));
  nnd2s1 _____0_448013(.DIN1 (________21294), .DIN2 (________21784), .Q
       (__9_0___26707));
  hi1s1 ___0__448014(.DIN (_____0__21783), .Q (___9____26163));
  nor2s1 ____0__448015(.DIN1 (________21312), .DIN2 (____0___21813), .Q
       (________22249));
  nor2s1 ___0___448016(.DIN1 (_____9__21782), .DIN2 (_____9__25145), .Q
       (________22739));
  or2s1 ___0___448017(.DIN1 (________26125), .DIN2 (___0_0__21676), .Q
       (________26130));
  nor2s1 ___0_0_448018(.DIN1 (________21323), .DIN2 (________21781), .Q
       (__9__0__26449));
  or2s1 ___0___448019(.DIN1 (___00___20701), .DIN2 (________21780), .Q
       (____00__24886));
  hi1s1 ___0___448020(.DIN (________21779), .Q (__9_9___26414));
  nnd2s1 ___0___448021(.DIN1 (________21132), .DIN2 (________21778), .Q
       (________24865));
  nnd2s1 ____0__448022(.DIN1 (___0____21687), .DIN2 (________21777), .Q
       (____9___23794));
  nor2s1 _______448023(.DIN1 (________22017), .DIN2 (________21101), .Q
       (________22189));
  nor2s1 ___0_9_448024(.DIN1 (________22113), .DIN2 (____9___21252), .Q
       (__90_0__26318));
  nnd2s1 ___0___448025(.DIN1 (________21088), .DIN2 (________22341), .Q
       (________25672));
  nnd2s1 _______448026(.DIN1 (________21177), .DIN2 (________21776), .Q
       (_________28294));
  nnd2s1 ___0_448027(.DIN1 (________21775), .DIN2 (________21774), .Q
       (________25774));
  nnd2s1 ______448028(.DIN1 (________21277), .DIN2 (________21378), .Q
       (__9__0__26494));
  and2s1 ___0___448029(.DIN1 (________21295), .DIN2 (________21824), .Q
       (________25478));
  nnd2s1 _______448030(.DIN1 (_____0__21773), .DIN2 (________21216), .Q
       (___0_0__23500));
  nor2s1 ___0__448031(.DIN1 (_____9__21772), .DIN2 (________21771), .Q
       (____99__22894));
  nnd2s1 ___0__448032(.DIN1 (________21309), .DIN2 (___9_9__20643), .Q
       (______0__31325));
  nnd2s1 _______448033(.DIN1 (____99__21165), .DIN2
       (_____________________18662), .Q (________21770));
  nnd2s1 ___00__448034(.DIN1 (____0___21262), .DIN2 (________20435), .Q
       (________21769));
  hi1s1 _______448035(.DIN (________21767), .Q (________21768));
  hi1s1 _______448036(.DIN (________21765), .Q (________21766));
  hi1s1 _______448037(.DIN (___9____22482), .Q (________21764));
  hi1s1 _____9_448038(.DIN (________21925), .Q (_____0__21763));
  nnd2s1 ___00__448039(.DIN1 (____0___21169), .DIN2
       (____0_________________18658), .Q (________21762));
  or2s1 ___00__448040(.DIN1 (_____________0___18697), .DIN2
       (________21760), .Q (________21761));
  nnd2s1 ___0___448041(.DIN1 (________22425), .DIN2 (________23814), .Q
       (________21759));
  or2s1 _______448042(.DIN1 (_____9__21756), .DIN2 (________21755), .Q
       (_____0__21757));
  nor2s1 ___009_448043(.DIN1 (________20347), .DIN2 (____9___21807), .Q
       (________21754));
  nnd2s1 ______448044(.DIN1 (____9___21164), .DIN2 (_____9__21278), .Q
       (________21753));
  nnd2s1 _______448045(.DIN1 (________21273), .DIN2
       (_____________________18662), .Q (________21752));
  nnd2s1 _______448046(.DIN1 (____9___21163), .DIN2 (_____0__21821), .Q
       (________21751));
  nor2s1 _____448047(.DIN1 (___90___21546), .DIN2 (________21135), .Q
       (_____0__21749));
  nnd2s1 _____9_448048(.DIN1 (_____9__21112), .DIN2 (________22332), .Q
       (_____9__21748));
  nor2s1 _____0_448049(.DIN1 (________20389), .DIN2 (________21746), .Q
       (________21747));
  nor2s1 _____0_448050(.DIN1 (________19652), .DIN2 (_________32487),
       .Q (________21745));
  nor2s1 _______448051(.DIN1 (________21198), .DIN2 (________21746), .Q
       (________21744));
  nor2s1 _______448052(.DIN1 (________21742), .DIN2 (________21741), .Q
       (________21743));
  and2s1 ______448053(.DIN1 (_____0__21739), .DIN2 (____0___21360), .Q
       (________21740));
  nor2s1 _______448054(.DIN1 (_______18991), .DIN2 (_________34116), .Q
       (_____9__21738));
  nnd2s1 ___0___448055(.DIN1 (__9_____26456), .DIN2 (_____9__19648), .Q
       (________21737));
  nor2s1 _______448056(.DIN1 (________20841), .DIN2 (________22132), .Q
       (________21736));
  nor2s1 ___0___448057(.DIN1 (________25015), .DIN2 (___0____21682), .Q
       (________21735));
  and2s1 _______448058(.DIN1 (________21733), .DIN2 (________21109), .Q
       (________21734));
  nor2s1 _______448059(.DIN1 (________21114), .DIN2 (________21741), .Q
       (________21732));
  nor2s1 ___0___448060(.DIN1 (________21730), .DIN2 (_____0__21729), .Q
       (________21731));
  nnd2s1 ___0___448061(.DIN1 (____0___22812), .DIN2 (___0____23448), .Q
       (____09__21728));
  nnd2s1 ___0___448062(.DIN1 (________21290), .DIN2 (________19480), .Q
       (____0___21727));
  nnd2s1 ___0___448063(.DIN1 (________22412), .DIN2 (________23814), .Q
       (____0___21726));
  nor2s1 ___0___448064(.DIN1 (____0___21724), .DIN2 (____9___21258), .Q
       (____0___21725));
  nnd2s1 ___0___448065(.DIN1 (________21336), .DIN2 (__900_), .Q
       (____0___21723));
  or2s1 ___0___448066(.DIN1 (___9____23389), .DIN2 (__9_____26456), .Q
       (____0___21722));
  xor2s1 ___0___448067(.DIN1 (________21942), .DIN2 (____9____30874),
       .Q (____0___21721));
  hi1s1 ___0___448068(.DIN (____00__21719), .Q (____0___21720));
  nor2s1 ___0__448069(.DIN1 (____0___24888), .DIN2 (____0___21992), .Q
       (___099__21718));
  nnd2s1 ___009_448070(.DIN1 (____9___21439), .DIN2 (___09___21716), .Q
       (___09___21717));
  nnd2s1 ___0___448071(.DIN1 (_____0__21308), .DIN2 (________21777), .Q
       (___09___21715));
  hi1s1 ___0___448072(.DIN (___0_____27804), .Q (___09___21714));
  hi1s1 ___0___448073(.DIN (___09___21712), .Q (___09___21713));
  hi1s1 ___0__448074(.DIN (___0____21709), .Q (___0____21710));
  nnd2s1 ___09__448075(.DIN1 (____0___21172), .DIN2 (___0____21690), .Q
       (___0____21707));
  hi1s1 ___000_448076(.DIN (__9_____26784), .Q (___0____21706));
  hi1s1 _____9_448077(.DIN (________23273), .Q (___0_0__21705));
  hi1s1 _______448078(.DIN (___0____21703), .Q (___0____21704));
  hi1s1 _____9_448079(.DIN (________25887), .Q (___0____21702));
  nor2s1 ___0___448080(.DIN1 (________21228), .DIN2 (___0____21701), .Q
       (________22210));
  nnd2s1 _____0_448081(.DIN1 (___0____21681), .DIN2 (________20917), .Q
       (________22133));
  nor2s1 _____0_448082(.DIN1 (___0____21700), .DIN2 (________21092), .Q
       (_____9__21933));
  nor2s1 ___0__448083(.DIN1 (___0____21699), .DIN2 (________21110), .Q
       (________22159));
  hi1s1 ___0___448084(.DIN (___9____23394), .Q (________22194));
  nnd2s1 ___0_448085(.DIN1 (________21302), .DIN2 (___0____21698), .Q
       (________21888));
  nnd2s1 _____448086(.DIN1 (___0____21697), .DIN2 (___9____19721), .Q
       (________21935));
  nor2s1 ___0__448087(.DIN1 (___0_0__21696), .DIN2 (___0_9__21695), .Q
       (____9___21896));
  hi1s1 ___0__448088(.DIN (____9___25170), .Q (____9___22257));
  hi1s1 ___0___448089(.DIN (__9_0___26517), .Q (________23700));
  nor2s1 _______448090(.DIN1 (________21501), .DIN2 (________21117), .Q
       (_____9__21884));
  nnd2s1 ______448091(.DIN1 (___0____21697), .DIN2 (___0____21694), .Q
       (____09__22181));
  nor2s1 _______448092(.DIN1 (________21495), .DIN2 (________21411), .Q
       (________22114));
  and2s1 _______448093(.DIN1 (___0____21693), .DIN2 (________21785), .Q
       (________22135));
  hi1s1 ___0___448094(.DIN (__90_9__26308), .Q (________22955));
  hi1s1 _____0_448095(.DIN (________25392), .Q (_____0__22700));
  or2s1 _______448096(.DIN1 (___0____21692), .DIN2 (___0____21691), .Q
       (________22125));
  nnd2s1 ______448097(.DIN1 (________21137), .DIN2 (___0____21690), .Q
       (________21937));
  hi1s1 _______448098(.DIN (________22967), .Q (________22218));
  hi1s1 _______448099(.DIN (________25158), .Q (________22144));
  xor2s1 ___0__448100(.DIN1 (___0____21689), .DIN2 (______9__33856), .Q
       (_________30231));
  hi1s1 _______448101(.DIN (________22185), .Q (________22882));
  hi1s1 _______448102(.DIN (_________34159), .Q (________22244));
  hi1s1 ___99__448103(.DIN (___0____21688), .Q (___900__22446));
  nor2s1 ___0___448104(.DIN1 (________21221), .DIN2 (________25064), .Q
       (________22140));
  nnd2s1 _______448105(.DIN1 (___0____21687), .DIN2 (_____0__20156), .Q
       (________21921));
  hi1s1 _______448106(.DIN (__9_____26779), .Q (__9__9__26757));
  nnd2s1 ______448107(.DIN1 (________21330), .DIN2 (________22341), .Q
       (____90__21895));
  hi1s1 _______448108(.DIN (___0_0__21686), .Q (________22134));
  hi1s1 _______448109(.DIN (__9_9___26791), .Q (____9___22170));
  hi1s1 _____9_448110(.DIN (________24724), .Q (________22130));
  hi1s1 _____448111(.DIN (________22685), .Q (__90____26273));
  hi1s1 ___0___448112(.DIN (________25734), .Q (____9___22441));
  hi1s1 _______448113(.DIN (________21957), .Q (_____9__22884));
  hi1s1 _______448114(.DIN (___0__0__27287), .Q (____9___22349));
  hi1s1 _____9_448115(.DIN (___0_9__21685), .Q (___0____23498));
  hi1s1 _____0_448116(.DIN (_____0__23028), .Q (________22126));
  hi1s1 _______448117(.DIN (_________35056), .Q (___9_0__25184));
  hi1s1 ______448118(.DIN (____00__21904), .Q (___90___26154));
  and2s1 ___0___448119(.DIN1 (_____9__21146), .DIN2 (___0____21684), .Q
       (________22222));
  hi1s1 _____448120(.DIN (___0____21683), .Q (___0____24403));
  nor2s1 ___0_448121(.DIN1 (___0____21682), .DIN2 (________25782), .Q
       (________22143));
  nor2s1 _______448122(.DIN1 (_____0__20207), .DIN2 (________21293), .Q
       (________24642));
  hi1s1 ___0___448123(.DIN (________22152), .Q (________26084));
  and2s1 _______448124(.DIN1 (___0____21681), .DIN2 (________21511), .Q
       (_____0__24772));
  nor2s1 ___0___448125(.DIN1 (________23757), .DIN2 (________23875), .Q
       (__90____26262));
  nnd2s1 _______448126(.DIN1 (________21099), .DIN2 (________21776), .Q
       (________21886));
  or2s1 _______448127(.DIN1 (___0____21680), .DIN2 (_________34116), .Q
       (______9__34084));
  nor2s1 ______448128(.DIN1 (________21788), .DIN2 (________21274), .Q
       (________22212));
  hi1s1 ___99__448129(.DIN (___0____21679), .Q (____00__24701));
  nor2s1 _______448130(.DIN1 (____9___21898), .DIN2 (______0__35068),
       .Q (_____0__22216));
  nnd2s1 _______448131(.DIN1 (_____0__21240), .DIN2 (________20872), .Q
       (____9___21899));
  hi1s1 _____9_448132(.DIN (___0____21678), .Q (___90___24242));
  hi1s1 _______448133(.DIN (______0__30591), .Q (_________31164));
  hi1s1 ___0___448134(.DIN (________22392), .Q (____0___22814));
  and2s1 _______448135(.DIN1 (________21305), .DIN2 (___0____21677), .Q
       (________22221));
  hi1s1 _______448136(.DIN (_____0__22108), .Q (_____0__22242));
  and2s1 ___0___448137(.DIN1 (________21320), .DIN2 (___0____21698), .Q
       (___0____22592));
  nor2s1 ___0___448138(.DIN1 (________21148), .DIN2 (___0_0__21676), .Q
       (________25058));
  and2s1 ___0_9_448139(.DIN1 (____0___24705), .DIN2 (________23295), .Q
       (________22276));
  nnd2s1 ______448140(.DIN1 (___0____21644), .DIN2 (___0_0__21658), .Q
       (_____0__22148));
  nnd2s1 ___0___448141(.DIN1 (____0___25661), .DIN2 (___0_9__21675), .Q
       (________23853));
  nnd2s1 ___0___448142(.DIN1 (________25604), .DIN2 (___0____21674), .Q
       (________25483));
  nnd2s1 ___0___448143(.DIN1 (___0____21673), .DIN2 (___9_9__21589), .Q
       (________22316));
  or2s1 ___0___448144(.DIN1 (____9___19945), .DIN2 (___0____21672), .Q
       (________23109));
  xnr2s1 ___0___448145(.DIN1 (________19160), .DIN2 (____9____32728),
       .Q (_____0__23958));
  nnd2s1 _______448146(.DIN1 (________21324), .DIN2 (________22332), .Q
       (__9__0__26664));
  hi1s1 ___0___448147(.DIN (____9___21901), .Q (____00__22356));
  nor2s1 _______448148(.DIN1 (___0____21671), .DIN2 (________21108), .Q
       (____9___26144));
  nnd2s1 ___0___448149(.DIN1 (________21321), .DIN2 (________19257), .Q
       (_____0__26077));
  or2s1 _______448150(.DIN1 (________24855), .DIN2 (___0____21670), .Q
       (___9____25249));
  hi1s1 ___0_9_448151(.DIN (___0____21669), .Q (___00____27196));
  and2s1 _______448152(.DIN1 (________21395), .DIN2 (_____9__22147), .Q
       (___9____24314));
  or2s1 ___0__448153(.DIN1 (___0____21668), .DIN2 (___99___23435), .Q
       (___9_0__23413));
  and2s1 _______448154(.DIN1 (________25052), .DIN2 (________21322), .Q
       (____9___25742));
  hi1s1 _______448155(.DIN (___0_0__21667), .Q (__90____26258));
  nnd2s1 _____0_448156(.DIN1 (___0____21665), .DIN2 (_____0__21821), .Q
       (________24557));
  nor2s1 ______448157(.DIN1 (________21213), .DIN2 (________21095), .Q
       (________22410));
  nnd2s1 ______448158(.DIN1 (________21292), .DIN2 (___0____21663), .Q
       (________24824));
  nnd2s1 _____0_448159(.DIN1 (___0____21687), .DIN2 (_____0__21821), .Q
       (________22369));
  hi1s1 _______448160(.DIN (_____0__22366), .Q (__9_____26548));
  hi1s1 ___0_448161(.DIN (___0_9__21666), .Q (__9_____26583));
  nor2s1 _______448162(.DIN1 (____0___21357), .DIN2 (_____0__21327), .Q
       (___00___24334));
  nnd2s1 _______448163(.DIN1 (___0____21665), .DIN2 (___0____21664), .Q
       (_____9__25674));
  nnd2s1 _______448164(.DIN1 (________21311), .DIN2 (___0____21663), .Q
       (________25836));
  hi1s1 ___0___448165(.DIN (___0____21662), .Q (__9_____27037));
  nor2s1 ____09_448166(.DIN1 (________21506), .DIN2 (___0____21655), .Q
       (________25437));
  hi1s1 ___0__448167(.DIN (________22678), .Q (________23919));
  nor2s1 _____9_448168(.DIN1 (_____0__20198), .DIN2 (________21741), .Q
       (____0___22359));
  hi1s1 ___00__448169(.DIN (_________33103), .Q (_________31618));
  nor2s1 _______448170(.DIN1 (________20062), .DIN2 (___0____21661), .Q
       (________25513));
  nor2s1 ___0_9_448171(.DIN1 (___0____21660), .DIN2 (________21318), .Q
       (___9_9__23395));
  hi1s1 _______448172(.DIN (____9___22078), .Q (________24440));
  nor2s1 _____0_448173(.DIN1 (________21145), .DIN2 (___0____21661), .Q
       (__9_____26381));
  nor2s1 ___0_0_448174(.DIN1 (___0____21660), .DIN2 (________21282), .Q
       (________23101));
  nor2s1 ___0__448175(.DIN1 (___0____21659), .DIN2 (_____0__21729), .Q
       (____9___23255));
  nnd2s1 ______448176(.DIN1 (____0___21171), .DIN2 (___0_0__21658), .Q
       (________23140));
  nnd2s1 ____0_448177(.DIN1 (________21866), .DIN2 (___0_9__21657), .Q
       (________22246));
  and2s1 ___0___448178(.DIN1 (________21795), .DIN2 (________21481), .Q
       (_____9__24828));
  nnd2s1 _______448179(.DIN1 (_____9__21119), .DIN2 (________21794), .Q
       (__9_____26623));
  nnd2s1 ___0_9_448180(.DIN1 (_____0__21288), .DIN2 (___9____20669), .Q
       (________26032));
  nor2s1 _______448181(.DIN1 (___0____21651), .DIN2 (___0____21655), .Q
       (___99___23432));
  nnd2s1 ___0__448182(.DIN1 (________21795), .DIN2 (________20970), .Q
       (___00____27182));
  nor2s1 _______448183(.DIN1 (____0____29098), .DIN2 (________21303),
       .Q (____9____32697));
  hi1s1 ______448184(.DIN (___0____21654), .Q (___0_____27696));
  nnd2s1 ___09__448185(.DIN1 (________20956), .DIN2 (________20574), .Q
       (___0____21653));
  or2s1 ______448186(.DIN1 (___0____21651), .DIN2 (____0___20795), .Q
       (___0____21652));
  nnd2s1 ___0___448187(.DIN1 (___9____21566), .DIN2 (___0____20756), .Q
       (___0____21650));
  nor2s1 ______448188(.DIN1 (________21115), .DIN2 (________21733), .Q
       (___0_0__21649));
  nnd2s1 _______448189(.DIN1 (_________31648), .DIN2 (____9__18955), .Q
       (___0_9__21648));
  nor2s1 _______448190(.DIN1 (________19613), .DIN2 (________20915), .Q
       (___0____21647));
  nor2s1 _______448191(.DIN1 (_____9__20030), .DIN2 (________21004), .Q
       (___0____21646));
  nor2s1 _______448192(.DIN1 (________21319), .DIN2 (_____0__20991), .Q
       (___0____21645));
  nnd2s1 _______448193(.DIN1 (________21150), .DIN2 (________21497), .Q
       (___0____21643));
  nnd2s1 ______448194(.DIN1 (___9____20674), .DIN2 (________20249), .Q
       (___0____21642));
  nnd2s1 _______448195(.DIN1 (____99__21354), .DIN2 (____0___20791), .Q
       (___0_0__21641));
  nnd2s1 _______448196(.DIN1 (________19873), .DIN2 (________21011), .Q
       (___00___21640));
  nor2s1 ___0___448197(.DIN1 (_____9__21493), .DIN2 (________21176), .Q
       (___00___21639));
  nnd2s1 ___09__448198(.DIN1 (___0____20721), .DIN2 (____9___20596), .Q
       (___00___21638));
  nnd2s1 ___09_448199(.DIN1 (________21027), .DIN2 (___09___19848), .Q
       (___00___21637));
  or2s1 _______448200(.DIN1 (________21730), .DIN2 (________21512), .Q
       (___00___21636));
  nor2s1 _______448201(.DIN1 (________21730), .DIN2 (________21371), .Q
       (___00___21635));
  nnd2s1 ___0_9_448202(.DIN1 (____99__20981), .DIN2 (____0___21816), .Q
       (___00___21634));
  or2s1 ___0___448203(.DIN1 (___999__21632), .DIN2 (________20862), .Q
       (___000__21633));
  nnd2s1 _______448204(.DIN1 (_____9__21400), .DIN2 (________21470), .Q
       (___99___21631));
  or2s1 _______448205(.DIN1 (________20470), .DIN2 (___9____21620), .Q
       (___99___21630));
  hi1s1 ____0__448206(.DIN (___99___21628), .Q (___99___21629));
  and2s1 ___0___448207(.DIN1 (________20929), .DIN2 (________19962), .Q
       (___99___21627));
  hi1s1 ____0__448208(.DIN (___0____21697), .Q (___99___21626));
  nor2s1 ___0_9_448209(.DIN1 (_____0___34426), .DIN2 (________21949),
       .Q (___990));
  or2s1 _____0_448210(.DIN1 (___9____21624), .DIN2 (_____9__20971), .Q
       (___9_9__21625));
  nor2s1 ___00__448211(.DIN1 (___9____24300), .DIN2 (_________30341),
       .Q (___9____21623));
  nnd2s1 _______448212(.DIN1 (___9____21614), .DIN2 (___00___20703), .Q
       (___9____21622));
  or2s1 _____0_448213(.DIN1 (________20998), .DIN2 (___9____21620), .Q
       (___9____21621));
  nor2s1 _____9_448214(.DIN1 (___9____21618), .DIN2 (________20953), .Q
       (___9____21619));
  nnd2s1 _______448215(.DIN1 (________21477), .DIN2 (________20809), .Q
       (___9_0__21617));
  nor2s1 _____9_448216(.DIN1 (________20930), .DIN2 (________21389), .Q
       (___9_9__21616));
  nor2s1 ______448217(.DIN1 (_____9__20856), .DIN2 (___9____21614), .Q
       (___9____21615));
  nor2s1 _______448218(.DIN1 (________19664), .DIN2 (___009__20707), .Q
       (___9____21613));
  nnd2s1 ___0___448219(.DIN1 (________20966), .DIN2 (________21974), .Q
       (___9____21612));
  nor2s1 ___0__448220(.DIN1 (___9____21610), .DIN2 (_____9__20875), .Q
       (___9____21611));
  xor2s1 ___0_0_448221(.DIN1 (_________31479), .DIN2 (_________30104),
       .Q (___9____21609));
  xor2s1 ___0___448222(.DIN1 (_________34447), .DIN2 (____0____30981),
       .Q (___9_0__21608));
  xor2s1 ___0___448223(.DIN1 (_____________18898), .DIN2
       (_________31479), .Q (___9_9__21607));
  nnd2s1 _______448224(.DIN1 (_____0__21485), .DIN2 (________20934), .Q
       (___9____21606));
  nor2s1 _______448225(.DIN1 (________21086), .DIN2 (________20968), .Q
       (___9____21605));
  nnd2s1 _______448226(.DIN1 (____9___20974), .DIN2 (_____0__19525), .Q
       (___9____21604));
  nor2s1 ______448227(.DIN1 (____0___20427), .DIN2 (_____9__20961), .Q
       (___9____21603));
  and2s1 _______448228(.DIN1 (________21456), .DIN2 (___0_0__21658), .Q
       (___9____21602));
  nnd2s1 _______448229(.DIN1 (___9____20690), .DIN2 (________21489), .Q
       (___9____21601));
  hi1s1 ___0___448230(.DIN (_____9__21800), .Q (___9____21600));
  nnd2s1 _______448231(.DIN1 (___9____20642), .DIN2 (________21367), .Q
       (___9_0__21599));
  nnd2s1 ___0_9_448232(.DIN1 (____0___20792), .DIN2 (________19575), .Q
       (___9_9__21598));
  nnd2s1 ___0_9_448233(.DIN1 (________20808), .DIN2 (___0_0__21658), .Q
       (___9____21597));
  nor2s1 ___0_9_448234(.DIN1 (_____9__21038), .DIN2 (________20948), .Q
       (___9____21596));
  nnd2s1 ___0_448235(.DIN1 (________21491), .DIN2 (_____0__21335), .Q
       (___9____21594));
  nor2s1 ___0_0_448236(.DIN1 (___9____21592), .DIN2 (________21022), .Q
       (___9____21593));
  nnd2s1 ___0_0_448237(.DIN1 (___9_0__21580), .DIN2 (inData[30]), .Q
       (___9____21591));
  nnd2s1 ___0_0_448238(.DIN1 (________21057), .DIN2 (___9_9__21589), .Q
       (___9_0__21590));
  nnd2s1 ___0_0_448239(.DIN1 (________21035), .DIN2 (___90___21549), .Q
       (___9____21588));
  nnd2s1 ___0__448240(.DIN1 (_________35082), .DIN2 (________19962), .Q
       (___9____21587));
  nnd2s1 ___0___448241(.DIN1 (___000__20699), .DIN2 (____0___20327), .Q
       (___9____21586));
  nor2s1 ___0___448242(.DIN1 (____0________________18591), .DIN2
       (________20864), .Q (___9____21585));
  nnd2s1 ___0__448243(.DIN1 (____00__20324), .DIN2 (___9____21583), .Q
       (___9____21584));
  nor2s1 ___0___448244(.DIN1 (_________29585), .DIN2 (____0____30080),
       .Q (___9____21582));
  nnd2s1 ___0___448245(.DIN1 (___9_0__21580), .DIN2 (inData[28]), .Q
       (___9____21581));
  nor2s1 ___0___448246(.DIN1 (________19912), .DIN2 (________20818), .Q
       (___9_9__21579));
  nor2s1 ___0___448247(.DIN1 (______9__28578), .DIN2 (____0____30080),
       .Q (___9____21578));
  nnd2s1 ___0___448248(.DIN1 (_____9__20865), .DIN2 (____0___20045), .Q
       (___9____21577));
  nor2s1 ___0__448249(.DIN1 (___9____21575), .DIN2 (___999__20698), .Q
       (___9____21576));
  nnd2s1 ___0__448250(.DIN1 (________20999), .DIN2 (___9_9__21589), .Q
       (___9____21574));
  nor2s1 ___0___448251(.DIN1 (____0___21991), .DIN2 (________21028), .Q
       (___9____21573));
  nor2s1 ___0___448252(.DIN1 (____0___20330), .DIN2 (___0_0__20724), .Q
       (___9____21572));
  nnd2s1 ___0___448253(.DIN1 (___0____20764), .DIN2
       (__________________0___18628), .Q (___9_0__21571));
  nor2s1 ___0___448254(.DIN1 (________21425), .DIN2 (________21300), .Q
       (___9_9__21570));
  nor2s1 ___0__448255(.DIN1 (___9____21568), .DIN2 (________21507), .Q
       (___9____21569));
  nnd2s1 ___0___448256(.DIN1 (___9____21566), .DIN2 (___0____20748), .Q
       (___9____21567));
  nnd2s1 ___0__448257(.DIN1 (________21017), .DIN2 (____0___20042), .Q
       (___9____21565));
  nnd2s1 ___0___448258(.DIN1 (________20863), .DIN2 (________20099), .Q
       (___9____21564));
  nnd2s1 ___0___448259(.DIN1 (___9_0__21580), .DIN2 (inData[31]), .Q
       (___9____21563));
  nnd2s1 ___0___448260(.DIN1 (_____9__20806), .DIN2 (___9_0__21561), .Q
       (___9____21562));
  nor2s1 ___0___448261(.DIN1 (___0____20726), .DIN2 (________20437), .Q
       (___9_9__21560));
  nor2s1 ___0___448262(.DIN1 (________20084), .DIN2 (_____9__21474), .Q
       (___9____21559));
  nor2s1 ___0__448263(.DIN1 (___0____20753), .DIN2 (________20810), .Q
       (___9____21558));
  or2s1 ___0___448264(.DIN1 (___9____21556), .DIN2 (_________28837), .Q
       (___9____21557));
  nor2s1 ___0_448265(.DIN1 (____0___21080), .DIN2 (___0____20729), .Q
       (___9____21555));
  nor2s1 ___0_9_448266(.DIN1 (_____9__19668), .DIN2 (________21026), .Q
       (___9____21554));
  nor2s1 ___0_9_448267(.DIN1 (____0___20234), .DIN2 (____9___20979), .Q
       (___9_0__21553));
  nnd2s1 ___0_9_448268(.DIN1 (________20928), .DIN2 (____0___21988), .Q
       (___909__21552));
  nnd2s1 ___0_448269(.DIN1 (___0____20728), .DIN2 (________22037), .Q
       (___90___21551));
  nnd2s1 ___090_448270(.DIN1 (________21519), .DIN2 (___90___21549), .Q
       (___90___21550));
  nnd2s1 ___090_448271(.DIN1 (________20963), .DIN2 (inData[26]), .Q
       (___90___21548));
  nor2s1 ___090_448272(.DIN1 (___90___21546), .DIN2 (________21033), .Q
       (___90___21547));
  nor2s1 ___09__448273(.DIN1 (___90___21544), .DIN2 (____9___21535), .Q
       (___90___21545));
  nor2s1 ___09__448274(.DIN1 (________21174), .DIN2 (____99__21542), .Q
       (___900__21543));
  and2s1 ___09__448275(.DIN1 (_________31648), .DIN2 (________20122),
       .Q (____9___21541));
  nor2s1 _______448276(.DIN1 (___9____20683), .DIN2 (________20451), .Q
       (____9___21540));
  nnd2s1 ___09__448277(.DIN1 (________20967), .DIN2 (________19675), .Q
       (____9___21539));
  nor2s1 ___09__448278(.DIN1 (________20854), .DIN2 (____9___21537), .Q
       (____9___21538));
  nor2s1 ___09__448279(.DIN1 (________21021), .DIN2 (____9___21535), .Q
       (____9___21536));
  nnd2s1 ___09__448280(.DIN1 (___0____20760), .DIN2 (____90__21533), .Q
       (____9___21534));
  or2s1 ___09__448281(.DIN1 (________19459), .DIN2 (________20939), .Q
       (_____9__21532));
  nnd2s1 ___09__448282(.DIN1 (________21525), .DIN2 (________21530), .Q
       (________21531));
  nnd2s1 ___09__448283(.DIN1 (________20536), .DIN2 (___9____20670), .Q
       (________21529));
  and2s1 ___09__448284(.DIN1 (________21005), .DIN2 (_____0__19862), .Q
       (________21528));
  and2s1 ___09__448285(.DIN1 (_________31648), .DIN2 (______18941), .Q
       (________21527));
  nnd2s1 ___09_448286(.DIN1 (________21525), .DIN2 (________21518), .Q
       (________21526));
  nnd2s1 ___09_448287(.DIN1 (________21525), .DIN2 (___0_0__20771), .Q
       (________21524));
  nor2s1 ___09__448288(.DIN1 (_____9__21522), .DIN2 (___9____21620), .Q
       (_____0__21523));
  nnd2s1 ___09__448289(.DIN1 (________20908), .DIN2 (inData[28]), .Q
       (________21521));
  nnd2s1 _______448290(.DIN1 (________21519), .DIN2 (________21518), .Q
       (________21520));
  nnd2s1 _______448291(.DIN1 (___0_0__20708), .DIN2 (____0___21988), .Q
       (________21517));
  nor2s1 _______448292(.DIN1 (___0_9__20751), .DIN2 (________21372), .Q
       (________21516));
  or2s1 _______448293(.DIN1 (________21032), .DIN2 (____9___21537), .Q
       (________21515));
  nor2s1 _______448294(.DIN1 (_____0__20942), .DIN2 (____9___20601), .Q
       (_____0__21514));
  hi1s1 ______448295(.DIN (________22425), .Q (________21999));
  nnd2s1 ____00_448296(.DIN1 (___0____20709), .DIN2 (_____0__20274), .Q
       (________21836));
  nnd2s1 ____00_448297(.DIN1 (________21100), .DIN2 (_____9__21513), .Q
       (___0____21709));
  nor2s1 ____0__448298(.DIN1 (___0____21659), .DIN2 (________21512), .Q
       (________21838));
  nor2s1 ____0__448299(.DIN1 (______18933), .DIN2 (___9____20687), .Q
       (_____0__21840));
  nnd2s1 ____0__448300(.DIN1 (_____0__20807), .DIN2 (___09___20787), .Q
       (________22302));
  and2s1 ____00_448301(.DIN1 (________20921), .DIN2 (________21511), .Q
       (____0___21987));
  hi1s1 _______448302(.DIN (____0___21992), .Q (____0___21993));
  hi1s1 ____0__448303(.DIN (________23236), .Q (____0___22357));
  nor2s1 ___0___448304(.DIN1 (________21206), .DIN2 (___9_0__20672), .Q
       (___0____21656));
  nnd2s1 ___0___448305(.DIN1 (________21490), .DIN2 (________21510), .Q
       (___0____21708));
  nnd2s1 ___0__448306(.DIN1 (_____9__21484), .DIN2 (________21510), .Q
       (___0____21688));
  nnd2s1 ___0___448307(.DIN1 (________20815), .DIN2 (________21509), .Q
       (___0____21662));
  nnd2s1 ___0_9_448308(.DIN1 (____90__20876), .DIN2 (________21785), .Q
       (___0_9__21666));
  nor2s1 ___0_9_448309(.DIN1 (________21508), .DIN2 (____99__20885), .Q
       (___0____21669));
  nor2s1 ___0___448310(.DIN1 (________21976), .DIN2 (_____0__20933), .Q
       (___0____21679));
  nor2s1 ___09_448311(.DIN1 (____0____________0_), .DIN2
       (________20867), .Q (________21967));
  nnd2s1 ___09__448312(.DIN1 (____0___20985), .DIN2 (________21776), .Q
       (____00__21985));
  nnd2s1 ___099_448313(.DIN1 (___0____22589), .DIN2 (________19570), .Q
       (________24000));
  nor2s1 ___099_448314(.DIN1 (________21488), .DIN2 (________20918), .Q
       (____0___21989));
  nor2s1 ___448315(.DIN1 (___9____19725), .DIN2 (________21013), .Q
       (___09___21712));
  nor2s1 ____00_448316(.DIN1 (___9_9__20662), .DIN2 (________21500), .Q
       (____9___21981));
  nor2s1 ____00_448317(.DIN1 (________19269), .DIN2 (________21507), .Q
       (____0___21906));
  nor2s1 _______448318(.DIN1 (___9____21592), .DIN2 (________21482), .Q
       (_____0__21783));
  nnd2s1 ____09_448319(.DIN1 (________21015), .DIN2 (________20394), .Q
       (________21779));
  nor2s1 _____0_448320(.DIN1 (________21506), .DIN2 (____09__21364), .Q
       (________22392));
  nor2s1 _______448321(.DIN1 (________21505), .DIN2 (___0____20741), .Q
       (________22122));
  nnd2s1 ____0_448322(.DIN1 (________20927), .DIN2 (________21976), .Q
       (________21977));
  nnd2s1 ____0__448323(.DIN1 (________20902), .DIN2 (___0__18931), .Q
       (________22035));
  nnd2s1 ____0__448324(.DIN1 (________21340), .DIN2 (_____0__21504), .Q
       (___0_____27289));
  nor2s1 ____0__448325(.DIN1 (____0___21363), .DIN2 (_____0__20904), .Q
       (_____0__22670));
  hi1s1 _______448326(.DIN (___0_0__22608), .Q (_____0__23591));
  or2s1 ____0__448327(.DIN1 (________21492), .DIN2 (________21478), .Q
       (________21998));
  nor2s1 ____0__448328(.DIN1 (________21483), .DIN2 (_____9__21503), .Q
       (___0____24389));
  nor2s1 ____448329(.DIN1 (________19613), .DIN2 (________21037), .Q
       (________22152));
  or2s1 ____0__448330(.DIN1 (________19631), .DIN2 (___9_0__21580), .Q
       (________22048));
  nor2s1 ___0_0_448331(.DIN1 (________21487), .DIN2 (________21473), .Q
       (___9_0__22491));
  and2s1 ____0__448332(.DIN1 (__9_____26370), .DIN2 (________21377), .Q
       (________24571));
  nor2s1 ____0__448333(.DIN1 (___9____21592), .DIN2 (_____9__21503), .Q
       (_____9__22743));
  nor2s1 _______448334(.DIN1 (________21502), .DIN2 (___0_0__20762), .Q
       (____0___22358));
  nnd2s1 ___0__448335(.DIN1 (________21124), .DIN2 (____90__21801), .Q
       (________22766));
  nnd2s1 ____0__448336(.DIN1 (________20824), .DIN2 (___0__18931), .Q
       (_____9__21970));
  nor2s1 ____0__448337(.DIN1 (________21060), .DIN2 (_____9__20951), .Q
       (________24749));
  nor2s1 ____0__448338(.DIN1 (________21502), .DIN2 (_____0__21494), .Q
       (____9___22348));
  nor2s1 ____0__448339(.DIN1 (________21479), .DIN2 (________21376), .Q
       (_____0__26117));
  nor2s1 ____0__448340(.DIN1 (________21501), .DIN2 (________21500), .Q
       (___0____22603));
  nnd2s1 _______448341(.DIN1 (________21498), .DIN2 (________21499), .Q
       (________22678));
  nnd2s1 ____0__448342(.DIN1 (________20994), .DIN2 (________19884), .Q
       (____09__24992));
  nnd2s1 ____0__448343(.DIN1 (________21498), .DIN2 (________21497), .Q
       (________23005));
  hi1s1 _____0_448344(.DIN (________21496), .Q (_____9__23161));
  or2s1 ____0__448345(.DIN1 (________21495), .DIN2 (_____0__21494), .Q
       (___9____26235));
  nor2s1 ____0_448346(.DIN1 (_____9__21493), .DIN2 (________20832), .Q
       (___9_0__26207));
  nor2s1 ____0__448347(.DIN1 (____0___20889), .DIN2 (________20801), .Q
       (________22112));
  nor2s1 ____0_448348(.DIN1 (________20277), .DIN2 (___0____20739), .Q
       (___0____22559));
  or2s1 ____0_448349(.DIN1 (________21492), .DIN2 (____9___21350), .Q
       (________22026));
  hi1s1 ___0___448350(.DIN (_________29496), .Q (_________33541));
  nor2s1 ____0__448351(.DIN1 (___9____20665), .DIN2 (________21235), .Q
       (________23136));
  nor2s1 ____0__448352(.DIN1 (___0____21659), .DIN2 (___0____20720), .Q
       (___9____22458));
  nnd2s1 ____0__448353(.DIN1 (________21491), .DIN2 (____00__20510), .Q
       (____09__22815));
  nor2s1 ____0__448354(.DIN1 (____9___21351), .DIN2 (_____0__21494), .Q
       (________24105));
  nor2s1 ______448355(.DIN1 (___9____20641), .DIN2 (________20931), .Q
       (__9_____26350));
  nor2s1 ___0__448356(.DIN1 (________21889), .DIN2 (_________35080), .Q
       (____9___25943));
  nor2s1 ___0___448357(.DIN1 (___9____19725), .DIN2 (________20907), .Q
       (_________28636));
  nnd2s1 ___0___448358(.DIN1 (________21490), .DIN2 (________21489), .Q
       (___9____23397));
  nor2s1 ___0___448359(.DIN1 (___9____19725), .DIN2 (___9____20686), .Q
       (____0___25853));
  nor2s1 ____0_448360(.DIN1 (________21488), .DIN2 (________20938), .Q
       (___9____25206));
  nor2s1 ____0_448361(.DIN1 (________21487), .DIN2 (________21338), .Q
       (________22123));
  nnd2s1 ____09_448362(.DIN1 (________21231), .DIN2 (___9_9__21589), .Q
       (___9____23394));
  nnd2s1 _____0_448363(.DIN1 (________20820), .DIN2 (________21486), .Q
       (____9___25170));
  nor2s1 ______448364(.DIN1 (________21495), .DIN2 (________21118), .Q
       (___0____24378));
  nnd2s1 ____0__448365(.DIN1 (________21382), .DIN2 (________21976), .Q
       (________22002));
  nnd2s1 ____0__448366(.DIN1 (_____0__21120), .DIN2 (_____0__21485), .Q
       (_____0__22014));
  nnd2s1 ___0___448367(.DIN1 (_____9__21484), .DIN2 (________21489), .Q
       (___99___22533));
  nor2s1 ____0__448368(.DIN1 (________21483), .DIN2 (________21482), .Q
       (___9____24260));
  nnd2s1 _____0_448369(.DIN1 (________21007), .DIN2 (________21481), .Q
       (________23145));
  nnd2s1 _______448370(.DIN1 (___09___20786), .DIN2 (________21480), .Q
       (________22289));
  nor2s1 ____0__448371(.DIN1 (________21479), .DIN2 (________21478), .Q
       (____0___26053));
  nor2s1 ______448372(.DIN1 (____09__20990), .DIN2 (_____9__21326), .Q
       (__9_0___26897));
  nnd2s1 ___0___448373(.DIN1 (________21332), .DIN2 (___0____21663), .Q
       (___00____27220));
  nor2s1 ___0_9_448374(.DIN1 (________21887), .DIN2 (_____0__20817), .Q
       (___0_0___27370));
  nnd2s1 _______448375(.DIN1 (_____9__20922), .DIN2 (________21468), .Q
       (______9__33828));
  nnd2s1 _______448376(.DIN1 (________21008), .DIN2 (________21477), .Q
       (__9_0___26517));
  nor2s1 _______448377(.DIN1 (________21476), .DIN2 (________20869), .Q
       (__90_9__26308));
  nor2s1 ____09_448378(.DIN1 (_____0__21475), .DIN2 (_____0__21030), .Q
       (___0_____27804));
  nor2s1 _______448379(.DIN1 (________21508), .DIN2 (_____9__21474), .Q
       (___0_____27291));
  nor2s1 ___0___448380(.DIN1 (________21472), .DIN2 (________21473), .Q
       (__9_____26784));
  or2s1 _______448381(.DIN1 (________21472), .DIN2 (________20870), .Q
       (__9_____26828));
  or2s1 _______448382(.DIN1 (________21471), .DIN2 (_____9__21503), .Q
       (___9_0__26177));
  nor2s1 _______448383(.DIN1 (________21508), .DIN2 (___9____20689), .Q
       (________25913));
  nnd2s1 _______448384(.DIN1 (_____0__20799), .DIN2 (________20825), .Q
       (_________31486));
  nor2s1 ___0___448385(.DIN1 (________21470), .DIN2 (___0____20712), .Q
       (_________31956));
  nnd2s1 _______448386(.DIN1 (____9___20973), .DIN2 (________21468), .Q
       (____0____32823));
  nor2s1 ______448387(.DIN1 (___0____19828), .DIN2 (________20945), .Q
       (_____9___30624));
  nnd2s1 ___0_0_448388(.DIN1 (________21463), .DIN2 (________21510), .Q
       (________21467));
  nor2s1 _______448389(.DIN1 (_____9__21019), .DIN2 (________21512), .Q
       (________21466));
  nnd2s1 _______448390(.DIN1 (________20955), .DIN2 (____9___21808), .Q
       (_____0__21465));
  nnd2s1 ______448391(.DIN1 (________21463), .DIN2 (________21518), .Q
       (_____9__21464));
  nnd2s1 ______448392(.DIN1 (___9_0__20682), .DIN2 (________21461), .Q
       (________21462));
  and2s1 _______448393(.DIN1 (________20919), .DIN2 (___0____21677), .Q
       (________21460));
  nnd2s1 _______448394(.DIN1 (___09___20781), .DIN2 (________21458), .Q
       (________21459));
  nnd2s1 _____448395(.DIN1 (________21456), .DIN2 (________20593), .Q
       (________21457));
  nnd2s1 _______448396(.DIN1 (___0____20711), .DIN2 (_____9__20932), .Q
       (_____0__21455));
  nnd2s1 ___00__448397(.DIN1 (____0___21447), .DIN2 (____0___21453), .Q
       (____09__21454));
  nor2s1 _______448398(.DIN1 (_____0__20304), .DIN2 (________21406), .Q
       (____0___21452));
  xor2s1 ___0_9_448399(.DIN1 (_________18847), .DIN2 (_________34362),
       .Q (____0___21451));
  xor2s1 ___0_448400(.DIN1 (____0___21449), .DIN2 (____009__31815), .Q
       (____0___21450));
  nnd2s1 ___0___448401(.DIN1 (____0___21447), .DIN2 (____0___19600), .Q
       (____0___21448));
  nnd2s1 _______448402(.DIN1 (___090__20780), .DIN2 (________21387), .Q
       (____00__21446));
  xor2s1 ___0___448403(.DIN1 (_________34489), .DIN2 (_________34077),
       .Q (____99__21445));
  nnd2s1 ___09__448404(.DIN1 (________20995), .DIN2 (________19957), .Q
       (____9___21444));
  nnd2s1 ___448405(.DIN1 (____0___20986), .DIN2 (________21098), .Q
       (____9___21443));
  nnd2s1 ___0___448406(.DIN1 (____0___21356), .DIN2 (____9___21441), .Q
       (____9___21442));
  hi1s1 ___0___448407(.DIN (____9___21439), .Q (____9___21440));
  and2s1 ___0___448408(.DIN1 (___0____22589), .DIN2 (________23757), .Q
       (____90__21438));
  nnd2s1 ___0___448409(.DIN1 (____0___20890), .DIN2 (________21776), .Q
       (_____9__21437));
  nor2s1 ___090_448410(.DIN1 (________21978), .DIN2 (____9___21535), .Q
       (________21436));
  nnd2s1 ___0___448411(.DIN1 (________21031), .DIN2 (_____9__20283), .Q
       (________21434));
  hi1s1 ___0___448412(.DIN (___009__23445), .Q (________21433));
  and2s1 ___09__448413(.DIN1 (____9___20980), .DIN2 (________21458), .Q
       (________21432));
  nnd2s1 ___090_448414(.DIN1 (___0____20747), .DIN2 (________21368), .Q
       (________21431));
  nor2s1 ___0___448415(.DIN1 (_____0__21429), .DIN2 (________21507), .Q
       (________21430));
  nnd2s1 ___09__448416(.DIN1 (________20898), .DIN2 (____0___21988), .Q
       (_____9__21428));
  and2s1 ___0___448417(.DIN1 (____0____30080), .DIN2 (______18938), .Q
       (________21427));
  nor2s1 ___09__448418(.DIN1 (________21425), .DIN2 (________21424), .Q
       (________21426));
  nnd2s1 ___0___448419(.DIN1 (___9____21566), .DIN2 (________21477), .Q
       (________21423));
  nnd2s1 ___09_448420(.DIN1 (________20434), .DIN2 (____00__20982), .Q
       (________21422));
  hi1s1 _______448421(.DIN (________21420), .Q (________21421));
  nnd2s1 ___09__448422(.DIN1 (___00___20706), .DIN2 (_____0__20439), .Q
       (_____0__21419));
  hi1s1 ______448423(.DIN (________21417), .Q (________21418));
  hi1s1 _______448424(.DIN (________21415), .Q (________21416));
  and2s1 _____448425(.DIN1 (_____9__21029), .DIN2 (________21458), .Q
       (________21414));
  hi1s1 _______448426(.DIN (__9_____26555), .Q (________21413));
  hi1s1 ____0__448427(.DIN (________21411), .Q (________21412));
  nnd2s1 _______448428(.DIN1 (________20997), .DIN2 (________19981), .Q
       (_____0__21410));
  or2s1 _______448429(.DIN1 (________21407), .DIN2 (________21406), .Q
       (________21408));
  nor2s1 _____9_448430(.DIN1 (________21061), .DIN2 (________25782), .Q
       (________21405));
  or2s1 _______448431(.DIN1 (____0___21724), .DIN2 (____00__20790), .Q
       (________21404));
  nor2s1 ______448432(.DIN1 (____9___20218), .DIN2 (________21402), .Q
       (________21403));
  nnd2s1 ______448433(.DIN1 (_____9__21400), .DIN2 (________20946), .Q
       (_____0__21401));
  xor2s1 _______448434(.DIN1 (_________18861), .DIN2 (_________31578),
       .Q (________21399));
  and2s1 _______448435(.DIN1 (___9____21614), .DIN2 (________21397), .Q
       (________21398));
  hi1s1 ____0__448436(.DIN (________21395), .Q (________21396));
  nnd2s1 _______448437(.DIN1 (________21733), .DIN2 (________20405), .Q
       (________21394));
  nor2s1 _______448438(.DIN1 (_________18862), .DIN2 (___0____20740),
       .Q (_____0__21393));
  hi1s1 _______448439(.DIN (________21041), .Q (_____9__21392));
  hi1s1 _______448440(.DIN (________21390), .Q (________21391));
  nor2s1 _____9_448441(.DIN1 (________21310), .DIN2 (________21389), .Q
       (________21767));
  nor2s1 ______448442(.DIN1 (________21506), .DIN2 (________20947), .Q
       (___0____21683));
  nnd2s1 _____9_448443(.DIN1 (________20812), .DIN2 (________20802), .Q
       (________21765));
  nor2s1 _____448444(.DIN1 (________20935), .DIN2 (________21388), .Q
       (________21918));
  or2s1 _____448445(.DIN1 (________21750), .DIN2 (________20992), .Q
       (____0___21909));
  and2s1 _____0_448446(.DIN1 (___0____20755), .DIN2 (___0____21663), .Q
       (____0___21907));
  nnd2s1 _______448447(.DIN1 (________20969), .DIN2 (______18933), .Q
       (________21915));
  nor2s1 _______448448(.DIN1 (________19613), .DIN2 (_____9__21383), .Q
       (________23103));
  nnd2s1 _______448449(.DIN1 (_____0__21384), .DIN2 (________21387), .Q
       (________21950));
  nnd2s1 ___0___448450(.DIN1 (____9___21349), .DIN2 (________21480), .Q
       (____00__21719));
  hi1s1 _______448451(.DIN (________21386), .Q (___0_____27778));
  nnd2s1 _______448452(.DIN1 (________21343), .DIN2 (________21385), .Q
       (________21786));
  nnd2s1 _____448453(.DIN1 (_____0__21384), .DIN2 (___0_0__21658), .Q
       (___0_0__21667));
  nnd2s1 _______448454(.DIN1 (___0____20766), .DIN2 (____0___21905), .Q
       (___0_9__21685));
  nnd2s1 ___0___448455(.DIN1 (________20905), .DIN2 (____90__21801), .Q
       (___90___22448));
  nor2s1 _______448456(.DIN1 (___0____21659), .DIN2 (_____9__21383), .Q
       (___90___22453));
  nor2s1 _____9_448457(.DIN1 (________21730), .DIN2 (_____9__21383), .Q
       (_____9__22933));
  hi1s1 ___0___448458(.DIN (___0____24393), .Q (________24908));
  nnd2s1 _______448459(.DIN1 (________21382), .DIN2 (________21381), .Q
       (________21975));
  hi1s1 ___0__448460(.DIN (___09___23526), .Q (__9_0___26521));
  hi1s1 ___0___448461(.DIN (________21380), .Q (____0___21986));
  nor2s1 ___09__448462(.DIN1 (________19989), .DIN2 (________21379), .Q
       (___090__21711));
  nnd2s1 _______448463(.DIN1 (___09___20788), .DIN2 (________22674), .Q
       (___0_0__21686));
  nnd2s1 ____0__448464(.DIN1 (___9____20676), .DIN2 (____0___21816), .Q
       (____9___21805));
  hi1s1 _____9_448465(.DIN (___0____21682), .Q (________25044));
  hi1s1 _______448466(.DIN (________24660), .Q (________22069));
  hi1s1 _______448467(.DIN (___90___23350), .Q (________21997));
  hi1s1 ______448468(.DIN (__9_9___26695), .Q (____0___21912));
  nnd2s1 _______448469(.DIN1 (________21063), .DIN2 (________21378), .Q
       (___0____21654));
  nor2s1 _______448470(.DIN1 (________22136), .DIN2 (________20944), .Q
       (________21798));
  hi1s1 _______448471(.DIN (__9_____26717), .Q (__9_____26964));
  nor2s1 _______448472(.DIN1 (___90___20608), .DIN2 (________21370), .Q
       (____0___21908));
  hi1s1 ____0__448473(.DIN (________21845), .Q (________21928));
  and2s1 _____0_448474(.DIN1 (________21377), .DIN2 (________21214), .Q
       (________21920));
  nnd2s1 ______448475(.DIN1 (________20937), .DIN2 (____0___21359), .Q
       (_____0__22023));
  nnd2s1 ______448476(.DIN1 (___9____21614), .DIN2 (________21203), .Q
       (____9___21806));
  nnd2s1 _______448477(.DIN1 (___9____21614), .DIN2 (____9___21070), .Q
       (________22054));
  nor2s1 _____0_448478(.DIN1 (________21495), .DIN2 (________21376), .Q
       (___0____21703));
  hi1s1 _____0_448479(.DIN (__9_00__26798), .Q (_____9__22127));
  nnd2s1 _______448480(.DIN1 (___9____21614), .DIN2 (________21053), .Q
       (_____0__21995));
  nnd2s1 ____00_448481(.DIN1 (________21519), .DIN2 (____0___21267), .Q
       (____9___21983));
  nor2s1 _______448482(.DIN1 (______18933), .DIN2 (________20805), .Q
       (_____9__22223));
  nor2s1 _______448483(.DIN1 (________21978), .DIN2 (___0____20777), .Q
       (___0____21678));
  nnd2s1 ____90_448484(.DIN1 (___0____20736), .DIN2 (____9___21256), .Q
       (________21892));
  nnd2s1 ___0_448485(.DIN1 (________20936), .DIN2 (________21375), .Q
       (___90___22451));
  nor2s1 _______448486(.DIN1 (___99___19764), .DIN2 (________21402), .Q
       (_____0__22855));
  hi1s1 ____0__448487(.DIN (_____0__21374), .Q (________24563));
  nnd2s1 ___0___448488(.DIN1 (___0____20725), .DIN2
       (____0____________0_), .Q (_____0__22138));
  nnd2s1 _______448489(.DIN1 (____0___20796), .DIN2 (________21477), .Q
       (_____0__22108));
  nor2s1 _____9_448490(.DIN1 (________21409), .DIN2 (___9____20679), .Q
       (____0___22363));
  nnd2s1 _______448491(.DIN1 (____9___20975), .DIN2 (________21373), .Q
       (________21916));
  nnd2s1 _____9_448492(.DIN1 (________20940), .DIN2 (_____9__21199), .Q
       (____00__21904));
  nor2s1 _____9_448493(.DIN1 (___0____21651), .DIN2 (____0___21170), .Q
       (________21957));
  nor2s1 ___0___448494(.DIN1 (________21472), .DIN2 (___99___20696), .Q
       (_____0__22099));
  nnd2s1 _______448495(.DIN1 (____9___20977), .DIN2 (________21372), .Q
       (_____0__23028));
  nnd2s1 ______448496(.DIN1 (___0____20776), .DIN2 (____9___21897), .Q
       (________25158));
  nor2s1 _______448497(.DIN1 (________19613), .DIN2 (________21371), .Q
       (________22381));
  nnd2s1 _____9_448498(.DIN1 (_____0__21020), .DIN2 (________20210), .Q
       (________24682));
  or2s1 _______448499(.DIN1 (________21495), .DIN2 (________21024), .Q
       (________24216));
  nor2s1 _______448500(.DIN1 (____99__20509), .DIN2 (________21370), .Q
       (________24680));
  or2s1 _______448501(.DIN1 (___9____21610), .DIN2 (________21406), .Q
       (____9___21902));
  hi1s1 ___0___448502(.DIN (___9____26174), .Q (___9____23399));
  and2s1 ______448503(.DIN1 (________20926), .DIN2 (___0____21690), .Q
       (____9___22799));
  or2s1 _______448504(.DIN1 (________22136), .DIN2 (________21512), .Q
       (________21996));
  or2s1 ______448505(.DIN1 (____0____29098), .DIN2 (____9___20878), .Q
       (________21973));
  nor2s1 _______448506(.DIN1 (____9____30882), .DIN2 (________20804),
       .Q (_____9__25918));
  nnd2s1 _______448507(.DIN1 (________20958), .DIN2 (________21368), .Q
       (___9____22482));
  or2s1 _______448508(.DIN1 (____9___21353), .DIN2 (________21402), .Q
       (________23938));
  nor2s1 ______448509(.DIN1 (________21234), .DIN2 (________21367), .Q
       (________24724));
  nor2s1 _______448510(.DIN1 (________21488), .DIN2 (___0____20717), .Q
       (____0___22362));
  and2s1 _______448511(.DIN1 (_________31648), .DIN2 (________21366),
       .Q (_________29668));
  and2s1 ___0___448512(.DIN1 (_____9__21484), .DIN2 (_____0__21365), .Q
       (________22093));
  nnd2s1 _______448513(.DIN1 (___9____20630), .DIN2 (___0____21663), .Q
       (________23539));
  nor2s1 _______448514(.DIN1 (___0____21659), .DIN2 (________21371), .Q
       (________22343));
  nor2s1 ____0__448515(.DIN1 (________21409), .DIN2 (____09__21364), .Q
       (________22387));
  nnd2s1 _______448516(.DIN1 (___9____20688), .DIN2 (____9___21346), .Q
       (________22370));
  nor2s1 _______448517(.DIN1 (____0___21363), .DIN2 (___0____20772), .Q
       (____9___22078));
  nnd2s1 ____09_448518(.DIN1 (____0___20987), .DIN2 (________22341), .Q
       (____9___21901));
  hi1s1 ______448519(.DIN (___0____23502), .Q (____0___22263));
  nnd2s1 _____0_448520(.DIN1 (________21051), .DIN2 (___0____21663), .Q
       (________22967));
  or2s1 _______448521(.DIN1 (____0___21362), .DIN2 (________21367), .Q
       (________22150));
  nnd2s1 _______448522(.DIN1 (_____9__21334), .DIN2 (____0___21361), .Q
       (____0___21910));
  nor2s1 _______448523(.DIN1 (________20369), .DIN2 (___9____21620), .Q
       (________21959));
  nnd2s1 _______448524(.DIN1 (________20896), .DIN2 (____0___21988), .Q
       (________23698));
  nnd2s1 _____0_448525(.DIN1 (___9_9__20671), .DIN2 (________21893), .Q
       (_____0__22366));
  nnd2s1 ____0__448526(.DIN1 (_____0__20952), .DIN2 (____0___21360), .Q
       (___9____22461));
  nnd2s1 ____0__448527(.DIN1 (_____0__22690), .DIN2 (________20861), .Q
       (________23642));
  and2s1 _____448528(.DIN1 (________21456), .DIN2 (________21387), .Q
       (_____9__21923));
  nnd2s1 ______448529(.DIN1 (____0___21359), .DIN2 (___0_9__20761), .Q
       (________23922));
  nor2s1 ___0_0_448530(.DIN1 (___0____21660), .DIN2 (___99___20693), .Q
       (________22220));
  nnd2s1 ___0___448531(.DIN1 (____9___20880), .DIN2 (____0___21816), .Q
       (________26074));
  nnd2s1 ______448532(.DIN1 (____0___20793), .DIN2 (____0___21988), .Q
       (___9____26223));
  nnd2s1 ______448533(.DIN1 (___9____21614), .DIN2 (________21211), .Q
       (____0___25560));
  nnd2s1 _____9_448534(.DIN1 (________25726), .DIN2 (____0___21358), .Q
       (___0____23488));
  nor2s1 ____0_448535(.DIN1 (___9____19725), .DIN2 (____0___20989), .Q
       (____99__24517));
  nnd2s1 ____0__448536(.DIN1 (________21491), .DIN2 (________21470), .Q
       (____9___25168));
  nor2s1 ______448537(.DIN1 (____0___21357), .DIN2 (________20811), .Q
       (________25715));
  nnd2s1 ______448538(.DIN1 (____0___21356), .DIN2 (________20312), .Q
       (____9___23800));
  and2s1 _____9_448539(.DIN1 (___0____20749), .DIN2 (________22341), .Q
       (________23233));
  nor2s1 _____9_448540(.DIN1 (____00__21355), .DIN2 (___9____20673), .Q
       (_____9__25001));
  nnd2s1 _____0_448541(.DIN1 (________20545), .DIN2 (___0____21663), .Q
       (___0____25333));
  hi1s1 _______448542(.DIN (___99___23429), .Q (__9_____26655));
  and2s1 _____448543(.DIN1 (____9___21257), .DIN2 (____99__21354), .Q
       (___9____26213));
  nor2s1 _______448544(.DIN1 (________21341), .DIN2 (___9____21620), .Q
       (________22965));
  nnd2s1 _______448545(.DIN1 (___0____20769), .DIN2 (____0___21988), .Q
       (________21925));
  nor2s1 _______448546(.DIN1 (____0___21362), .DIN2 (___0_0__20733), .Q
       (__9_____26650));
  nor2s1 ______448547(.DIN1 (____9___21353), .DIN2 (________21370), .Q
       (_____0__24173));
  nnd2s1 _______448548(.DIN1 (_____9__21000), .DIN2 (_____0__22118), .Q
       (________25419));
  nor2s1 _______448549(.DIN1 (____9___21352), .DIN2 (___0____25354), .Q
       (__90_0__26291));
  nor2s1 ___0__448550(.DIN1 (___0____21660), .DIN2 (________20873), .Q
       (____0___24798));
  and2s1 _______448551(.DIN1 (_____0__21010), .DIN2 (________21458), .Q
       (___9_0__26167));
  or2s1 ___0___448552(.DIN1 (_____9__21894), .DIN2 (________20871), .Q
       (__9_____26875));
  nor2s1 _____448553(.DIN1 (________21502), .DIN2 (____9___21347), .Q
       (________25980));
  nor2s1 _______448554(.DIN1 (_____0__21046), .DIN2 (________21402), .Q
       (________23273));
  nnd2s1 _______448555(.DIN1 (___0____20738), .DIN2 (____9___19200), .Q
       (________25035));
  nnd2s1 _______448556(.DIN1 (_____0__21001), .DIN2 (____9___19200), .Q
       (____9___23707));
  nor2s1 _______448557(.DIN1 (___9____19725), .DIN2 (___0____20778), .Q
       (___0____25303));
  or2s1 _______448558(.DIN1 (____9___21351), .DIN2 (____9___21350), .Q
       (_____9__25928));
  nnd2s1 _______448559(.DIN1 (________21002), .DIN2 (________21238), .Q
       (___909__22454));
  nnd2s1 ___0___448560(.DIN1 (____9___21349), .DIN2 (___99___20695), .Q
       (________22091));
  hi1s1 ___0___448561(.DIN (____9___21348), .Q (________22859));
  nor2s1 _______448562(.DIN1 (________21495), .DIN2 (____9___21347), .Q
       (________25887));
  nnd2s1 _______448563(.DIN1 (____9___21346), .DIN2 (___0____20759), .Q
       (___9____22463));
  nor2s1 _______448564(.DIN1 (________21333), .DIN2 (________20964), .Q
       (____0___23085));
  nor2s1 _______448565(.DIN1 (________21506), .DIN2 (____9___20882), .Q
       (_____0__22924));
  hi1s1 ___0___448566(.DIN (____90__21345), .Q (__9_____26387));
  nor2s1 _____9_448567(.DIN1 (________21409), .DIN2 (_____0__20913), .Q
       (________22185));
  nnd2s1 ___0___448568(.DIN1 (___0_9__20723), .DIN2 (________21373), .Q
       (________25734));
  nnd2s1 ___0__448569(.DIN1 (________21342), .DIN2 (____90__21801), .Q
       (________22677));
  nnd2s1 _______448570(.DIN1 (_________31648), .DIN2 (_____9__21344),
       .Q (____90___32662));
  nnd2s1 ______448571(.DIN1 (________21343), .DIN2 (________21477), .Q
       (___0_____27600));
  nnd2s1 ___0___448572(.DIN1 (________21342), .DIN2 (_____0__21365), .Q
       (___9____22495));
  nnd2s1 _____0_448573(.DIN1 (___0____20735), .DIN2 (________21458), .Q
       (________22818));
  nor2s1 ______448574(.DIN1 (____0___21363), .DIN2 (________21341), .Q
       (________22685));
  nnd2s1 ___0___448575(.DIN1 (________20906), .DIN2 (________22341), .Q
       (_____0__22952));
  nnd2s1 ______448576(.DIN1 (________21340), .DIN2 (________21486), .Q
       (________25392));
  nnd2s1 _______448577(.DIN1 (________21040), .DIN2 (________21378), .Q
       (________22946));
  nor2s1 _______448578(.DIN1 (________21339), .DIN2 (___0____20768), .Q
       (________25722));
  nnd2s1 _____0_448579(.DIN1 (____00__20886), .DIN2 (________21373), .Q
       (__9_____26779));
  nor2s1 ____0__448580(.DIN1 (________21472), .DIN2 (________21338), .Q
       (________25524));
  and2s1 _____9_448581(.DIN1 (________20822), .DIN2 (________21337), .Q
       (___0_0__23481));
  hi1s1 ___0___448582(.DIN (________21336), .Q (___9_0__26157));
  nor2s1 _______448583(.DIN1 (________21505), .DIN2 (___0____20754), .Q
       (______0__28751));
  nnd2s1 _______448584(.DIN1 (___0____20757), .DIN2 (________20380), .Q
       (___0__0__27287));
  nnd2s1 _____9_448585(.DIN1 (_____9__21400), .DIN2 (_____0__21335), .Q
       (________23119));
  and2s1 _____9_448586(.DIN1 (___9____21614), .DIN2 (_____9__21287), .Q
       (__9_____26472));
  nnd2s1 _______448587(.DIN1 (____09__20428), .DIN2 (___0____21663), .Q
       (__9_____26358));
  nnd2s1 ______448588(.DIN1 (________20950), .DIN2 (____0___19948), .Q
       (______0__30591));
  nnd2s1 _______448589(.DIN1 (_____9__21334), .DIN2 (___0____21663), .Q
       (______0__28974));
  nor2s1 _____448590(.DIN1 (_____9__21894), .DIN2 (____0___20797), .Q
       (____09__22365));
  nor2s1 _____0_448591(.DIN1 (________21333), .DIN2 (________20916), .Q
       (__9_____26553));
  nnd2s1 ______448592(.DIN1 (________21094), .DIN2 (________20843), .Q
       (___00___23438));
  nnd2s1 _______448593(.DIN1 (____09__20798), .DIN2 (____9___21346), .Q
       (__9_9___26791));
  nnd2s1 ___0_0_448594(.DIN1 (________21332), .DIN2 (________21373), .Q
       (__9_____26877));
  nnd2s1 _____448595(.DIN1 (________21477), .DIN2 (________21509), .Q
       (________21930));
  nor2s1 _______448596(.DIN1 (________21508), .DIN2 (________20960), .Q
       (___0_____27430));
  ib1s1 _______448597(.DIN (________21469), .Q (________21758));
  nor2s1 ______448598(.DIN1 (______9__33436), .DIN2 (_________33797),
       .Q (_________34159));
  nor2s1 ___0___448599(.DIN1 (___9____20622), .DIN2 (____9___20884), .Q
       (_________33103));
  nor2s1 _______448600(.DIN1 (________22050), .DIN2 (___9____20621), .Q
       (________21331));
  and2s1 _______448601(.DIN1 (____0___20421), .DIN2 (________22109), .Q
       (________21330));
  nor2s1 _______448602(.DIN1 (________19929), .DIN2 (________20494), .Q
       (________21329));
  nor2s1 ______448603(.DIN1 (____9___20412), .DIN2 (____9___20883), .Q
       (________21328));
  or2s1 _______448604(.DIN1 (________21180), .DIN2 (_____9__21326), .Q
       (_____0__21327));
  nnd2s1 _______448605(.DIN1 (_____0__21279), .DIN2 (____9___19297), .Q
       (________21325));
  nor2s1 _____448606(.DIN1 (________21323), .DIN2 (________20993), .Q
       (________21324));
  nnd2s1 _______448607(.DIN1 (____90__21066), .DIN2 (________20459), .Q
       (________21322));
  nor2s1 _______448608(.DIN1 (________21505), .DIN2 (___9____20631), .Q
       (________21321));
  nor2s1 _______448609(.DIN1 (________21319), .DIN2 (________21424), .Q
       (________21320));
  nnd2s1 _______448610(.DIN1 (________21281), .DIN2 (________20076), .Q
       (________21318));
  hi1s1 ____0_448611(.DIN (________21376), .Q (_____0__21317));
  nnd2s1 ___0__448612(.DIN1 (________21315), .DIN2 (____0___20229), .Q
       (_____9__21316));
  nnd2s1 ___09__448613(.DIN1 (________21313), .DIN2 (________20490), .Q
       (________21314));
  nnd2s1 ______448614(.DIN1 (________20472), .DIN2 (_____9__19476), .Q
       (________21312));
  nor2s1 _______448615(.DIN1 (________21310), .DIN2 (_____9__21326), .Q
       (________21311));
  nor2s1 ___09__448616(.DIN1 (____9___20319), .DIN2 (________20480), .Q
       (________21309));
  nor2s1 _____0_448617(.DIN1 (________21059), .DIN2 (____9___21162), .Q
       (_____0__21308));
  nor2s1 ___090_448618(.DIN1 (________21306), .DIN2 (________21104), .Q
       (_____9__21307));
  nor2s1 _______448619(.DIN1 (________21153), .DIN2 (________21291), .Q
       (________21305));
  nor2s1 _______448620(.DIN1 (____9___20322), .DIN2 (________20449), .Q
       (________21304));
  or2s1 _______448621(.DIN1 (____99__19685), .DIN2 (_____0__21173), .Q
       (________21303));
  nor2s1 _______448622(.DIN1 (________21310), .DIN2 (________21424), .Q
       (________21302));
  nor2s1 ___0___448623(.DIN1 (____0___21265), .DIN2 (________21300), .Q
       (________21301));
  nor2s1 _______448624(.DIN1 (_____0__21298), .DIN2 (________20496), .Q
       (________21299));
  nnd2s1 _______448625(.DIN1 (_____0__20465), .DIN2 (________20213), .Q
       (_____9__21297));
  nnd2s1 ___0___448626(.DIN1 (____9___20414), .DIN2 (________21372), .Q
       (________21296));
  nor2s1 _______448627(.DIN1 (____0___21357), .DIN2 (____0___20424), .Q
       (________21295));
  hi1s1 _______448628(.DIN (________21478), .Q (________21294));
  nnd2s1 ______448629(.DIN1 (________20458), .DIN2 (________21778), .Q
       (________21293));
  nor2s1 _______448630(.DIN1 (________21276), .DIN2 (________21291), .Q
       (________21292));
  or2s1 ___0___448631(.DIN1 (________22050), .DIN2 (_____9__20483), .Q
       (________21290));
  nor2s1 ___0__448632(.DIN1 (________20195), .DIN2 (________20541), .Q
       (________21289));
  nnd2s1 _______448633(.DIN1 (________21212), .DIN2 (_____9__21287), .Q
       (_____0__21288));
  hi1s1 _______448634(.DIN (_____0__21494), .Q (________21286));
  nnd2s1 _______448635(.DIN1 (________21189), .DIN2 (_____0__21821), .Q
       (________21285));
  or2s1 ___0_9_448636(.DIN1 (________21283), .DIN2 (________20004), .Q
       (________21284));
  nnd2s1 _____448637(.DIN1 (________21281), .DIN2 (________21006), .Q
       (________21282));
  nnd2s1 _______448638(.DIN1 (_____0__21279), .DIN2 (_____9__21278), .Q
       (________21280));
  nor2s1 _______448639(.DIN1 (________21276), .DIN2 (_____9__21326), .Q
       (________21277));
  and2s1 ______448640(.DIN1 (________21236), .DIN2 (___0____21684), .Q
       (________21275));
  hi1s1 ____0_448641(.DIN (_____9__21334), .Q (________21274));
  nnd2s1 ______448642(.DIN1 (_____9__21182), .DIN2 (_______19050), .Q
       (________21273));
  or2s1 ___0_9_448643(.DIN1 (________20280), .DIN2 (___9____20640), .Q
       (________21272));
  nnd2s1 ___0___448644(.DIN1 (________20488), .DIN2 (___0____20773), .Q
       (________21271));
  or2s1 ___0__448645(.DIN1 (inData[29]), .DIN2 (____9___21158), .Q
       (_____0__21270));
  nnd2s1 ___0___448646(.DIN1 (________20577), .DIN2 (________22131), .Q
       (____09__21269));
  nnd2s1 ___0__448647(.DIN1 (____90__20595), .DIN2 (____0___21267), .Q
       (____0___21268));
  nor2s1 ___0___448648(.DIN1 (____0___21265), .DIN2 (________21424), .Q
       (____0___21266));
  nor2s1 ___0__448649(.DIN1 (____0___21263), .DIN2 (_____9__21093), .Q
       (____0___21264));
  nor2s1 ___0_9_448650(.DIN1 (________20407), .DIN2 (________20093), .Q
       (____0___21262));
  nor2s1 ___0_9_448651(.DIN1 (____00__21260), .DIN2 (________21217), .Q
       (____0___21261));
  or2s1 ___448652(.DIN1 (_________9_______18809), .DIN2
       (_____00__33954), .Q (____99__21259));
  nnd2s1 ___09__448653(.DIN1 (____9___21257), .DIN2 (____9___21256), .Q
       (____9___21258));
  nor2s1 ___09__448654(.DIN1 (________20453), .DIN2 (________20161), .Q
       (____9___21255));
  nor2s1 ___09__448655(.DIN1 (________20333), .DIN2 (____9___21253), .Q
       (____9___21254));
  nnd2s1 ___09_448656(.DIN1 (________21373), .DIN2 (_____0__20567), .Q
       (____9___21252));
  and2s1 ___09__448657(.DIN1 (________22312), .DIN2 (________20578), .Q
       (____9___21251));
  nor2s1 ___09__448658(.DIN1 (___90___21546), .DIN2 (________20527), .Q
       (____90__21250));
  nnd2s1 ___09__448659(.DIN1 (________20350), .DIN2 (________20432), .Q
       (_____9__21249));
  nor2s1 ___09__448660(.DIN1 (________20477), .DIN2 (________21224), .Q
       (________21248));
  and2s1 ___09__448661(.DIN1 (________20526), .DIN2 (________21489), .Q
       (________21247));
  or2s1 ___09__448662(.DIN1 (________21245), .DIN2 (_____0__20576), .Q
       (________21246));
  nor2s1 _______448663(.DIN1 (________20563), .DIN2 (_____9__20529), .Q
       (________21244));
  nnd2s1 _______448664(.DIN1 (___000___27171), .DIN2 (_________29585),
       .Q (________21243));
  nnd2s1 ______448665(.DIN1 (___9____20618), .DIN2 (________21241), .Q
       (________21242));
  hi1s1 _______448666(.DIN (________21338), .Q (_____0__21240));
  nor2s1 _______448667(.DIN1 (________21495), .DIN2 (_____0__20585), .Q
       (________21415));
  nor2s1 ____0__448668(.DIN1 (_____9__21239), .DIN2 (________20553), .Q
       (_____0__21831));
  nnd2s1 ____90_448669(.DIN1 (___9____20645), .DIN2 (____9___21069), .Q
       (____0___21814));
  nnd2s1 ____448670(.DIN1 (_____9__21219), .DIN2 (___0____21694), .Q
       (________22024));
  nnd2s1 ____00_448671(.DIN1 (________20535), .DIN2 (________21238), .Q
       (________21799));
  nnd2s1 ___099_448672(.DIN1 (________21223), .DIN2 (________21205), .Q
       (________21791));
  nnd2s1 ___09__448673(.DIN1 (________21237), .DIN2 (_____9__22435), .Q
       (________23100));
  nnd2s1 _____9_448674(.DIN1 (________21236), .DIN2 (________20543), .Q
       (___0_9__21695));
  nor2s1 _______448675(.DIN1 (____0___19953), .DIN2 (________20447), .Q
       (___0____21693));
  hi1s1 _______448676(.DIN (________21235), .Q (_____0__21773));
  nnd2s1 _______448677(.DIN1 (________21215), .DIN2 (________21238), .Q
       (___0_9__21675));
  nor2s1 _______448678(.DIN1 (________21234), .DIN2 (________21047), .Q
       (________21926));
  and2s1 ______448679(.DIN1 (_____0__21279), .DIN2 (________21233), .Q
       (________21919));
  or2s1 ___09__448680(.DIN1 (________20258), .DIN2 (________23052), .Q
       (____0___21817));
  nnd2s1 _______448681(.DIN1 (________21232), .DIN2 (________20468), .Q
       (________21496));
  nnd2s1 ___09_448682(.DIN1 (________21231), .DIN2 (___9_0__21561), .Q
       (____9___21439));
  nor2s1 ___09__448683(.DIN1 (_____0__21230), .DIN2 (________21062), .Q
       (___0____21673));
  nnd2s1 ___09__448684(.DIN1 (_____9__20455), .DIN2 (___9_0__21561), .Q
       (___09___21716));
  nor2s1 ___099_448685(.DIN1 (_____9__21229), .DIN2 (________21227), .Q
       (_____9__21792));
  nor2s1 ___09__448686(.DIN1 (________21228), .DIN2 (________21227), .Q
       (________21775));
  nnd2s1 ____0_448687(.DIN1 (___90___20609), .DIN2 (________21226), .Q
       (________21435));
  nnd2s1 ____0__448688(.DIN1 (_____0__20429), .DIN2 (________20954), .Q
       (___0____21672));
  or2s1 ____0_448689(.DIN1 (____0________________18647), .DIN2
       (___90___20610), .Q (___0____21701));
  nnd2s1 _______448690(.DIN1 (___9____20627), .DIN2 (____9___21897), .Q
       (________21781));
  nnd2s1 _______448691(.DIN1 (________21044), .DIN2 (________21776), .Q
       (____9___21348));
  nnd2s1 _______448692(.DIN1 (________21281), .DIN2 (_____0__20827), .Q
       (________21336));
  nnd2s1 ____0_448693(.DIN1 (_____9__20539), .DIN2 (________21226), .Q
       (________21380));
  nor2s1 _____0_448694(.DIN1 (________21323), .DIN2 (________21196), .Q
       (____90__21345));
  hi1s1 _______448695(.DIN (_________35076), .Q (____0_0__30932));
  nor2s1 _______448696(.DIN1 (________21234), .DIN2 (________21064), .Q
       (________22132));
  nnd2s1 _______448697(.DIN1 (________21281), .DIN2 (___9____20668), .Q
       (___0_0__22608));
  hi1s1 _______448698(.DIN (________21225), .Q (___0____24368));
  nor2s1 ____9_448699(.DIN1 (________21224), .DIN2 (________20214), .Q
       (________21871));
  nnd2s1 ____0_448700(.DIN1 (________21223), .DIN2 (________21222), .Q
       (___009__23445));
  nnd2s1 ____0_448701(.DIN1 (________21042), .DIN2 (________21222), .Q
       (________21850));
  nnd2s1 _______448702(.DIN1 (________21232), .DIN2 (___9_0__20654), .Q
       (___9____23379));
  nor2s1 ______448703(.DIN1 (____0___21363), .DIN2 (________20571), .Q
       (___0____24398));
  nnd2s1 _____0_448704(.DIN1 (________21034), .DIN2 (____90__21156), .Q
       (___90___23350));
  nnd2s1 _______448705(.DIN1 (________21281), .DIN2 (________20838), .Q
       (___0____23502));
  nor2s1 ____0__448706(.DIN1 (________20840), .DIN2 (________21221), .Q
       (________24632));
  nnd2s1 ____0__448707(.DIN1 (________21223), .DIN2 (________21201), .Q
       (___9____22505));
  nnd2s1 ____0__448708(.DIN1 (________20487), .DIN2 (___9__18934), .Q
       (_____9__21800));
  nor2s1 _______448709(.DIN1 (___9____20666), .DIN2 (_____0__21210), .Q
       (________24132));
  hi1s1 _______448710(.DIN (_____0__21220), .Q (________24821));
  nor2s1 ______448711(.DIN1 (____9____30882), .DIN2 (___0____20737), .Q
       (________24475));
  nnd2s1 _______448712(.DIN1 (_____9__21219), .DIN2 (________21218), .Q
       (____0___24705));
  nnd2s1 _______448713(.DIN1 (________21232), .DIN2 (________20335), .Q
       (________22149));
  xnr2s1 _______448714(.DIN1 (_____0__19153), .DIN2 (_____99__29264),
       .Q (____000__28138));
  and2s1 _______448715(.DIN1 (________21281), .DIN2 (________20828), .Q
       (_____0__24616));
  or2s1 _______448716(.DIN1 (________20215), .DIN2 (________21217), .Q
       (_____0__23933));
  and2s1 _______448717(.DIN1 (________21194), .DIN2 (________21216), .Q
       (___99___23435));
  nnd2s1 ______448718(.DIN1 (________21215), .DIN2 (________21511), .Q
       (____90__23792));
  hi1s1 ____0_448719(.DIN (________21214), .Q (__9_____26440));
  nnd2s1 ____0__448720(.DIN1 (________21223), .DIN2 (________21023), .Q
       (________25803));
  nor2s1 _____0_448721(.DIN1 (________21213), .DIN2 (________20443), .Q
       (____0___24888));
  nor2s1 _______448722(.DIN1 (________21501), .DIN2 (________20462), .Q
       (__9_____26660));
  nor2s1 _______448723(.DIN1 (____9___21067), .DIN2 (_____0__20484), .Q
       (________24902));
  nnd2s1 ____0__448724(.DIN1 (____0___20422), .DIN2 (________21373), .Q
       (________25704));
  nnd2s1 _______448725(.DIN1 (________21212), .DIN2 (________21211), .Q
       (____00__24792));
  nor2s1 _______448726(.DIN1 (___9____20656), .DIN2 (_____0__21210), .Q
       (___09___24420));
  nor2s1 _______448727(.DIN1 (_____9__20557), .DIN2 (________21207), .Q
       (________24183));
  nnd2s1 _______448728(.DIN1 (________21204), .DIN2 (________21211), .Q
       (________23236));
  hi1s1 ____0__448729(.DIN (_____9__21209), .Q (________22688));
  and2s1 ____0__448730(.DIN1 (_____9__21045), .DIN2 (________21043), .Q
       (________22730));
  nnd2s1 _______448731(.DIN1 (________20556), .DIN2 (________21208), .Q
       (__9_00__26798));
  nor2s1 _______448732(.DIN1 (________20199), .DIN2 (________20591), .Q
       (________24659));
  nor2s1 _______448733(.DIN1 (___9____20615), .DIN2 (________21207), .Q
       (________25064));
  nnd2s1 _______448734(.DIN1 (___9____20616), .DIN2 (____9___19200), .Q
       (__9_____26871));
  nnd2s1 _______448735(.DIN1 (_____0__21200), .DIN2 (________21206), .Q
       (__9_____26631));
  hi1s1 _______448736(.DIN (____0___21356), .Q (________21741));
  nnd2s1 ____0__448737(.DIN1 (_____9__21065), .DIN2 (________21205), .Q
       (____0___25661));
  nnd2s1 _____448738(.DIN1 (________21202), .DIN2 (________21222), .Q
       (___09___23526));
  and2s1 _____0_448739(.DIN1 (________20554), .DIN2 (________21226), .Q
       (__90_0__26281));
  nnd2s1 _______448740(.DIN1 (________20457), .DIN2 (________20080), .Q
       (_________29496));
  nnd2s1 _______448741(.DIN1 (________20568), .DIN2 (______0__28643),
       .Q (________21469));
  nnd2s1 _______448742(.DIN1 (________21204), .DIN2 (________21203), .Q
       (________23222));
  nnd2s1 ____0__448743(.DIN1 (________21202), .DIN2 (________21201), .Q
       (_____0__23695));
  hi1s1 ____0__448744(.DIN (____0___21358), .Q (__9__9__26921));
  nnd2s1 _______448745(.DIN1 (_____0__21200), .DIN2 (_____9__21199), .Q
       (___0____22601));
  nnd2s1 _______448746(.DIN1 (________21232), .DIN2 (________20168), .Q
       (___99___23429));
  nor2s1 _____448747(.DIN1 (________21333), .DIN2 (________20440), .Q
       (________22106));
  nnd2s1 _______448748(.DIN1 (________20528), .DIN2 (____9___21346), .Q
       (___0____24393));
  nor2s1 _____0_448749(.DIN1 (________21198), .DIN2 (___9____20637), .Q
       (____0___22812));
  nor2s1 _____0_448750(.DIN1 (________21197), .DIN2 (________20409), .Q
       (________26101));
  nor2s1 _______448751(.DIN1 (________21506), .DIN2 (________21195), .Q
       (_____9__25145));
  nnd2s1 _______448752(.DIN1 (___9____20629), .DIN2 (___9__18934), .Q
       (________25604));
  nor2s1 ____09_448753(.DIN1 (________21788), .DIN2 (________21196), .Q
       (__9_____26499));
  nnd2s1 _______448754(.DIN1 (____9___20600), .DIN2 (_____9__19965), .Q
       (____0____30044));
  or2s1 _____0_448755(.DIN1 (________21409), .DIN2 (________21195), .Q
       (___99___26242));
  nnd2s1 _______448756(.DIN1 (________21194), .DIN2 (________21193), .Q
       (________24660));
  nnd2s1 _______448757(.DIN1 (______0__35088), .DIN2 (________20309),
       .Q (_________28737));
  nor2s1 _______448758(.DIN1 (____0___20233), .DIN2 (________21192), .Q
       (_____0___31450));
  nnd2s1 _______448759(.DIN1 (_____0__20456), .DIN2 (________20831), .Q
       (_________32606));
  nor2s1 _______448760(.DIN1 (___0____19831), .DIN2 (________20397), .Q
       (____9____31798));
  nor2s1 _______448761(.DIN1 (________19607), .DIN2 (________21192), .Q
       (____99___31805));
  nnd2s1 _______448762(.DIN1 (___9_0__20624), .DIN2 (_____0__21191), .Q
       (_________33925));
  nor2s1 ____448763(.DIN1 (____9___20501), .DIN2 (________20489), .Q
       (_________34116));
  and2s1 _______448764(.DIN1 (________21189), .DIN2 (________21188), .Q
       (_____9__21190));
  and2s1 _______448765(.DIN1 (________21141), .DIN2 (________20241), .Q
       (________21187));
  nnd2s1 _______448766(.DIN1 (____9___20418), .DIN2 (inData[6]), .Q
       (________21186));
  nnd2s1 ______448767(.DIN1 (____0___19854), .DIN2 (________20473), .Q
       (________21185));
  xor2s1 _____9_448768(.DIN1 (_________31376), .DIN2 (____0____31818),
       .Q (________21184));
  nnd2s1 _______448769(.DIN1 (_____9__21182), .DIN2
       (_________________18693), .Q (_____0__21183));
  nor2s1 ______448770(.DIN1 (________21180), .DIN2 (________21424), .Q
       (________21181));
  nor2s1 _______448771(.DIN1 (_____9__20125), .DIN2 (________21133), .Q
       (________21179));
  hi1s1 _______448772(.DIN (________26099), .Q (________21178));
  nor2s1 ______448773(.DIN1 (________20845), .DIN2 (________21176), .Q
       (________21177));
  or2s1 _______448774(.DIN1 (________21174), .DIN2 (_____0__21173), .Q
       (________21175));
  and2s1 _______448775(.DIN1 (________21136), .DIN2 (________19433), .Q
       (____0___21172));
  hi1s1 ____0__448776(.DIN (____0___21170), .Q (____0___21171));
  nor2s1 _______448777(.DIN1 (___9____21610), .DIN2 (___9_9__20633), .Q
       (____0___21169));
  nor2s1 _______448778(.DIN1 (____0___21167), .DIN2 (________20498), .Q
       (____0___21168));
  xor2s1 ___0___448779(.DIN1 (____________18893), .DIN2
       (_________31505), .Q (____00__21166));
  nnd2s1 _______448780(.DIN1 (________20486), .DIN2 (inData[4]), .Q
       (____99__21165));
  nor2s1 _______448781(.DIN1 (___9____20625), .DIN2 (________21113), .Q
       (____9___21164));
  nor2s1 _____0_448782(.DIN1 (________20292), .DIN2 (____9___21162), .Q
       (____9___21163));
  nnd2s1 ______448783(.DIN1 (___9____20619), .DIN2 (inData[10]), .Q
       (____9___21161));
  and2s1 _______448784(.DIN1 (____9___21257), .DIN2 (____0___20516), .Q
       (____9___21160));
  nnd2s1 ___0_9_448785(.DIN1 (____9___21158), .DIN2 (________20285), .Q
       (____9___21159));
  nnd2s1 ______448786(.DIN1 (____9___21257), .DIN2 (____90__21156), .Q
       (____9___21157));
  nor2s1 ___0___448787(.DIN1 (________19999), .DIN2 (________20560), .Q
       (_____9__21155));
  or2s1 _______448788(.DIN1 (________21153), .DIN2 (________21300), .Q
       (________21154));
  or2s1 ___0___448789(.DIN1 (____0___19859), .DIN2 (___90___20611), .Q
       (________21152));
  nnd2s1 ______448790(.DIN1 (________20452), .DIN2 (____9___21897), .Q
       (________21151));
  hi1s1 ____0__448791(.DIN (________21148), .Q (________21149));
  nnd2s1 _______448792(.DIN1 (________21212), .DIN2 (________21397), .Q
       (_____0__21147));
  nor2s1 ______448793(.DIN1 (________21145), .DIN2 (________21144), .Q
       (_____9__21146));
  hi1s1 ____0__448794(.DIN (________25864), .Q (________21143));
  nnd2s1 ____0__448795(.DIN1 (________19916), .DIN2 (________20475), .Q
       (________21142));
  nnd2s1 ____09_448796(.DIN1 (___0____20710), .DIN2 (________19560), .Q
       (_____0__21140));
  nnd2s1 ___09_448797(.DIN1 (_____0__21279), .DIN2 (________19568), .Q
       (_____9__21139));
  nor2s1 ___09__448798(.DIN1 (____0___20047), .DIN2 (________20589), .Q
       (________21138));
  and2s1 ______448799(.DIN1 (________21136), .DIN2 (________21025), .Q
       (________21137));
  or2s1 _______448800(.DIN1 (________21134), .DIN2 (________21133), .Q
       (________21135));
  nor2s1 ___0___448801(.DIN1 (________21131), .DIN2 (________21227), .Q
       (________21132));
  nor2s1 _______448802(.DIN1 (________19441), .DIN2 (_____9__21129), .Q
       (_____0__21130));
  nor2s1 ___09__448803(.DIN1 (________21127), .DIN2 (_____9__20438), .Q
       (________21128));
  and2s1 _______448804(.DIN1 (_____9__21129), .DIN2 (_________28734),
       .Q (________21126));
  hi1s1 ___0___448805(.DIN (________21124), .Q (________21125));
  nnd2s1 _______448806(.DIN1 (________20531), .DIN2 (________21122), .Q
       (________21123));
  nnd2s1 ___09_448807(.DIN1 (_____0__21120), .DIN2 (________21372), .Q
       (________21121));
  hi1s1 ____0__448808(.DIN (________21118), .Q (_____9__21119));
  or2s1 _______448809(.DIN1 (________21502), .DIN2 (________21058), .Q
       (________21117));
  and2s1 ______448810(.DIN1 (________20406), .DIN2 (________21115), .Q
       (________21116));
  nor2s1 _____9_448811(.DIN1 (________21750), .DIN2 (________21323), .Q
       (_____9__21112));
  nor2s1 _______448812(.DIN1 (_____0__20895), .DIN2 (________21133), .Q
       (________21111));
  nnd2s1 ___0___448813(.DIN1 (________21189), .DIN2 (________21777), .Q
       (________21110));
  nor2s1 _______448814(.DIN1 (___0____19803), .DIN2 (________20400), .Q
       (________21109));
  or2s1 _______448815(.DIN1 (___9_9__20681), .DIN2 (_____9__21326), .Q
       (________21108));
  nnd2s1 _______448816(.DIN1 (________21232), .DIN2 (________20150), .Q
       (________21107));
  nnd2s1 ___0___448817(.DIN1 (_____0__21056), .DIN2 (____0___21360), .Q
       (________21106));
  nor2s1 ___09__448818(.DIN1 (________21104), .DIN2 (________20191), .Q
       (________21105));
  nnd2s1 ___09__448819(.DIN1 (___9____20626), .DIN2 (________21136), .Q
       (_____0__21103));
  nnd2s1 ___09__448820(.DIN1 (_____0__20530), .DIN2 (________19877), .Q
       (_____9__21102));
  hi1s1 _______448821(.DIN (________21100), .Q (________21101));
  and2s1 _______448822(.DIN1 (_____9__21055), .DIN2 (________21098), .Q
       (________21099));
  nor2s1 ___0___448823(.DIN1 (________20190), .DIN2 (________20565), .Q
       (________21097));
  and2s1 _____0_448824(.DIN1 (_____9__21219), .DIN2 (_____9__20401), .Q
       (________21096));
  hi1s1 ____0_448825(.DIN (________21094), .Q (________21095));
  hi1s1 ____0__448826(.DIN (__9_____26639), .Q (________21092));
  hi1s1 _______448827(.DIN (____0___21447), .Q (________21091));
  nor2s1 _______448828(.DIN1 (________20850), .DIN2 (________21089), .Q
       (________21090));
  nor2s1 ______448829(.DIN1 (____00__21355), .DIN2 (_____9__21093), .Q
       (________21088));
  nor2s1 _______448830(.DIN1 (________21086), .DIN2 (_____9__20594), .Q
       (________21087));
  xor2s1 _______448831(.DIN1 (____09__21084), .DIN2 (____0___21083), .Q
       (_____0__21085));
  hi1s1 _______448832(.DIN (________25115), .Q (____0___21082));
  nor2s1 _____448833(.DIN1 (____0___21080), .DIN2 (________20573), .Q
       (____0___21081));
  xor2s1 _______448834(.DIN1 (_____99__29264), .DIN2 (outData[31]), .Q
       (____0___21079));
  nnd2s1 _______448835(.DIN1 (________19644), .DIN2 (________20592), .Q
       (____0___21078));
  or2s1 _______448836(.DIN1 (________23682), .DIN2 (________20495), .Q
       (____0___21077));
  xor2s1 _____0_448837(.DIN1 (______________18868), .DIN2
       (_____99__29264), .Q (____0___21076));
  nor2s1 _______448838(.DIN1 (________20158), .DIN2 (________21217), .Q
       (____00__21075));
  nnd2s1 _______448839(.DIN1 (________21232), .DIN2 (________20463), .Q
       (____99__21074));
  nnd2s1 _______448840(.DIN1 (________20533), .DIN2 (______18933), .Q
       (____9___21073));
  nor2s1 ___0___448841(.DIN1 (____9___21071), .DIN2 (____9___20411), .Q
       (____9___21072));
  hi1s1 ____0__448842(.DIN (________21371), .Q (___0____21665));
  and2s1 _______448843(.DIN1 (_____0__21279), .DIN2 (________21368), .Q
       (___9____22459));
  nnd2s1 ______448844(.DIN1 (________21204), .DIN2 (____9___21070), .Q
       (_____0__21374));
  nnd2s1 ______448845(.DIN1 (________21212), .DIN2 (________21203), .Q
       (________21417));
  nnd2s1 ____9__448846(.DIN1 (________20858), .DIN2 (____9___21069), .Q
       (________21386));
  hi1s1 _______448847(.DIN (____9___21068), .Q (____00__21811));
  nor2s1 _____0_448848(.DIN1 (________21488), .DIN2 (________21217), .Q
       (________21796));
  nor2s1 _____9_448849(.DIN1 (________20821), .DIN2 (________20481), .Q
       (___0____21644));
  hi1s1 ____0__448850(.DIN (________25973), .Q (___0____21670));
  nnd2s1 ____9_448851(.DIN1 (___9_0__20614), .DIN2 (____9___20223), .Q
       (_____0__22206));
  nor2s1 ____9__448852(.DIN1 (_____9__21229), .DIN2 (____9___21067), .Q
       (________21420));
  nnd2s1 _____9_448853(.DIN1 (________20445), .DIN2 (____9___20881), .Q
       (___0____21655));
  nnd2s1 _______448854(.DIN1 (________21232), .DIN2 (________20176), .Q
       (________21760));
  or2s1 _______448855(.DIN1 (________20479), .DIN2 (________21054), .Q
       (____0___22180));
  nor2s1 ______448856(.DIN1 (________20830), .DIN2 (________20476), .Q
       (_____9__21782));
  nnd2s1 ___09_448857(.DIN1 (_____9__21065), .DIN2 (________21222), .Q
       (___0____21674));
  nor2s1 _____0_448858(.DIN1 (____0___21362), .DIN2 (________21064), .Q
       (________21755));
  nnd2s1 _____9_448859(.DIN1 (___9____20664), .DIN2 (____9___21069), .Q
       (________21390));
  hi1s1 ____0__448860(.DIN (________21063), .Q (___0____21661));
  nor2s1 ___09__448861(.DIN1 (_____9__20846), .DIN2 (________21062), .Q
       (________21787));
  hi1s1 ____0__448862(.DIN (________21061), .Q (________21790));
  hi1s1 ____0_448863(.DIN (_____0__21485), .Q (___0____21691));
  nor2s1 _____0_448864(.DIN1 (___9_0__20663), .DIN2 (________21060), .Q
       (___99___21628));
  and2s1 _______448865(.DIN1 (_____0__21279), .DIN2 (________21381), .Q
       (____9___22163));
  and2s1 ___099_448866(.DIN1 (________21202), .DIN2 (________21205), .Q
       (________21780));
  nor2s1 _______448867(.DIN1 (________21059), .DIN2 (________21113), .Q
       (________21395));
  and2s1 _______448868(.DIN1 (________21136), .DIN2 (________22141), .Q
       (_____0__21739));
  nor2s1 ______448869(.DIN1 (____9___20219), .DIN2 (________21217), .Q
       (___0_0__21676));
  nor2s1 _______448870(.DIN1 (________21058), .DIN2 (___9____20647), .Q
       (____0___21990));
  nnd2s1 _____0_448871(.DIN1 (____90__21066), .DIN2 (________21205), .Q
       (________21411));
  hi1s1 ____0__448872(.DIN (________21370), .Q (___0____21681));
  nnd2s1 ______448873(.DIN1 (________21057), .DIN2 (_____0__20866), .Q
       (________21771));
  nor2s1 _______448874(.DIN1 (________21922), .DIN2 (_____0__20492), .Q
       (________21866));
  nor2s1 _______448875(.DIN1 (________21197), .DIN2 (_____0__20558), .Q
       (____9___22986));
  nnd2s1 ____0_448876(.DIN1 (_____0__21056), .DIN2 (________22131), .Q
       (_____0__21729));
  nor2s1 _______448877(.DIN1 (________20829), .DIN2 (_____0__21210), .Q
       (___0____21682));
  hi1s1 ___0___448878(.DIN (_________30341), .Q (____9___22073));
  nor2s1 ____9__448879(.DIN1 (____9___20415), .DIN2 (________21052), .Q
       (____0___21815));
  nor2s1 ______448880(.DIN1 (____9___21984), .DIN2 (________20471), .Q
       (________22412));
  hi1s1 ___0___448881(.DIN (_________31134), .Q (___0_____27735));
  nor2s1 _______448882(.DIN1 (_____9__20836), .DIN2 (_____9__20448), .Q
       (_____0__22089));
  nor2s1 _______448883(.DIN1 (________20083), .DIN2 (________20572), .Q
       (___0_0__24352));
  nor2s1 ____9__448884(.DIN1 (________21049), .DIN2 (________21048), .Q
       (___0____21700));
  nnd2s1 _______448885(.DIN1 (________20941), .DIN2 (____0___20143), .Q
       (________22665));
  nnd2s1 ______448886(.DIN1 (_____9__21055), .DIN2 (______18933), .Q
       (________21746));
  or2s1 _______448887(.DIN1 (_____0__20402), .DIN2 (________21054), .Q
       (________23295));
  nnd2s1 _______448888(.DIN1 (________21053), .DIN2 (________21204), .Q
       (________23219));
  and2s1 _______448889(.DIN1 (________20431), .DIN2 (___9____20657), .Q
       (___0____21687));
  nnd2s1 ____9__448890(.DIN1 (____90__21066), .DIN2 (________19887), .Q
       (________23007));
  nor2s1 _______448891(.DIN1 (____90__19937), .DIN2 (________21052), .Q
       (________21845));
  and2s1 _______448892(.DIN1 (_____0__20549), .DIN2 (________21373), .Q
       (________25148));
  nnd2s1 ____0_448893(.DIN1 (___90___20607), .DIN2 (________19580), .Q
       (____9___21807));
  hi1s1 ___0___448894(.DIN (_________31478), .Q (______0__31254));
  nor2s1 _______448895(.DIN1 (________20384), .DIN2 (________21207), .Q
       (_____9__24181));
  nnd2s1 ____0__448896(.DIN1 (________20874), .DIN2 (________21141), .Q
       (___9____24323));
  hi1s1 ___0___448897(.DIN (_________33174), .Q (__9_____26456));
  nnd2s1 _______448898(.DIN1 (________21051), .DIN2 (________21050), .Q
       (___9____26174));
  nor2s1 _______448899(.DIN1 (________21049), .DIN2 (________20163), .Q
       (________24855));
  nor2s1 ____448900(.DIN1 (________21052), .DIN2 (________21048), .Q
       (____0___21992));
  nor2s1 _______448901(.DIN1 (____9___20316), .DIN2 (________21058), .Q
       (________26125));
  nor2s1 _______448902(.DIN1 (____0___21362), .DIN2 (________21047), .Q
       (___0____24412));
  nor2s1 _______448903(.DIN1 (_____0__21046), .DIN2 (________21058), .Q
       (___0____21697));
  nnd2s1 ____0__448904(.DIN1 (_____9__21045), .DIN2 (________21776), .Q
       (________26059));
  and2s1 _______448905(.DIN1 (________21281), .DIN2 (___09___20784), .Q
       (________21795));
  hi1s1 ______448906(.DIN (______0__35078), .Q (_________31295));
  nnd2s1 ____0__448907(.DIN1 (________21044), .DIN2 (________21043), .Q
       (_____0__23811));
  nnd2s1 _______448908(.DIN1 (________21204), .DIN2 (_____9__21287), .Q
       (__90_0__26271));
  or2s1 _______448909(.DIN1 (________20460), .DIN2 (________21054), .Q
       (__9_____26489));
  nnd2s1 ____0__448910(.DIN1 (________21042), .DIN2 (________21205), .Q
       (________25380));
  nor2s1 _____448911(.DIN1 (________20849), .DIN2 (____9___20976), .Q
       (________22425));
  nor2s1 ____9__448912(.DIN1 (________21174), .DIN2 (_____9__20206), .Q
       (_________32487));
  nnd2s1 ____99_448913(.DIN1 (____90__21066), .DIN2 (_____9__19936), .Q
       (__9_____26717));
  nnd2s1 _______448914(.DIN1 (___909__20613), .DIN2 (________21373), .Q
       (__9_____26555));
  nnd2s1 ____0__448915(.DIN1 (________20562), .DIN2 (___9_0__21561), .Q
       (________23770));
  nnd2s1 ____9__448916(.DIN1 (________20404), .DIN2 (_________35092),
       .Q (________23917));
  nnd2s1 _____0_448917(.DIN1 (________20399), .DIN2 (______18933), .Q
       (________23875));
  nor2s1 _______448918(.DIN1 (________21505), .DIN2 (____99__20604), .Q
       (__9_9___26695));
  nor2s1 _______448919(.DIN1 (________22037), .DIN2 (_____9__21009), .Q
       (________21040));
  nnd2s1 ____0_448920(.DIN1 (________20914), .DIN2 (____0___21905), .Q
       (________21037));
  nnd2s1 _______448921(.DIN1 (____9___20133), .DIN2 (________19514), .Q
       (________21036));
  nor2s1 _______448922(.DIN1 (____0___20984), .DIN2 (________20800), .Q
       (________21035));
  or2s1 _______448923(.DIN1 (________21032), .DIN2 (________21018), .Q
       (________21033));
  nor2s1 _______448924(.DIN1 (________19385), .DIN2 (________20949), .Q
       (________21031));
  nnd2s1 ______448925(.DIN1 (________21098), .DIN2 (____9___21808), .Q
       (_____0__21030));
  nor2s1 _______448926(.DIN1 (________21310), .DIN2 (___0____20734), .Q
       (_____9__21029));
  nnd2s1 _______448927(.DIN1 (________20957), .DIN2 (_____9__20293), .Q
       (________21028));
  nor2s1 _______448928(.DIN1 (________20090), .DIN2 (_____0__20332), .Q
       (________21027));
  nnd2s1 _______448929(.DIN1 (_____9__20391), .DIN2 (________21025), .Q
       (________21026));
  nnd2s1 _______448930(.DIN1 (___9____20648), .DIN2 (________21023), .Q
       (________21024));
  or2s1 _______448931(.DIN1 (________21021), .DIN2 (________20925), .Q
       (________21022));
  nor2s1 _______448932(.DIN1 (_____9__21019), .DIN2 (________21018), .Q
       (_____0__21020));
  and2s1 _______448933(.DIN1 (________21016), .DIN2 (___0____19786), .Q
       (________21017));
  nor2s1 _______448934(.DIN1 (________21276), .DIN2 (________21014), .Q
       (________21015));
  nnd2s1 _______448935(.DIN1 (____0___20988), .DIN2 (________21012), .Q
       (________21013));
  nnd2s1 _______448936(.DIN1 (________20240), .DIN2
       (_____________________18668), .Q (________21011));
  nor2s1 _____0_448937(.DIN1 (___0____21671), .DIN2 (_____9__21009), .Q
       (_____0__21010));
  nor2s1 _______448938(.DIN1 (____0___21263), .DIN2 (___9____20660), .Q
       (________21008));
  and2s1 _______448939(.DIN1 (___09___20785), .DIN2 (________21006), .Q
       (________21007));
  nnd2s1 _______448940(.DIN1 (________20346), .DIN2 (________21003), .Q
       (________21005));
  nor2s1 _______448941(.DIN1 (________21003), .DIN2 (____0___20139), .Q
       (________21004));
  nor2s1 _____0_448942(.DIN1 (________20534), .DIN2 (________20920), .Q
       (________21002));
  and2s1 _____448943(.DIN1 (________20803), .DIN2 (____9___20503), .Q
       (_____0__21001));
  and2s1 _______448944(.DIN1 (____0___20325), .DIN2 (___0____21698), .Q
       (_____9__21000));
  nor2s1 _____448945(.DIN1 (________20454), .DIN2 (________20998), .Q
       (________20999));
  nor2s1 _______448946(.DIN1 (________19522), .DIN2 (________20089), .Q
       (________20997));
  and2s1 _______448947(.DIN1 (________20848), .DIN2 (____9___21070), .Q
       (________20996));
  nor2s1 _______448948(.DIN1 (____0___20231), .DIN2 (________19974), .Q
       (________20995));
  nor2s1 _______448949(.DIN1 (________21014), .DIN2 (________20993), .Q
       (________20994));
  nnd2s1 _______448950(.DIN1 (________20446), .DIN2 (____0___21361), .Q
       (________20992));
  nnd2s1 ______448951(.DIN1 (________21378), .DIN2 (________19879), .Q
       (_____0__20991));
  nnd2s1 _______448952(.DIN1 (____0___21361), .DIN2 (________20393), .Q
       (____09__20990));
  nnd2s1 _______448953(.DIN1 (____0___20988), .DIN2 (________20109), .Q
       (____0___20989));
  and2s1 _____0_448954(.DIN1 (________20819), .DIN2 (____9___21441), .Q
       (____0___20987));
  nor2s1 ______448955(.DIN1 (_____0__19419), .DIN2 (___0____20750), .Q
       (____0___20986));
  nor2s1 _______448956(.DIN1 (____0___20984), .DIN2 (____0___21363), .Q
       (____0___20985));
  nor2s1 ______448957(.DIN1 (____9___19494), .DIN2 (_____0__20294), .Q
       (____00__20982));
  nor2s1 ______448958(.DIN1 (________21131), .DIN2 (___9____20650), .Q
       (____99__20981));
  nor2s1 ______448959(.DIN1 (____0___21265), .DIN2 (___0_0__21696), .Q
       (____9___20980));
  or2s1 _______448960(.DIN1 (____9___20978), .DIN2 (________20334), .Q
       (____9___20979));
  hi1s1 ____0__448961(.DIN (____9___20976), .Q (____9___20977));
  nor2s1 ______448962(.DIN1 (____0___21265), .DIN2 (________20852), .Q
       (____9___20975));
  or2s1 _______448963(.DIN1 (________20564), .DIN2 (________20152), .Q
       (____9___20974));
  nor2s1 _______448964(.DIN1 (____90__20972), .DIN2 (_____0__20372), .Q
       (____9___20973));
  or2s1 _____9_448965(.DIN1 (________20162), .DIN2 (________20970), .Q
       (_____9__20971));
  nor2s1 ____0__448966(.DIN1 (____9___21984), .DIN2 (_____0__20189), .Q
       (________20969));
  nnd2s1 ____0_448967(.DIN1 (________20842), .DIN2 (________20175), .Q
       (________20968));
  nor2s1 _______448968(.DIN1 (________19921), .DIN2 (_____9__20371), .Q
       (________20967));
  nor2s1 _____9_448969(.DIN1 (________20965), .DIN2 (_____0__20284), .Q
       (________20966));
  nnd2s1 _______448970(.DIN1 (________20844), .DIN2 (________20208), .Q
       (________20964));
  nor2s1 _______448971(.DIN1 (_____0__20962), .DIN2 (________20104), .Q
       (________20963));
  nor2s1 ______448972(.DIN1 (________20160), .DIN2 (________20339), .Q
       (_____9__20961));
  nnd2s1 _______448973(.DIN1 (________20851), .DIN2 (________22211), .Q
       (________20960));
  nnd2s1 _____9_448974(.DIN1 (_____0__20116), .DIN2 (inData[24]), .Q
       (________20959));
  and2s1 _______448975(.DIN1 (________20957), .DIN2 (___0____21690), .Q
       (________20958));
  nor2s1 _____0_448976(.DIN1 (___09___20782), .DIN2 (___00___20704), .Q
       (________20956));
  and2s1 ______448977(.DIN1 (________20954), .DIN2 (________20368), .Q
       (________20955));
  or2s1 _____0_448978(.DIN1 (________21750), .DIN2 (___0____21671), .Q
       (________20953));
  nor2s1 _______448979(.DIN1 (________21483), .DIN2 (____0___20887), .Q
       (_____0__20952));
  nor2s1 _____448980(.DIN1 (________20159), .DIN2 (________20478), .Q
       (_____9__20951));
  nor2s1 _______448981(.DIN1 (________19245), .DIN2 (________20949), .Q
       (________20950));
  nnd2s1 _______448982(.DIN1 (____90__20314), .DIN2 (____0___19856), .Q
       (________20948));
  nnd2s1 _______448983(.DIN1 (_____9__20912), .DIN2 (________20946), .Q
       (________20947));
  nnd2s1 _______448984(.DIN1 (_____0__20245), .DIN2 (________19565), .Q
       (________20945));
  nnd2s1 _______448985(.DIN1 (_____9__20096), .DIN2 (____0___21905), .Q
       (________20944));
  nor2s1 _______448986(.DIN1 (outData[9]), .DIN2 (_________33817), .Q
       (________20943));
  nnd2s1 _______448987(.DIN1 (________20360), .DIN2 (_____0__19562), .Q
       (_____0__20942));
  hi1s1 ____0__448988(.DIN (_____0__21210), .Q (________20940));
  and2s1 _______448989(.DIN1 (________20149), .DIN2
       (_____________________18624), .Q (________20939));
  nnd2s1 ____448990(.DIN1 (________20937), .DIN2 (________21511), .Q
       (________20938));
  nor2s1 ___0__448991(.DIN1 (________21978), .DIN2 (________20098), .Q
       (________20936));
  nnd2s1 ______448992(.DIN1 (___9____20667), .DIN2 (________20934), .Q
       (________20935));
  nnd2s1 ___0___448993(.DIN1 (________20157), .DIN2 (_____9__20932), .Q
       (_____0__20933));
  or2s1 _____0_448994(.DIN1 (________20930), .DIN2 (___9____20652), .Q
       (________20931));
  nnd2s1 ___0___448995(.DIN1 (____9___20318), .DIN2 (inData[10]), .Q
       (________20929));
  nor2s1 _______448996(.DIN1 (___9____21592), .DIN2 (________20853), .Q
       (________20928));
  and2s1 ______448997(.DIN1 (___0____20765), .DIN2 (________19905), .Q
       (________20927));
  nor2s1 _______448998(.DIN1 (_____9__21019), .DIN2 (________20925), .Q
       (________20926));
  or2s1 ___0__448999(.DIN1 (________19647), .DIN2 (_____0__20923), .Q
       (________20924));
  nor2s1 _______449000(.DIN1 (___9____19763), .DIN2 (________20344), .Q
       (_____9__20922));
  nor2s1 _____9_449001(.DIN1 (____09__20519), .DIN2 (________20920), .Q
       (________20921));
  and2s1 _______449002(.DIN1 (____0___21361), .DIN2 (___0____21684), .Q
       (________20919));
  nnd2s1 ______449003(.DIN1 (________20937), .DIN2 (________20917), .Q
       (________20918));
  hi1s1 ____0__449004(.DIN (________21194), .Q (________20916));
  nnd2s1 _______449005(.DIN1 (________20914), .DIN2 (_____9__19611), .Q
       (________20915));
  nnd2s1 _______449006(.DIN1 (_____9__20912), .DIN2 (_____0__21335), .Q
       (_____0__20913));
  nnd2s1 _______449007(.DIN1 (________20910), .DIN2 (________20521), .Q
       (________20911));
  or2s1 ___0_9_449008(.DIN1 (_________34439), .DIN2 (_________33186),
       .Q (________20909));
  nor2s1 _______449009(.DIN1 (___0____19792), .DIN2 (________20897), .Q
       (________20908));
  nnd2s1 ___0__449010(.DIN1 (___9____20685), .DIN2 (________20813), .Q
       (________20907));
  nor2s1 ___0___449011(.DIN1 (____00__20420), .DIN2 (____0___20232), .Q
       (________20906));
  nor2s1 ___0___449012(.DIN1 (________21862), .DIN2 (_____0__20847), .Q
       (________20905));
  nnd2s1 ______449013(.DIN1 (____9___21808), .DIN2 (________21497), .Q
       (_____0__20904));
  nnd2s1 ___09_449014(.DIN1 (________20281), .DIN2 (inData[28]), .Q
       (_____9__20903));
  nor2s1 _______449015(.DIN1 (________20901), .DIN2 (________20823), .Q
       (________20902));
  nor2s1 ______449016(.DIN1 (________20899), .DIN2 (_____9__20155), .Q
       (________20900));
  nor2s1 ____0__449017(.DIN1 (_____9__21979), .DIN2 (________20925), .Q
       (________20898));
  nor2s1 ____0__449018(.DIN1 (_____0__20895), .DIN2 (________20925), .Q
       (________20896));
  nor2s1 _____9_449019(.DIN1 (____0___20893), .DIN2 (________20174), .Q
       (____09__20894));
  nor2s1 _____0_449020(.DIN1 (________20183), .DIN2 (________19865), .Q
       (____0___20892));
  nnd2s1 _______449021(.DIN1 (____09__20145), .DIN2 (____0___19501), .Q
       (____0___20891));
  nor2s1 _______449022(.DIN1 (____0___20889), .DIN2 (____0___20888), .Q
       (____0___20890));
  nor2s1 _______449023(.DIN1 (___9____21618), .DIN2 (________20993), .Q
       (____00__20886));
  nnd2s1 _______449024(.DIN1 (________20814), .DIN2 (________22109), .Q
       (____99__20885));
  nor2s1 _______449025(.DIN1 (________20275), .DIN2 (____9___20883), .Q
       (____9___20884));
  nnd2s1 _______449026(.DIN1 (_____9__20912), .DIN2 (____9___20881), .Q
       (____9___20882));
  and2s1 _____0_449027(.DIN1 (________20299), .DIN2 (____9___21441), .Q
       (____9___20880));
  nor2s1 _______449028(.DIN1 (___099), .DIN2 (_________33817), .Q
       (____9___20879));
  nnd2s1 _______449029(.DIN1 (___0_9__21657), .DIN2 (____9___20877), .Q
       (____9___20878));
  nor2s1 ______449030(.DIN1 (________20930), .DIN2 (________20523), .Q
       (____90__20876));
  nnd2s1 _______449031(.DIN1 (________20874), .DIN2 (___9____20684), .Q
       (_____9__20875));
  nnd2s1 _______449032(.DIN1 (_____0__20857), .DIN2 (________20872), .Q
       (________20873));
  nnd2s1 _______449033(.DIN1 (________20279), .DIN2 (________21486), .Q
       (________20871));
  nnd2s1 _____9_449034(.DIN1 (________20835), .DIN2 (________20970), .Q
       (________20870));
  or2s1 _____9_449035(.DIN1 (________20868), .DIN2 (________20348), .Q
       (________20869));
  nnd2s1 _____449036(.DIN1 (________21510), .DIN2 (_____0__20866), .Q
       (________20867));
  or2s1 _______449037(.DIN1 (______________________18630), .DIN2
       (________20855), .Q (_____9__20865));
  nor2s1 _______449038(.DIN1 (_____0__19468), .DIN2 (________21372), .Q
       (________20864));
  nnd2s1 _______449039(.DIN1 (_____9__20361), .DIN2 (inData[0]), .Q
       (________20863));
  or2s1 _______449040(.DIN1 (_____9__20164), .DIN2 (________20008), .Q
       (________20862));
  hi1s1 ______449041(.DIN (________20860), .Q (________20861));
  nor2s1 _______449042(.DIN1 (____9___20222), .DIN2 (____9___20034), .Q
       (________20859));
  nnd2s1 ____9__449043(.DIN1 (________20858), .DIN2 (________20257), .Q
       (________21225));
  xor2s1 _______449044(.DIN1 (_______19000), .DIN2 (_________34023), .Q
       (____90___29908));
  and2s1 _______449045(.DIN1 (_____0__20857), .DIN2 (________20196), .Q
       (____9___21349));
  nnd2s1 _____9_449046(.DIN1 (_____9__20856), .DIN2 (________21211), .Q
       (____9___21809));
  or2s1 _____9_449047(.DIN1 (______________________18629), .DIN2
       (________20855), .Q (________21855));
  nor2s1 ____449048(.DIN1 (________20854), .DIN2 (________20853), .Q
       (________21382));
  nor2s1 _______449049(.DIN1 (________21750), .DIN2 (________20852), .Q
       (________21063));
  nnd2s1 _____9_449050(.DIN1 (________20379), .DIN2 (________20833), .Q
       (____9___21350));
  nnd2s1 ____9__449051(.DIN1 (________20834), .DIN2 (________21794), .Q
       (________21500));
  hi1s1 ____0__449052(.DIN (________21062), .Q (________21463));
  nnd2s1 ____9__449053(.DIN1 (________20851), .DIN2 (________22109), .Q
       (_____9__21474));
  nor2s1 ______449054(.DIN1 (________20850), .DIN2 (________20849), .Q
       (________21150));
  nor2s1 _____449055(.DIN1 (________20153), .DIN2 (________21060), .Q
       (________22342));
  and2s1 _____9_449056(.DIN1 (________20848), .DIN2 (________21397), .Q
       (_____9__21756));
  nor2s1 ___09__449057(.DIN1 (________20398), .DIN2 (_____0__20847), .Q
       (________21490));
  nor2s1 ___099_449058(.DIN1 (_____9__20846), .DIN2 (_____0__20847), .Q
       (________21342));
  nor2s1 ____0__449059(.DIN1 (_____0__21230), .DIN2 (________20450), .Q
       (________21124));
  nnd2s1 ____0__449060(.DIN1 (_____0__20857), .DIN2 (________20970), .Q
       (________21473));
  nnd2s1 ____9__449061(.DIN1 (___0____20719), .DIN2 (________21375), .Q
       (________21482));
  nnd2s1 ____9__449062(.DIN1 (_____0__20181), .DIN2 (inData[24]), .Q
       (____9___21068));
  nor2s1 ____9__449063(.DIN1 (________20849), .DIN2 (________20845), .Q
       (________21498));
  nnd2s1 ____9_449064(.DIN1 (________20269), .DIN2 (________19509), .Q
       (________22183));
  nor2s1 ____90_449065(.DIN1 (___0____20746), .DIN2 (________20853), .Q
       (________21100));
  nnd2s1 ____9_449066(.DIN1 (________20954), .DIN2 (___90___21549), .Q
       (_____9__21493));
  nnd2s1 ____9_449067(.DIN1 (________20844), .DIN2 (________20843), .Q
       (________21235));
  nnd2s1 ____9__449068(.DIN1 (________20842), .DIN2 (___0_9__20779), .Q
       (____09__21364));
  nnd2s1 ____9__449069(.DIN1 (________20858), .DIN2 (________20202), .Q
       (___9____21583));
  nnd2s1 ______449070(.DIN1 (___0____20716), .DIN2 (________21023), .Q
       (________21118));
  nor2s1 _______449071(.DIN1 (____0___20043), .DIN2 (________21060), .Q
       (________21148));
  hi1s1 ____0__449072(.DIN (________20841), .Q (____99__21903));
  or2s1 ____9__449073(.DIN1 (_____________________18668), .DIN2
       (________20114), .Q (____9___21537));
  nnd2s1 _____9_449074(.DIN1 (________20848), .DIN2 (________20290), .Q
       (___09___23522));
  nor2s1 _______449075(.DIN1 (_____0__21429), .DIN2 (___9____20646), .Q
       (____0___21447));
  nnd2s1 ____9__449076(.DIN1 (________20957), .DIN2 (____0___21991), .Q
       (____9___21535));
  nor2s1 _______449077(.DIN1 (____0____________0_), .DIN2
       (________20849), .Q (_____0__21485));
  nnd2s1 ____9__449078(.DIN1 (________20858), .DIN2 (________20839), .Q
       (_____0__22690));
  hi1s1 ______449079(.DIN (_________30472), .Q (____90___28993));
  hi1s1 ______449080(.DIN (___0____22597), .Q (__99____27157));
  hi1s1 ____0_449081(.DIN (________20840), .Q (________22139));
  nnd2s1 ____9__449082(.DIN1 (________20364), .DIN2 (________20839), .Q
       (____0___21911));
  nnd2s1 _____0_449083(.DIN1 (________20838), .DIN2 (_____9__20826), .Q
       (____0___21358));
  nor2s1 ____9__449084(.DIN1 (_____0__19282), .DIN2 (____9___20315), .Q
       (___9____21566));
  nnd2s1 ____9__449085(.DIN1 (_____0__20837), .DIN2 (________22131), .Q
       (________21507));
  nor2s1 ____9__449086(.DIN1 (___0____21651), .DIN2 (_____9__20836), .Q
       (________21491));
  nnd2s1 ____9__449087(.DIN1 (________20835), .DIN2 (________21481), .Q
       (________21338));
  nnd2s1 _______449088(.DIN1 (________20937), .DIN2 (____9___20128), .Q
       (________25052));
  and2s1 _______449089(.DIN1 (____0___20794), .DIN2 (________21337), .Q
       (_____9__21400));
  nor2s1 ____9__449090(.DIN1 (________20920), .DIN2 (___9____20628), .Q
       (________24909));
  hi1s1 _______449091(.DIN (_____00__33954), .Q (_________33797));
  hi1s1 _______449092(.DIN (____9___21158), .Q (___9_0__21580));
  nnd2s1 ____9__449093(.DIN1 (________20834), .DIN2 (________20833), .Q
       (_____0__21494));
  nnd2s1 ____0__449094(.DIN1 (_____9__20856), .DIN2 (________21397), .Q
       (________22783));
  hi1s1 _______449095(.DIN (______9__33247), .Q (_________33268));
  nor2s1 ____9__449096(.DIN1 (____9___20506), .DIN2 (____9___20502), .Q
       (________25639));
  nor2s1 ____9__449097(.DIN1 (________20262), .DIN2 (___9____20649), .Q
       (________23104));
  nnd2s1 _____9_449098(.DIN1 (_____9__20856), .DIN2 (________21053), .Q
       (________25115));
  nnd2s1 ____9__449099(.DIN1 (________20937), .DIN2 (________20308), .Q
       (________25817));
  nor2s1 ____9_449100(.DIN1 (________20113), .DIN2 (________20832), .Q
       (___0____22589));
  nnd2s1 _______449101(.DIN1 (________20957), .DIN2 (___0_0__19810), .Q
       (________21512));
  nnd2s1 _______449102(.DIN1 (____0___20326), .DIN2 (________20831), .Q
       (_________30341));
  nor2s1 _____9_449103(.DIN1 (________20830), .DIN2 (___9____20677), .Q
       (________25901));
  nnd2s1 _____9_449104(.DIN1 (________20291), .DIN2 (____9___19200), .Q
       (___900__26147));
  hi1s1 ______449105(.DIN (___000___27171), .Q (_____90__31526));
  nnd2s1 ____9__449106(.DIN1 (________20835), .DIN2 (________20828), .Q
       (________26018));
  nnd2s1 ____9__449107(.DIN1 (____0___19857), .DIN2 (_________35090),
       .Q (___9____26159));
  nor2s1 _______449108(.DIN1 (_____9__20499), .DIN2 (________20187), .Q
       (_________31478));
  nor2s1 _______449109(.DIN1 (________21387), .DIN2 (________20266), .Q
       (_________31326));
  nor2s1 _______449110(.DIN1 (_____0__21335), .DIN2 (________20310), .Q
       (______0__30607));
  nor2s1 ______449111(.DIN1 (________20467), .DIN2 (________20112), .Q
       (_________32554));
  nnd2s1 _______449112(.DIN1 (________20874), .DIN2 (________20566), .Q
       (__9_____26496));
  nnd2s1 ____99_449113(.DIN1 (_____0__20827), .DIN2 (_____9__20826), .Q
       (__9_____26937));
  nnd2s1 ______449114(.DIN1 (________20253), .DIN2 (________20825), .Q
       (_________33144));
  nnd2s1 _______449115(.DIN1 (________20184), .DIN2 (________21472), .Q
       (____099__30093));
  nor2s1 _______449116(.DIN1 (________21470), .DIN2 (_____9__20188), .Q
       (_________29500));
  nnd2s1 ______449117(.DIN1 (________20270), .DIN2 (_____9__20932), .Q
       (____99__25750));
  nor2s1 _______449118(.DIN1 (____9___20599), .DIN2 (________20267), .Q
       (______0__29851));
  nnd2s1 ______449119(.DIN1 (____9___20129), .DIN2 (________21487), .Q
       (____9____32728));
  nor2s1 ______449120(.DIN1 (____0___20514), .DIN2 (________20185), .Q
       (_________33564));
  nor2s1 ______449121(.DIN1 (________19544), .DIN2 (________20265), .Q
       (_________31134));
  nnd2s1 _______449122(.DIN1 (________20357), .DIN2 (___0____19815), .Q
       (______9__33856));
  nor2s1 _____449123(.DIN1 (________21889), .DIN2 (________20823), .Q
       (________20824));
  nor2s1 _______449124(.DIN1 (________20821), .DIN2 (________20444), .Q
       (________20822));
  and2s1 _______449125(.DIN1 (________20819), .DIN2 (_____9__20816), .Q
       (________20820));
  and2s1 _______449126(.DIN1 (____9___20134), .DIN2
       (_____________________18637), .Q (________20818));
  nnd2s1 ___0_449127(.DIN1 (________20305), .DIN2 (_____9__20816), .Q
       (_____0__20817));
  and2s1 _____9_449128(.DIN1 (________20814), .DIN2 (________20813), .Q
       (________20815));
  hi1s1 ____0__449129(.DIN (________21207), .Q (________20812));
  nnd2s1 _______449130(.DIN1 (____90__21156), .DIN2 (____0___20423), .Q
       (________20811));
  nnd2s1 ____0__449131(.DIN1 (___0____20767), .DIN2 (________20809), .Q
       (________20810));
  nor2s1 ____0__449132(.DIN1 (____9___19588), .DIN2 (_____9__20836), .Q
       (________20808));
  nnd2s1 ____0_449133(.DIN1 (___9_9__20653), .DIN2 (________21397), .Q
       (_____0__20807));
  nor2s1 ____09_449134(.DIN1 (____9___21980), .DIN2 (________20998), .Q
       (_____9__20806));
  nnd2s1 _______449135(.DIN1 (________21530), .DIN2 (_____9__20263), .Q
       (________20805));
  nnd2s1 _______449136(.DIN1 (________20803), .DIN2 (________20802), .Q
       (________20804));
  or2s1 _______449137(.DIN1 (________20800), .DIN2 (________20469), .Q
       (________20801));
  nor2s1 _______449138(.DIN1 (________20343), .DIN2 (________20170), .Q
       (_____0__20799));
  nor2s1 _______449139(.DIN1 (____9___21900), .DIN2 (___0____20758), .Q
       (____09__20798));
  nnd2s1 _______449140(.DIN1 (________20851), .DIN2 (________21486), .Q
       (____0___20797));
  nor2s1 _______449141(.DIN1 (________21114), .DIN2 (___0_0__20752), .Q
       (____0___20796));
  nnd2s1 _______449142(.DIN1 (____0___20794), .DIN2 (________20946), .Q
       (____0___20795));
  nor2s1 _______449143(.DIN1 (________21471), .DIN2 (____0___20329), .Q
       (____0___20793));
  and2s1 _______449144(.DIN1 (________20544), .DIN2 (____0___20791), .Q
       (____0___20792));
  nnd2s1 _______449145(.DIN1 (________20385), .DIN2 (____0___20791), .Q
       (____00__20790));
  nor2s1 _______449146(.DIN1 (____0___19115), .DIN2 (_________33817),
       .Q (___099__20789));
  and2s1 _______449147(.DIN1 (___0____20731), .DIN2 (____09__20331), .Q
       (___09___20788));
  nnd2s1 _______449148(.DIN1 (___9____20659), .DIN2 (________21203), .Q
       (___09___20787));
  and2s1 ______449149(.DIN1 (___09___20785), .DIN2 (___09___20784), .Q
       (___09___20786));
  nor2s1 _______449150(.DIN1 (___09___20782), .DIN2 (________20171), .Q
       (___09___20783));
  nor2s1 _____449151(.DIN1 (________21319), .DIN2 (________21153), .Q
       (___09___20781));
  and2s1 _____9_449152(.DIN1 (____0___20794), .DIN2 (___0_9__20779), .Q
       (___090__20780));
  or2s1 _____9_449153(.DIN1 (________21407), .DIN2 (____0___20144), .Q
       (___0____20778));
  nnd2s1 _______449154(.DIN1 (________20914), .DIN2 (________20493), .Q
       (___0____20777));
  and2s1 _______449155(.DIN1 (____0___20141), .DIN2 (___0____21698), .Q
       (___0____20776));
  nnd2s1 _______449156(.DIN1 (________20014), .DIN2 (________20259), .Q
       (___0____20775));
  nnd2s1 _______449157(.DIN1 (___0____20773), .DIN2 (________19924), .Q
       (___0____20774));
  nnd2s1 _______449158(.DIN1 (____9___21808), .DIN2 (___0_0__20771), .Q
       (___0____20772));
  and2s1 _______449159(.DIN1 (________20848), .DIN2 (________21211), .Q
       (___0_9__20770));
  and2s1 _______449160(.DIN1 (________20957), .DIN2 (_____9__21278), .Q
       (___0____20769));
  nnd2s1 _______449161(.DIN1 (___0____20767), .DIN2 (________21774), .Q
       (___0____20768));
  and2s1 _______449162(.DIN1 (___0____20765), .DIN2 (_____9__21278), .Q
       (___0____20766));
  nnd2s1 _______449163(.DIN1 (________20340), .DIN2 (___0____20763), .Q
       (___0____20764));
  nnd2s1 ______449164(.DIN1 (___0_9__20761), .DIN2 (________19886), .Q
       (___0_0__20762));
  nor2s1 _______449165(.DIN1 (________20248), .DIN2 (________20239), .Q
       (___0____20760));
  nor2s1 _______449166(.DIN1 (________21862), .DIN2 (___0____20758), .Q
       (___0____20759));
  and2s1 _______449167(.DIN1 (___0____20767), .DIN2 (___0____20756), .Q
       (___0____20757));
  nor2s1 _______449168(.DIN1 (________22113), .DIN2 (_____0__20146), .Q
       (___0____20755));
  or2s1 ______449169(.DIN1 (___0____20753), .DIN2 (___0_0__20752), .Q
       (___0____20754));
  nnd2s1 _______449170(.DIN1 (___0____20750), .DIN2 (________20525), .Q
       (___0_9__20751));
  and2s1 _______449171(.DIN1 (____0___20988), .DIN2 (___0____20748), .Q
       (___0____20749));
  nor2s1 _______449172(.DIN1 (___0____20746), .DIN2 (____9___20127), .Q
       (___0____20747));
  nnd2s1 _______449173(.DIN1 (____9___20220), .DIN2 (inData[16]), .Q
       (___0____20745));
  nor2s1 ___09__449174(.DIN1 (___0_0__20743), .DIN2 (_________33186),
       .Q (___0____20744));
  nnd2s1 ______449175(.DIN1 (________20147), .DIN2 (____9____31759), .Q
       (___0_9__20742));
  nnd2s1 _____0_449176(.DIN1 (___9____20658), .DIN2 (___90___20606), .Q
       (___0____20741));
  hi1s1 _______449177(.DIN (_____9__21182), .Q (___0____20740));
  or2s1 _______449178(.DIN1 (____0___21263), .DIN2 (___0_0__20752), .Q
       (___0____20739));
  hi1s1 ____0_449179(.DIN (___0____20737), .Q (___0____20738));
  hi1s1 _____9_449180(.DIN (________21145), .Q (___0____20736));
  nor2s1 _______449181(.DIN1 (___0____20734), .DIN2 (________20993), .Q
       (___0____20735));
  hi1s1 _____0_449182(.DIN (________21204), .Q (___0_0__20733));
  nnd2s1 _____0_449183(.DIN1 (___0____20731), .DIN2 (___0____20730), .Q
       (___0_9__20732));
  nnd2s1 ______449184(.DIN1 (________21012), .DIN2 (____90__20410), .Q
       (___0____20729));
  or2s1 ______449185(.DIN1 (______________________18629), .DIN2
       (___0____20727), .Q (___0____20728));
  nor2s1 _______449186(.DIN1 (________19355), .DIN2 (_________31047),
       .Q (___0____20726));
  and2s1 ______449187(.DIN1 (________20238), .DIN2 (________21372), .Q
       (___0____20725));
  nnd2s1 _______449188(.DIN1 (________22187), .DIN2 (________19995), .Q
       (___0_0__20724));
  nor2s1 _______449189(.DIN1 (___0____20722), .DIN2 (________20255), .Q
       (___0_9__20723));
  nnd2s1 _______449190(.DIN1 (________20287), .DIN2 (________22050), .Q
       (___0____20721));
  nnd2s1 ______449191(.DIN1 (___0____20719), .DIN2 (____0___21905), .Q
       (___0____20720));
  nnd2s1 ___09__449192(.DIN1 (________20119), .DIN2 (________20151), .Q
       (___0____20718));
  nnd2s1 ______449193(.DIN1 (___0____20716), .DIN2 (___9_0__19698), .Q
       (___0____20717));
  nor2s1 _______449194(.DIN1 (_______19013), .DIN2 (_________33186), .Q
       (___0____20714));
  nnd2s1 ___0__449195(.DIN1 (________20298), .DIN2 (inData[2]), .Q
       (___0____20713));
  or2s1 _______449196(.DIN1 (________20872), .DIN2 (________20282), .Q
       (___0____20712));
  nor2s1 ____0__449197(.DIN1 (________22017), .DIN2 (________20276), .Q
       (___0____20711));
  nor2s1 _______449198(.DIN1 (___0____19784), .DIN2 (_____0__20342), .Q
       (___0____20709));
  and2s1 _____0_449199(.DIN1 (________20957), .DIN2 (________22131), .Q
       (___0_0__20708));
  nnd2s1 _______449200(.DIN1 (________20186), .DIN2 (____9___20132), .Q
       (___009__20707));
  nor2s1 _____0_449201(.DIN1 (___00___20705), .DIN2 (___00___20704), .Q
       (___00___20706));
  hi1s1 _______449202(.DIN (___00___20701), .Q (___00___20702));
  xor2s1 _______449203(.DIN1 (______0__18865), .DIN2 (______9__32232),
       .Q (___00___20700));
  nnd2s1 _______449204(.DIN1 (________20358), .DIN2 (_____0__19956), .Q
       (___000__20699));
  nnd2s1 _____0_449205(.DIN1 (____9___21803), .DIN2 (________20124), .Q
       (___999__20698));
  nnd2s1 ___09__449206(.DIN1 (________20095), .DIN2 (inData[2]), .Q
       (___99___20697));
  nnd2s1 _______449207(.DIN1 (_____0__20857), .DIN2 (___99___20695), .Q
       (___99___20696));
  nor2s1 _____9_449208(.DIN1 (________20082), .DIN2 (____0___20230), .Q
       (___99___20694));
  nnd2s1 _______449209(.DIN1 (_____0__20857), .DIN2 (___09___20784), .Q
       (___99___20693));
  nor2s1 ___09_449210(.DIN1 (___99___20691), .DIN2 (_____0__20923), .Q
       (___99___20692));
  nor2s1 _______449211(.DIN1 (___0____21692), .DIN2 (________20998), .Q
       (___9____20690));
  nnd2s1 _______449212(.DIN1 (________20105), .DIN2 (_____0__21504), .Q
       (___9____20689));
  nor2s1 _______449213(.DIN1 (____0___21167), .DIN2 (________20998), .Q
       (___9____20688));
  nnd2s1 _____9_449214(.DIN1 (____0___20227), .DIN2 (_____0__20069), .Q
       (___9____20687));
  nnd2s1 ___0__449215(.DIN1 (___9____20685), .DIN2 (___9____20684), .Q
       (___9____20686));
  nor2s1 ______449216(.DIN1 (________19657), .DIN2 (_________31047), .Q
       (___9____20683));
  nor2s1 _______449217(.DIN1 (___9_9__20681), .DIN2 (___0_0__21696), .Q
       (___9_0__20682));
  xor2s1 _______449218(.DIN1 (outData[27]), .DIN2 (_________31154), .Q
       (___9____20680));
  nnd2s1 ____0__449219(.DIN1 (________20842), .DIN2 (________20946), .Q
       (___9____20679));
  nor2s1 ______449220(.DIN1 (________20297), .DIN2 (___9____20677), .Q
       (___9____20678));
  and2s1 _____9_449221(.DIN1 (________20111), .DIN2 (________22109), .Q
       (___9____20676));
  or2s1 _______449222(.DIN1 (________19970), .DIN2 (_____9__20351), .Q
       (___9____20675));
  nor2s1 _____449223(.DIN1 (________19466), .DIN2 (________20236), .Q
       (___9____20674));
  nnd2s1 _____0_449224(.DIN1 (________20301), .DIN2 (_____9__20816), .Q
       (___9____20673));
  nnd2s1 ___09__449225(.DIN1 (____9___20320), .DIN2 (________20053), .Q
       (___9_0__20672));
  nor2s1 _______449226(.DIN1 (________20868), .DIN2 (________20302), .Q
       (___9_9__20671));
  or2s1 _______449227(.DIN1 (____0________________18589), .DIN2
       (_____9__20115), .Q (___9____20670));
  nnd2s1 _______449228(.DIN1 (________20848), .DIN2 (________21203), .Q
       (___9____20669));
  and2s1 _______449229(.DIN1 (________20937), .DIN2 (________20148), .Q
       (____9___21352));
  nnd2s1 _____9_449230(.DIN1 (_____9__20856), .DIN2 (____9___21070), .Q
       (____0___21819));
  nnd2s1 _____9_449231(.DIN1 (________20260), .DIN2 (_____0__21885), .Q
       (________21425));
  nnd2s1 _____0_449232(.DIN1 (___9____20668), .DIN2 (_____9__20826), .Q
       (_____9__21209));
  nnd2s1 ____9__449233(.DIN1 (___9____20667), .DIN2 (____0___21267), .Q
       (________21341));
  nor2s1 ____9__449234(.DIN1 (_____9__20491), .DIN2 (________20365), .Q
       (____99__21542));
  nnd2s1 ____9__449235(.DIN1 (_____0__19892), .DIN2 (________20367), .Q
       (________21379));
  nor2s1 ____0_449236(.DIN1 (_____9__20244), .DIN2 (________21481), .Q
       (________21041));
  nor2s1 _______449237(.DIN1 (___9____20666), .DIN2 (___9____20655), .Q
       (________21061));
  and2s1 _______449238(.DIN1 (___9____20661), .DIN2 (_________35092),
       .Q (________21793));
  nnd2s1 _____9_449239(.DIN1 (________20848), .DIN2 (___00___20703), .Q
       (________21214));
  nnd2s1 _______449240(.DIN1 (________20848), .DIN2 (_____9__21287), .Q
       (________22378));
  nor2s1 _____9_449241(.DIN1 (___9____20665), .DIN2 (________20182), .Q
       (________21094));
  nnd2s1 _______449242(.DIN1 (_____9__20856), .DIN2 (________21203), .Q
       (____09__21994));
  nnd2s1 ____9__449243(.DIN1 (___9____20664), .DIN2 (________20839), .Q
       (_____0__21220));
  nnd2s1 _______449244(.DIN1 (________21378), .DIN2 (____9___21897), .Q
       (________21389));
  hi1s1 _____9_449245(.DIN (___9_0__20663), .Q (____0___21359));
  nor2s1 _______449246(.DIN1 (_____0__20088), .DIN2 (___9____21618), .Q
       (____99__21354));
  or2s1 _______449247(.DIN1 (___9_9__20662), .DIN2 (________21060), .Q
       (____9___21347));
  and2s1 ______449248(.DIN1 (___9____20661), .DIN2 (_________35090), .Q
       (___0____21668));
  nor2s1 _____449249(.DIN1 (___0____20753), .DIN2 (___9____20660), .Q
       (________21340));
  nnd2s1 _____449250(.DIN1 (___9____20659), .DIN2 (________21397), .Q
       (________21377));
  nor2s1 _____9_449251(.DIN1 (________20060), .DIN2 (_____9__20836), .Q
       (_____0__21384));
  and2s1 _____9_449252(.DIN1 (___9____20658), .DIN2 (_____0__21504), .Q
       (________21343));
  nnd2s1 _______449253(.DIN1 (_____9__20912), .DIN2 (___0_9__20779), .Q
       (____0___21170));
  nnd2s1 _______449254(.DIN1 (________22674), .DIN2 (________19512), .Q
       (________22056));
  dffacs1 __________________449255(.CLRB (reset), .CLK (clk), .DIN
       (____0___20140), .QN (_________34497));
  nor2s1 ____0__449256(.DIN1 (____0___20425), .DIN2 (___9____20632), .Q
       (____9___22347));
  nnd2s1 ____9__449257(.DIN1 (________20897), .DIN2 (_________31587),
       .Q (____0____31816));
  or2s1 ______449258(.DIN1 (___0____21680), .DIN2 (_________33186), .Q
       (_____0___31454));
  nor2s1 ____9_449259(.DIN1 (______18933), .DIN2 (_____9__21522), .Q
       (________21519));
  hi1s1 ____0__449260(.DIN (________21195), .Q (________21456));
  nnd2s1 _______449261(.DIN1 (________20957), .DIN2 (___9____20657), .Q
       (_____9__21383));
  nnd2s1 ______449262(.DIN1 (____9___20130), .DIN2 (_____0__20520), .Q
       (____0___21813));
  nor2s1 _______449263(.DIN1 (___9____20656), .DIN2 (___9____20655), .Q
       (___0____24408));
  nnd2s1 _______449264(.DIN1 (________20354), .DIN2 (____9___19587), .Q
       (________21406));
  nnd2s1 ______449265(.DIN1 (___9_0__20654), .DIN2 (_____9__20912), .Q
       (________21949));
  and2s1 _______449266(.DIN1 (___9____20659), .DIN2 (________21211), .Q
       (___9_0__22472));
  and2s1 _______449267(.DIN1 (___9_9__20653), .DIN2 (________21211), .Q
       (________23729));
  nor2s1 _______449268(.DIN1 (___0____20763), .DIN2 (___9____20652), .Q
       (_____9__21334));
  nnd2s1 _______449269(.DIN1 (________20306), .DIN2 (_________35090),
       .Q (________22029));
  nnd2s1 ____9__449270(.DIN1 (________20834), .DIN2 (________20569), .Q
       (________21478));
  nnd2s1 _______449271(.DIN1 (___0____20716), .DIN2 (___99_), .Q
       (________21376));
  hi1s1 ____0_449272(.DIN (_________31153), .Q (_________29280));
  nnd2s1 ____9_449273(.DIN1 (___0____20765), .DIN2 (________20201), .Q
       (_____9__21503));
  nnd2s1 ____9__449274(.DIN1 (___0____20716), .DIN2 (____9___19943), .Q
       (________22275));
  hi1s1 ____0__449275(.DIN (________21212), .Q (________21367));
  nor2s1 _______449276(.DIN1 (___9____20651), .DIN2 (________21144), .Q
       (________21332));
  nor2s1 ____0__449277(.DIN1 (____9___21980), .DIN2 (_____0__20847), .Q
       (_____9__21484));
  nor2s1 ____99_449278(.DIN1 (________21476), .DIN2 (___9____20650), .Q
       (____0___21356));
  nor2s1 ____9__449279(.DIN1 (____9___20508), .DIN2 (___9____20649), .Q
       (________22001));
  and2s1 _______449280(.DIN1 (_____9__20826), .DIN2 (_____9__20197), .Q
       (________23284));
  and2s1 _______449281(.DIN1 (___9_9__20653), .DIN2 (____9___21070), .Q
       (________25782));
  nnd2s1 _____449282(.DIN1 (___9____20648), .DIN2 (___9_0__20644), .Q
       (________21370));
  nor2s1 _______449283(.DIN1 (___9____20647), .DIN2 (___9____20649), .Q
       (________26000));
  nor2s1 _______449284(.DIN1 (___9____20647), .DIN2 (________21054), .Q
       (___0____25354));
  nnd2s1 ______449285(.DIN1 (________20570), .DIN2 (____0___20138), .Q
       (________26068));
  nnd2s1 _____0_449286(.DIN1 (___0____20765), .DIN2 (________21375), .Q
       (________21371));
  or2s1 ____9__449287(.DIN1 (____0___20512), .DIN2 (________21048), .Q
       (________23321));
  and2s1 _______449288(.DIN1 (___0____20731), .DIN2 (____9___20037), .Q
       (________21733));
  nnd2s1 _______449289(.DIN1 (___9____20659), .DIN2 (____9___21070), .Q
       (___00____27222));
  nor2s1 ____9__449290(.DIN1 (____0____________0_), .DIN2
       (_____9__21522), .Q (________21525));
  nor2s1 _______449291(.DIN1 (___0____21659), .DIN2 (___9____20646), .Q
       (____9___25458));
  hi1s1 ______449292(.DIN (________21974), .Q (___9_9__21589));
  nor2s1 _______449293(.DIN1 (____9____30882), .DIN2 (____9___20321),
       .Q (________25015));
  nnd2s1 ____9_449294(.DIN1 (___9____20645), .DIN2 (________20839), .Q
       (____0___25470));
  nnd2s1 ____9_449295(.DIN1 (____99__20135), .DIN2 (____9___19200), .Q
       (____0___23620));
  nnd2s1 _____449296(.DIN1 (___9____20661), .DIN2 (________20442), .Q
       (________25973));
  nnd2s1 ____9_449297(.DIN1 (_____0__20827), .DIN2 (___09___20785), .Q
       (________25726));
  nnd2s1 _____0_449298(.DIN1 (___9_9__20653), .DIN2 (________21203), .Q
       (________25864));
  or2s1 _____0_449299(.DIN1 (____0____________0_), .DIN2
       (________20800), .Q (___9____21620));
  nnd2s1 ____9__449300(.DIN1 (________20356), .DIN2 (_________35092),
       .Q (___9____23416));
  nnd2s1 _______449301(.DIN1 (___09___20785), .DIN2 (___9____20668), .Q
       (____9___22886));
  nnd2s1 ____9__449302(.DIN1 (________20937), .DIN2 (___9_0__20644), .Q
       (________21402));
  or2s1 _____9_449303(.DIN1 (___9____20655), .DIN2 (________20829), .Q
       (_____0__25790));
  nnd2s1 ____9__449304(.DIN1 (____9___20603), .DIN2 (________20118), .Q
       (________26099));
  hi1s1 ______449305(.DIN (__9_00__26989), .Q (_________33204));
  nnd2s1 _____9_449306(.DIN1 (___9_9__20653), .DIN2 (_____9__21287), .Q
       (__9_____26370));
  nnd2s1 _____9_449307(.DIN1 (________20848), .DIN2 (________21053), .Q
       (_________28837));
  nnd2s1 _____0_449308(.DIN1 (________20838), .DIN2 (___09___20785), .Q
       (__9_____26639));
  or2s1 _______449309(.DIN1 (___0_0__21658), .DIN2 (________20165), .Q
       (_________33007));
  nor2s1 _______449310(.DIN1 (________21470), .DIN2 (________20167), .Q
       (____0_0__31861));
  nnd2s1 ____0__449311(.DIN1 (___9_9__20643), .DIN2 (________20373), .Q
       (____90___33582));
  hi1s1 _______449312(.DIN (________21339), .Q (________21477));
  nnd2s1 ____99_449313(.DIN1 (___9____20661), .DIN2 (________20844), .Q
       (__900_));
  hi1s1 _______449314(.DIN (_________28365), .Q (____0_0__31851));
  hi1s1 ____0_449315(.DIN (_________32639), .Q (_________31648));
  nnd2s1 ____0__449316(.DIN1 (____99__20225), .DIN2 (________20825), .Q
       (____9____30874));
  hi1s1 _______449317(.DIN (________24923), .Q (_________33278));
  hi1s1 _______449318(.DIN (___9____20642), .Q (___9____21614));
  nor2s1 ____0_449319(.DIN1 (________20178), .DIN2 (________20965), .Q
       (_________30496));
  nnd2s1 _______449320(.DIN1 (_____9___30173), .DIN2 (_________29858),
       .Q (____0____30080));
  hi1s1 _______449321(.DIN (___9____20641), .Q (___0____21663));
  nor2s1 _______449322(.DIN1 (________19461), .DIN2 (________20179), .Q
       (_________33174));
  xor2s1 ____09_449323(.DIN1 (_____9__19085), .DIN2 (_________29330),
       .Q (___9____20640));
  nnd2s1 _______449324(.DIN1 (________20029), .DIN2 (___9____20638), .Q
       (___9____20639));
  or2s1 _______449325(.DIN1 (___0____21692), .DIN2 (________20522), .Q
       (___9____20637));
  nnd2s1 _______449326(.DIN1 (___9____20635), .DIN2 (___9_0__20634), .Q
       (___9____20636));
  or2s1 _______449327(.DIN1 (______9__33899), .DIN2 (___9____20632), .Q
       (___9_9__20633));
  nnd2s1 _____0_449328(.DIN1 (________21385), .DIN2 (________22339), .Q
       (___9____20631));
  and2s1 _____0_449329(.DIN1 (_____9__20548), .DIN2 (___0____21684), .Q
       (___9____20630));
  nor2s1 _____0_449330(.DIN1 (________20247), .DIN2 (___9____20628), .Q
       (___9____20629));
  nor2s1 ______449331(.DIN1 (____0___19860), .DIN2 (________19880), .Q
       (___9____20627));
  nor2s1 ______449332(.DIN1 (___9____20625), .DIN2 (_____0__20895), .Q
       (___9____20626));
  nor2s1 _______449333(.DIN1 (___9_9__20623), .DIN2 (________19914), .Q
       (___9_0__20624));
  and2s1 _______449334(.DIN1 (________22227), .DIN2
       (____0________________18651), .Q (___9____20622));
  nor2s1 _______449335(.DIN1 (____0___19595), .DIN2 (________19895), .Q
       (___9____20621));
  nor2s1 _______449336(.DIN1 (________19933), .DIN2 (________19903), .Q
       (___9____20620));
  nor2s1 _______449337(.DIN1
       (____________________________________18836), .DIN2
       (______9__33899), .Q (___9____20619));
  nor2s1 ______449338(.DIN1 (________20123), .DIN2 (___9____20617), .Q
       (___9____20618));
  nor2s1 ______449339(.DIN1 (___9____20656), .DIN2 (___9____20615), .Q
       (___9____20616));
  nnd2s1 ____00_449340(.DIN1 (________19931), .DIN2 (________20901), .Q
       (___9_0__20614));
  and2s1 _______449341(.DIN1 (________19885), .DIN2 (_____0__22118), .Q
       (___909__20613));
  nnd2s1 _______449342(.DIN1 (___09___19849), .DIN2 (_____0__20392), .Q
       (___90___20612));
  nor2s1 _______449343(.DIN1 (________20007), .DIN2 (________20022), .Q
       (___90___20611));
  nnd2s1 _______449344(.DIN1 (____0___20517), .DIN2 (___900__20605), .Q
       (___90___20610));
  nor2s1 ______449345(.DIN1 (___90___20608), .DIN2 (________20538), .Q
       (___90___20609));
  and2s1 ______449346(.DIN1 (___90___20606), .DIN2 (___900__20605), .Q
       (___90___20607));
  nnd2s1 ______449347(.DIN1 (____9___20603), .DIN2 (________20242), .Q
       (____99__20604));
  and2s1 _______449348(.DIN1 (________19994), .DIN2 (___9____22524), .Q
       (____9___20602));
  nnd2s1 _____0_449349(.DIN1 (____9___19939), .DIN2 (________19315), .Q
       (____9___20601));
  nor2s1 _______449350(.DIN1 (____9___20599), .DIN2 (________19932), .Q
       (____9___20600));
  and2s1 ______449351(.DIN1 (____9___20597), .DIN2 (________19517), .Q
       (____9___20598));
  nnd2s1 _______449352(.DIN1 (____0___20044), .DIN2
       (____0________________18591), .Q (____9___20596));
  nor2s1 ______449353(.DIN1 (________20071), .DIN2 (____0___20889), .Q
       (____90__20595));
  nnd2s1 _____0_449354(.DIN1 (____0___20511), .DIN2 (________20593), .Q
       (_____9__20594));
  or2s1 _______449355(.DIN1 (____0________________18649), .DIN2
       (____0___20426), .Q (________20592));
  nnd2s1 ____449356(.DIN1 (________19971), .DIN2 (________21368), .Q
       (________20591));
  nnd2s1 _____0_449357(.DIN1 (________20055), .DIN2 (inData[6]), .Q
       (________20590));
  nor2s1 _____0_449358(.DIN1 (_________28828), .DIN2 (____9___20036),
       .Q (________20589));
  nor2s1 _______449359(.DIN1 (________20587), .DIN2 (________20250), .Q
       (________20588));
  nnd2s1 ___09_449360(.DIN1 (________19869), .DIN2 (inData[0]), .Q
       (________20586));
  or2s1 ____0__449361(.DIN1 (________20261), .DIN2 (________21054), .Q
       (_____0__20585));
  and2s1 _____9_449362(.DIN1 (________20583), .DIN2 (_____0__19992), .Q
       (_____9__20584));
  and2s1 ___09__449363(.DIN1 (________19890), .DIN2 (_________33370),
       .Q (________20582));
  nnd2s1 _____0_449364(.DIN1 (________20580), .DIN2 (_____0__19882), .Q
       (________20581));
  nnd2s1 _______449365(.DIN1 (____00__20040), .DIN2
       (_____________________18662), .Q (________20579));
  nor2s1 _______449366(.DIN1 (________19372), .DIN2 (________20028), .Q
       (________20578));
  nor2s1 _______449367(.DIN1 (___9____21592), .DIN2 (____9___20035), .Q
       (________20577));
  nnd2s1 ______449368(.DIN1 (_____9__20575), .DIN2 (________20574), .Q
       (_____0__20576));
  nnd2s1 _______449369(.DIN1 (___0____20756), .DIN2 (________20388), .Q
       (________20573));
  nnd2s1 _____9_449370(.DIN1 (________20555), .DIN2 (________21050), .Q
       (________20572));
  or2s1 _______449371(.DIN1 (________21862), .DIN2 (________20532), .Q
       (________20571));
  nor2s1 _______449372(.DIN1 (___9____20615), .DIN2 (________20829), .Q
       (________20568));
  nor2s1 _______449373(.DIN1 (_____0__21298), .DIN2 (________19863), .Q
       (_____0__20567));
  nor2s1 _______449374(.DIN1 (________20564), .DIN2 (________19883), .Q
       (________20565));
  nnd2s1 ______449375(.DIN1 (________20006), .DIN2 (________19384), .Q
       (________20563));
  nor2s1 _______449376(.DIN1 (________20561), .DIN2 (________20832), .Q
       (________20562));
  nor2s1 _______449377(.DIN1 (________20559), .DIN2 (________20052), .Q
       (________20560));
  or2s1 _____0_449378(.DIN1 (_____9__20557), .DIN2 (________20829), .Q
       (_____0__20558));
  and2s1 _____9_449379(.DIN1 (________20555), .DIN2 (___0____21684), .Q
       (________20556));
  nor2s1 _______449380(.DIN1 (___9_9__20662), .DIN2 (____0___20515), .Q
       (________20554));
  nor2s1 _____9_449381(.DIN1 (________19606), .DIN2 (_____9__20001), .Q
       (________20553));
  nor2s1 _____9_449382(.DIN1 (________20085), .DIN2 (________20551), .Q
       (________20552));
  nnd2s1 ___090_449383(.DIN1 (________19969), .DIN2 (inData[26]), .Q
       (________20550));
  and2s1 _____0_449384(.DIN1 (_____9__20548), .DIN2 (________22332), .Q
       (_____0__20549));
  nnd2s1 _______449385(.DIN1 (________20546), .DIN2 (___09___19845), .Q
       (________20547));
  and2s1 _______449386(.DIN1 (________20544), .DIN2 (________20543), .Q
       (________20545));
  nnd2s1 ______449387(.DIN1 (________19993), .DIN2 (inData[0]), .Q
       (________20542));
  nor2s1 _______449388(.DIN1 (_____________________18626), .DIN2
       (____9___19941), .Q (________20541));
  nnd2s1 _______449389(.DIN1 (________20024), .DIN2 (inData[10]), .Q
       (_____0__20540));
  nor2s1 _____9_449390(.DIN1 (___9_9__20662), .DIN2 (________20538), .Q
       (_____9__20539));
  or2s1 _____449391(.DIN1 (_____09__31192), .DIN2 (________20050), .Q
       (________20537));
  nnd2s1 _______449392(.DIN1 (________19972), .DIN2 (______18933), .Q
       (________20536));
  nor2s1 ______449393(.DIN1 (________20534), .DIN2 (____0___20518), .Q
       (________20535));
  nor2s1 _______449394(.DIN1 (________20009), .DIN2 (________20532), .Q
       (________20533));
  nor2s1 ______449395(.DIN1 (________19618), .DIN2 (____990__34521), .Q
       (________20531));
  nnd2s1 _______449396(.DIN1 (________19920), .DIN2 (________22050), .Q
       (_____0__20530));
  nnd2s1 ______449397(.DIN1 (___090), .DIN2 (________19342), .Q
       (_____9__20529));
  nor2s1 _______449398(.DIN1 (____9___21900), .DIN2 (____0___20889), .Q
       (________20528));
  or2s1 _______449399(.DIN1 (_____0__19669), .DIN2 (____0___20513), .Q
       (________20527));
  nor2s1 _____9_449400(.DIN1 (_____9__20846), .DIN2 (________20525), .Q
       (________20526));
  nnd2s1 _____9_449401(.DIN1 (________19928), .DIN2 (inData[4]), .Q
       (________20524));
  hi1s1 _______449402(.DIN (____9___21808), .Q (________21176));
  nor2s1 _____9_449403(.DIN1 (________21879), .DIN2 (________20832), .Q
       (________21044));
  nor2s1 ____9__449404(.DIN1 (________19329), .DIN2 (___09___19847), .Q
       (____90__21533));
  nor2s1 ____9__449405(.DIN1 (________20386), .DIN2 (________20538), .Q
       (_____9__21065));
  nor2s1 ______449406(.DIN1 (___9____21575), .DIN2 (_____9__20172), .Q
       (________21051));
  and2s1 ______449407(.DIN1 (________20482), .DIN2 (______18933), .Q
       (________21057));
  nnd2s1 _______449408(.DIN1 (_____9__21199), .DIN2 (________19998), .Q
       (___0____20737));
  hi1s1 ____0__449409(.DIN (________20523), .Q (________21236));
  nor2s1 ____9_449410(.DIN1 (________20561), .DIN2 (________20522), .Q
       (________21231));
  nor2s1 _______449411(.DIN1 (____9____30882), .DIN2 (________19896),
       .Q (________20840));
  nor2s1 _______449412(.DIN1 (________20868), .DIN2 (___9____20632), .Q
       (________20941));
  hi1s1 ____0__449413(.DIN (_________33186), .Q (________21315));
  hi1s1 _______449414(.DIN (________20521), .Q (_____0__21173));
  nnd2s1 ____90_449415(.DIN1 (________19973), .DIN2 (________19469), .Q
       (________21245));
  nnd2s1 ____449416(.DIN1 (_____0__20520), .DIN2 (________22110), .Q
       (____9___21253));
  nnd2s1 ____9__449417(.DIN1 (________20166), .DIN2 (________19913), .Q
       (________21192));
  nor2s1 _____0_449418(.DIN1 (________21180), .DIN2 (___9____20617), .Q
       (________21034));
  nor2s1 ______449419(.DIN1 (___0____19836), .DIN2 (____9___20505), .Q
       (________20841));
  nnd2s1 ______449420(.DIN1 (________21499), .DIN2 (________21098), .Q
       (____9___20976));
  nor2s1 _____0_449421(.DIN1 (____09__20519), .DIN2 (____0___20518), .Q
       (________21215));
  nor2s1 ____9__449422(.DIN1 (_____________________18636), .DIN2
       (_____9__22679), .Q (________22434));
  nnd2s1 ____9__449423(.DIN1 (____0___20517), .DIN2 (____0___21816), .Q
       (________21227));
  nnd2s1 _______449424(.DIN1 (________20396), .DIN2 (________20802), .Q
       (____9___21802));
  nnd2s1 _______449425(.DIN1 (____0___20516), .DIN2 (________21241), .Q
       (________21300));
  nor2s1 _______449426(.DIN1 (________19980), .DIN2 (____0___20515), .Q
       (________23239));
  nor2s1 ____9__449427(.DIN1 (________19935), .DIN2 (________21054), .Q
       (___0____22597));
  nor2s1 ____00_449428(.DIN1 (___09___19851), .DIN2 (____0___20514), .Q
       (__9_00__26989));
  nor2s1 _______449429(.DIN1 (____90__20126), .DIN2 (____0___20513), .Q
       (________21189));
  nor2s1 ____9_449430(.DIN1 (___90___21546), .DIN2 (________19906), .Q
       (_____0__21056));
  nnd2s1 ____9__449431(.DIN1 (________21043), .DIN2 (______18933), .Q
       (________21089));
  nor2s1 ____9_449432(.DIN1 (________20387), .DIN2 (________20375), .Q
       (________23052));
  nnd2s1 _______449433(.DIN1 (____9___20597), .DIN2 (___99___19769), .Q
       (________22067));
  nor2s1 _______449434(.DIN1 (________21213), .DIN2 (____0___20512), .Q
       (________21194));
  nnd2s1 ____0__449435(.DIN1 (_____0__19927), .DIN2 (_____9__19908), .Q
       (________24923));
  nnd2s1 _____9_449436(.DIN1 (____0___20511), .DIN2 (____00__20510), .Q
       (________21195));
  nor2s1 _______449437(.DIN1 (____99__20509), .DIN2 (____9___20507), .Q
       (_____9__21219));
  nor2s1 _______449438(.DIN1 (____9___20508), .DIN2 (____9___20507), .Q
       (________25622));
  hi1s1 ______449439(.DIN (____9___20506), .Q (____9___21069));
  nor2s1 ____9__449440(.DIN1 (____9___20504), .DIN2 (________20538), .Q
       (________21202));
  or2s1 _______449441(.DIN1 (___9____20615), .DIN2 (____9___20505), .Q
       (________24822));
  nor2s1 ____0__449442(.DIN1 (_____9__19926), .DIN2 (____90__20500), .Q
       (_________28365));
  nnd2s1 _______449443(.DIN1 (________21206), .DIN2 (______0__28643),
       .Q (________21207));
  nor2s1 ____9__449444(.DIN1 (____9___20504), .DIN2 (____0___20515), .Q
       (________21223));
  nnd2s1 ______449445(.DIN1 (____9___20503), .DIN2 (______0__28643), .Q
       (_____0__21210));
  nor2s1 ____9_449446(.DIN1 (________20376), .DIN2 (____9___20502), .Q
       (___9____26215));
  nor2s1 ____0__449447(.DIN1 (________19189), .DIN2 (________19878), .Q
       (______9__33247));
  nor2s1 ____0__449448(.DIN1 (___9____19722), .DIN2 (____90__20031), .Q
       (______0__33107));
  nor2s1 _______449449(.DIN1 (____9___20501), .DIN2 (_________32919),
       .Q (_________32639));
  nor2s1 ____00_449450(.DIN1 (________19541), .DIN2 (____90__20500), .Q
       (____009__31815));
  nor2s1 ____00_449451(.DIN1 (____00__19852), .DIN2 (____9___20033), .Q
       (____0____30981));
  hi1s1 _______449452(.DIN (___9____20646), .Q (_____0__21279));
  or2s1 _____0_449453(.DIN1 (_____0__21298), .DIN2 (________19979), .Q
       (________21424));
  nor2s1 ____99_449454(.DIN1 (_____0___33866), .DIN2 (________20408),
       .Q (________21281));
  nor2s1 ____0__449455(.DIN1 (___0____19788), .DIN2 (________20026), .Q
       (_________30472));
  nor2s1 ____00_449456(.DIN1 (_____9__20499), .DIN2 (________19870), .Q
       (_________32410));
  nor2s1 ____00_449457(.DIN1 (________19420), .DIN2 (________19889), .Q
       (_________34077));
  nnd2s1 _______449458(.DIN1 (________19904), .DIN2 (________19577), .Q
       (____00___31810));
  nor2s1 ____00_449459(.DIN1 (_________33989), .DIN2 (___0____19830),
       .Q (_____00__33954));
  nor2s1 ____00_449460(.DIN1 (________19620), .DIN2 (________19930), .Q
       (_____0___32851));
  nnd2s1 _____449461(.DIN1 (________21530), .DIN2 (________20497), .Q
       (________20498));
  nnd2s1 ______449462(.DIN1 (_____9__20087), .DIN2 (________19978), .Q
       (________20496));
  nnd2s1 _______449463(.DIN1 (________20383), .DIN2
       (_________________18783), .Q (________20495));
  and2s1 _____9_449464(.DIN1 (___9____19692), .DIN2
       (__________0___0___18823), .Q (________20494));
  nor2s1 _______449465(.DIN1 (_____9__20491), .DIN2 (________21508), .Q
       (_____0__20492));
  and2s1 ______449466(.DIN1 (_____9__19900), .DIN2 (inData[12]), .Q
       (________20490));
  nor2s1 _______449467(.DIN1 (____0___19401), .DIN2 (____9___20417), .Q
       (________20489));
  nnd2s1 _______449468(.DIN1 (________19901), .DIN2 (inData[30]), .Q
       (________20488));
  nor2s1 _______449469(.DIN1 (________20461), .DIN2 (___9____20628), .Q
       (________20487));
  nor2s1 ______449470(.DIN1 (_____________0___18679), .DIN2
       (________20485), .Q (________20486));
  hi1s1 ____0__449471(.DIN (________20814), .Q (_____0__20484));
  nor2s1 _______449472(.DIN1 (________19519), .DIN2 (________20482), .Q
       (_____9__20483));
  hi1s1 _____0_449473(.DIN (_____9__20912), .Q (________20481));
  nnd2s1 _______449474(.DIN1 (________20377), .DIN2 (________19471), .Q
       (________20480));
  hi1s1 _______449475(.DIN (________20478), .Q (________20479));
  nor2s1 _____449476(.DIN1 (_____0__19449), .DIN2 (____9___19942), .Q
       (________20477));
  hi1s1 _____9_449477(.DIN (____0___20794), .Q (________20476));
  nnd2s1 _______449478(.DIN1 (_____0__20474), .DIN2
       (_____________________18667), .Q (________20475));
  nnd2s1 _______449479(.DIN1 (_____0__20474), .DIN2 (________21976), .Q
       (________20473));
  or2s1 ______449480(.DIN1 (_____________________18664), .DIN2
       (________22000), .Q (________20472));
  or2s1 ____0__449481(.DIN1 (________20470), .DIN2 (________20469), .Q
       (________20471));
  and2s1 ____9__449482(.DIN1 (________20467), .DIN2 (____00__20510), .Q
       (________20468));
  nor2s1 _______449483(.DIN1 (________19662), .DIN2 (________20485), .Q
       (________20466));
  or2s1 ____9__449484(.DIN1 (___0____19822), .DIN2 (_____9__20464), .Q
       (_____0__20465));
  and2s1 ____9__449485(.DIN1 (____9___20881), .DIN2 (________21387), .Q
       (________20463));
  or2s1 _______449486(.DIN1 (________20461), .DIN2 (____0___20515), .Q
       (________20462));
  hi1s1 ______449487(.DIN (________20459), .Q (________20460));
  and2s1 ____00_449488(.DIN1 (________21774), .DIN2 (___0____20748), .Q
       (________20458));
  nor2s1 _______449489(.DIN1 (___9_0), .DIN2 (________19899), .Q
       (________20457));
  nor2s1 _______449490(.DIN1 (_____0__19371), .DIN2 (________20016), .Q
       (_____0__20456));
  nor2s1 _______449491(.DIN1 (________20454), .DIN2 (________20522), .Q
       (_____9__20455));
  nnd2s1 ______449492(.DIN1 (_____0__20012), .DIN2 (___9____19757), .Q
       (________20453));
  and2s1 _______449493(.DIN1 (___0____21698), .DIN2 (________20543), .Q
       (________20452));
  nor2s1 ____09_449494(.DIN1
       (______________________________________0_____________18891),
       .DIN2 (____9___20597), .Q (________20451));
  nnd2s1 _______449495(.DIN1 (________19888), .DIN2 (________19507), .Q
       (________20449));
  hi1s1 _______449496(.DIN (___9_0__20654), .Q (_____9__20448));
  hi1s1 _______449497(.DIN (________20446), .Q (________20447));
  hi1s1 _______449498(.DIN (________20444), .Q (________20445));
  nnd2s1 _______449499(.DIN1 (________20442), .DIN2 (________21193), .Q
       (________20443));
  nnd2s1 _______449500(.DIN1 (____09__20048), .DIN2 (___0____19823), .Q
       (________20441));
  nnd2s1 _______449501(.DIN1 (________20442), .DIN2 (________20843), .Q
       (________20440));
  nor2s1 _______449502(.DIN1 (____9___19391), .DIN2 (____0___19855), .Q
       (_____0__20439));
  nnd2s1 ______449503(.DIN1 (________20056), .DIN2 (________19868), .Q
       (_____9__20438));
  nor2s1 _______449504(.DIN1 (_________33835), .DIN2 (____9___20597),
       .Q (________20437));
  and2s1 _______449505(.DIN1 (________19925), .DIN2 (________20435), .Q
       (________20436));
  nor2s1 _______449506(.DIN1 (________19656), .DIN2 (________19988), .Q
       (________20434));
  xor2s1 _____449507(.DIN1 (_____9__19658), .DIN2 (_________28939), .Q
       (________20433));
  nnd2s1 _______449508(.DIN1 (________20013), .DIN2 (___9____20638), .Q
       (________20432));
  hi1s1 _______449509(.DIN (________20925), .Q (________20431));
  or2s1 _____449510(.DIN1 (____00__19496), .DIN2 (____9___20038), .Q
       (________20430));
  nor2s1 ______449511(.DIN1 (____0___20984), .DIN2 (________20469), .Q
       (_____0__20429));
  and2s1 _______449512(.DIN1 (________20555), .DIN2 (________22332), .Q
       (____09__20428));
  nor2s1 _______449513(.DIN1 (____0________________18652), .DIN2
       (____0___20426), .Q (____0___20427));
  nnd2s1 _______449514(.DIN1 (____0___20516), .DIN2 (____0___20423), .Q
       (____0___20424));
  and2s1 _______449515(.DIN1 (________20544), .DIN2 (____9___21256), .Q
       (____0___20422));
  nor2s1 _______449516(.DIN1 (________21407), .DIN2 (____00__20420), .Q
       (____0___20421));
  nor2s1 _____449517(.DIN1 (____9__19015), .DIN2 (________20061), .Q
       (____99__20419));
  nor2s1 ____9__449518(.DIN1 (________19176), .DIN2 (____9___20417), .Q
       (____9___20418));
  nor2s1 _______449519(.DIN1 (_________31220), .DIN2 (_________30592),
       .Q (____9___20416));
  nnd2s1 _______449520(.DIN1 (________20403), .DIN2 (________20355), .Q
       (____9___20415));
  nor2s1 _______449521(.DIN1 (____9___20413), .DIN2 (________21198), .Q
       (____9___20414));
  nor2s1 ____9_449522(.DIN1 (_____9__19984), .DIN2 (________20003), .Q
       (____9___20412));
  nnd2s1 _______449523(.DIN1 (____9___20603), .DIN2 (____90__20410), .Q
       (____9___20411));
  nnd2s1 ______449524(.DIN1 (_____9__21199), .DIN2 (____9___20503), .Q
       (________20409));
  nor2s1 _______449525(.DIN1 (___0____20730), .DIN2 (________20015), .Q
       (________20407));
  nnd2s1 ____9__449526(.DIN1 (________22000), .DIN2 (________20405), .Q
       (________20406));
  and2s1 ____9__449527(.DIN1 (________20843), .DIN2 (________20403), .Q
       (________20404));
  nnd2s1 ____9__449528(.DIN1 (________20917), .DIN2 (_____9__20401), .Q
       (_____0__20402));
  nor2s1 ____449529(.DIN1 (________21115), .DIN2 (________22000), .Q
       (________20400));
  nor2s1 ____09_449530(.DIN1 (________20398), .DIN2 (_____9__20058), .Q
       (________20399));
  or2s1 _______449531(.DIN1 (____0___19853), .DIN2 (____0___20328), .Q
       (________20397));
  nnd2s1 _____0_449532(.DIN1 (________20396), .DIN2 (________20065), .Q
       (________21789));
  nnd2s1 _______449533(.DIN1 (________19982), .DIN2 (____9___20599), .Q
       (___9____20642));
  nor2s1 _______449534(.DIN1 (________20395), .DIN2 (________20378), .Q
       (___0____20710));
  nor2s1 _____9_449535(.DIN1 (_____9__20846), .DIN2 (________21198), .Q
       (_____0__21120));
  nor2s1 _____9_449536(.DIN1 (________19968), .DIN2 (_____9__19676), .Q
       (________21237));
  nnd2s1 ____9__449537(.DIN1 (________20394), .DIN2 (________20393), .Q
       (________21196));
  nnd2s1 _______449538(.DIN1 (_____9__20464), .DIN2 (_____0__20392), .Q
       (___9____20641));
  hi1s1 _______449539(.DIN (___9_9__20653), .Q (________21064));
  hi1s1 ______449540(.DIN (_____9__20391), .Q (____9___21162));
  hi1s1 _____0_449541(.DIN (___9____20659), .Q (________21047));
  nor2s1 ____9_449542(.DIN1 (____9___19202), .DIN2 (____0___20426), .Q
       (________21104));
  nnd2s1 ____9__449543(.DIN1 (________20017), .DIN2 (________20390), .Q
       (___0_9__20715));
  nor2s1 ____9__449544(.DIN1 (____0___20518), .DIN2 (___9____20628), .Q
       (___00___20701));
  hi1s1 _______449545(.DIN (_________35092), .Q (________21049));
  nor2s1 _______449546(.DIN1 (________20389), .DIN2 (________20832), .Q
       (_____9__21045));
  hi1s1 _____9_449547(.DIN (___0____20750), .Q (_____9__21055));
  nnd2s1 ____0__449548(.DIN1 (________20388), .DIN2 (________22341), .Q
       (____9___21067));
  nnd2s1 ____0__449549(.DIN1 (________21201), .DIN2 (________21218), .Q
       (___9_0__20663));
  nor2s1 ____90_449550(.DIN1 (____0________________18651), .DIN2
       (________19894), .Q (________21283));
  nor2s1 ____90_449551(.DIN1 (________20387), .DIN2 (____9___20502), .Q
       (________20860));
  hi1s1 _____0_449552(.DIN (___9____20655), .Q (_____0__21200));
  nor2s1 _____449553(.DIN1 (________20386), .DIN2 (____0___20515), .Q
       (________21042));
  nor2s1 ____90_449554(.DIN1 (____0________________18651), .DIN2
       (________19934), .Q (_____9__21038));
  hi1s1 _____449555(.DIN (________20385), .Q (________21291));
  nor2s1 ____9__449556(.DIN1 (________20384), .DIN2 (____9___20505), .Q
       (________21221));
  hi1s1 _____0_449557(.DIN (_________35090), .Q (________21052));
  nnd2s1 _______449558(.DIN1 (________20383), .DIN2 (_____0__20382), .Q
       (________21339));
  nnd2s1 ____0_449559(.DIN1 (____0___21905), .DIN2 (____0___21988), .Q
       (________21133));
  nor2s1 _____449560(.DIN1 (_____9__20491), .DIN2 (_____9__21894), .Q
       (________21224));
  nnd2s1 ____0__449561(.DIN1 (_____0__19985), .DIN2 (_____9__20381), .Q
       (_____9__21129));
  nor2s1 ____0__449562(.DIN1 (________19661), .DIN2 (________20485), .Q
       (_____9__21182));
  or2s1 _____9_449563(.DIN1 (_____________________18667), .DIN2
       (________22000), .Q (________22312));
  nnd2s1 ______449564(.DIN1 (________20482), .DIN2
       (____0____________0_), .Q (________21062));
  nnd2s1 ______449565(.DIN1 (________21385), .DIN2 (________20380), .Q
       (_____9__21093));
  nor2s1 ____99_449566(.DIN1 (_____0__19534), .DIN2 (____0___19858), .Q
       (____9___21158));
  nnd2s1 ____0__449567(.DIN1 (_____9__20464), .DIN2
       (__________________0___18628), .Q (________21145));
  nor2s1 _______449568(.DIN1 (____0________________18648), .DIN2
       (_____9__21894), .Q (________21174));
  nor2s1 ____0__449569(.DIN1 (________21114), .DIN2 (____00__20420), .Q
       (________21141));
  hi1s1 ______449570(.DIN (_________35094), .Q (_________31336));
  hi1s1 _______449571(.DIN (____0___21363), .Q (____9___21346));
  hi1s1 ______449572(.DIN (____9___21803), .Q (________21323));
  nnd2s1 ____0__449573(.DIN1 (________21375), .DIN2 (________20200), .Q
       (________21113));
  hi1s1 ______449574(.DIN (________20379), .Q (________21058));
  hi1s1 _______449575(.DIN (___0____20734), .Q (________21785));
  nnd2s1 _______449576(.DIN1 (________20378), .DIN2
       (____0_________________18596), .Q (________21974));
  and2s1 ____0_449577(.DIN1 (________21375), .DIN2 (____0___21812), .Q
       (________21136));
  nor2s1 _____9_449578(.DIN1 (________21889), .DIN2 (________21788), .Q
       (____9___21257));
  hi1s1 ______449579(.DIN (_________30428), .Q (_________31578));
  nor2s1 ______449580(.DIN1 (________20374), .DIN2 (________20377), .Q
       (________21212));
  nor2s1 ____0__449581(.DIN1 (________20018), .DIN2 (____00__20510), .Q
       (___000___27171));
  or2s1 _____9_449582(.DIN1 (_____0__21046), .DIN2 (____9___20507), .Q
       (________21217));
  nor2s1 _____0_449583(.DIN1 (________20376), .DIN2 (________20375), .Q
       (__9_____26632));
  or2s1 _____449584(.DIN1 (___9____21575), .DIN2 (________20930), .Q
       (_____9__21326));
  hi1s1 _______449585(.DIN (___9____20649), .Q (____90__21066));
  hi1s1 _______449586(.DIN (_________31376), .Q (______0__33983));
  nor2s1 _____0_449587(.DIN1 (________20374), .DIN2 (________19867), .Q
       (________21204));
  nor2s1 ______449588(.DIN1 (________19484), .DIN2 (________20025), .Q
       (_____0___30999));
  nor2s1 _______449589(.DIN1 (____9___20599), .DIN2 (________20054), .Q
       (_________31479));
  nor2s1 _______449590(.DIN1 (____09__20235), .DIN2 (_____9__21199), .Q
       (_________31153));
  nor2s1 ____449591(.DIN1 (___0_0__19835), .DIN2 (_____0__19909), .Q
       (_________33384));
  hi1s1 _______449592(.DIN (___9____20677), .Q (________21232));
  nor2s1 ____0__449593(.DIN1 (___9__), .DIN2 (________19876), .Q
       (_________34362));
  nor2s1 _______449594(.DIN1 (________19387), .DIN2 (___0____19794), .Q
       (________20373));
  or2s1 _______449595(.DIN1 (___9____19743), .DIN2 (____9___20224), .Q
       (_____0__20372));
  nor2s1 ____00_449596(.DIN1 (________19673), .DIN2 (________20390), .Q
       (_____9__20371));
  nor2s1 ______449597(.DIN1 (_____09__31192), .DIN2 (____9___19684), .Q
       (________20370));
  nnd2s1 _______449598(.DIN1 (________20497), .DIN2 (________20368), .Q
       (________20369));
  nnd2s1 _______449599(.DIN1 (_____9__20216), .DIN2 (_____0__20002), .Q
       (________20367));
  and2s1 _______449600(.DIN1 (________20349), .DIN2
       (_________________18709), .Q (________20366));
  nor2s1 _____9_449601(.DIN1 (________21509), .DIN2 (________22341), .Q
       (________20365));
  hi1s1 _______449602(.DIN (____9___20502), .Q (________20364));
  nor2s1 _______449603(.DIN1 (___00___19776), .DIN2 (_____0__20362), .Q
       (________20363));
  and2s1 ____9__449604(.DIN1 (________21313), .DIN2 (_______19024), .Q
       (_____9__20361));
  nnd2s1 _______449605(.DIN1 (________20359), .DIN2 (_____0__20392), .Q
       (________20360));
  nnd2s1 _______449606(.DIN1 (_____9__20341), .DIN2 (________19674), .Q
       (________20358));
  nor2s1 _____9_449607(.DIN1 (________19364), .DIN2 (___0_9), .Q
       (________20357));
  and2s1 _______449608(.DIN1 (________21193), .DIN2 (________20355), .Q
       (________20356));
  nor2s1 ____99_449609(.DIN1 (________20353), .DIN2 (_____0__20352), .Q
       (________20354));
  nor2s1 ____99_449610(.DIN1 (________20901), .DIN2 (________19672), .Q
       (_____9__20351));
  nnd2s1 ______449611(.DIN1 (________20349), .DIN2 (________19535), .Q
       (________20350));
  or2s1 _______449612(.DIN1 (________21131), .DIN2 (________20347), .Q
       (________20348));
  nnd2s1 ______449613(.DIN1 (________20286), .DIN2 (_____0__19439), .Q
       (________20346));
  nnd2s1 ____9__449614(.DIN1 (________20110), .DIN2 (________20813), .Q
       (________20345));
  or2s1 ______449615(.DIN1 (________20343), .DIN2 (___9____19738), .Q
       (________20344));
  nor2s1 ____449616(.DIN1 (___9____19739), .DIN2 (_____9__20341), .Q
       (_____0__20342));
  and2s1 ____449617(.DIN1 (________22037), .DIN2 (___9____20651), .Q
       (________20340));
  nor2s1 ____99_449618(.DIN1 (___9____19752), .DIN2 (________20338), .Q
       (________20339));
  and2s1 ____9__449619(.DIN1 (____90__25071), .DIN2 (________20336), .Q
       (________20337));
  and2s1 ____9__449620(.DIN1 (________21470), .DIN2 (___0_0__21658), .Q
       (________20335));
  nor2s1 _______449621(.DIN1 (_____________________18638), .DIN2
       (________20386), .Q (________20334));
  and2s1 ____9__449622(.DIN1 (________20268), .DIN2 (________21115), .Q
       (________20333));
  nor2s1 ____9__449623(.DIN1 (_____0__20392), .DIN2 (________19642), .Q
       (_____0__20332));
  nnd2s1 ____9__449624(.DIN1 (________19654), .DIN2 (____0___20330), .Q
       (____09__20331));
  nnd2s1 ____9_449625(.DIN1 (___9____19715), .DIN2 (________20493), .Q
       (____0___20329));
  nnd2s1 ____9__449626(.DIN1 (________20338), .DIN2 (___9____19756), .Q
       (____0___20327));
  nor2s1 _______449627(.DIN1 (____9___19392), .DIN2 (________19635), .Q
       (____0___20326));
  nor2s1 ____9__449628(.DIN1 (_____0__21971), .DIN2 (________21310), .Q
       (____0___20325));
  nnd2s1 ______449629(.DIN1 (___9____20645), .DIN2 (________20081), .Q
       (____00__20324));
  nnd2s1 ____9__449630(.DIN1 (________20120), .DIN2 (________19228), .Q
       (____99__20323));
  nor2s1 ____9__449631(.DIN1 (__________________0___18628), .DIN2
       (________19625), .Q (____9___20322));
  or2s1 ____9_449632(.DIN1 (___9____20666), .DIN2 (________20384), .Q
       (____9___20321));
  nor2s1 _____9_449633(.DIN1 (____9___20319), .DIN2 (________19623), .Q
       (____9___20320));
  xor2s1 ____09_449634(.DIN1 (_______19028), .DIN2 (_________30524), .Q
       (____9___20318));
  nor2s1 _______449635(.DIN1 (_________31702), .DIN2 (___9____19747),
       .Q (____9___20317));
  or2s1 ____9__449636(.DIN1 (___0____19842), .DIN2 (____99__20509), .Q
       (____9___20316));
  or2s1 ______449637(.DIN1 (___9_0__19717), .DIN2 (________21228), .Q
       (____9___20315));
  nnd2s1 ____99_449638(.DIN1 (________20338), .DIN2 (_____9__20313), .Q
       (____90__20314));
  nor2s1 ____9__449639(.DIN1 (________20311), .DIN2 (________20117), .Q
       (________20312));
  nnd2s1 _______449640(.DIN1 (____9___19678), .DIN2 (________20309), .Q
       (________20310));
  nor2s1 _____9_449641(.DIN1 (________20307), .DIN2 (_____0__21046), .Q
       (________20308));
  nor2s1 ____9__449642(.DIN1 (________21333), .DIN2 (________21213), .Q
       (________20306));
  nor2s1 _______449643(.DIN1 (________20300), .DIN2 (_____0__20304), .Q
       (________20305));
  nor2s1 ____9_449644(.DIN1 (____0___19497), .DIN2 (___0____19779), .Q
       (_____9__20303));
  nnd2s1 ____90_449645(.DIN1 (________22211), .DIN2 (________19578), .Q
       (________20302));
  nor2s1 _____9_449646(.DIN1 (________21407), .DIN2 (________20300), .Q
       (________20301));
  and2s1 _______449647(.DIN1 (___0____20756), .DIN2 (________20809), .Q
       (________20299));
  and2s1 _____449648(.DIN1 (________21313), .DIN2 (___9____19759), .Q
       (________20298));
  nnd2s1 ____9__449649(.DIN1 (_____0__21335), .DIN2 (________21337), .Q
       (________20297));
  xor2s1 _______449650(.DIN1 (____99___35108), .DIN2 (________20295),
       .Q (________20296));
  nnd2s1 ______449651(.DIN1 (___9____19740), .DIN2 (____9___19491), .Q
       (_____0__20294));
  nor2s1 ____9_449652(.DIN1 (________20292), .DIN2 (___90___21544), .Q
       (_____9__20293));
  nor2s1 _______449653(.DIN1 (_____9__20557), .DIN2 (___0____19832), .Q
       (________20291));
  or2s1 _____0_449654(.DIN1 (____9___21070), .DIN2 (________21211), .Q
       (________20290));
  nor2s1 _______449655(.DIN1 (________20288), .DIN2 (____9___19683), .Q
       (________20289));
  nnd2s1 _______449656(.DIN1 (___00___19774), .DIN2 (________20286), .Q
       (________20287));
  nnd2s1 ____0__449657(.DIN1 (________19632), .DIN2 (_________30612),
       .Q (________20285));
  nnd2s1 _______449658(.DIN1 (________20389), .DIN2 (_____9__20283), .Q
       (_____0__20284));
  or2s1 _______449659(.DIN1 (____9___20881), .DIN2 (___9_9__19736), .Q
       (________20282));
  nor2s1 _______449660(.DIN1 (________20280), .DIN2 (___009), .Q
       (________20281));
  nor2s1 _____0_449661(.DIN1 (________20278), .DIN2 (________20277), .Q
       (________20279));
  nnd2s1 _______449662(.DIN1 (_____9__21278), .DIN2 (_______18973), .Q
       (________20276));
  and2s1 _____449663(.DIN1 (____9___19680), .DIN2 (_____0__20274), .Q
       (________20275));
  and2s1 ____90_449664(.DIN1 (________19962), .DIN2 (______0__30345),
       .Q (_____9__20273));
  or2s1 ______449665(.DIN1 (_____________________18665), .DIN2
       (________20271), .Q (________20272));
  and2s1 _____0_449666(.DIN1 (________19967), .DIN2 (_____9__21278), .Q
       (________20270));
  nnd2s1 _______449667(.DIN1 (________20268), .DIN2 (___0____20730), .Q
       (________20269));
  nnd2s1 _______449668(.DIN1 (___9_9__20643), .DIN2 (________19363), .Q
       (________20267));
  nnd2s1 _______449669(.DIN1 (________19616), .DIN2 (___0____19808), .Q
       (________20266));
  nnd2s1 _______449670(.DIN1 (___0____19814), .DIN2 (________19898), .Q
       (________20265));
  or2s1 _______449671(.DIN1 (_____________18898), .DIN2
       (________20154), .Q (_____0__20264));
  nor2s1 _______449672(.DIN1 (_____0__21230), .DIN2 (________20470), .Q
       (_____9__20263));
  or2s1 _______449673(.DIN1 (________21502), .DIN2 (________20261), .Q
       (________20262));
  nor2s1 ______449674(.DIN1 (___9_0__19727), .DIN2 (___9____19734), .Q
       (________20260));
  nnd2s1 _______449675(.DIN1 (___9_0__19745), .DIN2 (___0_9__19825), .Q
       (________20259));
  and2s1 _______449676(.DIN1 (___9____20645), .DIN2 (________20257), .Q
       (________20258));
  nor2s1 ______449677(.DIN1 (________19264), .DIN2 (___0_0__19785), .Q
       (________20256));
  nnd2s1 _______449678(.DIN1 (_____0__20254), .DIN2 (___0____19833), .Q
       (________20255));
  nor2s1 ______449679(.DIN1 (___9____19750), .DIN2 (________20252), .Q
       (________20253));
  hi1s1 _______449680(.DIN (________20250), .Q (________20251));
  nnd2s1 _______449681(.DIN1 (___9____19760), .DIN2 (_____0__22063), .Q
       (________20249));
  nor2s1 ______449682(.DIN1 (________19061), .DIN2 (________20247), .Q
       (________20248));
  and2s1 _______449683(.DIN1 (________21313), .DIN2 (_________34477),
       .Q (________20246));
  or2s1 _____9_449684(.DIN1 (_____________________18620), .DIN2
       (_____9__19621), .Q (_____0__20245));
  nnd2s1 _____449685(.DIN1 (________20831), .DIN2 (________19174), .Q
       (_____9__20244));
  and2s1 _______449686(.DIN1 (________20242), .DIN2 (________20241), .Q
       (________20243));
  nnd2s1 _______449687(.DIN1 (___0____19795), .DIN2 (________20027), .Q
       (________20240));
  nor2s1 ______449688(.DIN1 (________19437), .DIN2 (____9___20221), .Q
       (________20239));
  nor2s1 _______449689(.DIN1 (________20237), .DIN2 (________20389), .Q
       (________20238));
  nor2s1 ______449690(.DIN1 (_____9__21513), .DIN2 (________20271), .Q
       (________20236));
  nor2s1 _______449691(.DIN1 (________20091), .DIN2 (___9____19731), .Q
       (____0___20234));
  nnd2s1 _______449692(.DIN1 (____9___19394), .DIN2 (________19660), .Q
       (____0___20233));
  nnd2s1 _____0_449693(.DIN1 (________20077), .DIN2 (________20813), .Q
       (____0___20232));
  nnd2s1 _____0_449694(.DIN1 (________19548), .DIN2 (___0____19790), .Q
       (____0___20231));
  nnd2s1 _____449695(.DIN1 (________20169), .DIN2 (___90___19687), .Q
       (____0___20230));
  and2s1 _______449696(.DIN1 (___0____21680), .DIN2 (_________34447),
       .Q (____0___20229));
  nnd2s1 _______449697(.DIN1 (________19671), .DIN2 (inData[0]), .Q
       (____0___20228));
  and2s1 ______449698(.DIN1 (____90__21801), .DIN2 (____00__20226), .Q
       (____0___20227));
  nor2s1 _______449699(.DIN1 (___0____19816), .DIN2 (____9___20224), .Q
       (____99__20225));
  nnd2s1 _______449700(.DIN1 (________20075), .DIN2 (________20194), .Q
       (____9___20223));
  nor2s1 _______449701(.DIN1 (________19343), .DIN2 (____9___20221), .Q
       (____9___20222));
  and2s1 _____449702(.DIN1 (_____9__20106), .DIN2 (____________9_), .Q
       (____9___20220));
  hi1s1 _______449703(.DIN (____9_9__33643), .Q (____0___21083));
  nor2s1 ____0_449704(.DIN1 (____9___20219), .DIN2 (____9___20218), .Q
       (________20478));
  hi1s1 _____9_449705(.DIN (____90__20217), .Q (_____9__22156));
  and2s1 _______449706(.DIN1 (_____9__20216), .DIN2
       (____0________________18652), .Q (___00___20705));
  nor2s1 ____0__449707(.DIN1 (________20215), .DIN2 (____99__20509), .Q
       (________20459));
  nor2s1 ____0_449708(.DIN1 (________22113), .DIN2 (___0____20763), .Q
       (________20385));
  hi1s1 _______449709(.DIN (________20214), .Q (________20910));
  nnd2s1 ______449710(.DIN1 (_____0__20254), .DIN2 (________20213), .Q
       (________20523));
  nor2s1 ____0__449711(.DIN1 (___0____21699), .DIN2 (____9___19944), .Q
       (_____9__20391));
  nnd2s1 _____0_449712(.DIN1 (_____9__20816), .DIN2
       (____0________________18648), .Q (________20521));
  hi1s1 _______449713(.DIN (________21530), .Q (____0___20888));
  nnd2s1 ____9__449714(.DIN1 (_____9__20068), .DIN2 (______18933), .Q
       (________20450));
  hi1s1 _______449715(.DIN (________20829), .Q (________20803));
  xor2s1 _____0_449716(.DIN1 (________20212), .DIN2 (______0__28643),
       .Q (_________28556));
  or2s1 ______449717(.DIN1 (___9____19729), .DIN2 (________20211), .Q
       (________21016));
  hi1s1 _____0_449718(.DIN (________20482), .Q (___0____20758));
  and2s1 _______449719(.DIN1 (________20210), .DIN2 (____0___21360), .Q
       (___0____20719));
  nnd2s1 _______449720(.DIN1 (_____9__20932), .DIN2 (________20209), .Q
       (____0___20887));
  nnd2s1 _______449721(.DIN1 (________19633), .DIN2 (________21797), .Q
       (________21144));
  or2s1 _______449722(.DIN1 (____0_________________18596), .DIN2
       (________20177), .Q (________20800));
  nor2s1 _______449723(.DIN1 (_____0__20382), .DIN2 (_____9__21344), .Q
       (________21012));
  nnd2s1 _____449724(.DIN1 (_____9__20216), .DIN2 (_____9__20011), .Q
       (________22672));
  nor2s1 _____9_449725(.DIN1 (____9___19296), .DIN2 (________20203), .Q
       (________20842));
  nnd2s1 _____9_449726(.DIN1 (________19670), .DIN2 (________21976), .Q
       (________21018));
  nor2s1 ____0__449727(.DIN1 (________19653), .DIN2 (________22037), .Q
       (____90__21156));
  nnd2s1 ____0__449728(.DIN1 (________22339), .DIN2 (________20070), .Q
       (___0_0__20752));
  nor2s1 _______449729(.DIN1 (____0___21080), .DIN2 (________20277), .Q
       (________20814));
  nor2s1 ____9__449730(.DIN1 (________21131), .DIN2 (_____0__20304), .Q
       (___9____20685));
  nor2s1 _______449731(.DIN1 (________19866), .DIN2 (________20063), .Q
       (_________30428));
  nnd2s1 ____449732(.DIN1 (___0____19781), .DIN2
       (_________________0___18607), .Q (___9____20677));
  nnd2s1 ____0__449733(.DIN1 (________21193), .DIN2 (________20208), .Q
       (________21048));
  or2s1 ____0__449734(.DIN1 (_____________________18668), .DIN2
       (________22110), .Q (________22187));
  nor2s1 ____0__449735(.DIN1 (___9____19725), .DIN2 (________21887), .Q
       (___0____20767));
  nor2s1 _______449736(.DIN1 (_____0__20207), .DIN2 (_____0__20304), .Q
       (________20874));
  hi1s1 _______449737(.DIN (_____9__20206), .Q (___0_9__21657));
  nnd2s1 ____0_449738(.DIN1 (________20205), .DIN2
       (____0________________18592), .Q (___0____20750));
  hi1s1 _______449739(.DIN (____0___21357), .Q (____0___20791));
  and2s1 ____0__449740(.DIN1 (____9___20224), .DIN2
       (_________________0___18607), .Q (_____9__20826));
  and2s1 ____0__449741(.DIN1 (________20210), .DIN2 (________20204), .Q
       (___0____20765));
  nnd2s1 ______449742(.DIN1 (________20074), .DIN2
       (_________________0___18633), .Q (___9____20649));
  nor2s1 ____0__449743(.DIN1 (___0____19789), .DIN2 (________20203), .Q
       (____0___20794));
  hi1s1 _____449744(.DIN (________21208), .Q (___0____21671));
  or2s1 ____449745(.DIN1 (___9_0__19737), .DIN2 (________20203), .Q
       (_____9__20836));
  nor2s1 _____0_449746(.DIN1 (___0____19807), .DIN2 (________20831), .Q
       (________20970));
  and2s1 _______449747(.DIN1 (___9____20645), .DIN2 (________20202), .Q
       (________25582));
  nnd2s1 ____0__449748(.DIN1 (________20066), .DIN2
       (____0________________18592), .Q (________20849));
  nnd2s1 ______449749(.DIN1 (________20268), .DIN2 (___9____19694), .Q
       (________22674));
  nnd2s1 _______449750(.DIN1 (________20201), .DIN2 (________20200), .Q
       (________20925));
  and2s1 _____449751(.DIN1 (________20252), .DIN2
       (_________________0___18607), .Q (_____0__20857));
  or2s1 _____0_449752(.DIN1 (__________________0___18628), .DIN2
       (________20390), .Q (___0_0__21696));
  nor2s1 _____0_449753(.DIN1 (_____0__20392), .DIN2 (________20390), .Q
       (________21378));
  nor2s1 _____0_449754(.DIN1 (_____0___33866), .DIN2 (___9____19751),
       .Q (_____9__20912));
  and2s1 ____99_449755(.DIN1 (___0____19813), .DIN2
       (_____________________18601), .Q (_____9__20856));
  nor2s1 _______449756(.DIN1 (___0____21699), .DIN2 (________20199), .Q
       (________20957));
  nor2s1 ______449757(.DIN1 (____9___19203), .DIN2 (________19962), .Q
       (_________33817));
  nor2s1 _______449758(.DIN1 (___0_9__19844), .DIN2 (___0____19824), .Q
       (_________33186));
  or2s1 ____9__449759(.DIN1 (________20311), .DIN2 (________20300), .Q
       (_____0__20198));
  and2s1 ____9__449760(.DIN1 (________20196), .DIN2 (___9____21624), .Q
       (_____9__20197));
  nor2s1 ______449761(.DIN1 (________20194), .DIN2 (___99___19766), .Q
       (________20195));
  nnd2s1 _____9_449762(.DIN1 (________20192), .DIN2
       (_________________18695), .Q (________20193));
  nor2s1 _______449763(.DIN1 (________20010), .DIN2 (____9___20883), .Q
       (________20191));
  nor2s1 _______449764(.DIN1 (___9____19728), .DIN2 (____9___20221), .Q
       (________20190));
  or2s1 _______449765(.DIN1 (________20237), .DIN2 (________20470), .Q
       (_____0__20189));
  nnd2s1 _____9_449766(.DIN1 (___0____19827), .DIN2 (________20309), .Q
       (_____9__20188));
  nnd2s1 _____0_449767(.DIN1 (___909), .DIN2 (________19564), .Q
       (________20187));
  or2s1 ______449768(.DIN1 (____0________________18649), .DIN2
       (________19983), .Q (________20186));
  nnd2s1 ______449769(.DIN1 (___9____19748), .DIN2 (________19362), .Q
       (________20185));
  nor2s1 ______449770(.DIN1 (________19556), .DIN2 (___00_), .Q
       (________20184));
  nor2s1 ____9__449771(.DIN1 (________20564), .DIN2 (________20247), .Q
       (________20183));
  hi1s1 _____9_449772(.DIN (________20442), .Q (________20182));
  nnd2s1 _______449773(.DIN1 (________20280), .DIN2 (_____9__20180), .Q
       (_____0__20181));
  nnd2s1 _______449774(.DIN1 (________19626), .DIN2 (___0____19821), .Q
       (________20179));
  nnd2s1 ______449775(.DIN1 (________20177), .DIN2 (_____0__19649), .Q
       (________20178));
  and2s1 ____9_449776(.DIN1 (________20175), .DIN2 (___0_9__20779), .Q
       (________20176));
  hi1s1 _______449777(.DIN (________20173), .Q (________20174));
  nor2s1 ____00_449778(.DIN1 (________19643), .DIN2 (_____9__20341), .Q
       (________20171));
  nnd2s1 _______449779(.DIN1 (________20169), .DIN2 (_____9__19360), .Q
       (________20170));
  and2s1 ____00_449780(.DIN1 (___0_0__21658), .DIN2 (____00__20510), .Q
       (________20168));
  or2s1 ____00_449781(.DIN1 (________20196), .DIN2 (________20872), .Q
       (________20167));
  or2s1 ____0_449782(.DIN1 (________20593), .DIN2 (________20175), .Q
       (________20165));
  nor2s1 _______449783(.DIN1 (________19077), .DIN2 (________20247), .Q
       (_____9__20164));
  nnd2s1 ____99_449784(.DIN1 (________20843), .DIN2 (________21216), .Q
       (________20163));
  or2s1 ______449785(.DIN1 (________19641), .DIN2 (___09___19850), .Q
       (________20162));
  nor2s1 ____9_449786(.DIN1 (________20160), .DIN2 (_____9__20341), .Q
       (________20161));
  nor2s1 ____9__449787(.DIN1 (________20158), .DIN2 (____9___21353), .Q
       (________20159));
  and2s1 _______449788(.DIN1 (___0____21690), .DIN2 (_____0__20156), .Q
       (________20157));
  or2s1 _______449789(.DIN1 (_______19014), .DIN2 (________20154), .Q
       (_____9__20155));
  or2s1 ____99_449790(.DIN1 (________20158), .DIN2 (_____0__21046), .Q
       (________20153));
  nor2s1 ____9_449791(.DIN1 (_____0__20021), .DIN2 (________21226), .Q
       (________20152));
  nnd2s1 _______449792(.DIN1 (___90_), .DIN2 (____0___20330), .Q
       (________20151));
  and2s1 ____9__449793(.DIN1 (________20946), .DIN2 (________21337), .Q
       (________20150));
  nnd2s1 ____9__449794(.DIN1 (___0____19829), .DIN2 (____0___19950), .Q
       (________20149));
  and2s1 ____9__449795(.DIN1 (________21201), .DIN2 (___9____19708), .Q
       (________20148));
  nnd2s1 _______449796(.DIN1 (________21313), .DIN2 (________19066), .Q
       (________20147));
  nnd2s1 ____9__449797(.DIN1 (___0____21677), .DIN2 (________21458), .Q
       (_____0__20146));
  or2s1 _____449798(.DIN1 (________20194), .DIN2 (________22333), .Q
       (____09__20145));
  nnd2s1 ____00_449799(.DIN1 (___9____20684), .DIN2 (____0___20143), .Q
       (____0___20144));
  nnd2s1 ____9__449800(.DIN1 (___0_9__20779), .DIN2 (________19259), .Q
       (____0___20142));
  nor2s1 ____9__449801(.DIN1 (________21180), .DIN2 (___0____20763), .Q
       (____0___20141));
  or2s1 _______449802(.DIN1 (_________30104), .DIN2 (_________30374),
       .Q (____0___20140));
  nor2s1 ____9__449803(.DIN1 (________19919), .DIN2 (________20205), .Q
       (____0___20139));
  nor2s1 ____449804(.DIN1 (________20307), .DIN2 (____9___21353), .Q
       (____0___20138));
  or2s1 _____9_449805(.DIN1 (________19232), .DIN2 (________20280), .Q
       (____0___20137));
  nnd2s1 ____9__449806(.DIN1 (________21774), .DIN2 (________20813), .Q
       (____00__20136));
  nor2s1 _______449807(.DIN1 (________20384), .DIN2 (___9____20656), .Q
       (____99__20135));
  nnd2s1 ____90_449808(.DIN1 (________20461), .DIN2 (___9____19758), .Q
       (____9___20134));
  or2s1 _______449809(.DIN1 (_____________________18624), .DIN2
       (________20390), .Q (____9___20133));
  nnd2s1 ____9__449810(.DIN1 (____90__19677), .DIN2 (___0____19783), .Q
       (____9___20132));
  nnd2s1 ____9__449811(.DIN1 (________22211), .DIN2 (________20380), .Q
       (____9___20131));
  or2s1 ____90_449812(.DIN1 (_____9__21513), .DIN2 (___0____22552), .Q
       (____9___20130));
  nor2s1 ____90_449813(.DIN1 (____9___19493), .DIN2 (________19646), .Q
       (____9___20129));
  nor2s1 _____9_449814(.DIN1 (____9___20219), .DIN2 (____9___21353), .Q
       (____9___20128));
  or2s1 _____449815(.DIN1 (____90__20126), .DIN2 (_____9__20125), .Q
       (____9___20127));
  nor2s1 ____449816(.DIN1 (________20123), .DIN2 (________21276), .Q
       (________20124));
  nnd2s1 _____9_449817(.DIN1 (___900), .DIN2 (inData[14]), .Q
       (________20122));
  nnd2s1 _______449818(.DIN1 (________20120), .DIN2 (outData[13]), .Q
       (________20121));
  nnd2s1 ____0__449819(.DIN1 (____99__19946), .DIN2 (________21115), .Q
       (________20119));
  nor2s1 _____449820(.DIN1 (________20117), .DIN2 (________20347), .Q
       (________20118));
  and2s1 _______449821(.DIN1 (________20192), .DIN2 (_________34478),
       .Q (_____0__20116));
  nor2s1 _______449822(.DIN1 (________19553), .DIN2 (___0_9__19809), .Q
       (_____9__20115));
  nnd2s1 ______449823(.DIN1 (________20201), .DIN2 (_____0__20097), .Q
       (________20114));
  nnd2s1 _______449824(.DIN1 (____0___19951), .DIN2 (____09__19955), .Q
       (________20113));
  nnd2s1 ______449825(.DIN1 (_____0__19639), .DIN2 (________19255), .Q
       (________20112));
  and2s1 _____9_449826(.DIN1 (________20110), .DIN2 (________20109), .Q
       (________20111));
  nor2s1 _______449827(.DIN1 (_______18958), .DIN2 (________20101), .Q
       (________20108));
  nnd2s1 _____0_449828(.DIN1 (_____9__20106), .DIN2 (_____0__19341), .Q
       (_____0__20107));
  and2s1 _____9_449829(.DIN1 (________20809), .DIN2 (________20109), .Q
       (________20105));
  nnd2s1 _______449830(.DIN1 (___0____21680), .DIN2 (____0__18959), .Q
       (________20104));
  or2s1 _______449831(.DIN1 (_____________18900), .DIN2
       (________20154), .Q (________20103));
  nor2s1 _______449832(.DIN1 (____0), .DIN2 (________20101), .Q
       (________20102));
  nnd2s1 _______449833(.DIN1 (___90___19690), .DIN2 (inData[16]), .Q
       (________20100));
  or2s1 _______449834(.DIN1 (_____00__30456), .DIN2 (____9____31759),
       .Q (________20099));
  nnd2s1 _____9_449835(.DIN1 (___9____20657), .DIN2 (_____0__20097), .Q
       (________20098));
  nor2s1 ______449836(.DIN1 (___0____19811), .DIN2 (________21032), .Q
       (_____9__20096));
  nor2s1 ______449837(.DIN1 (_____0__19659), .DIN2 (________20154), .Q
       (________20095));
  nor2s1 _______449838(.DIN1 (________20073), .DIN2 (___0__), .Q
       (________20093));
  nor2s1 _______449839(.DIN1 (________20091), .DIN2 (___0____19801), .Q
       (________20092));
  nnd2s1 _______449840(.DIN1 (___0_0__19826), .DIN2 (________19527), .Q
       (________20090));
  nor2s1 _______449841(.DIN1 (________22050), .DIN2 (________19666), .Q
       (________20089));
  hi1s1 ______449842(.DIN (_____9__20087), .Q (_____0__20088));
  hi1s1 _______449843(.DIN (________20085), .Q (________20086));
  nor2s1 ____0__449844(.DIN1 (________20084), .DIN2 (________20278), .Q
       (___9____20658));
  hi1s1 _______449845(.DIN (________21054), .Q (___9____20648));
  hi1s1 _____9_449846(.DIN (________20375), .Q (___9____20664));
  hi1s1 _______449847(.DIN (____0_9__33692), .Q (___0____20773));
  hi1s1 _____0_449848(.DIN (____9___20507), .Q (___0_9__20761));
  hi1s1 _______449849(.DIN (________20525), .Q (____0___20983));
  nor2s1 ____0__449850(.DIN1 (________20072), .DIN2 (_____9__20341), .Q
       (___00___20704));
  hi1s1 _____449851(.DIN (________20394), .Q (________20852));
  hi1s1 _____449852(.DIN (________20555), .Q (___9____20652));
  and2s1 ______449853(.DIN1 (____0___20143), .DIN2 (________20241), .Q
       (________20819));
  and2s1 ____0__449854(.DIN1 (________20872), .DIN2 (________21480), .Q
       (________20828));
  nor2s1 ____0__449855(.DIN1 (________20083), .DIN2 (________22113), .Q
       (________20446));
  nnd2s1 ____0__449856(.DIN1 (________20082), .DIN2
       (_________________0___18607), .Q (________20444));
  nnd2s1 _______449857(.DIN1 (________20081), .DIN2
       (_____________________18601), .Q (____9___20506));
  or2s1 _______449858(.DIN1 (_____________________18619), .DIN2
       (________20080), .Q (________20823));
  and2s1 _______449859(.DIN1 (___9_9__19744), .DIN2 (_____0__20079), .Q
       (___0____20727));
  nor2s1 ____0__449860(.DIN1 (____0________________18592), .DIN2
       (________20286), .Q (___9____20667));
  nnd2s1 ______449861(.DIN1 (___0____19819), .DIN2 (_____9__20078), .Q
       (________20949));
  hi1s1 _______449862(.DIN (___90___20606), .Q (___9____20650));
  and2s1 _______449863(.DIN1 (________20210), .DIN2 (____9___19589), .Q
       (_____0__20837));
  hi1s1 _____9_449864(.DIN (_____9__20548), .Q (_____9__21009));
  nor2s1 _______449865(.DIN1 (___9__18934), .DIN2 (________20386), .Q
       (________20379));
  nnd2s1 ____9__449866(.DIN1 (________20077), .DIN2 (____0___20143), .Q
       (____0___20425));
  nor2s1 _______449867(.DIN1 (________19374), .DIN2 (_____9__19630), .Q
       (________20855));
  nor2s1 _____449868(.DIN1 (_________35106), .DIN2 (____9___20504), .Q
       (________20834));
  nor2s1 ____0__449869(.DIN1 (____0___21080), .DIN2 (________21505), .Q
       (____0___20988));
  and2s1 ____0_449870(.DIN1 (________20076), .DIN2 (________21480), .Q
       (________20838));
  nnd2s1 _______449871(.DIN1 (________20075), .DIN2
       (__________________0___18628), .Q (___0____20734));
  nor2s1 _____9_449872(.DIN1 (_____0___33866), .DIN2 (________20825),
       .Q (________20835));
  nnd2s1 _____0_449873(.DIN1 (________20074), .DIN2 (_________35106),
       .Q (________20920));
  or2s1 ____0__449874(.DIN1 (________20073), .DIN2 (________20405), .Q
       (___0____20731));
  and2s1 ____0__449875(.DIN1 (________20338), .DIN2 (________20072), .Q
       (________21890));
  hi1s1 _______449876(.DIN (________20071), .Q (________20954));
  and2s1 ______449877(.DIN1 (________20380), .DIN2 (________20109), .Q
       (________20851));
  nor2s1 ____0__449878(.DIN1 (____0___19209), .DIN2 (_____9__20125), .Q
       (________20914));
  hi1s1 _______449879(.DIN (____0___20512), .Q (________20844));
  hi1s1 _______449880(.DIN (________21050), .Q (________21153));
  nnd2s1 ____99_449881(.DIN1 (___0_9__19802), .DIN2 (_____9__20932), .Q
       (___9____20646));
  xor2s1 ____0__449882(.DIN1 (________35107), .DIN2 (___09), .Q
       (________21039));
  nor2s1 ____9__449883(.DIN1 (____9___19587), .DIN2 (____9___19681), .Q
       (_____0__20923));
  and2s1 ____0__449884(.DIN1 (________20872), .DIN2 (___99___20695), .Q
       (_____0__20827));
  nnd2s1 ____0__449885(.DIN1 (___9____19753), .DIN2 (_____9__20313), .Q
       (_____9__22435));
  nor2s1 ____0__449886(.DIN1 (____00__19947), .DIN2 (________20821), .Q
       (___9_0__20654));
  or2s1 ____0__449887(.DIN1 (____9___20219), .DIN2 (___90___20608), .Q
       (___9____20647));
  nnd2s1 ____0_449888(.DIN1 (________20809), .DIN2 (________20070), .Q
       (___9____20660));
  nor2s1 ____0__449889(.DIN1 (_________35105), .DIN2 (________20247),
       .Q (___0____20716));
  nnd2s1 _______449890(.DIN1 (________19907), .DIN2 (_____0__22063), .Q
       (________20853));
  nor2s1 _______449891(.DIN1 (___0_9__19834), .DIN2 (___90___19689), .Q
       (________21510));
  nnd2s1 ______449892(.DIN1 (________20205), .DIN2 (_____0__20069), .Q
       (_____9__21522));
  nor2s1 _______449893(.DIN1 (__________________0___18628), .DIN2
       (________20067), .Q (____9___21803));
  nnd2s1 _______449894(.DIN1 (________20075), .DIN2 (_____0__20392), .Q
       (________21014));
  nor2s1 ______449895(.DIN1 (________19386), .DIN2 (___00___19773), .Q
       (________20839));
  nnd2s1 _______449896(.DIN1 (___99___19770), .DIN2 (________19381), .Q
       (_____9___30173));
  nnd2s1 ____9__449897(.DIN1 (_____9__20068), .DIN2
       (____0____________0_), .Q (_____0__20847));
  hi1s1 _______449898(.DIN (________21234), .Q (________21053));
  nor2s1 ____0__449899(.DIN1 (________19634), .DIN2 (___9____20665), .Q
       (___9____20661));
  nnd2s1 ____09_449900(.DIN1 (________20802), .DIN2 (____9___19200), .Q
       (___9____20655));
  nnd2s1 ____0__449901(.DIN1 (____0___20423), .DIN2 (____9___21897), .Q
       (________20993));
  nor2s1 ______449902(.DIN1 (___0____19782), .DIN2 (____90__19196), .Q
       (________20858));
  nor2s1 _______449903(.DIN1 (___0____19797), .DIN2 (________21397), .Q
       (_________31376));
  nor2s1 _______449904(.DIN1 (________19076), .DIN2 (________21313), .Q
       (________20897));
  nor2s1 _____0_449905(.DIN1 (___9____19723), .DIN2 (________20064), .Q
       (___9____20659));
  hi1s1 _______449906(.DIN (________20570), .Q (________21060));
  nor2s1 _______449907(.DIN1 (_____0__20392), .DIN2 (________20067), .Q
       (____0___21361));
  hi1s1 _______449908(.DIN (____9___20597), .Q (_________31047));
  hi1s1 ______449909(.DIN (_________32919), .Q (_________32407));
  nor2s1 ____09_449910(.DIN1 (___9____19749), .DIN2 (________20203), .Q
       (___09___20785));
  nnd2s1 ______449911(.DIN1 (________20066), .DIN2 (_____0__20069), .Q
       (________20998));
  nor2s1 _______449912(.DIN1 (________19181), .DIN2 (________20065), .Q
       (_____99__29264));
  nnd2s1 _______449913(.DIN1 (________19640), .DIN2 (______18933), .Q
       (____0___21363));
  hi1s1 _______449914(.DIN (________20532), .Q (________21372));
  nor2s1 ______449915(.DIN1 (________19470), .DIN2 (________20064), .Q
       (___9_9__20653));
  nor2s1 _______449916(.DIN1 (_____0__19170), .DIN2 (________20063), .Q
       (______0__32594));
  nor2s1 _______449917(.DIN1 (________19348), .DIN2 (________20965), .Q
       (_________33895));
  nor2s1 _______449918(.DIN1 (_____0__20069), .DIN2 (________20286), .Q
       (____9___21808));
  and2s1 _______449919(.DIN1 (________21226), .DIN2
       (_________________0___18633), .Q (________20937));
  nor2s1 _______449920(.DIN1 (________19610), .DIN2 (___0____19806), .Q
       (________20848));
  nnd2s1 ____0_449921(.DIN1 (___9____19730), .DIN2
       (_____________________18600), .Q (_________31505));
  hi1s1 _______449922(.DIN (________20062), .Q (________21373));
  hi1s1 _______449923(.DIN (________20061), .Q (______9__32927));
  hi1s1 ______449924(.DIN (_____0__21335), .Q (________20060));
  or2s1 ____9__449925(.DIN1 (________19168), .DIN2 (_____0__20362), .Q
       (_____0__20059));
  or2s1 ____9_449926(.DIN1 (________20057), .DIN2 (________20850), .Q
       (_____9__20058));
  nnd2s1 ____9__449927(.DIN1 (____0___20041), .DIN2 (___9____19733), .Q
       (________20056));
  nor2s1 ____9__449928(.DIN1 (________19090), .DIN2 (________20023), .Q
       (________20055));
  nnd2s1 _____0_449929(.DIN1 (________20053), .DIN2 (_____9__19169), .Q
       (________20054));
  nnd2s1 _______449930(.DIN1 (________19373), .DIN2 (___0___19042), .Q
       (________20052));
  and2s1 _____0_449931(.DIN1 (________19546), .DIN2
       (_____________________18662), .Q (________20051));
  nnd2s1 _____9_449932(.DIN1 (____0____29098), .DIN2 (_____0__20049),
       .Q (________20050));
  or2s1 _______449933(.DIN1 (_____________________18625), .DIN2
       (________19375), .Q (____09__20048));
  nor2s1 ____90_449934(.DIN1 (____90__19196), .DIN2 (____0___20046), .Q
       (____0___20047));
  nnd2s1 ____9__449935(.DIN1 (________19508), .DIN2
       (__________________0___18628), .Q (____0___20045));
  nnd2s1 _______449936(.DIN1 (________19249), .DIN2 (____0___19952), .Q
       (____0___20044));
  nnd2s1 ______449937(.DIN1 (________21222), .DIN2 (___9_0__20644), .Q
       (____0___20043));
  nnd2s1 ____9__449938(.DIN1 (____0___20041), .DIN2 (________19513), .Q
       (____0___20042));
  nnd2s1 _______449939(.DIN1 (_____0__19312), .DIN2 (inData[30]), .Q
       (____00__20040));
  nnd2s1 _______449940(.DIN1 (_____9__19486), .DIN2 (inData[28]), .Q
       (____99__20039));
  nor2s1 _______449941(.DIN1 (___0____20730), .DIN2 (____9___20037), .Q
       (____9___20038));
  nnd2s1 _______449942(.DIN1 (____0___20046), .DIN2 (_________31041),
       .Q (____9___20036));
  or2s1 _______449943(.DIN1 (___9____20625), .DIN2 (____9___19583), .Q
       (____9___20035));
  nor2s1 _______449944(.DIN1 (________19996), .DIN2 (____9___22438), .Q
       (____9___20034));
  nnd2s1 _______449945(.DIN1 (________19368), .DIN2 (________19179), .Q
       (____9___20033));
  and2s1 _______449946(.DIN1 (_________33370), .DIN2 (_____0__19134),
       .Q (____9___20032));
  nnd2s1 _______449947(.DIN1 (___0____19796), .DIN2 (________19326), .Q
       (____90__20031));
  and2s1 _______449948(.DIN1 (____0___19498), .DIN2
       (____0________________18592), .Q (_____9__20030));
  nor2s1 _______449949(.DIN1 (_________________18709), .DIN2
       (________19388), .Q (________20029));
  nor2s1 _______449950(.DIN1 (_____0__22063), .DIN2 (________20027), .Q
       (________20028));
  nnd2s1 _______449951(.DIN1 (____90__19487), .DIN2 (________19558), .Q
       (________20026));
  nnd2s1 _______449952(.DIN1 (________19554), .DIN2 (________19569), .Q
       (________20025));
  nor2s1 _____9_449953(.DIN1 (_________________18713), .DIN2
       (________20023), .Q (________20024));
  nor2s1 _______449954(.DIN1 (____0___19407), .DIN2 (_____0__20021), .Q
       (________20022));
  nor2s1 _____0_449955(.DIN1 (_________18852), .DIN2 (________20019),
       .Q (_____9__20020));
  nnd2s1 _____9_449956(.DIN1 (_____9__19458), .DIN2 (_____9__19370), .Q
       (________20018));
  nnd2s1 _____449957(.DIN1 (____0___20041), .DIN2
       (_____________________18623), .Q (________20017));
  nnd2s1 _______449958(.DIN1 (________19235), .DIN2 (________19473), .Q
       (________20016));
  nor2s1 _______449959(.DIN1 (_____0__19872), .DIN2 (________19902), .Q
       (________20015));
  or2s1 _______449960(.DIN1 (______________________18632), .DIN2
       (____9___19938), .Q (________20014));
  nor2s1 _______449961(.DIN1 (______________0___________________),
       .DIN2 (________19537), .Q (________20013));
  or2s1 _______449962(.DIN1 (_____9__20011), .DIN2 (________20010), .Q
       (_____0__20012));
  nnd2s1 _______449963(.DIN1 (________21518), .DIN2 (____0___21267), .Q
       (________20009));
  nor2s1 ____9__449964(.DIN1 (________20007), .DIN2 (________19864), .Q
       (________20008));
  nnd2s1 ____9__449965(.DIN1 (________21797), .DIN2 (________19338), .Q
       (________20006));
  nor2s1 _______449966(.DIN1 (________19334), .DIN2 (________20027), .Q
       (________20005));
  and2s1 ____9_449967(.DIN1 (________20003), .DIN2 (_____0__20002), .Q
       (________20004));
  nor2s1 ____9__449968(.DIN1 (________19655), .DIN2 (________20003), .Q
       (_____9__20001));
  nor2s1 _______449969(.DIN1 (________19999), .DIN2 (___9____19709), .Q
       (________20000));
  hi1s1 _______449970(.DIN (________20384), .Q (________19998));
  nnd2s1 _______449971(.DIN1 (________19344), .DIN2 (________19996), .Q
       (________19997));
  or2s1 _______449972(.DIN1 (_____________________18667), .DIN2
       (____9___20037), .Q (________19995));
  nnd2s1 _______449973(.DIN1 (________19915), .DIN2 (_____0__22063), .Q
       (________19994));
  nor2s1 _______449974(.DIN1 (________19167), .DIN2 (_____0__20362), .Q
       (________19993));
  or2s1 ____9__449975(.DIN1 (_____9__19991), .DIN2 (______9__28887), .Q
       (_____0__19992));
  or2s1 ____9__449976(.DIN1 (_____0__19086), .DIN2 (_____0__20362), .Q
       (________19990));
  nor2s1 _______449977(.DIN1 (____0________________18649), .DIN2
       (_____9__19330), .Q (________19989));
  and2s1 _______449978(.DIN1 (________19963), .DIN2 (_____9__20313), .Q
       (________19988));
  nnd2s1 _______449979(.DIN1 (______9__33436), .DIN2 (____0___19499),
       .Q (________19987));
  hi1s1 _______449980(.DIN (________19983), .Q (_____9__19984));
  hi1s1 _______449981(.DIN (________20064), .Q (________19982));
  nnd2s1 ______449982(.DIN1 (________19314), .DIN2 (_____0__20069), .Q
       (________19981));
  or2s1 ____9__449983(.DIN1 (____0___19954), .DIN2 (________20461), .Q
       (________19980));
  nnd2s1 ____9__449984(.DIN1 (_____0__22118), .DIN2 (________19978), .Q
       (________19979));
  nnd2s1 ____9__449985(.DIN1 (________19976), .DIN2 (_____0__19975), .Q
       (________19977));
  or2s1 _______449986(.DIN1 (____0________________18649), .DIN2
       (________20010), .Q (________19973));
  nnd2s1 _______449987(.DIN1 (_____0__21191), .DIN2 (___0____19787), .Q
       (________19972));
  nor2s1 _____9_449988(.DIN1 (____9___21898), .DIN2 (___9____19704), .Q
       (________19971));
  nor2s1 ______449989(.DIN1 (________19382), .DIN2 (________19349), .Q
       (________19970));
  and2s1 _______449990(.DIN1 (______9__33436), .DIN2 (________19359),
       .Q (________19969));
  nor2s1 ____9__449991(.DIN1 (_____0__20002), .DIN2 (________20010), .Q
       (________19968));
  hi1s1 _______449992(.DIN (________19967), .Q (____0___20513));
  nnd2s1 ____0__449993(.DIN1 (_____0__19966), .DIN2 (________19958), .Q
       (___9_0__20634));
  hi1s1 _____9_449994(.DIN (________21506), .Q (________20467));
  xor2s1 ____0__449995(.DIN1 (_________________0___18633), .DIN2
       (________19125), .Q (________20094));
  or2s1 _______449996(.DIN1 (_____________________18599), .DIN2
       (_____9__19965), .Q (________20377));
  and2s1 ______449997(.DIN1 (____0___19949), .DIN2 (________21797), .Q
       (________21127));
  nor2s1 ____0_449998(.DIN1 (________19959), .DIN2 (________19964), .Q
       (________20250));
  hi1s1 _______449999(.DIN (________20353), .Q (________20388));
  nnd2s1 _______450000(.DIN1 (________19963), .DIN2
       (____0________________18651), .Q (________20574));
  hi1s1 ______450001(.DIN (_____9__21344), .Q (________20383));
  hi1s1 ______450002(.DIN (________20561), .Q (_____0__20866));
  nnd2s1 _______450003(.DIN1 (___09_), .DIN2 (________19961), .Q
       (________20546));
  nnd2s1 _______450004(.DIN1 (________20003), .DIN2 (_____9__20011), .Q
       (_____9__20575));
  nnd2s1 _______450005(.DIN1 (_____9__19533), .DIN2 (________19327), .Q
       (____0___20328));
  nnd2s1 ____0__450006(.DIN1 (________19963), .DIN2 (________20072), .Q
       (____90__20217));
  hi1s1 _______450007(.DIN (________20177), .Q (________20378));
  nnd2s1 ____0_450008(.DIN1 (______9__28887), .DIN2 (_____9__19991), .Q
       (________20583));
  nnd2s1 _______450009(.DIN1 (___9_9__20623), .DIN2
       (____0______________), .Q (________20166));
  nor2s1 ____0__450010(.DIN1 (___0____19843), .DIN2 (________19960), .Q
       (________20085));
  nnd2s1 ____0__450011(.DIN1 (___0____21677), .DIN2 (________22332), .Q
       (_____9__20172));
  nnd2s1 _______450012(.DIN1 (________19335), .DIN2
       (_____________________18665), .Q (_____0__20520));
  and2s1 ____0_450013(.DIN1 (________19964), .DIN2 (________19959), .Q
       (________20587));
  hi1s1 _____0_450014(.DIN (____90__21801), .Q (_____9__21772));
  nor2s1 ____0__450015(.DIN1 (____9____30882), .DIN2 (___9____20656),
       .Q (________20396));
  or2s1 ____0__450016(.DIN1 (________19958), .DIN2 (_____0__19966), .Q
       (___9____20635));
  hi1s1 _______450017(.DIN (________20307), .Q (_____9__20401));
  hi1s1 _______450018(.DIN (________20242), .Q (____00__20420));
  hi1s1 _____0_450019(.DIN (____0___21362), .Q (___00___20703));
  hi1s1 _____450020(.DIN (________21887), .Q (________21778));
  hi1s1 _______450021(.DIN (________21488), .Q (________21218));
  nor2s1 ____09_450022(.DIN1 (___9____21575), .DIN2 (___9____20651), .Q
       (________20394));
  nor2s1 ____0__450023(.DIN1 (_____0___33866), .DIN2 (________19957),
       .Q (____0___20511));
  nnd2s1 ____0__450024(.DIN1 (_________28828), .DIN2 (_____0__19477),
       .Q (________20375));
  nor2s1 ____0__450025(.DIN1 (___9_9__20681), .DIN2 (___9____19705), .Q
       (________20544));
  nnd2s1 ____0__450026(.DIN1 (________19893), .DIN2 (_____0__19956), .Q
       (____0___20426));
  nnd2s1 ____0__450027(.DIN1 (___9____20684), .DIN2 (________21893), .Q
       (___9____20632));
  nnd2s1 _____9_450028(.DIN1 (____09__19955), .DIN2
       (____0____________0_), .Q (________20845));
  and2s1 ____0_450029(.DIN1 (________21006), .DIN2 (___9____21624), .Q
       (___9____20668));
  nor2s1 _______450030(.DIN1 (_________35105), .DIN2 (________20461),
       .Q (________20570));
  nnd2s1 ____0__450031(.DIN1 (_____0__20021), .DIN2 (___9__18934), .Q
       (____0___20518));
  hi1s1 ______450032(.DIN (________20405), .Q (_____0__20474));
  hi1s1 _____0_450033(.DIN (_____9__20341), .Q (________22227));
  nnd2s1 _______450034(.DIN1 (________20497), .DIN2
       (____0____________0_), .Q (________20522));
  or2s1 ____0_450035(.DIN1 (________21197), .DIN2 (___9____20666), .Q
       (____9___20505));
  nor2s1 _______450036(.DIN1 (____0_________________18659), .DIN2
       (________19550), .Q (___90___20606));
  nnd2s1 ____450037(.DIN1 (_____0__20021), .DIN2
       (_________________0___18633), .Q (____9___20507));
  nnd2s1 _______450038(.DIN1 (_________28828), .DIN2 (____90__19390),
       .Q (____9___20502));
  or2s1 _____0_450039(.DIN1 (________20534), .DIN2 (____0___19954), .Q
       (___9____20628));
  nor2s1 ____09_450040(.DIN1 (___9____21575), .DIN2 (____0___19953), .Q
       (________20555));
  or2s1 _______450041(.DIN1 (_________________0___18633), .DIN2
       (________20534), .Q (________20538));
  nor2s1 ____09_450042(.DIN1 (____0________________18592), .DIN2
       (____0___19952), .Q (________20482));
  hi1s1 _______450043(.DIN (____0___19951), .Q (___0____21692));
  nor2s1 _______450044(.DIN1 (_____0__20392), .DIN2 (____0___19950), .Q
       (________21050));
  nnd2s1 _______450045(.DIN1 (____0___19949), .DIN2 (_____0__20392), .Q
       (____0___21357));
  nor2s1 ____0__450046(.DIN1 (_________________0___18607), .DIN2
       (________19323), .Q (________20442));
  hi1s1 _______450047(.DIN (_____0__19985), .Q (________19986));
  nor2s1 _______450048(.DIN1 (____0_________________18596), .DIN2
       (____0___19948), .Q (________21530));
  or2s1 _____0_450049(.DIN1 (_________________0___18633), .DIN2
       (____09__20519), .Q (____0___20515));
  hi1s1 _______450050(.DIN (____00__19947), .Q (________21387));
  hi1s1 _____9_450051(.DIN (____99__19946), .Q (________22000));
  nor2s1 _______450052(.DIN1 (_____9__19543), .DIN2 (________19567), .Q
       (_____9___33022));
  hi1s1 _____450053(.DIN (________21381), .Q (___9____21592));
  hi1s1 _______450054(.DIN (________21509), .Q (________21508));
  hi1s1 _____450055(.DIN (________21233), .Q (________21978));
  nnd2s1 _______450056(.DIN1 (________19333), .DIN2 (____0___19119), .Q
       (____0_9__33692));
  and2s1 _______450057(.DIN1 (____0___19949), .DIN2
       (__________________0___18628), .Q (___0____21698));
  hi1s1 _______450058(.DIN (____9___19944), .Q (____0___21905));
  hi1s1 _______450059(.DIN (____9___19945), .Q (____09__22634));
  nnd2s1 _______450060(.DIN1 (____9___19492), .DIN2 (________19566), .Q
       (_________30693));
  nnd2s1 _______450061(.DIN1 (_____9__20557), .DIN2 (____9___19489), .Q
       (_________31154));
  nor2s1 _______450062(.DIN1 (________19140), .DIN2 (___0_9__19817), .Q
       (____0____32762));
  nor2s1 _______450063(.DIN1 (________21492), .DIN2 (___9____19724), .Q
       (____9___19943));
  nor2s1 _____0_450064(.DIN1 (___900__20605), .DIN2 (________19538), .Q
       (____9___19942));
  and2s1 _______450065(.DIN1 (____9___19940), .DIN2 (______18940), .Q
       (____9___19941));
  or2s1 _______450066(.DIN1 (______________________18631), .DIN2
       (____9___19938), .Q (____9___19939));
  nnd2s1 ____9__450067(.DIN1 (________21216), .DIN2 (___9____19703), .Q
       (____90__19937));
  nor2s1 _______450068(.DIN1 (________21492), .DIN2 (________20261), .Q
       (_____9__19936));
  nnd2s1 ____90_450069(.DIN1 (________20917), .DIN2 (___0____21694), .Q
       (________19935));
  nor2s1 ______450070(.DIN1 (____9___19490), .DIN2 (________19316), .Q
       (________19934));
  nor2s1 ____90_450071(.DIN1 (_____________________18665), .DIN2
       (________19532), .Q (________19933));
  nnd2s1 _____9_450072(.DIN1 (________19482), .DIN2 (____9___19111), .Q
       (________19932));
  hi1s1 _____9_450073(.DIN (________20390), .Q (________19931));
  nnd2s1 _______450074(.DIN1 (________19244), .DIN2 (________19874), .Q
       (________19930));
  nor2s1 _______450075(.DIN1 (_________28581), .DIN2 (___0____19804),
       .Q (________19929));
  nor2s1 ______450076(.DIN1 (________19065), .DIN2 (_____0__20362), .Q
       (________19928));
  nor2s1 _____0_450077(.DIN1 (________19246), .DIN2 (_____9__19926), .Q
       (_____0__19927));
  or2s1 _______450078(.DIN1 (_____________________18666), .DIN2
       (________20027), .Q (________19925));
  nnd2s1 ____450079(.DIN1 (____9___19587), .DIN2 (________19365), .Q
       (________19924));
  and2s1 ____9__450080(.DIN1 (______0__30345), .DIN2 (________19922),
       .Q (________19923));
  nor2s1 ____9__450081(.DIN1 (________19510), .DIN2 (____9___19940), .Q
       (________19921));
  or2s1 ____99_450082(.DIN1 (________19919), .DIN2 (_____0__19918), .Q
       (________19920));
  nor2s1 ____99_450083(.DIN1 (________20073), .DIN2 (____9___20037), .Q
       (_____9__19917));
  nnd2s1 _______450084(.DIN1 (________19915), .DIN2
       (_____________________18666), .Q (________19916));
  nnd2s1 ____9__450085(.DIN1 (________19913), .DIN2 (________19528), .Q
       (________19914));
  and2s1 _______450086(.DIN1 (________19911), .DIN2
       (_____________________18638), .Q (________19912));
  nnd2s1 ____9__450087(.DIN1 (_____0__21504), .DIN2 (________21774), .Q
       (________19910));
  nnd2s1 _______450088(.DIN1 (________19318), .DIN2 (_____9__19908), .Q
       (_____0__19909));
  nnd2s1 _______450089(.DIN1 (________20209), .DIN2 (________19905), .Q
       (________19906));
  nor2s1 _______450090(.DIN1 (___0__18943), .DIN2 (____0___20514), .Q
       (________19904));
  and2s1 ____9_450091(.DIN1 (________19902), .DIN2 (___9____19710), .Q
       (________19903));
  nor2s1 _______450092(.DIN1 (____0__18967), .DIN2 (________20019), .Q
       (________19901));
  nnd2s1 _______450093(.DIN1 (________19352), .DIN2 (________19217), .Q
       (_____9__19900));
  nnd2s1 _______450094(.DIN1 (________19875), .DIN2 (________19898), .Q
       (________19899));
  nor2s1 ____9__450095(.DIN1 (________19922), .DIN2 (______0__30345),
       .Q (________19897));
  or2s1 ____9_450096(.DIN1 (___9____20666), .DIN2 (_____9__20557), .Q
       (________19896));
  or2s1 _______450097(.DIN1 (________19377), .DIN2 (_____0__19321), .Q
       (________19895));
  or2s1 ____9__450098(.DIN1 (_____9__19891), .DIN2 (________19893), .Q
       (________19894));
  or2s1 ____9_450099(.DIN1 (_____9__19891), .DIN2 (________20010), .Q
       (_____0__19892));
  nnd2s1 _____0_450100(.DIN1 (_____9__19320), .DIN2 (inData[2]), .Q
       (________19890));
  nnd2s1 _______450101(.DIN1 (________20053), .DIN2 (________19464), .Q
       (________19889));
  or2s1 _______450102(.DIN1 (_____0__20392), .DIN2 (_____9__19524), .Q
       (________19888));
  and2s1 ______450103(.DIN1 (________19886), .DIN2 (________21784), .Q
       (________19887));
  and2s1 _____9_450104(.DIN1 (___0____21677), .DIN2 (________19884), .Q
       (________19885));
  nor2s1 _______450105(.DIN1 (________19328), .DIN2 (_____9__19581), .Q
       (________19883));
  or2s1 _____9_450106(.DIN1 (_____9__19881), .DIN2 (_________30710), .Q
       (_____0__19882));
  nnd2s1 _____9_450107(.DIN1 (___0____21677), .DIN2 (________19879), .Q
       (________19880));
  nnd2s1 _____9_450108(.DIN1 (________19542), .DIN2 (________19070), .Q
       (________19878));
  or2s1 _____9_450109(.DIN1 (________21003), .DIN2 (____0___19598), .Q
       (________19877));
  nnd2s1 _______450110(.DIN1 (________19875), .DIN2 (________19874), .Q
       (________19876));
  nnd2s1 ______450111(.DIN1 (________19915), .DIN2 (_____0__19872), .Q
       (________19873));
  nnd2s1 _______450112(.DIN1 (_____0__19552), .DIN2 (_________28581),
       .Q (_____9__19871));
  nnd2s1 ______450113(.DIN1 (________19539), .DIN2 (________19185), .Q
       (________19870));
  xor2s1 ____09_450114(.DIN1 (________19192), .DIN2 (_______18951), .Q
       (________19869));
  nor2s1 _____0_450115(.DIN1 (________19332), .DIN2 (________19357), .Q
       (________19868));
  hi1s1 _______450116(.DIN (________19866), .Q (________19867));
  nor2s1 _______450117(.DIN1 (___9_9__19706), .DIN2 (________19864), .Q
       (________19865));
  or2s1 ______450118(.DIN1 (________19624), .DIN2 (____0___19953), .Q
       (________19863));
  nnd2s1 _____9_450119(.DIN1 (___0____19838), .DIN2
       (____0________________18591), .Q (_____0__19862));
  nor2s1 _____0_450120(.DIN1 (____0___19860), .DIN2 (____9___19938), .Q
       (____09__19861));
  nor2s1 _______450121(.DIN1 (___0____19800), .DIN2 (___09___19846), .Q
       (____0___19859));
  nnd2s1 _______450122(.DIN1 (________19346), .DIN2 (________19166), .Q
       (____0___19858));
  and2s1 _______450123(.DIN1 (________21216), .DIN2 (________20355), .Q
       (____0___19857));
  nnd2s1 ______450124(.DIN1 (________21306), .DIN2 (________19893), .Q
       (____0___19856));
  and2s1 _______450125(.DIN1 (________20003), .DIN2
       (____0________________18649), .Q (____0___19855));
  nnd2s1 _____450126(.DIN1 (________19915), .DIN2
       (_____________________18668), .Q (____0___19854));
  or2s1 ______450127(.DIN1 (____00__19852), .DIN2 (___9____19742), .Q
       (____0___19853));
  xor2s1 ____0__450128(.DIN1 (_________28979), .DIN2 (___9___19030), .Q
       (___099));
  or2s1 _____450129(.DIN1 (____0___19503), .DIN2 (___09___19850), .Q
       (___09___19851));
  nnd2s1 _______450130(.DIN1 (___09___19848), .DIN2 (________19324), .Q
       (___09___19849));
  nor2s1 ______450131(.DIN1 (________19445), .DIN2 (___09___19846), .Q
       (___09___19847));
  or2s1 _______450132(.DIN1 (________19961), .DIN2 (___09_), .Q
       (___09___19845));
  or2s1 ____9__450133(.DIN1 (___99___19765), .DIN2 (____9___19940), .Q
       (___090));
  nor2s1 ______450134(.DIN1 (___0_9__19844), .DIN2 (_________33370), .Q
       (________20061));
  and2s1 ____0__450135(.DIN1 (________19960), .DIN2 (___0____19843), .Q
       (________20551));
  or2s1 ____0_450136(.DIN1 (___0____19842), .DIN2 (___90___20608), .Q
       (____9___20508));
  hi1s1 ______450137(.DIN (________20257), .Q (________20376));
  hi1s1 _______450138(.DIN (_____9__21019), .Q (___0____21664));
  or2s1 ____0__450139(.DIN1 (________21409), .DIN2 (________21086), .Q
       (________20830));
  nor2s1 ____0__450140(.DIN1 (___0__18931), .DIN2 (________19313), .Q
       (_____9__20087));
  xor2s1 ____0__450141(.DIN1 (____90__19196), .DIN2 (______9__28578),
       .Q (________22920));
  nor2s1 _______450142(.DIN1 (___0____19839), .DIN2 (___0____19841), .Q
       (____0___20893));
  nor2s1 _______450143(.DIN1 (____0________________18648), .DIN2
       (___9____19725), .Q (________20214));
  hi1s1 _____9_450144(.DIN (___0____20763), .Q (________21461));
  nnd2s1 _______450145(.DIN1 (___0____19840), .DIN2 (___0____19780), .Q
       (________20408));
  hi1s1 _______450146(.DIN (________21032), .Q (________21188));
  nnd2s1 _______450147(.DIN1 (____0___20041), .DIN2
       (__________________0___18628), .Q (________20062));
  nor2s1 ______450148(.DIN1 (_____0__20069), .DIN2 (________19474), .Q
       (________22039));
  hi1s1 ______450149(.DIN (________20120), .Q (____9___20417));
  nnd2s1 ______450150(.DIN1 (_____9__20283), .DIN2 (________19559), .Q
       (____90__20500));
  hi1s1 _______450151(.DIN (________21333), .Q (________20403));
  and2s1 _______450152(.DIN1 (___9_9__19726), .DIN2 (____90__20410), .Q
       (________20566));
  nnd2s1 _____0_450153(.DIN1 (_________30710), .DIN2 (_____9__19881),
       .Q (________20580));
  nor2s1 _______450154(.DIN1 (__________________0___18628), .DIN2
       (________19485), .Q (_____9__22042));
  nor2s1 _____0_450155(.DIN1 (_____9__20491), .DIN2 (___9____19725), .Q
       (_____9__20206));
  nnd2s1 _______450156(.DIN1 (___0____19841), .DIN2 (___0____19839), .Q
       (________20173));
  nnd2s1 _____450157(.DIN1 (________19336), .DIN2
       (____0_______________), .Q (________20071));
  and2s1 ____0__450158(.DIN1 (_____0__22118), .DIN2 (________19879), .Q
       (____0___20516));
  nor2s1 _____9_450159(.DIN1 (________22050), .DIN2 (_____0__21191), .Q
       (________21043));
  nor2s1 _____0_450160(.DIN1 (__________________0___18628), .DIN2
       (____0___19950), .Q (________21208));
  nnd2s1 _____0_450161(.DIN1 (___0____19838), .DIN2
       (____0________________18592), .Q (________20525));
  nor2s1 ____0__450162(.DIN1 (_____0__20352), .DIN2 (________21407), .Q
       (____9___20603));
  nor2s1 _____9_450163(.DIN1 (_____0__20382), .DIN2 (________19354), .Q
       (____0___20517));
  hi1s1 _______450164(.DIN (___0____19837), .Q (_________30592));
  hi1s1 _______450165(.DIN (_____0__20156), .Q (________21483));
  nnd2s1 ____0__450166(.DIN1 (____0___20041), .DIN2 (_____0__20392), .Q
       (___9____20617));
  hi1s1 _______450167(.DIN (________21238), .Q (________21501));
  or2s1 ____0__450168(.DIN1 (______18933), .DIN2 (____9___21900), .Q
       (________20469));
  nnd2s1 _______450169(.DIN1 (_____0__19516), .DIN2 (_____0___33866),
       .Q (____0___20512));
  hi1s1 _______450170(.DIN (___0____19836), .Q (____9___20503));
  nnd2s1 ____0_450171(.DIN1 (_____9__22147), .DIN2 (________20204), .Q
       (_____0__20895));
  nnd2s1 _______450172(.DIN1 (_____0__19918), .DIN2
       (____0________________18593), .Q (________20532));
  nor2s1 ____0_450173(.DIN1 (___9____21575), .DIN2 (________21310), .Q
       (_____9__20548));
  hi1s1 _______450174(.DIN (___0____20753), .Q (___0____20748));
  hi1s1 _____0_450175(.DIN (________21388), .Q (________21499));
  nnd2s1 _______450176(.DIN1 (___0_0__19835), .DIN2
       (____0_______________), .Q (________21198));
  nor2s1 _______450177(.DIN1 (___0_9__19834), .DIN2 (________19531), .Q
       (_____0__21365));
  hi1s1 _______450178(.DIN (____9___21804), .Q (________21489));
  nnd2s1 _______450179(.DIN1 (_____0__19918), .DIN2 (________19665), .Q
       (____0___20889));
  hi1s1 _______450180(.DIN (___0____19833), .Q (________20930));
  hi1s1 ______450181(.DIN (___0____19832), .Q (________21206));
  hi1s1 _______450182(.DIN (________20277), .Q (________21385));
  nnd2s1 _______450183(.DIN1 (___0____19831), .DIN2 (____9___19488), .Q
       (________21234));
  nnd2s1 _______450184(.DIN1 (________19465), .DIN2 (____09__19505), .Q
       (_________33989));
  nnd2s1 _______450185(.DIN1 (________19563), .DIN2
       (_____________________18634), .Q (_____9__22679));
  nor2s1 _______450186(.DIN1 (______18933), .DIN2 (________21879), .Q
       (________21098));
  hi1s1 _______450187(.DIN (___0____19830), .Q (______9__33899));
  hi1s1 _______450188(.DIN (_____9__20106), .Q (________20485));
  hi1s1 ______450189(.DIN (___0____19829), .Q (_____9__20464));
  nnd2s1 _______450190(.DIN1 (___0____19838), .DIN2 (_____0__20069), .Q
       (____0___20984));
  or2s1 ____09_450191(.DIN1 (______18933), .DIN2 (________20057), .Q
       (________20832));
  hi1s1 _____0_450192(.DIN (____00__21355), .Q (________21486));
  nor2s1 ______450193(.DIN1 (________19463), .DIN2 (_____9__19965), .Q
       (_____9__21199));
  nnd2s1 _______450194(.DIN1 (___0____19831), .DIN2
       (_________________9___18606), .Q (___9____20615));
  nnd2s1 ______450195(.DIN1 (_________29858), .DIN2 (__99____27118), .Q
       (____9___20597));
  nnd2s1 _______450196(.DIN1 (________19481), .DIN2 (_____0__20392), .Q
       (________21788));
  nnd2s1 ______450197(.DIN1 (____9___20319), .DIN2
       (_____________________18601), .Q (________20829));
  nor2s1 _______450198(.DIN1 (________19223), .DIN2 (________19529), .Q
       (______9__32232));
  nor2s1 ______450199(.DIN1 (________19250), .DIN2 (___0____19840), .Q
       (____9_9__33643));
  hi1s1 _____0_450200(.DIN (________20199), .Q (________21375));
  hi1s1 _______450201(.DIN (________20070), .Q (_____9__21894));
  nnd2s1 _______450202(.DIN1 (________19460), .DIN2 (____9___19396), .Q
       (_________32919));
  nnd2s1 _______450203(.DIN1 (________19911), .DIN2
       (_________________0___18633), .Q (________21054));
  or2s1 _______450204(.DIN1 (_____9__19340), .DIN2 (___0____19828), .Q
       (_________34023));
  hi1s1 ______450205(.DIN (________19520), .Q (____0___23716));
  or2s1 ____9__450206(.DIN1 (___000), .DIN2 (___9____19735), .Q
       (___0____19827));
  nnd2s1 _______450207(.DIN1 (________21241), .DIN2 (___0_9__19825), .Q
       (___0_0__19826));
  nnd2s1 ____9_450208(.DIN1 (_________34295), .DIN2 (___9_0__19707), .Q
       (___0____19824));
  nnd2s1 _______450209(.DIN1 (___0____19822), .DIN2 (________20194), .Q
       (___0____19823));
  or2s1 _______450210(.DIN1 (_____________________18610), .DIN2
       (___9____19693), .Q (___0____19821));
  nnd2s1 ______450211(.DIN1 (_____0___33489), .DIN2
       (_________________18768), .Q (___0____19820));
  or2s1 _______450212(.DIN1 (____0____________9_), .DIN2
       (___9____19691), .Q (___0____19819));
  xor2s1 _______450213(.DIN1 (_____________9___18703), .DIN2
       (___0__18931), .Q (___0____19818));
  nor2s1 _______450214(.DIN1 (________19547), .DIN2 (___0____19815), .Q
       (___0____19816));
  or2s1 _____9_450215(.DIN1 (_____________________18620), .DIN2
       (________19339), .Q (___0____19814));
  and2s1 ____9__450216(.DIN1 (____09__20235), .DIN2 (___0____19805), .Q
       (___0____19813));
  xor2s1 _______450217(.DIN1 (_______19037), .DIN2
       (_____________0___18759), .Q (___0____19812));
  nnd2s1 _______450218(.DIN1 (____0___21812), .DIN2 (___0_0__19810), .Q
       (___0____19811));
  nor2s1 _______450219(.DIN1 (____9___19053), .DIN2 (____9___20413), .Q
       (___0_9__19809));
  nnd2s1 _______450220(.DIN1 (___9____19699), .DIN2 (___0____19807), .Q
       (___0____19808));
  nnd2s1 _____0_450221(.DIN1 (___0____19805), .DIN2 (____9___20599), .Q
       (___0____19806));
  and2s1 _______450222(.DIN1 (____0___20330), .DIN2 (________19511), .Q
       (___0____19803));
  nor2s1 _______450223(.DIN1 (___0____20746), .DIN2 (________20292), .Q
       (___0_9__19802));
  nnd2s1 _______450224(.DIN1 (________19274), .DIN2 (___0____19800), .Q
       (___0____19801));
  xnr2s1 _______450225(.DIN1 (___0____19798), .DIN2
       (_________________18726), .Q (___0____19799));
  hi1s1 _______450226(.DIN (___0____19796), .Q (___0____19797));
  nnd2s1 ______450227(.DIN1 (____0___20330), .DIN2 (_____9__21513), .Q
       (___0____19795));
  nor2s1 _______450228(.DIN1 (_____________________18601), .DIN2
       (___00___19772), .Q (___0____19794));
  nnd2s1 ______450229(.DIN1 (________19220), .DIN2 (inData[20]), .Q
       (___0_0__19793));
  xor2s1 _______450230(.DIN1 (_________________18681), .DIN2
       (___9____19746), .Q (___0____19792));
  nnd2s1 _______450231(.DIN1 (________19173), .DIN2 (inData[22]), .Q
       (___0____19791));
  or2s1 ______450232(.DIN1 (__________________0_), .DIN2
       (___0____19789), .Q (___0____19790));
  nor2s1 ______450233(.DIN1 (___0____19787), .DIN2 (____9___20413), .Q
       (___0____19788));
  nnd2s1 _______450234(.DIN1 (________20213), .DIN2 (___9____19732), .Q
       (___0____19786));
  xor2s1 _______450235(.DIN1 (_______19040), .DIN2
       (_______________0_____________________18830), .Q
       (___0_0__19785));
  nor2s1 _______450236(.DIN1 (_________________9___18616), .DIN2
       (___0____19789), .Q (___0_9));
  and2s1 _______450237(.DIN1 (___0____19783), .DIN2
       (____0________________18651), .Q (___0____19784));
  nnd2s1 ______450238(.DIN1 (___9____19702), .DIN2 (___9____19700), .Q
       (___0____19782));
  nor2s1 _______450239(.DIN1 (___0____19780), .DIN2 (________21468), .Q
       (___0____19781));
  nor2s1 _______450240(.DIN1 (___9____19696), .DIN2 (________19425), .Q
       (___0____19779));
  xor2s1 ____0__450241(.DIN1 (________19135), .DIN2 (________19079), .Q
       (___0____19778));
  and2s1 _______450242(.DIN1 (___0_0), .DIN2 (____9__18949), .Q
       (___0__));
  xor2s1 _______450243(.DIN1 (___________), .DIN2 (___00___19777), .Q
       (___009));
  xnr2s1 _______450244(.DIN1 (_________18851), .DIN2 (___00___19775),
       .Q (___00___19776));
  hi1s1 _______450245(.DIN (_____0__19918), .Q (___00___19774));
  or2s1 _______450246(.DIN1 (_____________________18602), .DIN2
       (___00___19772), .Q (___00___19773));
  nor2s1 _______450247(.DIN1 (___0____20730), .DIN2 (___0_0), .Q
       (___00___19771));
  nor2s1 ______450248(.DIN1 (_____________________18608), .DIN2
       (___000), .Q (___00_));
  xor2s1 _______450249(.DIN1 (________19097), .DIN2 (____0____31818),
       .Q (___999));
  nnd2s1 ______450250(.DIN1 (___99___19769), .DIN2 (____9___22253), .Q
       (___99___19770));
  hi1s1 ______450251(.DIN (___99___19767), .Q (___99___19768));
  or2s1 _____0_450252(.DIN1 (___99___19765), .DIN2 (____9___19585), .Q
       (___99___19766));
  hi1s1 _______450253(.DIN (________20917), .Q (___99___19764));
  hi1s1 _______450254(.DIN (________20261), .Q (___99_));
  nor2s1 _______450255(.DIN1 (___0____19789), .DIN2 (____9___19197), .Q
       (___9____19763));
  xnr2s1 _______450256(.DIN1 (___9____19761), .DIN2
       (_________________18732), .Q (___9____19762));
  and2s1 _______450257(.DIN1 (___9____19695), .DIN2 (___0____20730), .Q
       (___9____19760));
  xor2s1 ______450258(.DIN1 (_____________0___18715), .DIN2
       (_____0__19351), .Q (___9____19759));
  hi1s1 ______450259(.DIN (_____0__20021), .Q (___9____19758));
  nnd2s1 _______450260(.DIN1 (___9____19756), .DIN2 (_____0__20002), .Q
       (___9____19757));
  xor2s1 _______450261(.DIN1 (___9_9__19754), .DIN2 (____9____29052),
       .Q (___9_0__19755));
  or2s1 _____9_450262(.DIN1 (___9____19752), .DIN2 (___0____19783), .Q
       (___9____19753));
  or2s1 _______450263(.DIN1 (___9____19697), .DIN2 (___0____19789), .Q
       (___9____19751));
  nor2s1 ______450264(.DIN1 (___9____19749), .DIN2 (___0____19815), .Q
       (___9____19750));
  nnd2s1 _______450265(.DIN1 (_____9__19638), .DIN2
       (_____________________18613), .Q (___9____19748));
  xor2s1 _______450266(.DIN1 (_________________18682), .DIN2
       (___9____19746), .Q (___9____19747));
  hi1s1 _______450267(.DIN (___9_9__19744), .Q (___9_0__19745));
  nor2s1 ______450268(.DIN1 (___0____19789), .DIN2 (___0____19815), .Q
       (___9____19743));
  nnd2s1 ______450269(.DIN1 (______9__33436), .DIN2 (___00____27191),
       .Q (___9____19741));
  or2s1 _______450270(.DIN1 (___9____19739), .DIN2 (_____9__19891), .Q
       (___9____19740));
  nor2s1 _____9_450271(.DIN1 (___9_0__19737), .DIN2 (___0____19815), .Q
       (___9____19738));
  nor2s1 ____9_450272(.DIN1 (____09__19601), .DIN2 (___9____19735), .Q
       (___9_9__19736));
  nnd2s1 _______450273(.DIN1 (___9____19733), .DIN2 (___9____19732), .Q
       (___9____19734));
  or2s1 _____0_450274(.DIN1 (_____________________18636), .DIN2
       (________20007), .Q (___9____19731));
  nnd2s1 _____0_450275(.DIN1 (_____0__19622), .DIN2
       (_____________________18599), .Q (___9____19730));
  hi1s1 _______450276(.DIN (________20387), .Q (________20202));
  nnd2s1 _______450277(.DIN1 (___9____19719), .DIN2 (___9____19729), .Q
       (________20067));
  nnd2s1 ______450278(.DIN1 (___9____19732), .DIN2 (________20194), .Q
       (________21847));
  nor2s1 _______450279(.DIN1 (_____0__20382), .DIN2 (___9___18975), .Q
       (___0____19830));
  hi1s1 _______450280(.DIN (________21776), .Q (_____0__21475));
  and2s1 _______450281(.DIN1 (____00__19592), .DIN2 (___9____19728), .Q
       (____9___20978));
  nnd2s1 ______450282(.DIN1 (________20213), .DIN2 (___9_0__19727), .Q
       (________20211));
  hi1s1 _______450283(.DIN (________22113), .Q (________21369));
  hi1s1 ______450284(.DIN (_____9__20381), .Q (___090___28044));
  hi1s1 ______450285(.DIN (___9_9__19726), .Q (________20117));
  hi1s1 _______450286(.DIN (________21794), .Q (____9___21351));
  hi1s1 _______450287(.DIN (____9____29953), .Q (_________29513));
  hi1s1 ______450288(.DIN (_____9__20557), .Q (________20065));
  hi1s1 _______450289(.DIN (________20454), .Q (________20368));
  hi1s1 ______450290(.DIN (________21472), .Q (________20076));
  hi1s1 ______450291(.DIN (_____9__20499), .Q (________20080));
  hi1s1 _______450292(.DIN (___9____19724), .Q (________20569));
  and2s1 _______450293(.DIN1 (____00__20226), .DIN2
       (____0________________18592), .Q (_____9__20068));
  and2s1 ______450294(.DIN1 (___9_9__19716), .DIN2 (___9____19723), .Q
       (________20063));
  nnd2s1 ______450295(.DIN1 (___9____19722), .DIN2
       (_____________________18605), .Q (___0____19836));
  hi1s1 _______450296(.DIN (___9____19721), .Q (________20215));
  nnd2s1 ____9__450297(.DIN1 (___9____19714), .DIN2 (________19472), .Q
       (____00__19947));
  nnd2s1 _______450298(.DIN1 (____9___19200), .DIN2 (______18932), .Q
       (________20336));
  nnd2s1 _______450299(.DIN1 (________21241), .DIN2 (________19098), .Q
       (_____0__20079));
  hi1s1 _______450300(.DIN (____9___21980), .Q (___0_0__20771));
  nor2s1 _______450301(.DIN1 (_______18950), .DIN2 (___99___19769), .Q
       (________20349));
  hi1s1 _______450302(.DIN (___9____19720), .Q (________25579));
  nnd2s1 _______450303(.DIN1 (___9____19719), .DIN2
       (_____________________18625), .Q (___0____19829));
  hi1s1 _______450304(.DIN (________21006), .Q (________21487));
  hi1s1 _______450305(.DIN (________21319), .Q (____0___20423));
  hi1s1 _______450306(.DIN (___0____21694), .Q (________20158));
  hi1s1 _______450307(.DIN (___90___21549), .Q (____0___21167));
  nnd2s1 ______450308(.DIN1 (____0___20330), .DIN2 (___9____19718), .Q
       (________20271));
  hi1s1 _____9_450309(.DIN (___0____21651), .Q (________20175));
  hi1s1 _______450310(.DIN (________21497), .Q (________20237));
  nor2s1 _______450311(.DIN1 (_____0__19612), .DIN2 (________19663), .Q
       (_____9__20216));
  nor2s1 _______450312(.DIN1 (___9_0__19717), .DIN2 (___9___18975), .Q
       (________20242));
  nor2s1 ____90_450313(.DIN1 (_____________________18663), .DIN2
       (___99___19769), .Q (_____9__20106));
  hi1s1 _______450314(.DIN (________22129), .Q (________20278));
  nnd2s1 _______450315(.DIN1 (___0____19805), .DIN2 (___9_9__19716), .Q
       (________20064));
  hi1s1 _______450316(.DIN (___9____19715), .Q (_____9__20125));
  and2s1 _____9_450317(.DIN1 (____0___19405), .DIN2 (___9____19714), .Q
       (___99___20695));
  nor2s1 _____0_450318(.DIN1 (____________________), .DIN2
       (________21468), .Q (________20252));
  hi1s1 _______450319(.DIN (___9____19713), .Q (______0__29662));
  hi1s1 _______450320(.DIN (________20398), .Q (________22116));
  hi1s1 _______450321(.DIN (________19884), .Q (_____0__21971));
  nor2s1 ____9__450322(.DIN1 (___9____19712), .DIN2 (___9____21568), .Q
       (________21233));
  nnd2s1 _____9_450323(.DIN1 (_____9__20313), .DIN2 (________19608), .Q
       (________20347));
  nnd2s1 _______450324(.DIN1 (___90___19688), .DIN2 (___0_9__19834), .Q
       (________20177));
  or2s1 _______450325(.DIN1 (___9____19711), .DIN2 (___9____19710), .Q
       (___0____22552));
  nnd2s1 _____450326(.DIN1 (________21197), .DIN2
       (______________________________________0__________0), .Q
       (____90__25071));
  nnd2s1 _______450327(.DIN1 (___9____19728), .DIN2 (________19996), .Q
       (________20386));
  nnd2s1 ______450328(.DIN1 (____99__19591), .DIN2 (____0___19402), .Q
       (_____0__21230));
  nnd2s1 _______450329(.DIN1 (_____0___33489), .DIN2 (________19353),
       .Q (_____9__21344));
  hi1s1 _______450330(.DIN (____0___19948), .Q (________20965));
  or2s1 ____0__450331(.DIN1 (____0_________________18656), .DIN2
       (_________34295), .Q (_____0__20304));
  or2s1 _______450332(.DIN1 (_____0___33866), .DIN2 (___0____19815), .Q
       (________20203));
  hi1s1 _____9_450333(.DIN (___9____19709), .Q (_________31395));
  hi1s1 _______450334(.DIN (___0_09__27568), .Q (____9____29986));
  hi1s1 _______450335(.DIN (___9____19708), .Q (____9___20219));
  or2s1 _______450336(.DIN1 (____0_________________18659), .DIN2
       (___9_0__19707), .Q (________20280));
  nnd2s1 _______450337(.DIN1 (_____0__19602), .DIN2 (____9___19584), .Q
       (________20307));
  nnd2s1 ____450338(.DIN1 (_____0___33489), .DIN2 (________19412), .Q
       (___0____20753));
  nor2s1 ____9__450339(.DIN1 (____0___19594), .DIN2 (___9_9__19706), .Q
       (________21238));
  and2s1 _______450340(.DIN1 (_____0___33489), .DIN2 (________19549),
       .Q (________20109));
  nor2s1 ____0__450341(.DIN1 (________19442), .DIN2 (___9____19705), .Q
       (_____0__20254));
  hi1s1 _______450342(.DIN (___9____19704), .Q (________20210));
  hi1s1 _____9_450343(.DIN (________21471), .Q (________21368));
  hi1s1 _______450344(.DIN (___9____19703), .Q (________21213));
  and2s1 _______450345(.DIN1 (___9____19702), .DIN2 (___9____19701), .Q
       (________20802));
  nnd2s1 _______450346(.DIN1 (_____0__19572), .DIN2 (___9____19700), .Q
       (________20384));
  and2s1 _____9_450347(.DIN1 (___9____19699), .DIN2 (________19615), .Q
       (________21193));
  hi1s1 _______450348(.DIN (___9_0__19698), .Q (____9___21353));
  nor2s1 _______450349(.DIN1 (_____0__19234), .DIN2 (___9_9), .Q
       (_________29330));
  nor2s1 _______450350(.DIN1 (___9____19697), .DIN2 (___9_0__19737), .Q
       (________20843));
  nnd2s1 ______450351(.DIN1 (___9____19696), .DIN2 (________19518), .Q
       (________20286));
  nor2s1 ____09_450352(.DIN1 (________19230), .DIN2 (____90__19196), .Q
       (___9____20645));
  nnd2s1 _______450353(.DIN1 (___9____19695), .DIN2 (___9____19694), .Q
       (________22110));
  hi1s1 _____0_450354(.DIN (____9___21984), .Q (___9_0__21561));
  nnd2s1 ____9__450355(.DIN1 (_____9__20313), .DIN2 (________19603), .Q
       (________21887));
  nnd2s1 ____9_450356(.DIN1 (________21797), .DIN2 (____0___19597), .Q
       (________21750));
  nor2s1 ____90_450357(.DIN1 (___9____19693), .DIN2 (________19555), .Q
       (_____0__21335));
  nnd2s1 ____9__450358(.DIN1 (___9____19714), .DIN2 (___9____19699), .Q
       (________21506));
  hi1s1 _______450359(.DIN (___99___22527), .Q (___0____23448));
  nnd2s1 ____9__450360(.DIN1 (________21824), .DIN2 (________19978), .Q
       (___0____20763));
  hi1s1 _______450361(.DIN (________20084), .Q (____0___21816));
  nor2s1 ____90_450362(.DIN1 (________19545), .DIN2 (_________31702),
       .Q (_________30374));
  nor2s1 ____9__450363(.DIN1 (___9____19691), .DIN2 (________19273), .Q
       (____90__21801));
  nnd2s1 ____9__450364(.DIN1 (___0____19822), .DIN2 (___9____19729), .Q
       (________20390));
  hi1s1 _____9_450365(.DIN (_________33370), .Q (_________33279));
  nor2s1 _______450366(.DIN1 (___9__), .DIN2 (___9_0), .Q
       (____00___33677));
  hi1s1 _______450367(.DIN (_____0__20207), .Q (________22341));
  hi1s1 _______450368(.DIN (___9____19692), .Q (________19962));
  nor2s1 _____0_450369(.DIN1 (________19256), .DIN2 (________19526), .Q
       (___909));
  and2s1 ____00_450370(.DIN1 (___0_9__19844), .DIN2 (________19164), .Q
       (___90___19690));
  nnd2s1 _____9_450371(.DIN1 (___90___19688), .DIN2 (________19576), .Q
       (___90___19689));
  or2s1 _______450372(.DIN1 (__________________0_), .DIN2
       (___9_0__19737), .Q (___90___19687));
  nor2s1 _______450373(.DIN1 (____0___24155), .DIN2 (________19254), .Q
       (___90___19686));
  nnd2s1 _______450374(.DIN1 (___0_0), .DIN2 (___9____19718), .Q
       (___90_));
  xor2s1 _______450375(.DIN1 (_____9__19133), .DIN2 (___9____21556), .Q
       (___900));
  nor2s1 _____0_450376(.DIN1 (_____9__20491), .DIN2 (_____0__20352), .Q
       (____99__19685));
  xor2s1 _______450377(.DIN1 (_____________18895), .DIN2
       (___00___19777), .Q (____9___19684));
  nnd2s1 _______450378(.DIN1 (________19227), .DIN2 (_____0__19252), .Q
       (____9___19683));
  nor2s1 ______450379(.DIN1 (inData[18]), .DIN2 (_________31702), .Q
       (____9___19682));
  or2s1 _______450380(.DIN1 (_______19003), .DIN2 (______9__33436), .Q
       (____9___19681));
  nor2s1 _______450381(.DIN1 (_____0__19429), .DIN2 (________19180), .Q
       (____9___19680));
  xor2s1 _______450382(.DIN1 (____9___19110), .DIN2 (______0__34461),
       .Q (____9___19679));
  nnd2s1 _______450383(.DIN1 (___9____19735), .DIN2
       (_____________________18610), .Q (____9___19678));
  nnd2s1 _______450384(.DIN1 (________20160), .DIN2 (___9____19739), .Q
       (____90__19677));
  nor2s1 _______450385(.DIN1 (_____0__19956), .DIN2 (_____0__20274), .Q
       (_____9__19676));
  nnd2s1 ______450386(.DIN1 (________20213), .DIN2 (___9____19719), .Q
       (________19675));
  nnd2s1 _______450387(.DIN1 (_____0__20002), .DIN2 (________19617), .Q
       (________19674));
  nor2s1 _____9_450388(.DIN1 (________20213), .DIN2 (________21797), .Q
       (________19673));
  nor2s1 _______450389(.DIN1 (___0____19822), .DIN2 (___9____19732), .Q
       (________19672));
  nnd2s1 _______450390(.DIN1 (_____9__19251), .DIN2 (_________18845),
       .Q (________19671));
  nor2s1 ______450391(.DIN1 (_____0__19669), .DIN2 (_____9__19668), .Q
       (________19670));
  nor2s1 _______450392(.DIN1 (______18933), .DIN2 (________21857), .Q
       (________19667));
  nnd2s1 ______450393(.DIN1 (____0___19596), .DIN2 (________19665), .Q
       (________19666));
  nor2s1 _______450394(.DIN1 (________19663), .DIN2 (_____9__19891), .Q
       (________19664));
  nnd2s1 _____450395(.DIN1 (________19661), .DIN2 (_________18862), .Q
       (________19662));
  or2s1 _______450396(.DIN1 (____0________________18589), .DIN2
       (____9___20413), .Q (________19660));
  xor2s1 _______450397(.DIN1 (____9__19045), .DIN2 (outData[20]), .Q
       (_____0__19659));
  xor2s1 ______450398(.DIN1 (______18932), .DIN2 (___0__18931), .Q
       (_____9__19658));
  xor2s1 _______450399(.DIN1 (____09__19311), .DIN2
       (______________0___________________9), .Q (________19657));
  and2s1 _____450400(.DIN1 (___0____19783), .DIN2 (________19655), .Q
       (________19656));
  hi1s1 _______450401(.DIN (____9___20037), .Q (________19654));
  hi1s1 _____0_450402(.DIN (_____0__22118), .Q (________19653));
  xor2s1 _______450403(.DIN1 (______0__34451), .DIN2 (_______18993), .Q
       (________19652));
  xor2s1 _______450404(.DIN1 (____0___19122), .DIN2
       (______________0____________________), .Q (________19651));
  nnd2s1 _____450405(.DIN1 (_________31702), .DIN2 (_________31388), .Q
       (________19650));
  or2s1 _______450406(.DIN1 (____0_____________0_), .DIN2
       (___9____19691), .Q (_____0__19649));
  nor2s1 _______450407(.DIN1 (___0____22547), .DIN2 (________19423), .Q
       (_____9__19648));
  xor2s1 ____09_450408(.DIN1 (________19136), .DIN2 (_______18999), .Q
       (________19647));
  nor2s1 _______450409(.DIN1 (________19645), .DIN2 (___000), .Q
       (________19646));
  or2s1 ____9__450410(.DIN1 (________19643), .DIN2 (_____0__20274), .Q
       (________19644));
  nnd2s1 _______450411(.DIN1 (_____0__21298), .DIN2 (________19978), .Q
       (________19642));
  and2s1 _______450412(.DIN1 (___9____19714), .DIN2
       (_____________________18615), .Q (________19641));
  nor2s1 ______450413(.DIN1 (________19457), .DIN2 (___9____19691), .Q
       (________19640));
  nnd2s1 ____9__450414(.DIN1 (_____9__19638), .DIN2 (____90__19582), .Q
       (_____0__19639));
  xnr2s1 _______450415(.DIN1 (______0__18842), .DIN2 (________19636),
       .Q (________19637));
  and2s1 _______450416(.DIN1 (_____9__19638), .DIN2
       (_____________________18612), .Q (________19635));
  hi1s1 _______450417(.DIN (________20208), .Q (________19634));
  nor2s1 ____9__450418(.DIN1 (____0___21724), .DIN2 (___9____19705), .Q
       (________19633));
  nor2s1 _____0_450419(.DIN1 (____00__19114), .DIN2 (________19631), .Q
       (________19632));
  and2s1 _______450420(.DIN1 (________21241), .DIN2 (_____0__20392), .Q
       (_____9__19630));
  nnd2s1 _______450421(.DIN1 (_________31702), .DIN2
       (______________________________________0_____________18889), .Q
       (________19629));
  or2s1 _______450422(.DIN1 (_________9_______18807), .DIN2
       (___9___18975), .Q (________19628));
  nor2s1 _______450423(.DIN1 (________19092), .DIN2 (_____0___32299),
       .Q (________19627));
  nor2s1 _______450424(.DIN1 (________19142), .DIN2 (________19183), .Q
       (________19626));
  or2s1 _____9_450425(.DIN1 (________19624), .DIN2 (________21241), .Q
       (________19625));
  and2s1 ____9_450426(.DIN1 (_____0__19622), .DIN2 (___90), .Q
       (________19623));
  nor2s1 _______450427(.DIN1 (________19620), .DIN2 (_____0__21885), .Q
       (_____9__19621));
  nnd2s1 ______450428(.DIN1 (___9____19719), .DIN2 (________20194), .Q
       (________19619));
  nor2s1 _______450429(.DIN1 (________19617), .DIN2 (________19238), .Q
       (________19618));
  nnd2s1 ____9__450430(.DIN1 (_____9__19638), .DIN2 (________19615), .Q
       (________19616));
  hi1s1 ______450431(.DIN (________20543), .Q (________20083));
  and2s1 _______450432(.DIN1 (___9____19696), .DIN2
       (____0________________18595), .Q (________20066));
  nor2s1 _____450433(.DIN1 (________19614), .DIN2 (_____9__19242), .Q
       (___0____19837));
  hi1s1 _____9_450434(.DIN (________21222), .Q (____9___20218));
  nor2s1 _____9_450435(.DIN1 (___0____20746), .DIN2 (________21021), .Q
       (________19967));
  nor2s1 _______450436(.DIN1 (________20123), .DIN2 (_____0__21298), .Q
       (___0____19833));
  or2s1 _______450437(.DIN1 (______________________18617), .DIN2
       (___0____19815), .Q (________20169));
  nor2s1 _______450438(.DIN1 (_____0__19612), .DIN2 (_____0__20274), .Q
       (_____9__21239));
  nnd2s1 _______450439(.DIN1 (________19605), .DIN2
       (_____________________18599), .Q (___0____19832));
  nor2s1 _______450440(.DIN1 (___0____19780), .DIN2 (___0____19815), .Q
       (________19974));
  nor2s1 ____9_450441(.DIN1 (_____9__21513), .DIN2 (___9____19711), .Q
       (____99__19946));
  nnd2s1 ______450442(.DIN1 (_____9__19611), .DIN2 (________21976), .Q
       (____9___19944));
  hi1s1 ______450443(.DIN (________20850), .Q (________20934));
  nor2s1 ______450444(.DIN1 (_____________________18602), .DIN2
       (___9____19723), .Q (________20081));
  and2s1 _______450445(.DIN1 (________19978), .DIN2
       (______________________18631), .Q (________20359));
  nor2s1 _______450446(.DIN1 (________19417), .DIN2 (________21857), .Q
       (____0___19951));
  or2s1 _______450447(.DIN1 (_______18966), .DIN2 (________19178), .Q
       (________20101));
  nor2s1 _______450448(.DIN1 (________19610), .DIN2 (___00___19772), .Q
       (________19866));
  nnd2s1 _______450449(.DIN1 (________20072), .DIN2 (___0____19783), .Q
       (________21122));
  nor2s1 _______450450(.DIN1 (_____0__20382), .DIN2 (_________34295),
       .Q (________20077));
  nnd2s1 _______450451(.DIN1 (___9____19695), .DIN2
       (_____________________18664), .Q (________20435));
  hi1s1 _______450452(.DIN (________19609), .Q (____0___25857));
  nor2s1 ______450453(.DIN1 (________19604), .DIN2 (___0____21699), .Q
       (________19907));
  nor2s1 _______450454(.DIN1 (____9___19586), .DIN2 (___0____19789), .Q
       (________20082));
  nor2s1 _______450455(.DIN1 (________20091), .DIN2 (___0____19800), .Q
       (________20074));
  nnd2s1 _______450456(.DIN1 (________19655), .DIN2 (________19617), .Q
       (________19983));
  hi1s1 _______450457(.DIN (________22119), .Q (________20300));
  nnd2s1 _______450458(.DIN1 (________19655), .DIN2 (________19608), .Q
       (________21228));
  nnd2s1 ____9__450459(.DIN1 (_____9__19611), .DIN2
       (_____________________18664), .Q (________20199));
  nnd2s1 ____09_450460(.DIN1 (________19607), .DIN2 (________22050), .Q
       (________21388));
  nor2s1 _______450461(.DIN1 (________19610), .DIN2 (___9____19723), .Q
       (________20257));
  nor2s1 ______450462(.DIN1 (____0________________18647), .DIN2
       (________19579), .Q (________20070));
  nnd2s1 _____0_450463(.DIN1 (____0___19593), .DIN2 (________19655), .Q
       (________20311));
  nnd2s1 _______450464(.DIN1 (_____0___32299), .DIN2 (___9_0__19707),
       .Q (________20120));
  nor2s1 _____0_450465(.DIN1 (________19430), .DIN2 (___9_0__19737), .Q
       (____9___20224));
  and2s1 ____0__450466(.DIN1 (_____0__20274), .DIN2 (________19606), .Q
       (____9___20883));
  nor2s1 _______450467(.DIN1 (________19605), .DIN2 (________19171), .Q
       (___9_9__20643));
  hi1s1 _______450468(.DIN (____0___20046), .Q (______0__30418));
  or2s1 ______450469(.DIN1 (_____________________18634), .DIN2
       (________20007), .Q (____9___20221));
  nor2s1 _______450470(.DIN1 (________21976), .DIN2 (_____0__19669), .Q
       (________20201));
  hi1s1 _______450471(.DIN (________20023), .Q (________20192));
  nor2s1 ______450472(.DIN1 (_____________________18664), .DIN2
       (________19604), .Q (________20493));
  or2s1 _______450473(.DIN1 (_____________________18635), .DIN2
       (___0____19800), .Q (____9___20504));
  nnd2s1 ______450474(.DIN1 (________19655), .DIN2 (________19603), .Q
       (________20353));
  nnd2s1 _____450475(.DIN1 (_____0__19602), .DIN2 (________19573), .Q
       (________21479));
  and2s1 _____9_450476(.DIN1 (___0____19822), .DIN2
       (_____________________18625), .Q (________20075));
  nor2s1 _____0_450477(.DIN1 (_____________________18665), .DIN2
       (___9____19711), .Q (________20268));
  nor2s1 _______450478(.DIN1 (___9____19693), .DIN2 (____09__19601), .Q
       (________20196));
  nnd2s1 _____450479(.DIN1 (____0___20330), .DIN2 (___9____19695), .Q
       (___9____22524));
  nor2s1 ______450480(.DIN1 (____0___19600), .DIN2 (_____0__21429), .Q
       (_____0__20156));
  nnd2s1 _______450481(.DIN1 (___0_0__19810), .DIN2
       (_____________________18663), .Q (________20854));
  hi1s1 _______450482(.DIN (________21025), .Q (___90___21544));
  nnd2s1 _______450483(.DIN1 (____0___19599), .DIN2 (________19434), .Q
       (________21032));
  hi1s1 _______450484(.DIN (____0___19598), .Q (________20205));
  and2s1 _______450485(.DIN1 (_____9__19551), .DIN2 (_____0___32299),
       .Q (________20154));
  hi1s1 _____0_450486(.DIN (___0____21660), .Q (________21481));
  nnd2s1 _______450487(.DIN1 (________20213), .DIN2 (____0___19597), .Q
       (________21276));
  nnd2s1 _______450488(.DIN1 (____0___19596), .DIN2 (____0___19595), .Q
       (________20470));
  nnd2s1 ____9__450489(.DIN1 (________20072), .DIN2 (________19603), .Q
       (____00__21355));
  nor2s1 _______450490(.DIN1 (____0___19594), .DIN2 (________20007), .Q
       (________21023));
  nor2s1 ____9__450491(.DIN1 (___9____19712), .DIN2 (_____0__21429), .Q
       (________21381));
  nnd2s1 _______450492(.DIN1 (________20072), .DIN2 (____0___19593), .Q
       (________21114));
  and2s1 _______450493(.DIN1 (____9___19590), .DIN2
       (____0_________________18656), .Q (___0____20756));
  nnd2s1 ______450494(.DIN1 (____00__19592), .DIN2 (_____0__19243), .Q
       (____99__20509));
  or2s1 _______450495(.DIN1 (_____________________18612), .DIN2
       (_____9__19571), .Q (________20831));
  nnd2s1 _______450496(.DIN1 (____99__19591), .DIN2 (________19431), .Q
       (________20561));
  nnd2s1 ______450497(.DIN1 (____9___19590), .DIN2 (_____0__20382), .Q
       (________20277));
  nor2s1 ______450498(.DIN1 (________19260), .DIN2 (________20007), .Q
       (________21201));
  nnd2s1 ____9__450499(.DIN1 (________19219), .DIN2 (inData[30]), .Q
       (____9___19945));
  nnd2s1 _____9_450500(.DIN1 (____0___19599), .DIN2 (____9___19589), .Q
       (_____9__21019));
  nnd2s1 _______450501(.DIN1 (________19416), .DIN2 (___90___19688), .Q
       (____9___21804));
  hi1s1 _______450502(.DIN (____9___19588), .Q (____9___20881));
  and2s1 _______450503(.DIN1 (____9___19587), .DIN2 (___0____19783), .Q
       (____0___20143));
  hi1s1 ______450504(.DIN (________20110), .Q (____0___21080));
  or2s1 _______450505(.DIN1 (____9___19586), .DIN2 (___9_0__19737), .Q
       (________20825));
  nor2s1 _______450506(.DIN1 (____0___21991), .DIN2 (________21021), .Q
       (___9____20657));
  nnd2s1 _______450507(.DIN1 (___9____19719), .DIN2 (____9___19585), .Q
       (________22333));
  hi1s1 _______450508(.DIN (________21476), .Q (_____9__20816));
  nnd2s1 _______450509(.DIN1 (________20213), .DIN2 (_____0__21885), .Q
       (________21180));
  nnd2s1 ____90_450510(.DIN1 (___9____19695), .DIN2
       (_____________________18668), .Q (________20405));
  nnd2s1 _____0_450511(.DIN1 (________19574), .DIN2 (____9___19584), .Q
       (________21488));
  hi1s1 _______450512(.DIN (____9___19583), .Q (_____9__20932));
  nor2s1 _______450513(.DIN1 (____0___19210), .DIN2 (___9____19739), .Q
       (________22211));
  or2s1 _______450514(.DIN1 (________19444), .DIN2 (________20007), .Q
       (_____0__21046));
  nnd2s1 ____9__450515(.DIN1 (____90__19582), .DIN2 (___9____19699), .Q
       (________21333));
  nor2s1 _______450516(.DIN1 (_____9__19515), .DIN2 (___000), .Q
       (___0_9__20779));
  nnd2s1 _______450517(.DIN1 (____9___19397), .DIN2 (___9_0__19707), .Q
       (___0____21680));
  and2s1 ______450518(.DIN1 (___0____19783), .DIN2
       (____0________________18649), .Q (________20338));
  nor2s1 _______450519(.DIN1 (____0___19594), .DIN2 (________20564), .Q
       (________21205));
  hi1s1 _______450520(.DIN (_____9__19581), .Q (________20247));
  nor2s1 _______450521(.DIN1 (________19580), .DIN2 (________19579), .Q
       (________21509));
  hi1s1 ______450522(.DIN (________19578), .Q (________21131));
  nor2s1 _______450523(.DIN1 (________19182), .DIN2 (________19577), .Q
       (________21480));
  nnd2s1 _______450524(.DIN1 (________20395), .DIN2 (________19576), .Q
       (________20389));
  hi1s1 _______450525(.DIN (________19864), .Q (________21226));
  nor2s1 _____9_450526(.DIN1 (_____9__19261), .DIN2 (___9____19739), .Q
       (________20813));
  nnd2s1 _____9_450527(.DIN1 (________19575), .DIN2 (________21241), .Q
       (___9____21618));
  nor2s1 _______450528(.DIN1 (____09__19408), .DIN2 (___000), .Q
       (________20946));
  nor2s1 _____9_450529(.DIN1 (_____0__19409), .DIN2 (___9____19739), .Q
       (________22109));
  nor2s1 ____9__450530(.DIN1 (______0__28643), .DIN2 (____9___19200),
       .Q (_____0__19985));
  nnd2s1 _____9_450531(.DIN1 (________19574), .DIN2 (________19573), .Q
       (________21502));
  nor2s1 ____9_450532(.DIN1 (____0___19600), .DIN2 (___9____21568), .Q
       (_____9__21278));
  nor2s1 _____450533(.DIN1 (__________________0___18670), .DIN2
       (________20292), .Q (___0____21690));
  nnd2s1 ____9_450534(.DIN1 (___9____19701), .DIN2 (_____0__19572), .Q
       (____0___21362));
  nnd2s1 ____9__450535(.DIN1 (___0____19783), .DIN2 (____0___19059), .Q
       (_____9__20341));
  or2s1 ____90_450536(.DIN1 (________19523), .DIN2 (_____0__21298), .Q
       (________22037));
  nor2s1 ____9_450537(.DIN1 (____9___22253), .DIN2 (_________31702), .Q
       (____9____31759));
  nor2s1 _______450538(.DIN1 (____9___22253), .DIN2 (___99___19769), .Q
       (________21313));
  and2s1 ____9__450539(.DIN1 (________21241), .DIN2 (________19978), .Q
       (________21458));
  and2s1 _______450540(.DIN1 (____0___19594), .DIN2
       (_____________________18641), .Q (_________32901));
  or2s1 _______450541(.DIN1 (____0___19504), .DIN2 (______9__33436), .Q
       (______0__33373));
  and2s1 _______450542(.DIN1 (___9____19722), .DIN2 (________19436), .Q
       (________21211));
  nor2s1 ____9__450543(.DIN1 (_____9__19571), .DIN2 (________19410), .Q
       (___0_0__21658));
  hi1s1 _______450544(.DIN (________19570), .Q (________23757));
  nnd2s1 _______450545(.DIN1 (____9___19201), .DIN2
       (____0________________18589), .Q (________19569));
  nor2s1 _______450546(.DIN1 (________19062), .DIN2 (___9____19712), .Q
       (________19568));
  hi1s1 _______450547(.DIN (________19566), .Q (________19567));
  or2s1 _______450548(.DIN1 (_____________________18622), .DIN2
       (________19564), .Q (________19565));
  nor2s1 _______450549(.DIN1 (_____________________18635), .DIN2
       (___9_9__19706), .Q (________19563));
  or2s1 _______450550(.DIN1 (_____0__20392), .DIN2 (________19099), .Q
       (_____0__19562));
  nnd2s1 _____9_450551(.DIN1 (_____________________18662), .DIN2
       (________19137), .Q (_____9__19561));
  nnd2s1 _______450552(.DIN1 (________19530), .DIN2 (___0_9__19834), .Q
       (________19560));
  nnd2s1 _______450553(.DIN1 (________19540), .DIN2 (________19576), .Q
       (________19559));
  nnd2s1 _______450554(.DIN1 (________19557), .DIN2
       (____0______________), .Q (________19558));
  nor2s1 _______450555(.DIN1 (________19141), .DIN2 (________19555), .Q
       (________19556));
  nnd2s1 ______450556(.DIN1 (________19553), .DIN2 (________19557), .Q
       (________19554));
  nor2s1 _____450557(.DIN1 (_________28766), .DIN2 (_____9__19551), .Q
       (_____0__19552));
  nnd2s1 _______450558(.DIN1 (________19549), .DIN2 (____0___19309), .Q
       (________19550));
  nnd2s1 ______450559(.DIN1 (________19547), .DIN2
       (_________________9___18616), .Q (________19548));
  nnd2s1 _______450560(.DIN1 (________19545), .DIN2 (inData[20]), .Q
       (________19546));
  nor2s1 _______450561(.DIN1 (________19564), .DIN2 (________19620), .Q
       (________19544));
  or2s1 _______450562(.DIN1 (_____________________18609), .DIN2
       (____09__19601), .Q (________19542));
  nor2s1 _______450563(.DIN1 (____0_______________), .DIN2
       (________19540), .Q (________19541));
  or2s1 _______450564(.DIN1 (_____________________18620), .DIN2
       (_____9__22215), .Q (________19539));
  and2s1 _______450565(.DIN1 (________19424), .DIN2 (_____9__20491), .Q
       (________19538));
  and2s1 _______450566(.DIN1 (________19536), .DIN2 (________19535), .Q
       (________19537));
  nor2s1 _______450567(.DIN1 (______________________18671), .DIN2
       (________19345), .Q (_____0__19534));
  or2s1 _______450568(.DIN1 (________19325), .DIN2 (___9____19701), .Q
       (_____9__19533));
  or2s1 _______450569(.DIN1 (_____________________18668), .DIN2
       (________20073), .Q (________19532));
  nnd2s1 ______450570(.DIN1 (________19530), .DIN2 (________19576), .Q
       (________19531));
  and2s1 _______450571(.DIN1 (_____9__22215), .DIN2 (___9__), .Q
       (________19529));
  nnd2s1 _______450572(.DIN1 (____9___19393), .DIN2 (______18933), .Q
       (________19528));
  nnd2s1 _______450573(.DIN1 (_____0__19506), .DIN2 (_______18971), .Q
       (________19527));
  nnd2s1 _______450574(.DIN1 (____00__19592), .DIN2 (____0___19207), .Q
       (_____0__19525));
  or2s1 _______450575(.DIN1 (______________________18631), .DIN2
       (________19523), .Q (_____9__19524));
  and2s1 _______450576(.DIN1 (________21003), .DIN2 (____0___19595), .Q
       (________19522));
  xor2s1 ______450577(.DIN1 (________19378), .DIN2
       (_________________18794), .Q (________19521));
  nor2s1 ____9__450578(.DIN1 (inData[30]), .DIN2 (________19263), .Q
       (________19520));
  nor2s1 ______450579(.DIN1 (________19518), .DIN2 (____0___19403), .Q
       (________19519));
  nnd2s1 _____9_450580(.DIN1 (_______19008), .DIN2 (inData[2]), .Q
       (________19517));
  nor2s1 _______450581(.DIN1 (________19555), .DIN2 (_____9__19515), .Q
       (_____0__19516));
  or2s1 _______450582(.DIN1 (_____________________18626), .DIN2
       (________19513), .Q (________19514));
  nnd2s1 _______450583(.DIN1 (____00), .DIN2 (________19511), .Q
       (________19512));
  and2s1 _____450584(.DIN1 (________19383), .DIN2 (___99___19765), .Q
       (________19510));
  nnd2s1 _____0_450585(.DIN1 (________21115), .DIN2 (_____0__22063), .Q
       (________19509));
  and2s1 _____9_450586(.DIN1 (________21824), .DIN2 (________19624), .Q
       (________19508));
  nnd2s1 _______450587(.DIN1 (_____9__19291), .DIN2 (_____0__19506), .Q
       (________19507));
  nnd2s1 _______450588(.DIN1 (____0___19504), .DIN2 (_______19002), .Q
       (____09__19505));
  nor2s1 ______450589(.DIN1 (____90__19582), .DIN2 (________19577), .Q
       (____0___19503));
  nnd2s1 _______450590(.DIN1 (____0___19307), .DIN2
       (_____________________18603), .Q (____0___19502));
  nnd2s1 _______450591(.DIN1 (___9____19733), .DIN2 (____0___19404), .Q
       (____0___19501));
  and2s1 _______450592(.DIN1 (___9__18942), .DIN2 (___9_9__19754), .Q
       (____0___19500));
  xnr2s1 _______450593(.DIN1 (_________9______18799), .DIN2
       (________19358), .Q (____0___19499));
  nor2s1 _______450594(.DIN1 (________19063), .DIN2 (____0___19497), .Q
       (____0___19498));
  nor2s1 _____9_450595(.DIN1 (_____9__21513), .DIN2 (____9___19108), .Q
       (____00__19496));
  nor2s1 _______450596(.DIN1 (____0________________18651), .DIN2
       (________19606), .Q (____9___19494));
  nor2s1 _______450597(.DIN1 (________19369), .DIN2 (________19555), .Q
       (____9___19493));
  nnd2s1 _______450598(.DIN1 (_____9__19543), .DIN2 (________19139), .Q
       (____9___19492));
  nnd2s1 _______450599(.DIN1 (____9___19490), .DIN2
       (____0________________18651), .Q (____9___19491));
  nnd2s1 _______450600(.DIN1 (___9____19701), .DIN2 (____9___19488), .Q
       (____9___19489));
  nnd2s1 _______450601(.DIN1 (________19553), .DIN2 (________19483), .Q
       (____90__19487));
  xor2s1 _______450602(.DIN1 (______0__34471), .DIN2 (________19226),
       .Q (_____9__19486));
  nnd2s1 _______450603(.DIN1 (________21824), .DIN2
       (______________________18629), .Q (________19485));
  nor2s1 _______450604(.DIN1 (________19483), .DIN2 (________19553), .Q
       (________19484));
  nnd2s1 _______450605(.DIN1 (___9_9__19716), .DIN2
       (_____________________18600), .Q (________19482));
  nor2s1 ______450606(.DIN1 (___9_0__19727), .DIN2 (____0___19206), .Q
       (________19481));
  or2s1 _______450607(.DIN1 (_____9__19467), .DIN2 (____0___19497), .Q
       (________19480));
  xor2s1 ____0__450608(.DIN1 (_____0___29362), .DIN2 (______0__28643),
       .Q (________19479));
  nnd2s1 ______450609(.DIN1 (_______19004), .DIN2 (inData[22]), .Q
       (________19478));
  nor2s1 _______450610(.DIN1 (________19435), .DIN2 (____00__19302), .Q
       (_____0__19477));
  nnd2s1 _______450611(.DIN1 (____99__19204), .DIN2 (________21115), .Q
       (_____9__19476));
  xor2s1 _______450612(.DIN1 (_________28581), .DIN2 (______0__28643),
       .Q (________19475));
  nnd2s1 ______450613(.DIN1 (____0___19595), .DIN2 (________22050), .Q
       (________19474));
  nnd2s1 _______450614(.DIN1 (________19472), .DIN2 (___0____19807), .Q
       (________19473));
  nnd2s1 _______450615(.DIN1 (___9_9__19716), .DIN2 (________19470), .Q
       (________19471));
  nnd2s1 _______450616(.DIN1 (____9___19490), .DIN2 (_____0__19956), .Q
       (________19469));
  nor2s1 _______450617(.DIN1 (____0________________18593), .DIN2
       (_____9__19467), .Q (_____0__19468));
  and2s1 _____0_450618(.DIN1 (________19511), .DIN2 (___9____19694), .Q
       (________19466));
  or2s1 _______450619(.DIN1 (____0_________________18656), .DIN2
       (_____9__19271), .Q (________19465));
  nnd2s1 _______450620(.DIN1 (___9_9__19716), .DIN2 (________19463), .Q
       (________19464));
  and2s1 _______450621(.DIN1 (________19461), .DIN2
       (_____________________18608), .Q (________19462));
  nnd2s1 ______450622(.DIN1 (___0_9__19844), .DIN2
       (____0_________________18657), .Q (________19460));
  nor2s1 _____0_450623(.DIN1 (________19147), .DIN2 (________20901), .Q
       (________19459));
  nnd2s1 _____9_450624(.DIN1 (____0___19597), .DIN2 (________19278), .Q
       (________19875));
  nor2s1 _____9_450625(.DIN1 (________19455), .DIN2 (___9____21610), .Q
       (___9_9__19726));
  and2s1 _______450626(.DIN1 (________19415), .DIN2 (____9___19490), .Q
       (___09___20782));
  nor2s1 ______450627(.DIN1 (________19457), .DIN2 (________19456), .Q
       (____09__19955));
  nor2s1 _____450628(.DIN1 (________19455), .DIN2 (___9_0__19717), .Q
       (________19578));
  nnd2s1 _______450629(.DIN1 (________19159), .DIN2 (_____0___28711),
       .Q (____9____30893));
  nnd2s1 ______450630(.DIN1 (________19454), .DIN2 (________19453), .Q
       (________19609));
  or2s1 _______450631(.DIN1 (___9____19697), .DIN2 (___9____19749), .Q
       (________19957));
  nnd2s1 _______450632(.DIN1 (_____9__19448), .DIN2 (________19184), .Q
       (________19898));
  nor2s1 _______450633(.DIN1 (____9___19299), .DIN2 (________19411), .Q
       (___9____19708));
  nor2s1 _______450634(.DIN1 (________19452), .DIN2 (_______19010), .Q
       (___0____22549));
  nnd2s1 _____9_450635(.DIN1 (____0___19212), .DIN2 (____0___21812), .Q
       (____9___19583));
  nor2s1 ______450636(.DIN1 (________19451), .DIN2 (________19450), .Q
       (_________34189));
  nor2s1 _____450637(.DIN1 (____0___19054), .DIN2 (________19456), .Q
       (_____9__19926));
  nnd2s1 _______450638(.DIN1 (_____0__19449), .DIN2 (_____0__19215), .Q
       (____9___20877));
  nnd2s1 ______450639(.DIN1 (_____9__19448), .DIN2
       (_____________________18621), .Q (________19874));
  nor2s1 _____9_450640(.DIN1 (________19447), .DIN2 (________19446), .Q
       (___99___19767));
  nor2s1 _____9_450641(.DIN1 (________20091), .DIN2 (________19445), .Q
       (_____9__19581));
  nnd2s1 ______450642(.DIN1 (____0___19595), .DIN2
       (____0________________18594), .Q (____0___19598));
  or2s1 ____9__450643(.DIN1 (_______18962), .DIN2 (________19961), .Q
       (___9____19709));
  nor2s1 _____450644(.DIN1 (________19444), .DIN2 (________20564), .Q
       (___9_0__19698));
  nnd2s1 _______450645(.DIN1 (________19443), .DIN2 (____0___19305), .Q
       (________19976));
  nor2s1 _______450646(.DIN1 (________19442), .DIN2 (________19513), .Q
       (________20393));
  and2s1 ______450647(.DIN1 (________19441), .DIN2 (________19440), .Q
       (________20212));
  or2s1 _______450648(.DIN1 (________19455), .DIN2 (____9___21071), .Q
       (________21742));
  or2s1 _______450649(.DIN1 (____0________________18595), .DIN2
       (_____0__19439), .Q (____0___19952));
  nor2s1 ______450650(.DIN1 (_____9__19438), .DIN2 (________19188), .Q
       (________20295));
  nnd2s1 _______450651(.DIN1 (____0___21988), .DIN2 (_____0__20097), .Q
       (___9____19704));
  nor2s1 ______450652(.DIN1 (________19996), .DIN2 (________19437), .Q
       (________19911));
  nor2s1 _____9_450653(.DIN1 (________19436), .DIN2 (________19435), .Q
       (___0____19831));
  nor2s1 _____0_450654(.DIN1 (____9___19295), .DIN2 (________20564), .Q
       (________19886));
  nnd2s1 _______450655(.DIN1 (___900__20605), .DIN2
       (____0________________18647), .Q (________20084));
  nnd2s1 _______450656(.DIN1 (_____0__19602), .DIN2 (___0___18983), .Q
       (____09__20519));
  nor2s1 _______450657(.DIN1 (________19455), .DIN2 (_____9__19281), .Q
       (________22119));
  nor2s1 ______450658(.DIN1 (____0___19860), .DIN2 (________19624), .Q
       (________19884));
  nnd2s1 _______450659(.DIN1 (________19434), .DIN2 (________19433), .Q
       (________21134));
  nor2s1 ____9__450660(.DIN1 (____9___20501), .DIN2 (___0_9__19844), .Q
       (___9____19692));
  nnd2s1 ______450661(.DIN1 (________19432), .DIN2 (____9___19107), .Q
       (________19964));
  nnd2s1 _______450662(.DIN1 (________19557), .DIN2 (________19431), .Q
       (________20454));
  or2s1 ______450663(.DIN1 (________20901), .DIN2 (____0___21724), .Q
       (____0___19953));
  nor2s1 _____0_450664(.DIN1 (________19518), .DIN2 (____9___19294), .Q
       (___0____19838));
  nor2s1 _____9_450665(.DIN1 (_____0__19068), .DIN2 (________19430), .Q
       (___0____19840));
  or2s1 _______450666(.DIN1 (________19128), .DIN2 (_____0__19429), .Q
       (________19893));
  nnd2s1 ______450667(.DIN1 (_____9__19428), .DIN2 (_____0__19124), .Q
       (_____0__19966));
  nor2s1 _______450668(.DIN1 (________19427), .DIN2 (________19426), .Q
       (___0____19841));
  or2s1 _______450669(.DIN1 (_____________________18608), .DIN2
       (____09__19601), .Q (________20309));
  nnd2s1 _______450670(.DIN1 (____0___19595), .DIN2 (________19425), .Q
       (________20057));
  and2s1 _______450671(.DIN1 (________19615), .DIN2
       (_____________________18615), .Q (____0___20514));
  and2s1 _____9_450672(.DIN1 (________19414), .DIN2
       (_____________________18602), .Q (____9___20319));
  nnd2s1 _______450673(.DIN1 (________19424), .DIN2
       (____0________________18647), .Q (_____0__20207));
  hi1s1 _______450674(.DIN (________19423), .Q (___9____23389));
  or2s1 _______450675(.DIN1 (____9___19298), .DIN2 (________19157), .Q
       (________20534));
  nor2s1 ____9__450676(.DIN1 (____09__19601), .DIN2 (_____9__19515), .Q
       (________21006));
  nor2s1 ____9_450677(.DIN1 (________19422), .DIN2 (________19421), .Q
       (_________30524));
  nnd2s1 _______450678(.DIN1 (________19413), .DIN2 (________19420), .Q
       (_____9__19965));
  or2s1 _______450679(.DIN1 (_____________________18623), .DIN2
       (_____0__19163), .Q (____9___19940));
  nnd2s1 ______450680(.DIN1 (___9____19733), .DIN2 (____0___19597), .Q
       (____0___21265));
  nnd2s1 ____9__450681(.DIN1 (_______19052), .DIN2 (____0___19597), .Q
       (________21319));
  nnd2s1 _______450682(.DIN1 (_____0__19449), .DIN2 (________19158), .Q
       (________22663));
  nnd2s1 ____9__450683(.DIN1 (________19444), .DIN2 (________19072), .Q
       (___0_09__27568));
  hi1s1 _______450684(.DIN (____0___19954), .Q (________21511));
  nnd2s1 _____0_450685(.DIN1 (________19424), .DIN2 (________19580), .Q
       (________21476));
  nor2s1 _____9_450686(.DIN1 (_____0__19419), .DIN2 (________19483), .Q
       (___90___21549));
  nor2s1 _____9_450687(.DIN1 (_____0__19419), .DIN2 (___0____19787), .Q
       (________21497));
  nnd2s1 _______450688(.DIN1 (________19130), .DIN2 (_____9__19418), .Q
       (_________29873));
  nnd2s1 _______450689(.DIN1 (___9____19694), .DIN2
       (_____________________18665), .Q (________20027));
  nor2s1 _______450690(.DIN1 (________19417), .DIN2 (________19483), .Q
       (____0___21267));
  nnd2s1 _______450691(.DIN1 (________19540), .DIN2 (________19416), .Q
       (________21879));
  nnd2s1 _______450692(.DIN1 (________19415), .DIN2 (_____0__19612), .Q
       (________20010));
  nnd2s1 ____9__450693(.DIN1 (____0_), .DIN2 (________19530), .Q
       (____9___21984));
  nnd2s1 _______450694(.DIN1 (________19414), .DIN2 (________19413), .Q
       (___9____20656));
  nnd2s1 _______450695(.DIN1 (________19194), .DIN2 (________19412), .Q
       (________20868));
  nor2s1 ______450696(.DIN1 (_____________________18635), .DIN2
       (________19445), .Q (_____0__20021));
  nnd2s1 _______450697(.DIN1 (________19545), .DIN2 (__99____27118), .Q
       (_________29858));
  nor2s1 _______450698(.DIN1 (________19444), .DIN2 (___9_9__19706), .Q
       (________20917));
  nor2s1 _____450699(.DIN1 (________19284), .DIN2 (________19411), .Q
       (________21794));
  nor2s1 _______450700(.DIN1 (________19150), .DIN2 (________19410), .Q
       (________21337));
  nor2s1 _______450701(.DIN1 (_____0__19409), .DIN2 (________20160), .Q
       (____9___21441));
  nor2s1 _______450702(.DIN1 (____09__19408), .DIN2 (________19555), .Q
       (____00__20510));
  nnd2s1 _______450703(.DIN1 (____0___19407), .DIN2
       (_____________________18634), .Q (________20461));
  nor2s1 ____9__450704(.DIN1 (____0___19406), .DIN2 (________20559), .Q
       (______0__30345));
  nnd2s1 ______450705(.DIN1 (________19434), .DIN2
       (______________________18671), .Q (________21730));
  nnd2s1 ____9__450706(.DIN1 (____0___19405), .DIN2 (________19615), .Q
       (___0____21651));
  and2s1 _______450707(.DIN1 (____0___19404), .DIN2
       (_____________________18626), .Q (____0___20041));
  nor2s1 _______450708(.DIN1 (____0________________18595), .DIN2
       (____0___19403), .Q (_____0__19918));
  nnd2s1 _______450709(.DIN1 (________19557), .DIN2 (____0___19402), .Q
       (____9___21900));
  or2s1 _______450710(.DIN1 (________19610), .DIN2 (________19470), .Q
       (___9____20666));
  nnd2s1 _______450711(.DIN1 (________19511), .DIN2
       (_____________________18665), .Q (____9___20037));
  nor2s1 ____9__450712(.DIN1 (________19523), .DIN2 (__909), .Q
       (___0____21684));
  hi1s1 _______450713(.DIN (_____0__20352), .Q (________21893));
  hi1s1 ______450714(.DIN (________21086), .Q (________21470));
  or2s1 ____90_450715(.DIN1 (____0___19504), .DIN2 (____9___19587), .Q
       (_____99__30363));
  nnd2s1 _______450716(.DIN1 (_____9__19448), .DIN2 (___0__18931), .Q
       (___9____21575));
  nnd2s1 ____9__450717(.DIN1 (________19270), .DIN2 (________19434), .Q
       (___0____21659));
  nnd2s1 _______450718(.DIN1 (________19412), .DIN2 (____0___19401), .Q
       (________21407));
  nor2s1 ____9__450719(.DIN1 (____0___21724), .DIN2 (________19513), .Q
       (___0____21677));
  hi1s1 _____9_450720(.DIN (_____0__23199), .Q (________23154));
  nor2s1 ____9__450721(.DIN1 (________19523), .DIN2 (_____9__19195), .Q
       (________22332));
  hi1s1 _______450722(.DIN (___9____19705), .Q (____9___21897));
  nnd2s1 _______450723(.DIN1 (________19574), .DIN2 (____00__19205), .Q
       (________21495));
  nor2s1 ____9__450724(.DIN1 (____9__19006), .DIN2 (___0__18931), .Q
       (_____0__22118));
  nnd2s1 ____9_450725(.DIN1 (____99__19398), .DIN2 (___0__18931), .Q
       (________22113));
  nor2s1 _______450726(.DIN1 (___0____19787), .DIN2 (________19417), .Q
       (________21776));
  nnd2s1 ______450727(.DIN1 (____9___19397), .DIN2 (____9___19396), .Q
       (_________33370));
  hi1s1 _____0_450728(.DIN (____9___19395), .Q (________23814));
  nnd2s1 _______450729(.DIN1 (________19553), .DIN2 (____9___19393), .Q
       (____9___19394));
  nor2s1 _______450730(.DIN1 (_____________________18615), .DIN2
       (_____0__19361), .Q (____9___19392));
  nor2s1 _______450731(.DIN1 (________19606), .DIN2 (___9____19756), .Q
       (____9___19391));
  nor2s1 ______450732(.DIN1 (________19258), .DIN2 (________19367), .Q
       (____90__19390));
  nnd2s1 _______450733(.DIN1 (_______19012), .DIN2 (inData[30]), .Q
       (_____9__19389));
  and2s1 _____0_450734(.DIN1 (________19536), .DIN2
       (______________0___________________), .Q (________19388));
  nor2s1 _____9_450735(.DIN1 (________19386), .DIN2 (________19470), .Q
       (________19387));
  nor2s1 _____0_450736(.DIN1 (____90__19292), .DIN2 (________19456), .Q
       (________19385));
  or2s1 _______450737(.DIN1 (________19383), .DIN2 (________19382), .Q
       (________19384));
  or2s1 ______450738(.DIN1 (____9___22253), .DIN2 (____9____30867), .Q
       (________19381));
  or2s1 _______450739(.DIN1 (_____________________18610), .DIN2
       (____09__19408), .Q (_____0__19380));
  xor2s1 _______450740(.DIN1 (_________32074), .DIN2 (________19378),
       .Q (_____9__19379));
  nor2s1 _______450741(.DIN1 (_____0__20069), .DIN2 (________19376), .Q
       (________19377));
  nnd2s1 _______450742(.DIN1 (___9____19733), .DIN2 (___9_0__19727), .Q
       (________19375));
  nor2s1 _______450743(.DIN1 (_____0__20392), .DIN2 (____0___19860), .Q
       (________19374));
  nnd2s1 _______450744(.DIN1 (____0___19406), .DIN2 (outData[25]), .Q
       (________19373));
  nor2s1 _______450745(.DIN1 (___9____19718), .DIN2 (___9____19710), .Q
       (________19372));
  and2s1 ______450746(.DIN1 (____0___19405), .DIN2 (________19410), .Q
       (_____0__19371));
  nnd2s1 _______450747(.DIN1 (________19369), .DIN2 (________19555), .Q
       (_____9__19370));
  nnd2s1 ______450748(.DIN1 (___9____19701), .DIN2 (________19367), .Q
       (________19368));
  nnd2s1 _______450749(.DIN1 (___0_9__19844), .DIN2 (outData[29]), .Q
       (________19366));
  and2s1 _______450750(.DIN1 (____0____33753), .DIN2 (___99), .Q
       (________19365));
  nor2s1 _______450751(.DIN1 (____0___19058), .DIN2 (___9____19749), .Q
       (________19364));
  nnd2s1 _______450752(.DIN1 (___9_9__19716), .DIN2 (________19277), .Q
       (________19363));
  or2s1 _____0_450753(.DIN1 (_____________________18614), .DIN2
       (_____0__19361), .Q (________19362));
  nnd2s1 _______450754(.DIN1 (_____9__19143), .DIN2 (____9___19586), .Q
       (_____9__19360));
  xnr2s1 ______450755(.DIN1 (_________9______18802), .DIN2
       (________19358), .Q (________19359));
  nor2s1 _______450756(.DIN1 (________19382), .DIN2 (________19337), .Q
       (________19357));
  nnd2s1 ____0__450757(.DIN1 (___9____20638), .DIN2 (____9__19041), .Q
       (________19356));
  xor2s1 _______450758(.DIN1 (______9__34490), .DIN2 (_______18963), .Q
       (________19355));
  nnd2s1 _____0_450759(.DIN1 (____0___19401), .DIN2 (________19353), .Q
       (________19354));
  or2s1 _______450760(.DIN1 (_____________0___18715), .DIN2
       (_____0__19351), .Q (________19352));
  and2s1 _______450761(.DIN1 (_______19022), .DIN2
       (_____________________18635), .Q (_____9__19350));
  nor2s1 _______450762(.DIN1 (___9_0__19727), .DIN2 (_______19049), .Q
       (________19349));
  nnd2s1 _____9_450763(.DIN1 (_____9__20078), .DIN2 (_______19019), .Q
       (________19348));
  nnd2s1 _____0_450764(.DIN1 (____9___19587), .DIN2 (___9___18953), .Q
       (________19347));
  nnd2s1 _______450765(.DIN1 (________19345), .DIN2 (____0___21453), .Q
       (________19346));
  nor2s1 _______450766(.DIN1 (________19343), .DIN2 (___9_9__19706), .Q
       (________19344));
  nnd2s1 _______450767(.DIN1 (____0___19404), .DIN2 (_______19048), .Q
       (________19342));
  nor2s1 _______450768(.DIN1 (_________________18693), .DIN2
       (_____9__19162), .Q (_____0__19341));
  hi1s1 ______450769(.DIN (________19339), .Q (_____9__19340));
  nnd2s1 _______450770(.DIN1 (________19337), .DIN2 (___0___18985), .Q
       (________19338));
  nor2s1 _______450771(.DIN1 (____0____________9_), .DIN2
       (_____9__20078), .Q (________19336));
  nor2s1 _______450772(.DIN1 (________19334), .DIN2 (________20073), .Q
       (________19335));
  or2s1 _______450773(.DIN1 (____0____________9___18654), .DIN2
       (____0___19504), .Q (________19333));
  nor2s1 _______450774(.DIN1 (_____0), .DIN2 (________20901), .Q
       (________19332));
  xor2s1 _______450775(.DIN1 (________19253), .DIN2 (______0__18865),
       .Q (_____0__19331));
  nnd2s1 _____9_450776(.DIN1 (________20072), .DIN2 (________19617), .Q
       (_____9__19330));
  and2s1 _______450777(.DIN1 (____00__19592), .DIN2 (________19328), .Q
       (________19329));
  nnd2s1 ______450778(.DIN1 (___9____19701), .DIN2 (________19436), .Q
       (________19327));
  or2s1 _______450779(.DIN1 (_____________________18604), .DIN2
       (________19325), .Q (________19326));
  or2s1 _____450780(.DIN1 (______________________18632), .DIN2
       (________19523), .Q (________19324));
  nnd2s1 ______450781(.DIN1 (____9___19293), .DIN2 (________19322), .Q
       (________19323));
  nor2s1 _______450782(.DIN1 (________19665), .DIN2 (_____9__19467), .Q
       (_____0__19321));
  xnr2s1 ______450783(.DIN1 (_________18859), .DIN2 (_____0__20962), .Q
       (_____9__19320));
  nnd2s1 _______450784(.DIN1 (________19103), .DIN2 (inData[10]), .Q
       (________19319));
  or2s1 ______450785(.DIN1 (________19456), .DIN2 (________19540), .Q
       (________19318));
  nor2s1 _______450786(.DIN1 (________19145), .DIN2 (________20073), .Q
       (________19317));
  nor2s1 ______450787(.DIN1 (____0________________18650), .DIN2
       (____9___21071), .Q (________19316));
  nnd2s1 _______450788(.DIN1 (___0_9__19825), .DIN2
       (______________________18632), .Q (________19315));
  nor2s1 ______450789(.DIN1 (____0________________18591), .DIN2
       (____0___19208), .Q (________19314));
  nnd2s1 _____0_450790(.DIN1 (____0___19055), .DIN2 (____99__19398), .Q
       (________19313));
  and2s1 ______450791(.DIN1 (____09__19311), .DIN2 (_______19017), .Q
       (_____0__19312));
  or2s1 _____9_450792(.DIN1 (________19069), .DIN2 (____0___19310), .Q
       (_________28305));
  nnd2s1 _______450793(.DIN1 (________19575), .DIN2
       (______________________18632), .Q (___09___19848));
  nnd2s1 _______450794(.DIN1 (___0_9__19844), .DIN2 (____0___19309), .Q
       (_____9__20180));
  and2s1 _______450795(.DIN1 (____0___19308), .DIN2 (________19071), .Q
       (___9____19720));
  dffacs1 ________________0_450796(.CLRB (reset), .CLK (clk), .DIN
       (_______19018), .QN (____________0_));
  nnd2s1 _______450797(.DIN1 (____0___21988), .DIN2 (____9___19198), .Q
       (________21059));
  nnd2s1 ______450798(.DIN1 (____0___19307), .DIN2
       (_____________________18604), .Q (___0____19796));
  nnd2s1 ______450799(.DIN1 (_______18994), .DIN2 (____0___19306), .Q
       (___9____19713));
  or2s1 _______450800(.DIN1 (____0___19305), .DIN2 (________19443), .Q
       (_____0__19975));
  nnd2s1 _______450801(.DIN1 (________19553), .DIN2 (________19266), .Q
       (________19913));
  hi1s1 _______450802(.DIN (___9_0__20644), .Q (___0____19842));
  nor2s1 _______450803(.DIN1 (_________________9___18606), .DIN2
       (________19435), .Q (____00__19852));
  nnd2s1 _____0_450804(.DIN1 (____0___19304), .DIN2 (____0___19303), .Q
       (_________28451));
  nnd2s1 _______450805(.DIN1 (________22684), .DIN2 (_______19001), .Q
       (_____9__23791));
  and2s1 _______450806(.DIN1 (_________30444), .DIN2 (___0___19034), .Q
       (___0____21689));
  nor2s1 _______450807(.DIN1 (_____________________18604), .DIN2
       (____00__19302), .Q (___9____19742));
  or2s1 _______450808(.DIN1 (____99__19301), .DIN2 (____9___19300), .Q
       (_________34004));
  nor2s1 _____0_450809(.DIN1 (____9___19299), .DIN2 (____9___19298), .Q
       (___9____19721));
  nor2s1 ____9__450810(.DIN1 (inData[30]), .DIN2 (________19218), .Q
       (________19570));
  nnd2s1 _______450811(.DIN1 (___0_9__19844), .DIN2 (inData[24]), .Q
       (________19999));
  nnd2s1 ____9__450812(.DIN1 (________19434), .DIN2 (____9___19297), .Q
       (________19613));
  nor2s1 _______450813(.DIN1 (________19287), .DIN2 (____9___19296), .Q
       (________20343));
  nor2s1 ______450814(.DIN1 (____9___19295), .DIN2 (___9_9__19706), .Q
       (________20833));
  and2s1 _______450815(.DIN1 (____0___19405), .DIN2
       (_____________________18612), .Q (___09___19850));
  nor2s1 ______450816(.DIN1 (________19430), .DIN2 (___9____19749), .Q
       (___9____19703));
  nor2s1 _______450817(.DIN1 (____99__19398), .DIN2 (________19442), .Q
       (___0____19828));
  nor2s1 _______450818(.DIN1 (________19437), .DIN2 (___9_9__19706), .Q
       (___999__21632));
  nnd2s1 ______450819(.DIN1 (___0_9__19844), .DIN2 (_________28766), .Q
       (___0____19804));
  nnd2s1 _______450820(.DIN1 (________19416), .DIN2 (________19155), .Q
       (_____9__19908));
  nor2s1 _______450821(.DIN1 (____0________________18595), .DIN2
       (____9___19294), .Q (________19919));
  nor2s1 _______450822(.DIN1 (___0____21699), .DIN2 (________22136), .Q
       (___9____19715));
  nnd2s1 ______450823(.DIN1 (________19461), .DIN2 (____9___19293), .Q
       (____9___19588));
  nor2s1 _______450824(.DIN1 (____90__19292), .DIN2 (_____9__20078), .Q
       (___0_0__19835));
  hi1s1 _______450825(.DIN (_________30807), .Q (___09_));
  nnd2s1 ______450826(.DIN1 (_____9__19291), .DIN2
       (______________________18630), .Q (___9_9__19744));
  nnd2s1 _____0_450827(.DIN1 (____00__19592), .DIN2 (_____9__19543), .Q
       (___9____19724));
  nor2s1 _______450828(.DIN1 (________19078), .DIN2 (____00__19592), .Q
       (___09___19846));
  and2s1 _______450829(.DIN1 (________19102), .DIN2
       (_____________________18665), .Q (________19902));
  nor2s1 _______450830(.DIN1 (_____________________18641), .DIN2
       (________19444), .Q (___0_9__19817));
  dffacs1 __________________450831(.CLRB (reset), .CLK (clk), .DIN
       (____0__18989), .Q (________________18674));
  or2s1 _____450832(.DIN1 (____0___21724), .DIN2 (___0____20722), .Q
       (___9_9__20681));
  nor2s1 _______450833(.DIN1 (________19290), .DIN2 (________19289), .Q
       (________19960));
  nnd2s1 _____0_450834(.DIN1 (________19413), .DIN2
       (_____________________18599), .Q (________20053));
  and2s1 _____450835(.DIN1 (________19549), .DIN2 (____0___19401), .Q
       (________20241));
  nnd2s1 _______450836(.DIN1 (____9___19393), .DIN2 (____0___19402), .Q
       (________20398));
  nor2s1 _____9_450837(.DIN1 (____09__19408), .DIN2 (____09__19601), .Q
       (___09___20784));
  nnd2s1 _______450838(.DIN1 (____9__19035), .DIN2 (________19288), .Q
       (____9____29953));
  nor2s1 _____0_450839(.DIN1 (________19287), .DIN2 (___9____19749), .Q
       (____90__20972));
  nor2s1 _______450840(.DIN1 (_____0__19956), .DIN2 (________19606), .Q
       (________21306));
  nnd2s1 ______450841(.DIN1 (________19286), .DIN2 (________19285), .Q
       (_____9__20381));
  nor2s1 _______450842(.DIN1 (________19284), .DIN2 (____9___19298), .Q
       (________21784));
  nnd2s1 _____9_450843(.DIN1 (________19545), .DIN2
       (_____________________18662), .Q (________20023));
  dffacs1 __________________450844(.CLRB (reset), .CLK (clk), .DIN
       (____0___19118), .QN (________________18673));
  nnd2s1 ______450845(.DIN1 (____0___19407), .DIN2 (________19996), .Q
       (________19864));
  nnd2s1 _____0_450846(.DIN1 (____00__19592), .DIN2 (________20091), .Q
       (____9___22438));
  nnd2s1 _____0_450847(.DIN1 (____9___19587), .DIN2 (________19283), .Q
       (________20019));
  nor2s1 _______450848(.DIN1 (______________________18671), .DIN2
       (____0___19600), .Q (________22292));
  nnd2s1 _____9_450849(.DIN1 (____90__19582), .DIN2 (________19472), .Q
       (___9____20665));
  nor2s1 _______450850(.DIN1 (___9____19729), .DIN2 (___99___19765), .Q
       (____0___19949));
  or2s1 _____450851(.DIN1 (_____________________18625), .DIN2
       (___99___19765), .Q (____0___19950));
  nor2s1 ____9__450852(.DIN1 (_____0__19282), .DIN2 (_____9__19281), .Q
       (________20110));
  nor2s1 _____0_450853(.DIN1 (____0________________18653), .DIN2
       (________19606), .Q (________19963));
  nnd2s1 _____9_450854(.DIN1 (_____0__19506), .DIN2 (_____9), .Q
       (____9___19938));
  nor2s1 _______450855(.DIN1 (______18933), .DIN2 (________19483), .Q
       (___9_9__20623));
  nor2s1 _______450856(.DIN1 (___9____19712), .DIN2 (________19265), .Q
       (________21025));
  nor2s1 _____450857(.DIN1 (_____9__21513), .DIN2 (___0____20746), .Q
       (________20209));
  nor2s1 _____0_450858(.DIN1 (____9___19296), .DIN2 (___9____19697), .Q
       (________20208));
  nor2s1 _______450859(.DIN1 (_____0__19409), .DIN2 (_____0__19144), .Q
       (____90__20410));
  nor2s1 _____0_450860(.DIN1 (____9___19296), .DIN2 (________19430), .Q
       (________20355));
  nnd2s1 _______450861(.DIN1 (____9___19295), .DIN2 (___0___18988), .Q
       (_________28593));
  nor2s1 ______450862(.DIN1 (________19280), .DIN2 (________19279), .Q
       (_____0___29178));
  nor2s1 _______450863(.DIN1 (________19278), .DIN2 (________19442), .Q
       (_____9__20499));
  and2s1 _____9_450864(.DIN1 (_____0__19449), .DIN2 (________19424), .Q
       (________21922));
  nor2s1 _____0_450865(.DIN1 (________19577), .DIN2 (_____0__19361), .Q
       (________20593));
  nnd2s1 _______450866(.DIN1 (________19277), .DIN2 (________19413), .Q
       (________20387));
  nor2s1 _______450867(.DIN1 (________19276), .DIN2 (________19275), .Q
       (_________28601));
  nnd2s1 _____450868(.DIN1 (________19540), .DIN2
       (____0_______________), .Q (____0___19948));
  nnd2s1 _______450869(.DIN1 (________19274), .DIN2 (_____9__19543), .Q
       (________20261));
  nor2s1 ______450870(.DIN1 (________19523), .DIN2 (____0___19860), .Q
       (________20543));
  nnd2s1 _______450871(.DIN1 (___9____19756), .DIN2 (________19608), .Q
       (____0___21263));
  hi1s1 _______450872(.DIN (_________31702), .Q (_________31587));
  nor2s1 _______450873(.DIN1 (_____0__19282), .DIN2 (___9____21610), .Q
       (________20380));
  nor2s1 _______450874(.DIN1 (____0___19860), .DIN2 (____9___19199), .Q
       (____9___21256));
  nnd2s1 _______450875(.DIN1 (____00__19592), .DIN2 (________19151), .Q
       (___9_9__20662));
  nnd2s1 _______450876(.DIN1 (________19148), .DIN2 (________19530), .Q
       (________20850));
  nor2s1 _______450877(.DIN1 (_____9__21513), .DIN2 (___9____19710), .Q
       (________19915));
  nnd2s1 _______450878(.DIN1 (____9___19393), .DIN2 (________19431), .Q
       (_____9__20846));
  nor2s1 _______450879(.DIN1 (________19273), .DIN2 (________19456), .Q
       (________21518));
  nor2s1 _______450880(.DIN1 (________19376), .DIN2 (_____9__19467), .Q
       (________20497));
  hi1s1 _______450881(.DIN (________19607), .Q (_____0__21191));
  nnd2s1 ______450882(.DIN1 (________19461), .DIN2 (________19645), .Q
       (________20821));
  nnd2s1 _____0_450883(.DIN1 (_____0__19272), .DIN2 (___00__19033), .Q
       (____0___20046));
  or2s1 _______450884(.DIN1 (_____9__19271), .DIN2 (___9_0__19717), .Q
       (_____9__21229));
  nnd2s1 _______450885(.DIN1 (____00__19592), .DIN2 (________19161), .Q
       (___90___20608));
  nnd2s1 ____9__450886(.DIN1 (________19270), .DIN2 (____9___19589), .Q
       (________21471));
  nor2s1 _______450887(.DIN1 (___9____19712), .DIN2 (________19269), .Q
       (________21777));
  nnd2s1 _______450888(.DIN1 (________19268), .DIN2 (_______19044), .Q
       (___90___23353));
  nnd2s1 _______450889(.DIN1 (________19416), .DIN2
       (____0____________9_), .Q (_____9__20283));
  nor2s1 ____9__450890(.DIN1 (_____9__19271), .DIN2 (____9___21071), .Q
       (________22129));
  nor2s1 ______450891(.DIN1 (____0___19600), .DIN2 (________19269), .Q
       (_____9__22147));
  nor2s1 _______450892(.DIN1 (_____0__19282), .DIN2 (____9___21071), .Q
       (________20809));
  nnd2s1 ____9__450893(.DIN1 (________19267), .DIN2 (________19165), .Q
       (______9__28887));
  nnd2s1 _______450894(.DIN1 (________19575), .DIN2 (________21824), .Q
       (___9____20651));
  nnd2s1 ____9_450895(.DIN1 (____0___19405), .DIN2 (____90__19582), .Q
       (___0____21660));
  nnd2s1 ____90_450896(.DIN1 (________19431), .DIN2 (________19266), .Q
       (____9___21980));
  nor2s1 _____9_450897(.DIN1 (________19265), .DIN2 (____0___19600), .Q
       (________22141));
  nor2s1 ____9__450898(.DIN1 (________19264), .DIN2 (________19263), .Q
       (___99___22527));
  nor2s1 _____450899(.DIN1 (________19149), .DIN2 (____9___19298), .Q
       (___0____21694));
  nor2s1 _______450900(.DIN1 (________19617), .DIN2 (________20160), .Q
       (________20003));
  nnd2s1 _______450901(.DIN1 (_____0__19262), .DIN2 (_____9__19105), .Q
       (_________30710));
  nor2s1 _______450902(.DIN1 (_____9__19261), .DIN2 (________20160), .Q
       (___9____20684));
  nor2s1 _______450903(.DIN1 (________19435), .DIN2 (________19367), .Q
       (_____9__21287));
  nor2s1 _____0_450904(.DIN1 (________19060), .DIN2 (_____9__19515), .Q
       (________20872));
  nor2s1 ____9_450905(.DIN1 (_____9__19271), .DIN2 (___9____21610), .Q
       (________21774));
  or2s1 ____9__450906(.DIN1 (________20901), .DIN2 (_____9__22215), .Q
       (________21310));
  nnd2s1 _____0_450907(.DIN1 (____0___19307), .DIN2 (___9____19700), .Q
       (_____9__20557));
  nor2s1 ____9__450908(.DIN1 (________19260), .DIN2 (________20564), .Q
       (________21222));
  nor2s1 _______450909(.DIN1 (_____0__19409), .DIN2 (________19643), .Q
       (_____0__21504));
  and2s1 _____9_450910(.DIN1 (____9___19589), .DIN2 (________19433), .Q
       (_____0__21821));
  nnd2s1 _____9_450911(.DIN1 (____0___19504), .DIN2
       (____0____________9___18654), .Q (_____0__20362));
  nnd2s1 _____0_450912(.DIN1 (________19645), .DIN2 (________19322), .Q
       (________21472));
  and2s1 ____9__450913(.DIN1 (____0___19307), .DIN2 (___9____19701), .Q
       (____9___21070));
  nnd2s1 _____0_450914(.DIN1 (________20072), .DIN2 (________19608), .Q
       (________21505));
  hi1s1 _____450915(.DIN (________19259), .Q (________21409));
  and2s1 ____9__450916(.DIN1 (___9____19701), .DIN2 (________19229), .Q
       (________21203));
  nor2s1 ____9__450917(.DIN1 (_____9__19271), .DIN2 (_____9__19281), .Q
       (________22339));
  nor2s1 _______450918(.DIN1 (________19258), .DIN2 (________19325), .Q
       (________21397));
  hi1s1 _____9_450919(.DIN (________19257), .Q (___9____19725));
  and2s1 ____9_450920(.DIN1 (_____0__19449), .DIN2 (___900__20605), .Q
       (____0____29098));
  hi1s1 _____9_450921(.DIN (____0___19400), .Q (___00___22540));
  ib1s1 _____450922(.DIN (____00__19399), .Q (________24221));
  and2s1 _______450923(.DIN1 (___9__), .DIN2
       (_____________________18622), .Q (________19256));
  or2s1 _______450924(.DIN1 (_____________________18614), .DIN2
       (________19410), .Q (________19255));
  or2s1 _______450925(.DIN1 (___0_), .DIN2 (________19253), .Q
       (________19254));
  nnd2s1 _____9_450926(.DIN1 (______18937), .DIN2 (_________34472), .Q
       (_____0__19252));
  hi1s1 ______450927(.DIN (___0____22594), .Q (_____9__19251));
  nor2s1 _____9_450928(.DIN1 (____________________), .DIN2
       (____9___19586), .Q (________19250));
  nnd2s1 _____9_450929(.DIN1 (________19425), .DIN2
       (____0________________18595), .Q (________19249));
  hi1s1 _______450930(.DIN (________19247), .Q (________19248));
  and2s1 _______450931(.DIN1 (________19245), .DIN2 (________19576), .Q
       (________19246));
  nnd2s1 _______450932(.DIN1 (___9__), .DIN2 (________19156), .Q
       (________19244));
  hi1s1 ____00_450933(.DIN (________19444), .Q (_____0__19243));
  hi1s1 ____9__450934(.DIN (________19241), .Q (_____9__19242));
  xor2s1 _____0_450935(.DIN1 (________19239), .DIN2 (_________34444),
       .Q (________19240));
  nnd2s1 _______450936(.DIN1 (___9____19752), .DIN2 (_____0__19612), .Q
       (________19238));
  nor2s1 _______450937(.DIN1 (outData[6]), .DIN2 (___0__18935), .Q
       (________19237));
  or2s1 _______450938(.DIN1 (_____________________18615), .DIN2
       (________19410), .Q (________19235));
  hi1s1 _______450939(.DIN (_____9__19233), .Q (_____0__19234));
  xor2s1 _____9_450940(.DIN1 (outData[17]), .DIN2 (________19231), .Q
       (________19232));
  nnd2s1 _____450941(.DIN1 (________19229), .DIN2 (___9____19700), .Q
       (________19230));
  xor2s1 _______450942(.DIN1 (_____________18894), .DIN2
       (__99____27109), .Q (________19228));
  nnd2s1 _______450943(.DIN1 (________19226), .DIN2 (______18929), .Q
       (________19227));
  xor2s1 ______450944(.DIN1 (_____9__19224), .DIN2 (_____0___34424), .Q
       (_____0__19225));
  and2s1 _______450945(.DIN1 (________19620), .DIN2
       (_____________________18620), .Q (________19223));
  xor2s1 _______450946(.DIN1 (________19221), .DIN2
       (_________________18766), .Q (________19222));
  or2s1 _______450947(.DIN1 (_________18847), .DIN2 (________23232), .Q
       (________19220));
  hi1s1 ____9__450948(.DIN (________19218), .Q (________19219));
  or2s1 _______450949(.DIN1
       (______________0______________________18825), .DIN2
       (______18936), .Q (________19217));
  hi1s1 _______450950(.DIN (_____9__19261), .Q (____0___19593));
  hi1s1 ______450951(.DIN (________19216), .Q (___0_____28026));
  nnd2s1 ______450952(.DIN1 (____9_), .DIN2 (________19610), .Q
       (_____0__19622));
  and2s1 ______450953(.DIN1 (_____0__19215), .DIN2 (________19580), .Q
       (________19257));
  nnd2s1 _______450954(.DIN1 (________19264), .DIN2 (________19154), .Q
       (____9___19395));
  nnd2s1 ______450955(.DIN1 (____09__19214), .DIN2 (____0___19213), .Q
       (____9___19495));
  hi1s1 ____9__450956(.DIN (____00__19302), .Q (___9____19702));
  hi1s1 _______450957(.DIN (________19415), .Q (________19663));
  nor2s1 _______450958(.DIN1 (_____________________18621), .DIN2
       (___9___18977), .Q (________19526));
  hi1s1 ____9__450959(.DIN (____0___19212), .Q (________19604));
  hi1s1 ____9__450960(.DIN (________19284), .Q (________19573));
  hi1s1 ____9_450961(.DIN (____0___19403), .Q (____0___19596));
  hi1s1 ____9__450962(.DIN (____0___19211), .Q (________21917));
  nor2s1 ____9__450963(.DIN1 (________19577), .DIN2 (________19410), .Q
       (________19259));
  hi1s1 _______450964(.DIN (____0___19210), .Q (________19603));
  hi1s1 ____9_450965(.DIN (________19905), .Q (_____0__19669));
  hi1s1 ____99_450966(.DIN (____9___19293), .Q (___9____19693));
  nor2s1 _______450967(.DIN1 (____0________________18595), .DIN2
       (_______18961), .Q (____00__20226));
  hi1s1 _______450968(.DIN (____0___19209), .Q (___0_0__19810));
  or2s1 _______450969(.DIN1 (inData[30]), .DIN2 (________19193), .Q
       (____00__19399));
  hi1s1 ____00_450970(.DIN (________19437), .Q (___9____19728));
  hi1s1 ____9_450971(.DIN (____0___19208), .Q (___9____19696));
  hi1s1 ____00_450972(.DIN (________19441), .Q (_________28734));
  nor2s1 _____0_450973(.DIN1 (____0______________), .DIN2
       (____0___19057), .Q (________19607));
  and2s1 _____9_450974(.DIN1 (________19245), .DIN2
       (____0_______________), .Q (________20395));
  hi1s1 ____9__450975(.DIN (____0___19207), .Q (___0____19800));
  xor2s1 ____9__450976(.DIN1 (_________9___18903), .DIN2 (outData[31]),
       .Q (_________30807));
  or2s1 ______450977(.DIN1 (______________________18617), .DIN2
       (____9___19586), .Q (________21468));
  hi1s1 ____0__450978(.DIN (_____0__19361), .Q (___9____19714));
  hi1s1 ____99_450979(.DIN (____0___19206), .Q (___9____19732));
  nnd2s1 _______450980(.DIN1 (_____0__19602), .DIN2 (____00__19205), .Q
       (________21492));
  hi1s1 ____0__450981(.DIN (________19557), .Q (________21857));
  hi1s1 _____9_450982(.DIN (____99__19204), .Q (___9____19711));
  hi1s1 _____450983(.DIN (____9___19203), .Q (___9_0__19707));
  hi1s1 ____450984(.DIN (____9___19202), .Q (_____0__20002));
  hi1s1 ____0__450985(.DIN (_____9__22215), .Q (_____0__21885));
  hi1s1 ______450986(.DIN (____9___19200), .Q (________21197));
  hi1s1 _____450987(.DIN (____9___19201), .Q (____9___20413));
  hi1s1 ____0__450988(.DIN (________19337), .Q (___9____19719));
  hi1s1 _____450989(.DIN (____9___19199), .Q (________19978));
  hi1s1 _____0_450990(.DIN (____9___19198), .Q (____9___21898));
  hi1s1 _______450991(.DIN (________19547), .Q (___9_0__19737));
  hi1s1 ____0_450992(.DIN (________21889), .Q (________21797));
  hi1s1 ______450993(.DIN (___9____19710), .Q (____0___20330));
  hi1s1 ____0__450994(.DIN (_____9__19281), .Q (___0____19783));
  hi1s1 ____0__450995(.DIN (____9___19197), .Q (___0____19815));
  hi1s1 _______450996(.DIN (____90__19196), .Q (_________28828));
  nor2s1 _______450997(.DIN1 (_____0__20382), .DIN2 (_____0__19282), .Q
       (______9__33436));
  hi1s1 ____0__450998(.DIN (_____9__19195), .Q (________21241));
  hi1s1 ____0__450999(.DIN (________19194), .Q (_____0___32299));
  nor2s1 _______451000(.DIN1 (_____________________18661), .DIN2
       (_____________________18662), .Q (_________31702));
  nor2s1 _______451001(.DIN1 (________19193), .DIN2 (________19264), .Q
       (_____0__23199));
  nnd2s1 _______451002(.DIN1 (____9___20501), .DIN2 (____09), .Q
       (_________34295));
  xor2s1 _______451003(.DIN1 (________19191), .DIN2
       (________________18787), .Q (________19192));
  xor2s1 ______451004(.DIN1 (_________________18730), .DIN2
       (____0___21449), .Q (________19190));
  and2s1 _______451005(.DIN1 (________19369), .DIN2
       (_____________________18611), .Q (________19189));
  nor2s1 _______451006(.DIN1 (_____9__19186), .DIN2 (________21366), .Q
       (_____0__19187));
  nnd2s1 _______451007(.DIN1 (___9__), .DIN2 (________19184), .Q
       (________19185));
  and2s1 _______451008(.DIN1 (________19369), .DIN2
       (_____________________18610), .Q (________19183));
  hi1s1 ____99_451009(.DIN (________19615), .Q (________19182));
  nor2s1 _______451010(.DIN1 (________19436), .DIN2 (________19258), .Q
       (________19181));
  nor2s1 _______451011(.DIN1 (________19617), .DIN2 (________19643), .Q
       (________19180));
  or2s1 _______451012(.DIN1 (_____________________18603), .DIN2
       (_____9__19177), .Q (________19179));
  nor2s1 _______451013(.DIN1 (_____0___34426), .DIN2 (_____), .Q
       (________19178));
  xor2s1 _____451014(.DIN1 (outData[8]), .DIN2 (__909___26328), .Q
       (________19176));
  xor2s1 _______451015(.DIN1 (___________0___18883), .DIN2
       (____0____31818), .Q (________19175));
  or2s1 _______451016(.DIN1 (_____________________18613), .DIN2
       (________19577), .Q (________19174));
  xor2s1 _______451017(.DIN1 (________19172), .DIN2
       (_________________18792), .Q (________19173));
  nor2s1 _______451018(.DIN1 (________19463), .DIN2 (________19610), .Q
       (________19171));
  nor2s1 _______451019(.DIN1 (________19463), .DIN2 (_____9__19169), .Q
       (_____0__19170));
  xor2s1 _______451020(.DIN1 (________19167), .DIN2
       (_________9______18800), .Q (________19168));
  nnd2s1 _______451021(.DIN1 (______18944), .DIN2 (____0___21991), .Q
       (________19166));
  xor2s1 _______451022(.DIN1 (outData[23]), .DIN2 (outData[24]), .Q
       (________19164));
  hi1s1 ____9__451023(.DIN (_____0__19163), .Q (____9___19585));
  hi1s1 ____9__451024(.DIN (________19325), .Q (_____0__19572));
  hi1s1 ____9__451025(.DIN (_____9__19162), .Q (________19661));
  and2s1 _______451026(.DIN1 (________19620), .DIN2
       (_____________________18621), .Q (___9_0));
  nnd2s1 _______451027(.DIN1 (________19161), .DIN2
       (_____________________18641), .Q (________19566));
  nnd2s1 _______451028(.DIN1 (________19160), .DIN2 (_______18965), .Q
       (________19423));
  hi1s1 ____99_451029(.DIN (________19472), .Q (_____9__19571));
  hi1s1 ____0__451030(.DIN (________19483), .Q (____99__19591));
  hi1s1 _______451031(.DIN (________19159), .Q (_________28762));
  and2s1 _______451032(.DIN1 (____9___20501), .DIN2
       (____0_________________18659), .Q (____9___19590));
  nor2s1 _______451033(.DIN1 (____0___21991), .DIN2 (_______18964), .Q
       (________19631));
  nnd2s1 _______451034(.DIN1 (________19645), .DIN2
       (_____________________18610), .Q (_____9__19458));
  hi1s1 _______451035(.DIN (________19158), .Q (________19579));
  hi1s1 ____9__451036(.DIN (________19157), .Q (____9___19584));
  nor2s1 _______451037(.DIN1 (________19386), .DIN2 (_____9__19169), .Q
       (________19605));
  nnd2s1 _______451038(.DIN1 (________19620), .DIN2 (________19156), .Q
       (________19339));
  hi1s1 _____9_451039(.DIN (________19414), .Q (___00___19772));
  or2s1 _____9_451040(.DIN1 (________19369), .DIN2 (________19645), .Q
       (___9____19735));
  hi1s1 ____9__451041(.DIN (________19155), .Q (___90___19688));
  nnd2s1 ____451042(.DIN1 (_______18970), .DIN2 (________19161), .Q
       (____0___19954));
  hi1s1 ____99_451043(.DIN (________20123), .Q (________19879));
  hi1s1 ____451044(.DIN (________19269), .Q (____0___19599));
  hi1s1 _____9_451045(.DIN (____90__20126), .Q (_____9__19611));
  nnd2s1 _______451046(.DIN1 (________19154), .DIN2 (inData[30]), .Q
       (____0___19400));
  nor2s1 _______451047(.DIN1 (_____________________18599), .DIN2
       (_____9__19169), .Q (____09__20235));
  nnd2s1 _____9_451048(.DIN1 (_____0__19153), .DIN2 (_______18968), .Q
       (__9__0__26618));
  nor2s1 _______451049(.DIN1 (____9___19488), .DIN2 (________19258), .Q
       (___9____19722));
  hi1s1 _______451050(.DIN (________20374), .Q (___0____19805));
  nnd2s1 _______451051(.DIN1 (_____0__19872), .DIN2 (_____9__21513), .Q
       (___0_0));
  nnd2s1 ____9__451052(.DIN1 (___9__), .DIN2 (___0__18931), .Q
       (___9____19705));
  nnd2s1 _______451053(.DIN1 (_____9__19152), .DIN2 (_____0__22063), .Q
       (________20292));
  hi1s1 ____00_451054(.DIN (____9___19297), .Q (___9____21568));
  nor2s1 ______451055(.DIN1 (_______18972), .DIN2 (________19577), .Q
       (___9____21624));
  nnd2s1 ____9__451056(.DIN1 (________19645), .DIN2 (____99), .Q
       (________21086));
  hi1s1 ____451057(.DIN (________19277), .Q (___9____19723));
  hi1s1 ____9__451058(.DIN (________19151), .Q (____0___19594));
  hi1s1 ____99_451059(.DIN (________19150), .Q (___9____19699));
  nor2s1 _______451060(.DIN1 (________19149), .DIN2 (________19411), .Q
       (___9_0__20644));
  nnd2s1 _______451061(.DIN1 (_____9__19152), .DIN2
       (_____________________18668), .Q (________21021));
  hi1s1 ____99_451062(.DIN (________19148), .Q (___9____19691));
  nnd2s1 _______451063(.DIN1 (________19146), .DIN2 (________19577), .Q
       (_____9__19638));
  xor2s1 ____9_451064(.DIN1 (____________18893), .DIN2 (__909___26328),
       .Q (_________28979));
  hi1s1 ____00_451065(.DIN (________20200), .Q (___90___21546));
  hi1s1 ____0__451066(.DIN (________19461), .Q (___000));
  hi1s1 ____00_451067(.DIN (________19147), .Q (___0____19822));
  hi1s1 ____0__451068(.DIN (________19270), .Q (_____0__21429));
  nor2s1 _____9_451069(.DIN1 (________19410), .DIN2 (________19146), .Q
       (________21216));
  hi1s1 _____451070(.DIN (________19145), .Q (___9____19695));
  nnd2s1 _______451071(.DIN1 (____0___19402), .DIN2 (________19266), .Q
       (________21862));
  hi1s1 ____0__451072(.DIN (___9____20638), .Q (___99___19769));
  nnd2s1 _______451073(.DIN1 (_____0__19215), .DIN2
       (____0________________18647), .Q (_____0__20352));
  or2s1 ____90_451074(.DIN1 (________19617), .DIN2 (_____9__19891), .Q
       (_____0__20274));
  hi1s1 ____0__451075(.DIN (________20160), .Q (_____9__20313));
  hi1s1 _____0_451076(.DIN (_____0__19144), .Q (________19655));
  hi1s1 ____0__451077(.DIN (___9____19756), .Q (___9____19739));
  hi1s1 ____0__451078(.DIN (____9___19397), .Q (_____0___33489));
  hi1s1 ____0__451079(.DIN (_____9__19143), .Q (___0____19789));
  hi1s1 ____0__451080(.DIN (_____9__19291), .Q (_____0__21298));
  hi1s1 ____0_451081(.DIN (________19274), .Q (________20007));
  nnd2s1 _______451082(.DIN1 (_____0__19282), .DIN2 (_____0__20382), .Q
       (_________34071));
  hi1s1 ____0__451083(.DIN (________19513), .Q (________20213));
  hi1s1 _______451084(.DIN (_____9__19668), .Q (________22131));
  nor2s1 ____0__451085(.DIN1 (________19141), .DIN2
       (_____________________18611), .Q (________19142));
  nor2s1 ______451086(.DIN1 (________19067), .DIN2 (________19139), .Q
       (________19140));
  nor2s1 ______451087(.DIN1 (______9__30537), .DIN2 (_________31281),
       .Q (________19138));
  nnd2s1 _______451088(.DIN1 (____0____28155), .DIN2 (inData[28]), .Q
       (________19137));
  xor2s1 ______451089(.DIN1 (_________9_______18812), .DIN2
       (_________9_______18810), .Q (________19136));
  xor2s1 _______451090(.DIN1 (_____0___34429), .DIN2 (______0__18849),
       .Q (________19135));
  nnd2s1 _______451091(.DIN1 (_________33530), .DIN2 (inData[30]), .Q
       (_____0__19134));
  nnd2s1 _____0_451092(.DIN1 (______18925), .DIN2
       (_________________18783), .Q (_____9__19133));
  nor2s1 ____0__451093(.DIN1 (___9____25205), .DIN2 (outData[3]), .Q
       (________19132));
  hi1s1 _______451094(.DIN (________19130), .Q (________19131));
  xor2s1 _______451095(.DIN1 (_________18864), .DIN2
       (_________________18683), .Q (________19129));
  nor2s1 _______451096(.DIN1 (_____0__19612), .DIN2 (________19617), .Q
       (________19128));
  nnd2s1 ______451097(.DIN1 (____0____31818), .DIN2 (_________31388),
       .Q (________19127));
  xor2s1 ______451098(.DIN1
       (______________0______________________18824), .DIN2
       (_________34487), .Q (________19126));
  nnd2s1 ______451099(.DIN1 (_________33835), .DIN2 (_________31388),
       .Q (________19125));
  hi1s1 _______451100(.DIN (____09__19123), .Q (_____0__19124));
  and2s1 _____0_451101(.DIN1 (_________34477), .DIN2 (____09__21084),
       .Q (____0___19122));
  and2s1 ____0__451102(.DIN1 (outData[3]), .DIN2 (___9____25205), .Q
       (____0___19121));
  nor2s1 _______451103(.DIN1 (_________31388), .DIN2 (_________33835),
       .Q (____0___19120));
  or2s1 ____0__451104(.DIN1 (____0_____________0___18655), .DIN2
       (_____0__20382), .Q (____0___19119));
  nor2s1 _______451105(.DIN1 (______________18871), .DIN2
       (_________________0___18660), .Q (____0___19118));
  nor2s1 ____0__451106(.DIN1 (_________34496), .DIN2 (____0___19116),
       .Q (____0___19117));
  nor2s1 ____0__451107(.DIN1 (____00__19114), .DIN2 (____99__19113), .Q
       (____0___19115));
  nor2s1 _____0_451108(.DIN1 (outData[19]), .DIN2 (outData[21]), .Q
       (____9___19112));
  nnd2s1 ____0__451109(.DIN1 (_____________________18599), .DIN2
       (________19386), .Q (____9___19111));
  nnd2s1 _______451110(.DIN1 (______0__30564), .DIN2 (____9___19109),
       .Q (____9___19110));
  nnd2s1 ______451111(.DIN1 (_____________________18664), .DIN2
       (___9____19718), .Q (____9___19108));
  hi1s1 ______451112(.DIN (____9___19106), .Q (____9___19107));
  nnd2s1 _______451113(.DIN1 (___________0___18883), .DIN2
       (____0____31818), .Q (____90));
  hi1s1 ______451114(.DIN (________19104), .Q (_____9__19105));
  nnd2s1 _______451115(.DIN1 (_________29646), .DIN2
       (_______________0___________________), .Q (________19103));
  nor2s1 _______451116(.DIN1 (___9____19718), .DIN2 (_____0__22063), .Q
       (________19102));
  hi1s1 ____9__451117(.DIN (________19100), .Q (________19101));
  nnd2s1 ______451118(.DIN1 (________19064), .DIN2 (________19098), .Q
       (________19099));
  nnd2s1 _____9_451119(.DIN1
       (______________________________________0_____________18887),
       .DIN2 (_________30612), .Q (________19097));
  nor2s1 ______451120(.DIN1 (_________31388), .DIN2 (____0____31818),
       .Q (_____0__19096));
  nor2s1 _____451121(.DIN1 (____9____29052), .DIN2
       (______________________________________0__________0__18892), .Q
       (_____9__19095));
  nor2s1 ____0__451122(.DIN1 (outData[29]), .DIN2 (_____________18905),
       .Q (________19094));
  nnd2s1 _______451123(.DIN1 (_________31281), .DIN2
       (_________9_______18806), .Q (________19093));
  nnd2s1 ______451124(.DIN1 (_________30491), .DIN2 (inData[6]), .Q
       (________19092));
  nor2s1 _______451125(.DIN1
       (______________________________________0__________0), .DIN2
       (_________28939), .Q (________19091));
  xor2s1 _____0_451126(.DIN1 (_________34478), .DIN2
       (_________________18696), .Q (________19090));
  or2s1 _______451127(.DIN1 (_____09__31192), .DIN2
       (________________18787), .Q (________19089));
  xor2s1 _______451128(.DIN1 (_________________18727), .DIN2
       (______0__34461), .Q (________19088));
  nor2s1 _______451129(.DIN1 (outData[14]), .DIN2 (outData[16]), .Q
       (________19087));
  xor2s1 _____9_451130(.DIN1 (_________________18797), .DIN2
       (___________________________________), .Q (_____0__19086));
  nor2s1 _____0_451131(.DIN1 (________19231), .DIN2
       (_____________18897), .Q (_____9__19085));
  nor2s1 _______451132(.DIN1 (outData[6]), .DIN2 (outData[8]), .Q
       (________19084));
  nor2s1 _______451133(.DIN1 (inData[2]), .DIN2 (__99____27118), .Q
       (________19083));
  nnd2s1 ____0__451134(.DIN1 (_____________9___18751), .DIN2
       (______18916), .Q (________19082));
  nor2s1 _______451135(.DIN1 (____0____31818), .DIN2
       (___________0___18883), .Q (________19081));
  xnr2s1 _____0_451136(.DIN1 (_________34452), .DIN2 (______0__34451),
       .Q (________19080));
  nor2s1 _____0_451137(.DIN1 (_____9__23665), .DIN2
       (_________________18792), .Q (________19079));
  nor2s1 _______451138(.DIN1 (________19077), .DIN2 (________20091), .Q
       (________19078));
  and2s1 ____0_451139(.DIN1 (__99____27118), .DIN2
       (_____________________18661), .Q (________19076));
  nor2s1 _______451140(.DIN1 (outData[30]), .DIN2 (_____________18902),
       .Q (________19075));
  xor2s1 _______451141(.DIN1 (_________34445), .DIN2
       (_____________0___18759), .Q (________19074));
  nnd2s1 _______451142(.DIN1
       (______________________________________0_____________18889),
       .DIN2 (___9___18981), .Q (________19073));
  or2s1 ____0__451143(.DIN1 (________19139), .DIN2
       (_____________________18640), .Q (________19072));
  nnd2s1 _______451144(.DIN1 (_______________18880), .DIN2
       (_____00__30456), .Q (________19071));
  nnd2s1 ____0__451145(.DIN1 (_____________________18609), .DIN2
       (______18922), .Q (________19070));
  and2s1 ____0__451146(.DIN1 (outData[4]), .DIN2 (outData[6]), .Q
       (________19069));
  nnd2s1 _______451147(.DIN1 (outData[3]), .DIN2 (___99___20691), .Q
       (________19454));
  nor2s1 _______451148(.DIN1 (outData[28]), .DIN2 (_____________18901),
       .Q (________19614));
  nor2s1 _______451149(.DIN1 (_________9_____), .DIN2 (______9__30537),
       .Q (________19188));
  nor2s1 _______451150(.DIN1 (_____0__19068), .DIN2
       (____________________), .Q (_____9__19143));
  nor2s1 _____451151(.DIN1 (____________________________________18836),
       .DIN2 (____0____31818), .Q (________19450));
  nnd2s1 ______451152(.DIN1 (outData[5]), .DIN2 (outData[7]), .Q
       (________19440));
  nor2s1 _______451153(.DIN1 (outData[12]), .DIN2 (outData[10]), .Q
       (________19958));
  nor2s1 _____9_451154(.DIN1 (________19996), .DIN2
       (_____________________18636), .Q (____0___19207));
  nor2s1 _____0_451155(.DIN1 (_____0__22063), .DIN2
       (_____________________18666), .Q (____99__19204));
  nnd2s1 _______451156(.DIN1 (___0__18921), .DIN2 (inData[31]), .Q
       (____0___19211));
  nnd2s1 ____09_451157(.DIN1 (________19231), .DIN2 (outData[14]), .Q
       (____0___19306));
  nor2s1 _______451158(.DIN1 (______18924), .DIN2
       (_________________18696), .Q (___9____19746));
  nor2s1 ______451159(.DIN1 (_____________________18661), .DIN2
       (_________________0___18660), .Q (____0___19212));
  nnd2s1 ______451160(.DIN1 (________19098), .DIN2 (_____9), .Q
       (____9___19199));
  nnd2s1 _____0_451161(.DIN1 (______________18869), .DIN2
       (____9____29052), .Q (____0___19303));
  and2s1 _______451162(.DIN1 (____0____31818), .DIN2
       (____________________________________18836), .Q (________19451));
  nor2s1 _______451163(.DIN1 (_________28603), .DIN2 (____9____29052),
       .Q (___9____21595));
  nor2s1 _____451164(.DIN1 (________19067), .DIN2
       (_____________________18639), .Q (________19151));
  nnd2s1 _______451165(.DIN1 (________25995), .DIN2 (outData[6]), .Q
       (________19285));
  nor2s1 _______451166(.DIN1 (outData[6]), .DIN2 (outData[4]), .Q
       (____0___19310));
  and2s1 ____09_451167(.DIN1 (_________31388), .DIN2
       (_________9_______18807), .Q (____99__19301));
  nnd2s1 ______451168(.DIN1 (_____________________18626), .DIN2
       (___9_0__19727), .Q (________19147));
  nnd2s1 _______451169(.DIN1 (________19066), .DIN2
       (______________0______________________18825), .Q
       (_____0__19351));
  or2s1 _______451170(.DIN1 (___9____24300), .DIN2 (outData[4]), .Q
       (________22869));
  nnd2s1 _____0_451171(.DIN1 (______________18871), .DIN2
       (_________28866), .Q (____0___19304));
  nnd2s1 _______451172(.DIN1 (____0___21449), .DIN2 (_________31131),
       .Q (___9____19761));
  nnd2s1 _______451173(.DIN1 (____0________________18594), .DIN2
       (________19665), .Q (____0___19208));
  nnd2s1 _______451174(.DIN1 (_____________________18614), .DIN2
       (____0___19056), .Q (________19150));
  or2s1 _______451175(.DIN1 (___99___20691), .DIN2 (outData[3]), .Q
       (________19453));
  nnd2s1 _____451176(.DIN1 (_____________________18626), .DIN2
       (___9____19729), .Q (____0___19206));
  nnd2s1 _______451177(.DIN1 (_____________18905), .DIN2 (outData[30]),
       .Q (________19159));
  nnd2s1 ____09_451178(.DIN1 (______18912), .DIN2 (inData[9]), .Q
       (________19263));
  nnd2s1 _______451179(.DIN1 (_____________18899), .DIN2
       (________20899), .Q (___0____19843));
  or2s1 _______451180(.DIN1 (________19065), .DIN2
       (_________________18797), .Q (___00___19775));
  nnd2s1 _______451181(.DIN1 (______________________18631), .DIN2
       (________19064), .Q (_____9__19195));
  nnd2s1 ______451182(.DIN1 (outData[18]), .DIN2 (________19231), .Q
       (_____9__19418));
  nnd2s1 _______451183(.DIN1 (_____18907), .DIN2 (inData[7]), .Q
       (________19218));
  nnd2s1 _______451184(.DIN1 (____0________________18593), .DIN2
       (________19063), .Q (_____0__19439));
  hi1s1 _____9_451185(.DIN (________19245), .Q (________19457));
  nnd2s1 ______451186(.DIN1 (outData[19]), .DIN2 (_______18990), .Q
       (________19288));
  nor2s1 _______451187(.DIN1 (________19287), .DIN2
       (__________________0_), .Q (____9___19197));
  nnd2s1 _______451188(.DIN1 (_________34479), .DIN2 (_________30215),
       .Q (_____9__19162));
  nor2s1 _______451189(.DIN1 (__99____27109), .DIN2
       (_____________18894), .Q (___00___19777));
  nor2s1 _______451190(.DIN1 (________19062), .DIN2 (___0____20730), .Q
       (________19270));
  nnd2s1 _______451191(.DIN1 (_____________________18621), .DIN2
       (________19278), .Q (________19564));
  nor2s1 _______451192(.DIN1 (outData[26]), .DIN2 (_____________18899),
       .Q (____0___19406));
  nor2s1 _______451193(.DIN1 (________19061), .DIN2
       (_____________________18638), .Q (________19274));
  nor2s1 _______451194(.DIN1 (___9_0__19727), .DIN2 (___9____19729), .Q
       (____0___19404));
  or2s1 _______451195(.DIN1 (_________34492), .DIN2 (__99____27118), .Q
       (________19536));
  nor2s1 _______451196(.DIN1 (________19420), .DIN2
       (_____________________18599), .Q (________19277));
  nnd2s1 _____9_451197(.DIN1 (_____18911), .DIN2
       (_________________9___18642), .Q (________19284));
  nnd2s1 _______451198(.DIN1 (_____________18900), .DIN2
       (_________28581), .Q (_________31220));
  nnd2s1 _____9_451199(.DIN1 (_____________18900), .DIN2
       (___9___18978), .Q (________19922));
  nor2s1 ______451200(.DIN1 (outData[11]), .DIN2 (outData[13]), .Q
       (_____9__19991));
  nor2s1 _______451201(.DIN1 (_____0__19068), .DIN2 (___0____19780), .Q
       (________19547));
  nor2s1 _____451202(.DIN1 (outData[11]), .DIN2 (outData[9]), .Q
       (_________29370));
  nor2s1 _______451203(.DIN1 (________19353), .DIN2
       (____0_________________18656), .Q (________19412));
  nnd2s1 _______451204(.DIN1 (_________34448), .DIN2 (______18923), .Q
       (____99__21810));
  and2s1 _______451205(.DIN1 (_____________________18662), .DIN2
       (_________________9___18669), .Q (_____0__20097));
  nnd2s1 _______451206(.DIN1 (_____9__21513), .DIN2 (____0___21991), .Q
       (___9____20625));
  nor2s1 ______451207(.DIN1 (_________________9___18669), .DIN2
       (__99____27118), .Q (________20200));
  nnd2s1 _______451208(.DIN1 (____0________________18595), .DIN2
       (________22050), .Q (____0___19497));
  nor2s1 _______451209(.DIN1 (________19353), .DIN2 (_____0__20382), .Q
       (________19549));
  nor2s1 _______451210(.DIN1 (________19098), .DIN2
       (__________________0___18628), .Q (_____0__19506));
  nnd2s1 _______451211(.DIN1 (_________________0___18660), .DIN2
       (_____________________18661), .Q (____90__20126));
  xor2s1 _______451212(.DIN1 (_____________18896), .DIN2 (outData[13]),
       .Q (________19443));
  nnd2s1 _______451213(.DIN1 (_________________9___18606), .DIN2
       (________19436), .Q (____00__19302));
  hi1s1 _______451214(.DIN (________19060), .Q (________19322));
  nnd2s1 ______451215(.DIN1 (____0________________18592), .DIN2
       (________19063), .Q (____0___19403));
  nnd2s1 ______451216(.DIN1 (_________________9___18627), .DIN2
       (_____0), .Q (________19337));
  hi1s1 _______451217(.DIN (________22136), .Q (________20204));
  nnd2s1 _______451218(.DIN1 (________19996), .DIN2 (________19343), .Q
       (________19445));
  hi1s1 ____451219(.DIN (________19229), .Q (________19367));
  nnd2s1 _______451220(.DIN1 (____0_________________18657), .DIN2
       (____09), .Q (____9___19397));
  nor2s1 _______451221(.DIN1 (________19141), .DIN2
       (_____________________18609), .Q (____9___19293));
  nor2s1 _____9_451222(.DIN1 (outData[15]), .DIN2 (outData[17]), .Q
       (________21942));
  nor2s1 _______451223(.DIN1 (____0___19309), .DIN2 (____09), .Q
       (____0___19401));
  nnd2s1 ______451224(.DIN1 (________19139), .DIN2
       (______________________18644), .Q (____9___19298));
  hi1s1 ____0_451225(.DIN (________19425), .Q (_____9__19467));
  nnd2s1 ______451226(.DIN1 (____0___19059), .DIN2 (_____9__20491), .Q
       (_____0__19409));
  nnd2s1 _______451227(.DIN1 (____0___19058), .DIN2 (________19287), .Q
       (________19430));
  nnd2s1 _______451228(.DIN1 (_____________________18612), .DIN2
       (___0____19807), .Q (_____0__19361));
  and2s1 _______451229(.DIN1 (____9___22253), .DIN2
       (_____________________18661), .Q (________19545));
  nnd2s1 _______451230(.DIN1 (__________________0_), .DIN2
       (________19287), .Q (___9____19697));
  hi1s1 ____00_451231(.DIN (_____9__19177), .Q (____0___19307));
  nnd2s1 _______451232(.DIN1 (______________________18630), .DIN2
       (_____9), .Q (________20123));
  hi1s1 _______451233(.DIN (____0___19057), .Q (____9___19393));
  and2s1 _______451234(.DIN1 (_____________________18619), .DIN2
       (________19278), .Q (____99__19398));
  nor2s1 _____0_451235(.DIN1 (____0___19056), .DIN2
       (_____________________18614), .Q (________19472));
  hi1s1 ____0__451236(.DIN (________19624), .Q (________19575));
  hi1s1 ______451237(.DIN (____0___19055), .Q (________19442));
  and2s1 _______451238(.DIN1 (_____________________18602), .DIN2
       (________19386), .Q (________19413));
  nor2s1 _______451239(.DIN1 (_____9__20011), .DIN2
       (____0________________18649), .Q (____9___19490));
  nnd2s1 _______451240(.DIN1 (___0____19780), .DIN2 (_____0__19068), .Q
       (____9___19296));
  hi1s1 _____0_451241(.DIN (________19266), .Q (___0____19787));
  hi1s1 _______451242(.DIN (_________________0___18633), .Q
       (_________35105));
  nor2s1 _______451243(.DIN1 (___9____19718), .DIN2
       (______________________18672), .Q (____9___19589));
  nnd2s1 _____9_451244(.DIN1 (____0_________________18596), .DIN2
       (____0___19054), .Q (_____9__20078));
  nnd2s1 _______451245(.DIN1 (_____________________18624), .DIN2
       (________20194), .Q (________19513));
  nor2s1 _____9_451246(.DIN1 (____0________________18646), .DIN2
       (___9___18980), .Q (___900__20605));
  and2s1 _____9_451247(.DIN1 (__99____27118), .DIN2
       (_________________9___18669), .Q (____0___21812));
  nnd2s1 _____0_451248(.DIN1 (_____________________18609), .DIN2
       (________19141), .Q (____09__19408));
  hi1s1 _______451249(.DIN (___0____20722), .Q (___9____19733));
  nnd2s1 _____0_451250(.DIN1 (___9_0__19727), .DIN2 (_____0), .Q
       (___99___19765));
  nor2s1 _____0_451251(.DIN1 (___0____19807), .DIN2
       (_____________________18612), .Q (________19615));
  nor2s1 _____0_451252(.DIN1 (________19580), .DIN2
       (____0________________18648), .Q (_____0__19449));
  and2s1 _____0_451253(.DIN1 (_____________________18662), .DIN2
       (_____________________18661), .Q (____9____30867));
  hi1s1 _______451254(.DIN (____9___19295), .Q (_____9__19543));
  nor2s1 _______451255(.DIN1 (_______18969), .DIN2
       (_____________________18611), .Q (________19461));
  and2s1 ______451256(.DIN1 (_____0__20382), .DIN2
       (____0_____________0___18655), .Q (____0___19504));
  nnd2s1 _______451257(.DIN1 (___9____19718), .DIN2 (____0___21453), .Q
       (___9____19712));
  hi1s1 _______451258(.DIN (___9____19752), .Q (________19606));
  hi1s1 _____0_451259(.DIN (____0_), .Q (________19456));
  hi1s1 ____0__451260(.DIN (____00), .Q (________20073));
  hi1s1 ____0_451261(.DIN (____99), .Q (________19555));
  nor2s1 _______451262(.DIN1 (_____0__19612), .DIN2
       (____0________________18651), .Q (___9____19756));
  nor2s1 ______451263(.DIN1 (____9___19053), .DIN2
       (____0________________18589), .Q (________19557));
  nnd2s1 _______451264(.DIN1 (______________________18672), .DIN2
       (___9____19718), .Q (____0___19600));
  nnd2s1 _______451265(.DIN1 (____0________________18589), .DIN2
       (____9___19053), .Q (________19483));
  hi1s1 _____0_451266(.DIN (____9_), .Q (___9_9__19716));
  hi1s1 _____0_451267(.DIN (__9_0), .Q (____9___21071));
  nnd2s1 _______451268(.DIN1 (____________________), .DIN2
       (_____0__19068), .Q (___9____19749));
  nnd2s1 ______451269(.DIN1 (_____________________18622), .DIN2
       (________19156), .Q (_____9__22215));
  nnd2s1 _______451270(.DIN1 (____0________________18651), .DIN2
       (_____0__19612), .Q (________20160));
  hi1s1 _______451271(.DIN (__909), .Q (________21824));
  nnd2s1 ______451272(.DIN1 (_____________________18621), .DIN2
       (________19184), .Q (____0___21724));
  hi1s1 ____0_451273(.DIN (_______19052), .Q (________20901));
  hi1s1 _______451274(.DIN (________19643), .Q (________20072));
  nor2s1 ______451275(.DIN1 (________19061), .DIN2 (________19077), .Q
       (____00__19592));
  nor2s1 _______451276(.DIN1 (___9___18976), .DIN2
       (_____________________18604), .Q (___9____19701));
  hi1s1 _______451277(.DIN (___9___18975), .Q (____9___19587));
  nor2s1 ____0__451278(.DIN1 (_____09__31192), .DIN2 (_____0___34425),
       .Q (_______19051));
  or2s1 ____0_451279(.DIN1 (_________30215), .DIN2 (_________34479), .Q
       (_______19050));
  nor2s1 ____0__451280(.DIN1 (_______19048), .DIN2
       (_____________________18626), .Q (_______19049));
  nnd2s1 _______451281(.DIN1 (_____________18902), .DIN2 (outData[30]),
       .Q (_______19047));
  xor2s1 _______451282(.DIN1 (_______________18882), .DIN2
       (_______________18880), .Q (____0__19046));
  nnd2s1 _____9_451283(.DIN1 (outData[21]), .DIN2 (outData[19]), .Q
       (____9__19045));
  hi1s1 _______451284(.DIN (_______19043), .Q (_______19044));
  nnd2s1 ____0_451285(.DIN1 (_____________18900), .DIN2 (outData[26]),
       .Q (___0___19042));
  xnr2s1 _____451286(.DIN1 (______9__34490), .DIN2
       (_________________18712), .Q (____9__19041));
  and2s1 _____0_451287(.DIN1 (_______19039), .DIN2
       (_____________0___18779), .Q (_______19040));
  nnd2s1 _____9_451288(.DIN1 (______18932), .DIN2 (______9__28578), .Q
       (_______19038));
  nnd2s1 ______451289(.DIN1 (_________34445), .DIN2 (____9__19036), .Q
       (_______19037));
  nnd2s1 _______451290(.DIN1 (outData[20]), .DIN2 (outData[18]), .Q
       (___0___19034));
  hi1s1 _______451291(.DIN (___9___19032), .Q (___00__19033));
  xor2s1 _______451292(.DIN1
       (______________________________________0_____________18887),
       .DIN2 (___________0___18883), .Q (___9___19031));
  nor2s1 ______451293(.DIN1 (________25995), .DIN2 (____99__19113), .Q
       (___9___19030));
  nor2s1 ______451294(.DIN1 (______________0___________________0),
       .DIN2 (______18914), .Q (_______19029));
  nnd2s1 _______451295(.DIN1 (outData[21]), .DIN2 (outData[20]), .Q
       (_______19028));
  nor2s1 _______451296(.DIN1 (_________________18680), .DIN2
       (__99____27118), .Q (_______19027));
  nor2s1 ____09_451297(.DIN1 (_________34432), .DIN2 (_________29688),
       .Q (_______19026));
  nnd2s1 _______451298(.DIN1 (_________29585), .DIN2
       (_________9______18801), .Q (_______19025));
  xor2s1 ______451299(.DIN1 (_________________18698), .DIN2
       (______________0____________________), .Q (_______19024));
  nnd2s1 ____0__451300(.DIN1 (______18927), .DIN2 (inData[10]), .Q
       (_______19023));
  nor2s1 _______451301(.DIN1 (________19061), .DIN2 (________19996), .Q
       (_______19022));
  nor2s1 _______451302(.DIN1 (_____0___31003), .DIN2 (_____00__30456),
       .Q (_______19021));
  nor2s1 ____0__451303(.DIN1 (________20899), .DIN2 (outData[20]), .Q
       (_______19020));
  nnd2s1 ____0__451304(.DIN1 (___0_9__19834), .DIN2 (____90__19292), .Q
       (_______19019));
  nor2s1 _______451305(.DIN1 (______________18870), .DIN2
       (_________________0___18660), .Q (_______19018));
  or2s1 ____0__451306(.DIN1 (____0____28155), .DIN2 (______0__34491),
       .Q (_______19017));
  nnd2s1 ____0_451307(.DIN1 (____0___19116), .DIN2 (_________34496), .Q
       (____0__19016));
  nor2s1 ____0__451308(.DIN1 (_____09__31192), .DIN2 (_________31917),
       .Q (____9__19015));
  xor2s1 ______451309(.DIN1 (_________34447), .DIN2
       (________________18756), .Q (_______19013));
  xnr2s1 _______451310(.DIN1 (________________18787), .DIN2
       (_________34434), .Q (_______19012));
  nor2s1 _______451311(.DIN1 (_________9______18801), .DIN2
       (_________29585), .Q (_______19011));
  hi1s1 ____9_451312(.DIN (_______19009), .Q (_______19010));
  xor2s1 _______451313(.DIN1 (_________________18712), .DIN2
       (_________________18694), .Q (_______19008));
  nor2s1 ______451314(.DIN1 (_____00__30456), .DIN2 (_________31388),
       .Q (____0__19007));
  or2s1 ____0__451315(.DIN1 (________19278), .DIN2
       (_____________________18619), .Q (____9__19006));
  nor2s1 ____0__451316(.DIN1 (______________18870), .DIN2
       (______18932), .Q (_______19005));
  xor2s1 _____0_451317(.DIN1 (_________________18698), .DIN2
       (_____________0___18684), .Q (_______19004));
  nor2s1 ____0__451318(.DIN1 (_______19002), .DIN2
       (____0_________________18656), .Q (_______19003));
  nnd2s1 ____0_451319(.DIN1 (outData[22]), .DIN2 (outData[20]), .Q
       (_______19001));
  nnd2s1 _____0_451320(.DIN1 (_____________18897), .DIN2
       (________19231), .Q (_______19000));
  nnd2s1 _____0_451321(.DIN1 (_______18998), .DIN2
       (_________9_______18811), .Q (_______18999));
  nnd2s1 _____9_451322(.DIN1 (________________18756), .DIN2
       (___0_0__20743), .Q (____0__18997));
  xor2s1 _______451323(.DIN1
       (______________________________________0_____________18889),
       .DIN2
       (______________________________________0_____________18891), .Q
       (____9__18996));
  xnr2s1 _______451324(.DIN1 (_____________0___18779), .DIN2
       (_______________0_____________________18830), .Q (_______18995));
  nnd2s1 _______451325(.DIN1 (_________34452), .DIN2 (______18917), .Q
       (_______18993));
  xor2s1 _______451326(.DIN1 (_________34463), .DIN2 (_________34464),
       .Q (_______18992));
  nor2s1 ____0__451327(.DIN1 (____00__19114), .DIN2 (_______18990), .Q
       (_______18991));
  nor2s1 _______451328(.DIN1
       (______________________________________0__________0), .DIN2
       (_________________0___18660), .Q (____0__18989));
  nnd2s1 ______451329(.DIN1 (____9____29052), .DIN2 (_________28603),
       .Q (___09));
  or2s1 ____0__451330(.DIN1 (________19139), .DIN2
       (_____________________18639), .Q (___0___18988));
  xor2s1 _______451331(.DIN1 (________________18788), .DIN2
       (________________18789), .Q (___0___18987));
  nnd2s1 _______451332(.DIN1 (_________31926), .DIN2
       (_________9_______18809), .Q (___0___18986));
  nnd2s1 ____0__451333(.DIN1 (_____________________18625), .DIN2
       (_____0), .Q (___0___18985));
  or2s1 ____0__451334(.DIN1 (____00__19114), .DIN2
       (_________________18746), .Q (___0___18984));
  hi1s1 ____9__451335(.DIN (________19149), .Q (___0___18983));
  nnd2s1 ______451336(.DIN1 (___9__18930), .DIN2
       (_________________18680), .Q (___0___18982));
  nor2s1 _____0_451337(.DIN1 (outData[29]), .DIN2 (outData[27]), .Q
       (___00));
  nnd2s1 ____0_451338(.DIN1 (___9___18981), .DIN2
       (_________9_______18807), .Q (___99));
  nnd2s1 _______451339(.DIN1 (_____________18894), .DIN2 (outData[14]),
       .Q (________19165));
  nnd2s1 _______451340(.DIN1 (___), .DIN2
       (__________________0___18643), .Q (________19157));
  nor2s1 _______451341(.DIN1 (___9___18980), .DIN2 (_______18974), .Q
       (________19158));
  nor2s1 _______451342(.DIN1 (________25995), .DIN2 (outData[10]), .Q
       (________19279));
  nnd2s1 _______451343(.DIN1 (__________________0___18670), .DIN2
       (_____9__21513), .Q (____0___19209));
  hi1s1 ____9__451344(.DIN (____00__19205), .Q (____9___19299));
  nnd2s1 _______451345(.DIN1 (____0_____________0_), .DIN2
       (____90__19292), .Q (________19155));
  nor2s1 _______451346(.DIN1 (____09), .DIN2
       (____0_________________18657), .Q (________19194));
  nnd2s1 _______451347(.DIN1
       (______________________________________0_____________18885),
       .DIN2 (_________31388), .Q (____0___19308));
  nnd2s1 _______451348(.DIN1 (_______18990), .DIN2 (outData[15]), .Q
       (_____9__19233));
  nor2s1 _______451349(.DIN1 (outData[21]), .DIN2 (outData[23]), .Q
       (________19959));
  nor2s1 _______451350(.DIN1 (outData[11]), .DIN2 (__909___26328), .Q
       (________19426));
  nor2s1 _____0_451351(.DIN1 (____0___19309), .DIN2 (________19353), .Q
       (____9___19203));
  nor2s1 _____451352(.DIN1 (_________9_______18812), .DIN2 (____), .Q
       (________19447));
  nor2s1 _____0_451353(.DIN1 (________19343), .DIN2 (________19996), .Q
       (________19328));
  nor2s1 _______451354(.DIN1 (outData[21]), .DIN2 (_________9_), .Q
       (________19421));
  nor2s1 _______451355(.DIN1 (_________9_______18809), .DIN2
       (_________31926), .Q (________19247));
  nnd2s1 _______451356(.DIN1 (_____0__19956), .DIN2 (_____0__19612), .Q
       (_____0__19144));
  nnd2s1 _______451357(.DIN1 (_____________18895), .DIN2 (outData[12]),
       .Q (________19267));
  nnd2s1 _______451358(.DIN1 (____0________________18649), .DIN2
       (_____9__20011), .Q (____9___19202));
  and2s1 _______451359(.DIN1 (______9__30537), .DIN2 (_________9_____),
       .Q (_____9__19438));
  hi1s1 _____9_451360(.DIN (________19161), .Q (________19260));
  nnd2s1 _____9_451361(.DIN1 (____0________________18648), .DIN2
       (____0___19059), .Q (____0___19210));
  nnd2s1 _______451362(.DIN1 (_____________________18666), .DIN2
       (_____9__21513), .Q (________19145));
  nor2s1 ______451363(.DIN1 (outData[19]), .DIN2 (_____________18898),
       .Q (________19422));
  nor2s1 _______451364(.DIN1 (___9___18979), .DIN2 (______9__30169), .Q
       (___0____19798));
  and2s1 ______451365(.DIN1 (_________34444), .DIN2 (________19239), .Q
       (________19636));
  nnd2s1 _____0_451366(.DIN1
       (______________________________________0__________0__18892),
       .DIN2 (____9____29052), .Q (_____0__23115));
  nnd2s1 _____451367(.DIN1 (________19665), .DIN2 (________19063), .Q
       (____9___19294));
  nnd2s1 _______451368(.DIN1 (______0__34491), .DIN2 (____0____28155),
       .Q (____09__19311));
  nor2s1 _______451369(.DIN1 (____99__19113), .DIN2 (outData[12]), .Q
       (________19275));
  nor2s1 _______451370(.DIN1 (____0______________), .DIN2
       (______18933), .Q (____9___19201));
  nor2s1 _____9_451371(.DIN1 (_________30104), .DIN2
       (_______________18873), .Q (________19236));
  nor2s1 _____0_451372(.DIN1 (outData[15]), .DIN2 (_______18990), .Q
       (___9_9));
  hi1s1 _____9_451373(.DIN (________19433), .Q (________19265));
  nor2s1 ____09_451374(.DIN1 (_________31388), .DIN2
       (_________9_______18807), .Q (____9___19300));
  nor2s1 _______451375(.DIN1 (________19576), .DIN2
       (____0_______________), .Q (________19148));
  nnd2s1 _______451376(.DIN1 (___9____19729), .DIN2 (_______19048), .Q
       (_____0__19163));
  hi1s1 _____9_451377(.DIN (_____0__19872), .Q (________19334));
  nor2s1 _____0_451378(.DIN1 (___9___18978), .DIN2 (outData[25]), .Q
       (________19289));
  nnd2s1 _______451379(.DIN1 (____09), .DIN2 (________19353), .Q
       (____9___19396));
  nnd2s1 _____9_451380(.DIN1 (____99__19113), .DIN2 (________25995), .Q
       (___0____19839));
  hi1s1 _______451381(.DIN (_________________0___18633), .Q
       (________35107));
  nor2s1 ______451382(.DIN1 (_____0__22063), .DIN2
       (_____________________18663), .Q (____9___19198));
  nor2s1 _______451383(.DIN1 (_________9_______18811), .DIN2
       (___9__18926), .Q (________19446));
  nnd2s1 _______451384(.DIN1 (_____________18901), .DIN2 (outData[28]),
       .Q (________19241));
  nor2s1 _____0_451385(.DIN1 (____99__19113), .DIN2 (outData[8]), .Q
       (________19280));
  nor2s1 _______451386(.DIN1 (outData[7]), .DIN2 (outData[9]), .Q
       (________19216));
  nor2s1 _______451387(.DIN1 (____0___21991), .DIN2
       (_________________9___18669), .Q (________19345));
  nor2s1 ______451388(.DIN1 (outData[31]), .DIN2 (_________9___18903),
       .Q (_________31653));
  nnd2s1 _______451389(.DIN1 (____________18893), .DIN2
       (___9____25205), .Q (________19441));
  nnd2s1 ______451390(.DIN1 (_________28939), .DIN2 (_________28866),
       .Q (___9_9__19754));
  nor2s1 _______451391(.DIN1 (outData[24]), .DIN2 (_____________18901),
       .Q (________20559));
  nor2s1 _______451392(.DIN1 (________19064), .DIN2
       (______________________18631), .Q (_____9__19291));
  nnd2s1 _______451393(.DIN1 (______18928), .DIN2 (inData[27]), .Q
       (________22334));
  nor2s1 _______451394(.DIN1 (______________________18644), .DIN2
       (________19139), .Q (________19574));
  nnd2s1 _____9_451395(.DIN1 (_________9_), .DIN2 (_______18990), .Q
       (_________30213));
  nnd2s1 _______451396(.DIN1 (_________0_), .DIN2 (________20899), .Q
       (________22684));
  hi1s1 ____0_451397(.DIN (____0___21360), .Q (_____9__21979));
  nor2s1 _____0_451398(.DIN1 (_____________________18661), .DIN2
       (_________34365), .Q (________19905));
  nor2s1 _______451399(.DIN1 (_______________0___________________),
       .DIN2 (_________29646), .Q (___0____22594));
  nor2s1 _____9_451400(.DIN1 (outData[24]), .DIN2 (outData[26]), .Q
       (_________31041));
  or2s1 ______451401(.DIN1 (_________9_______18807), .DIN2
       (___9___18981), .Q (____0____33753));
  nor2s1 _______451402(.DIN1 (_____9), .DIN2 (_____0__20392), .Q
       (___0_9__19825));
  hi1s1 ____9__451403(.DIN (___9___18977), .Q (_____9__19448));
  nor2s1 _______451404(.DIN1 (________19617), .DIN2
       (____0________________18651), .Q (________19415));
  nnd2s1 _______451405(.DIN1 (_____________________18663), .DIN2
       (_____0__22063), .Q (_____9__19668));
  nor2s1 _______451406(.DIN1 (outData[15]), .DIN2 (outData[13]), .Q
       (_____0___29715));
  nor2s1 _______451407(.DIN1 (________19343), .DIN2 (________20091), .Q
       (____0___19407));
  nnd2s1 ______451408(.DIN1 (_____________________18598), .DIN2
       (_________32644), .Q (____90__19196));
  nnd2s1 _____9_451409(.DIN1 (____0________________18649), .DIN2
       (_____9__20491), .Q (_____9__19261));
  nor2s1 _______451410(.DIN1 (_________31983), .DIN2 (_________32644),
       .Q (____9___19200));
  or2s1 ______451411(.DIN1 (________22050), .DIN2
       (____0______________), .Q (________19417));
  nor2s1 ______451412(.DIN1 (outData[26]), .DIN2 (outData[28]), .Q
       (_____9__19881));
  nor2s1 _______451413(.DIN1 (________19062), .DIN2
       (_____________________18667), .Q (____9___19297));
  nnd2s1 _______451414(.DIN1 (___9____19729), .DIN2 (________20194), .Q
       (________19382));
  nnd2s1 _____451415(.DIN1 (_________________0___18597), .DIN2
       (_________31983), .Q (________20374));
  nnd2s1 _______451416(.DIN1 (_________0___18904), .DIN2 (outData[31]),
       .Q (_____0___28711));
  nnd2s1 _______451417(.DIN1 (________19518), .DIN2 (________19665), .Q
       (________19376));
  nor2s1 ______451418(.DIN1 (________19420), .DIN2 (________19463), .Q
       (________19414));
  and2s1 _______451419(.DIN1 (____0______________), .DIN2
       (________22050), .Q (________19431));
  nnd2s1 _____9_451420(.DIN1 (_____________________18605), .DIN2
       (____9___19488), .Q (________19325));
  nnd2s1 _______451421(.DIN1 (_____________________18667), .DIN2
       (________19062), .Q (________19269));
  nnd2s1 _______451422(.DIN1 (____0_____________0___18655), .DIN2
       (_______19002), .Q (________19455));
  nor2s1 _____9_451423(.DIN1 (_____9__20491), .DIN2 (____0___19059), .Q
       (________19608));
  nnd2s1 _______451424(.DIN1 (_____________________18604), .DIN2
       (___9___18976), .Q (________19435));
  nor2s1 _______451425(.DIN1 (________22050), .DIN2
       (____0________________18592), .Q (________21003));
  hi1s1 _____9_451426(.DIN (___90), .Q (________19470));
  nor2s1 ______451427(.DIN1 (___0____20730), .DIN2 (________21976), .Q
       (___9____19694));
  nor2s1 _______451428(.DIN1 (___9____19718), .DIN2
       (_____________________18668), .Q (________19511));
  hi1s1 ____0__451429(.DIN (________19369), .Q (_____9__19515));
  hi1s1 _______451430(.DIN (_________________0___18633), .Q
       (_________35106));
  nor2s1 _______451431(.DIN1 (____90__19292), .DIN2
       (____0_____________0_), .Q (________19530));
  nnd2s1 ______451432(.DIN1 (outData[29]), .DIN2 (outData[28]), .Q
       (_________28766));
  nor2s1 ______451433(.DIN1 (outData[28]), .DIN2 (outData[30]), .Q
       (________19961));
  nnd2s1 ______451434(.DIN1 (____0________________18652), .DIN2
       (________19617), .Q (_____9__19281));
  nnd2s1 _______451435(.DIN1 (_____________________18636), .DIN2
       (________20091), .Q (________19437));
  hi1s1 _______451436(.DIN (_________________0___18633), .Q
       (____99___35108));
  nor2s1 ______451437(.DIN1 (____0____________0___18645), .DIN2
       (_______18974), .Q (________19424));
  hi1s1 ____0__451438(.DIN (_____9__19152), .Q (________22017));
  nor2s1 _______451439(.DIN1 (___0_9__19834), .DIN2 (________19576), .Q
       (________19416));
  hi1s1 ____00_451440(.DIN (_______18973), .Q (___0____20746));
  nor2s1 _____451441(.DIN1 (________19463), .DIN2
       (_____________________18600), .Q (____9___20599));
  hi1s1 ____0__451442(.DIN (________19273), .Q (________19540));
  nor2s1 _______451443(.DIN1 (____0___21453), .DIN2 (___9____19718), .Q
       (________19434));
  hi1s1 _____0_451444(.DIN (_______18972), .Q (____90__19582));
  or2s1 _____0_451445(.DIN1 (_______19002), .DIN2
       (____0_____________0___18655), .Q (_____9__19271));
  nnd2s1 _______451446(.DIN1 (_____________________18664), .DIN2
       (___0____20730), .Q (___9____19710));
  hi1s1 ______451447(.DIN (________19146), .Q (____0___19405));
  nor2s1 _______451448(.DIN1 (________19156), .DIN2 (________19184), .Q
       (____0___19597));
  and2s1 _______451449(.DIN1 (______18933), .DIN2
       (____0______________), .Q (________19553));
  nnd2s1 _______451450(.DIN1 (_____________________18639), .DIN2
       (________19067), .Q (________19444));
  hi1s1 _____0_451451(.DIN (_______18971), .Q (____0___19860));
  nnd2s1 _______451452(.DIN1 (______________________18629), .DIN2
       (________19098), .Q (________19523));
  nor2s1 _______451453(.DIN1 (_____________________18661), .DIN2
       (__99____27118), .Q (___9____20638));
  nor2s1 ______451454(.DIN1 (________19665), .DIN2 (________19518), .Q
       (____0___19595));
  nnd2s1 _______451455(.DIN1 (_____________________18623), .DIN2
       (_______19048), .Q (________21889));
  hi1s1 _______451456(.DIN (_______18970), .Q (___9_9__19706));
  nnd2s1 _______451457(.DIN1 (_____________________18611), .DIN2
       (_______18969), .Q (____09__19601));
  nnd2s1 _______451458(.DIN1 (_____________________18638), .DIN2
       (________19061), .Q (________20564));
  or2s1 _______451459(.DIN1 (_________________9___18669), .DIN2
       (_____________________18662), .Q (___0____21699));
  nor2s1 _______451460(.DIN1 (___0____20730), .DIN2
       (_____________________18664), .Q (________21115));
  nnd2s1 _______451461(.DIN1 (____0________________18653), .DIN2
       (_____9__20011), .Q (___9____21610));
  hi1s1 _______451462(.DIN (______0__28643), .Q (____9____30882));
  hi1s1 ______451463(.DIN (_____9__19551), .Q (___0_9__19844));
  nor2s1 _______451464(.DIN1 (____0___21991), .DIN2 (_____9__21513), .Q
       (____0___21988));
  nnd2s1 _______451465(.DIN1 (outData[5]), .DIN2 (outData[3]), .Q
       (_______18968));
  nor2s1 _______451466(.DIN1 (_________9_____), .DIN2
       (_________9_______18804), .Q (____0__18967));
  and2s1 ____0__451467(.DIN1 (_____0___34427), .DIN2
       (_________________18793), .Q (_______18966));
  nnd2s1 _______451468(.DIN1 (outData[2]), .DIN2 (outData[4]), .Q
       (_______18965));
  and2s1 _______451469(.DIN1 (______________________18672), .DIN2
       (_________________9___18669), .Q (_______18964));
  nor2s1 _______451470(.DIN1
       (______________0___________________9__18827), .DIN2
       (_________________18712), .Q (_______18963));
  nor2s1 _______451471(.DIN1 (_____________18902), .DIN2
       (_________0___18904), .Q (_______18962));
  nnd2s1 ____0_451472(.DIN1 (____0________________18593), .DIN2
       (____0________________18594), .Q (_______18961));
  nor2s1 ____0__451473(.DIN1 (outData[22]), .DIN2 (_________0_), .Q
       (_______18960));
  or2s1 _______451474(.DIN1 (______9__34440), .DIN2 (_________34439),
       .Q (____0__18959));
  and2s1 ____0_451475(.DIN1 (_____0___34427), .DIN2 (_____0___34426),
       .Q (_______18958));
  nor2s1 _______451476(.DIN1 (____________0___18686), .DIN2
       (_________________18718), .Q (_______18957));
  nor2s1 _______451477(.DIN1 (_________9_______18812), .DIN2
       (_____________________________________18839), .Q (_______18956));
  nor2s1 ____0__451478(.DIN1 (________________18771), .DIN2
       (_______________0____________________18829), .Q (____9__18955));
  or2s1 ____0__451479(.DIN1 (______0__34431), .DIN2 (_____09__34430),
       .Q (_______18954));
  and2s1 _______451480(.DIN1 (_________9_______18804), .DIN2
       (inData[16]), .Q (___9___18953));
  nor2s1 _______451481(.DIN1
       (______________________________________0_____________18891),
       .DIN2
       (______________________________________0_____________18889), .Q
       (___9___18952));
  nor2s1 _______451482(.DIN1 (_________________18742), .DIN2
       (_________________18744), .Q (___9_));
  and2s1 ______451483(.DIN1 (_________34434), .DIN2 (_________34433),
       .Q (_______18951));
  nnd2s1 ____0__451484(.DIN1 (_________34492), .DIN2
       (______________0___________________), .Q (_______18950));
  or2s1 ______451485(.DIN1 (_____0___34427), .DIN2
       (_________________18793), .Q (_____));
  nnd2s1 _______451486(.DIN1 (_____________________18665), .DIN2
       (_____________________18668), .Q (____9__18949));
  nor2s1 _______451487(.DIN1 (___________), .DIN2 (outData[13]), .Q
       (____09__19123));
  nor2s1 ____451488(.DIN1 (_______________18873), .DIN2
       (______________________________________0_____________18890), .Q
       (________19452));
  nor2s1 _______451489(.DIN1 (_____________18900), .DIN2 (outData[27]),
       .Q (___9___19032));
  nnd2s1 _______451490(.DIN1 (_____________________18613), .DIN2
       (_____________________18612), .Q (_______18972));
  nnd2s1 _______451491(.DIN1 (_____________________18620), .DIN2
       (_____________________18619), .Q (___9___18977));
  nnd2s1 _______451492(.DIN1 (outData[17]), .DIN2 (_________9_), .Q
       (____9__19035));
  nor2s1 _______451493(.DIN1 (_________9___18903), .DIN2 (outData[27]),
       .Q (________19104));
  or2s1 _______451494(.DIN1 (outData[3]), .DIN2 (outData[5]), .Q
       (_____0__19153));
  or2s1 ____451495(.DIN1 (_________9_______18810), .DIN2
       (___________0___18883), .Q (____0___19213));
  nor2s1 ______451496(.DIN1 (outData[23]), .DIN2 (_____________18900),
       .Q (________19290));
  nnd2s1 ______451497(.DIN1 (_____________18895), .DIN2 (outData[16]),
       .Q (_______18994));
  nor2s1 _______451498(.DIN1 (____0________________18652), .DIN2
       (____0________________18653), .Q (__9_0));
  nnd2s1 _____9_451499(.DIN1 (_____________18900), .DIN2 (outData[27]),
       .Q (_____0__19272));
  or2s1 _______451500(.DIN1 (outData[4]), .DIN2 (__________), .Q
       (________22872));
  and2s1 _______451501(.DIN1 (_____0___34424), .DIN2
       (_________________18795), .Q (________19378));
  nor2s1 _______451502(.DIN1 (__________________0___18670), .DIN2
       (_____________________18664), .Q (_______18973));
  nnd2s1 _____451503(.DIN1 (_____________18898), .DIN2 (outData[23]),
       .Q (________19268));
  nnd2s1 ____09_451504(.DIN1 (inData[9]), .DIN2 (inData[7]), .Q
       (________19193));
  nnd2s1 _____451505(.DIN1 (outData[22]), .DIN2 (_____________18899),
       .Q (________19432));
  nnd2s1 _______451506(.DIN1 (_________9______18801), .DIN2
       (_________9______18800), .Q (________19358));
  nnd2s1 ____0_451507(.DIN1 (___________0___18883), .DIN2
       (_________9_______18810), .Q (____09__19214));
  nor2s1 ______451508(.DIN1 (____0_______________), .DIN2
       (____0_________________18596), .Q (____0_));
  nor2s1 _______451509(.DIN1 (____0________________18650), .DIN2
       (____0________________18653), .Q (_____0__19429));
  nor2s1 ______451510(.DIN1 (inData[7]), .DIN2 (inData[9]), .Q
       (________19154));
  nnd2s1 _______451511(.DIN1 (_____________18894), .DIN2
       (_____________18895), .Q (____0___19305));
  nnd2s1 _____9_451512(.DIN1 (outData[13]), .DIN2 (___________), .Q
       (_____9__19428));
  nnd2s1 _______451513(.DIN1 (_______________18873), .DIN2
       (______________________________________0_____________18890), .Q
       (_______19009));
  nnd2s1 _______451514(.DIN1 (_____________________18626), .DIN2
       (_________________9___18627), .Q (________19383));
  nor2s1 _______451515(.DIN1 (_____________________18667), .DIN2
       (_____________________18664), .Q (____00));
  nnd2s1 _______451516(.DIN1 (_____________________18601), .DIN2
       (_____________________18602), .Q (____9_));
  nor2s1 _______451517(.DIN1 (outData[23]), .DIN2 (_____________18898),
       .Q (_______19043));
  nor2s1 _______451518(.DIN1 (_____________________18637), .DIN2
       (_____________________18638), .Q (_______18970));
  nnd2s1 _______451519(.DIN1 (_____________18897), .DIN2 (_________0_),
       .Q (_________30444));
  nor2s1 _______451520(.DIN1 (inData[27]), .DIN2 (inData[31]), .Q
       (________22433));
  and2s1 ______451521(.DIN1 (_____09__34430), .DIN2 (______0__34431),
       .Q (________23232));
  nnd2s1 _______451522(.DIN1 (_____________________18641), .DIN2
       (______________________18644), .Q (________19411));
  nnd2s1 ______451523(.DIN1 (_________9_______18804), .DIN2
       (_________9_____), .Q (________19283));
  or2s1 _______451524(.DIN1 (____0______________), .DIN2
       (____0________________18591), .Q (_____0__19419));
  nor2s1 _______451525(.DIN1 (_________________9___18642), .DIN2
       (__________________0___18643), .Q (____00__19205));
  nor2s1 _____0_451526(.DIN1 (_____________________18639), .DIN2
       (_____________________18640), .Q (________19161));
  nor2s1 _____9_451527(.DIN1 (______________________18644), .DIN2
       (_____________________18641), .Q (_____0__19602));
  nnd2s1 _______451528(.DIN1 (_____________________18639), .DIN2
       (_____________________18640), .Q (____9___19295));
  nor2s1 ______451529(.DIN1 (____0________________18594), .DIN2
       (____0________________18592), .Q (________19425));
  nor2s1 _______451530(.DIN1 (____0________________18652), .DIN2
       (____0________________18649), .Q (___9____19752));
  nnd2s1 _______451531(.DIN1 (_____________________18623), .DIN2
       (_____________________18624), .Q (___0____20722));
  nnd2s1 _____9_451532(.DIN1 (____0________________18653), .DIN2
       (____0________________18652), .Q (___9_0__19717));
  and2s1 _____9_451533(.DIN1 (_____________________18604), .DIN2
       (_____________________18603), .Q (___9____19700));
  nnd2s1 _______451534(.DIN1 (______________________18629), .DIN2
       (______________________18630), .Q (________19624));
  nnd2s1 _______451535(.DIN1 (____0________________18649), .DIN2
       (____0________________18652), .Q (_____9__19891));
  nnd2s1 _____451536(.DIN1 (_________________9___18616), .DIN2
       (__________________0_), .Q (____9___19586));
  nor2s1 _______451537(.DIN1 (_____________________18663), .DIN2
       (_____________________18668), .Q (____0___21360));
  nnd2s1 _______451538(.DIN1 (____0________________18651), .DIN2
       (____0________________18650), .Q (________19643));
  and2s1 _______451539(.DIN1 (_____________________18622), .DIN2
       (_____________________18619), .Q (________19620));
  or2s1 _______451540(.DIN1 (_____________________18612), .DIN2
       (_____________________18613), .Q (________19410));
  nor2s1 _______451541(.DIN1 (_____________________18619), .DIN2
       (_____________________18620), .Q (___9__));
  nor2s1 ______451542(.DIN1 (_________________18749), .DIN2
       (________________18754), .Q (____9));
  and2s1 ____0__451543(.DIN1 (_________________18793), .DIN2
       (_____0___34426), .Q (____0));
  nor2s1 ______451544(.DIN1 (_________34487), .DIN2 (_________34474),
       .Q (___0_));
  and2s1 ____0__451545(.DIN1
       (_____________________________________18839), .DIN2
       (_________9_______18812), .Q (______18948));
  nor2s1 _______451546(.DIN1 (_______________18880), .DIN2
       (______________________________________0_____________18885), .Q
       (______18947));
  nnd2s1 _______451547(.DIN1 (_________________18795), .DIN2
       (inData[24]), .Q (______18946));
  nnd2s1 ____09_451548(.DIN1 (_______________18873), .DIN2
       (_________9______18802), .Q (______18945));
  or2s1 ____0__451549(.DIN1 (_________________9___18669), .DIN2
       (______________________18672), .Q (______18944));
  nor2s1 ____0__451550(.DIN1 (_____________________18612), .DIN2
       (_____________________18614), .Q (___0__18943));
  nnd2s1 _______451551(.DIN1 (______________18870), .DIN2
       (______________18869), .Q (___9__18942));
  nnd2s1 ____0__451552(.DIN1 (________________18771), .DIN2
       (inData[6]), .Q (______18941));
  nnd2s1 _______451553(.DIN1 (_____________________18625), .DIN2
       (_____________________18624), .Q (______18940));
  and2s1 ____0__451554(.DIN1 (_________34465), .DIN2 (inData[10]), .Q
       (______18939));
  nnd2s1 _______451555(.DIN1 (________________18690), .DIN2
       (inData[12]), .Q (______18938));
  or2s1 ____0__451556(.DIN1 (________________18722), .DIN2
       (______0__34471), .Q (______18937));
  nor2s1 _______451557(.DIN1 (_____________0___18715), .DIN2
       (_____________0___18697), .Q (______18936));
  or2s1 _______451558(.DIN1 (outData[3]), .DIN2 (outData[2]), .Q
       (___0__18935));
  nnd2s1 _______451559(.DIN1 (outData[27]), .DIN2 (_________9___18903),
       .Q (_____0__19262));
  nor2s1 _______451560(.DIN1 (___________), .DIN2 (outData[9]), .Q
       (________19427));
  nnd2s1 _______451561(.DIN1 (_____________________18610), .DIN2
       (_____________________18611), .Q (________19060));
  nor2s1 _______451562(.DIN1 (_____________________18611), .DIN2
       (_____________________18610), .Q (____99));
  or2s1 ______451563(.DIN1 (outData[4]), .DIN2 (outData[2]), .Q
       (________19160));
  nor2s1 _______451564(.DIN1 (outData[10]), .DIN2 (_____________18894),
       .Q (________19276));
  nor2s1 _______451565(.DIN1 (_____________________18624), .DIN2
       (_____________________18623), .Q (_______19052));
  nnd2s1 _____0_451566(.DIN1 (____0________________18589), .DIN2
       (____0________________18590), .Q (____0___19057));
  nnd2s1 _______451567(.DIN1 (______________________18632), .DIN2
       (______________________18631), .Q (__909));
  nnd2s1 _______451568(.DIN1 (outData[8]), .DIN2 (__________), .Q
       (________19286));
  nor2s1 _______451569(.DIN1 (_____________________18600), .DIN2
       (_____________________18599), .Q (___90));
  nor2s1 _______451570(.DIN1 (______________________18631), .DIN2
       (______________________18632), .Q (_______18971));
  nor2s1 ____09_451571(.DIN1 (_________9______18802), .DIN2
       (_______________18873), .Q (________19100));
  nnd2s1 _______451572(.DIN1 (outData[16]), .DIN2 (_____________18897),
       .Q (________19130));
  nor2s1 _______451573(.DIN1 (outData[22]), .DIN2 (_____________18899),
       .Q (____9___19106));
  nor2s1 _____0_451574(.DIN1 (_____________________18621), .DIN2
       (_____________________18622), .Q (____0___19055));
  nnd2s1 _______451575(.DIN1 (____0____________9___18654), .DIN2
       (____0_____________0___18655), .Q (___9___18975));
  nor2s1 ______451576(.DIN1 (_________34472), .DIN2
       (________________18722), .Q (________19226));
  and2s1 _______451577(.DIN1 (_________34474), .DIN2 (_________34487),
       .Q (________19253));
  and2s1 _____0_451578(.DIN1 (_________34439), .DIN2 (______9__34440),
       .Q (_____0__20962));
  nnd2s1 _______451579(.DIN1 (inData[31]), .DIN2 (inData[27]), .Q
       (____9___22437));
  nor2s1 _______451580(.DIN1 (____0____________0___18645), .DIN2
       (____0________________18646), .Q (_____0__19215));
  nor2s1 _____0_451581(.DIN1 (_____________________18605), .DIN2
       (_________________9___18606), .Q (________19229));
  nnd2s1 _______451582(.DIN1 (_____________________18605), .DIN2
       (_________________9___18606), .Q (_____9__19177));
  nnd2s1 _______451583(.DIN1 (_____________18902), .DIN2
       (_________9___18903), .Q (_________28604));
  nnd2s1 ______451584(.DIN1 (__________________0___18643), .DIN2
       (_________________9___18642), .Q (________19149));
  nnd2s1 _______451585(.DIN1 (_____________________18614), .DIN2
       (_____________________18615), .Q (________19146));
  and2s1 _______451586(.DIN1
       (_______________0____________________18829), .DIN2
       (________________18771), .Q (________21366));
  nnd2s1 _______451587(.DIN1 (____0_________________18658), .DIN2
       (____0_________________18659), .Q (_____9__19551));
  nnd2s1 _______451588(.DIN1 (____0____________9_), .DIN2
       (____0_____________0_), .Q (________19273));
  or2s1 _______451589(.DIN1 (outData[1]), .DIN2 (outData[3]), .Q
       (___0____22547));
  nor2s1 _______451590(.DIN1 (_____________________18663), .DIN2
       (_____________________18665), .Q (_____9__19152));
  ib1s1 _______451591(.DIN (___0__18931), .Q (_________31431));
  nor2s1 _____451592(.DIN1 (____0_____________0_), .DIN2
       (____0____________9_), .Q (________19245));
  hi1s1 _______451593(.DIN (___0__18931), .Q (_________35110));
  hi1s1 _______451594(.DIN (___0__18931), .Q (____9____30860));
  nor2s1 _______451595(.DIN1 (____0________________18590), .DIN2
       (____0________________18589), .Q (________19266));
  or2s1 _______451596(.DIN1 (_____________________18603), .DIN2
       (_____________________18604), .Q (________19258));
  and2s1 _____451597(.DIN1 (____0________________18591), .DIN2
       (____0______________), .Q (____0___19402));
  nor2s1 _______451598(.DIN1 (_____________________18666), .DIN2
       (_____________________18668), .Q (_____0__19872));
  nor2s1 _______451599(.DIN1 (______________________18671), .DIN2
       (_____________________18667), .Q (________19433));
  or2s1 _______451600(.DIN1 (_____________________18602), .DIN2
       (_____________________18600), .Q (_____9__19169));
  nor2s1 _____0_451601(.DIN1 (____0_________________18657), .DIN2
       (____0_________________18658), .Q (____9___20501));
  nor2s1 ______451602(.DIN1 (_____________________18609), .DIN2
       (_____________________18608), .Q (________19369));
  or2s1 _______451603(.DIN1 (____0_____________0___18655), .DIN2
       (____0____________9___18654), .Q (_____0__19282));
  or2s1 _______451604(.DIN1 (_____________________18602), .DIN2
       (_____________________18601), .Q (________19610));
  nnd2s1 ______451605(.DIN1 (_____________________18668), .DIN2
       (_____________________18663), .Q (________22136));
  and2s1 ______451606(.DIN1 (_____________________18608), .DIN2
       (_____________________18609), .Q (________19645));
  or2s1 _______451607(.DIN1 (_____________________18615), .DIN2
       (_____________________18614), .Q (________19577));
  nor2s1 _______451608(.DIN1 (_____________________18598), .DIN2
       (_________________0___18597), .Q (______0__28643));
  hi1s1 _______451609(.DIN (_________________18713), .Q (___9__18930));
  hi1s1 _______451610(.DIN (______0__34471), .Q (______18929));
  hi1s1 _______451611(.DIN (inData[31]), .Q (______18928));
  hi1s1 _______451612(.DIN (________________18722), .Q (______18927));
  hi1s1 ______451613(.DIN (_________9_______18812), .Q (___9__18926));
  hi1s1 _____0_451614(.DIN
       (_______________0_____________________18831), .Q (______18925));
  hi1s1 _____9_451615(.DIN (_________34478), .Q (______18924));
  hi1s1 _____0_451616(.DIN (_____________9___18751), .Q (______18923));
  hi1s1 _______451617(.DIN (_____________________18611), .Q
       (______18922));
  hi1s1 _______451618(.DIN (inData[27]), .Q (___0__18921));
  hi1s1 _______451619(.DIN (________________18706), .Q (______18920));
  hi1s1 _______451620(.DIN (_________________18765), .Q (______18919));
  hi1s1 _______451621(.DIN
       (_____________________________________18839), .Q (_______18998));
  hi1s1 _____0_451622(.DIN (_____________________18615), .Q
       (____0___19056));
  hi1s1 _____451623(.DIN (_________9______18801), .Q (________19167));
  hi1s1 ______451624(.DIN (outData[23]), .Q (___9___18978));
  ib1s1 _______451625(.DIN (_________________0___18618), .Q
       (___0__18931));
  hi1s1 ______451626(.DIN (_____0___34429), .Q (________19172));
  hi1s1 _______451627(.DIN (_________________18741), .Q
       (_________29696));
  hi1s1 ______451628(.DIN (_________________18728), .Q (____9___19109));
  hi1s1 _____0_451629(.DIN (____0________________18646), .Q
       (_______18974));
  hi1s1 ______451630(.DIN (_________________18709), .Q (________19535));
  hi1s1 _______451631(.DIN (________________18754), .Q (_____0__20049));
  hi1s1 _______451632(.DIN (_________34445), .Q (_________32626));
  hi1s1 _______451633(.DIN (_________________18701), .Q
       (____9___22074));
  hi1s1 _____9_451634(.DIN (____0_____________0_), .Q (____0___19054));
  hi1s1 _______451635(.DIN (_____________0___18697), .Q
       (________19066));
  hi1s1 _______451636(.DIN (inData[14]), .Q (________20288));
  hi1s1 _______451637(.DIN (_____________0___18684), .Q
       (_________31606));
  hi1s1 _____451638(.DIN (inData[6]), .Q (_______19014));
  hi1s1 _______451639(.DIN (______________________18632), .Q
       (________19064));
  hi1s1 _______451640(.DIN (_________34475), .Q (____0___19116));
  hi1s1 ______451641(.DIN (____________0___18769), .Q (___0__0__27481));
  hi1s1 _______451642(.DIN (_____________________18640), .Q
       (________19067));
  hi1s1 _____9_451643(.DIN (_________________0___18633), .Q
       (___9__18934));
  hi1s1 _____0_451644(.DIN (_________________18761), .Q
       (________19239));
  hi1s1 _______451645(.DIN (_________9_______18806), .Q (___9___18981));
  hi1s1 _______451646(.DIN (________________18757), .Q (___0_0__20743));
  hi1s1 _______451647(.DIN (_________________18782), .Q
       (___9____21556));
  hi1s1 _______451648(.DIN (_________________18730), .Q
       (_________31131));
  hi1s1 _____0_451649(.DIN (clk), .Q (_________32437));
  hi1s1 _______451650(.DIN (_________________18744), .Q
       (___0_9___27842));
  hi1s1 _______451651(.DIN (_________________18727), .Q
       (______0__30564));
  hi1s1 _______451652(.DIN (_____________18900), .Q (outData[25]));
  hi1s1 _____0_451653(.DIN (_________34463), .Q (______9__30169));
  hi1s1 _____0_451654(.DIN (_____________________18622), .Q
       (________19184));
  hi1s1 _______451655(.DIN (________________18789), .Q
       (_________29688));
  hi1s1 _____9_451656(.DIN (inData[30]), .Q (________19264));
  hi1s1 _______451657(.DIN (____0_________________18657), .Q
       (____0___19309));
  hi1s1 _______451658(.DIN (____0________________18594), .Q
       (________19063));
  hi1s1 _______451659(.DIN (_____________________18608), .Q
       (________19141));
  hi1s1 _______451660(.DIN (_____________________18621), .Q
       (________19156));
  hi1s1 _______451661(.DIN (outData[1]), .Q (___99___20691));
  hi1s1 _____451662(.DIN (____0____________9___18654), .Q
       (_______19002));
  hi1s1 _______451663(.DIN (_____________0___18679), .Q
       (_________30215));
  hi1s1 _______451664(.DIN
       (_______________0_____________________18833), .Q
       (_____0___29362));
  hi1s1 _______451665(.DIN (_________________18763), .Q
       (____90___29904));
  hi1s1 _______451666(.DIN (______________________18671), .Q
       (________19062));
  hi1s1 _______451667(.DIN (_____________________18636), .Q
       (________19343));
  hi1s1 _______451668(.DIN (outData[17]), .Q (_______18990));
  hi1s1 ______451669(.DIN (outData[22]), .Q (________20899));
  hi1s1 _______451670(.DIN (_________________9___18616), .Q
       (________19287));
  hi1s1 _______451671(.DIN (_____________________18601), .Q
       (________19386));
  hi1s1 _______451672(.DIN (_________________18768), .Q
       (_________33530));
  hi1s1 _______451673(.DIN (____0_________________18659), .Q (____09));
  hi1s1 ______451674(.DIN (_______________0__________________), .Q
       (_________29646));
  hi1s1 _______451675(.DIN (_____________________18605), .Q
       (________19436));
  hi1s1 _______451676(.DIN (______________________18672), .Q
       (____0___21453));
  hi1s1 _______451677(.DIN (____0____________9_), .Q (____90__19292));
  hi1s1 ______451678(.DIN (___________0___18883), .Q (_________30612));
  hi1s1 ______451679(.DIN (_________9_), .Q (outData[19]));
  hi1s1 _______451680(.DIN (____0________________18651), .Q
       (_____0__19956));
  hi1s1 _______451681(.DIN (outData[16]), .Q (________19231));
  hi1s1 _______451682(.DIN (_____________18899), .Q (outData[24]));
  hi1s1 _______451683(.DIN (____0_______________), .Q (___0_9__19834));
  hi1s1 _______451684(.DIN (_________34474), .Q (_____9___32185));
  hi1s1 _______451685(.DIN (outData[8]), .Q (________25995));
  hi1s1 _______451686(.DIN (____0_________________18596), .Q
       (________19576));
  hi1s1 _______451687(.DIN (_____________18896), .Q (outData[15]));
  hi1s1 _______451688(.DIN (outData[27]), .Q (_________28581));
  hi1s1 _______451689(.DIN (_____________18902), .Q (outData[28]));
  hi1s1 _______451690(.DIN (____0________________18650), .Q
       (_____0__19612));
  hi1s1 _______451691(.DIN (_____________________18598), .Q
       (_________31983));
  hi1s1 _______451692(.DIN (inData[26]), .Q (_____09__31192));
  hi1s1 _______451693(.DIN (__________), .Q (outData[6]));
  hi1s1 ______451694(.DIN (_________________18718), .Q
       (______9__32271));
  hi1s1 _______451695(.DIN (____0________________18592), .Q
       (_____0__20069));
  hi1s1 _______451696(.DIN
       (______________________________________0_____________18885), .Q
       (_____00__30456));
  hi1s1 _______451697(.DIN (_____________18897), .Q (outData[18]));
  hi1s1 _______451698(.DIN (_____________18898), .Q (outData[21]));
  hi1s1 _______451699(.DIN
       (______________0______________________18828), .Q
       (___0_____27914));
  hi1s1 ______451700(.DIN (_________0___18904), .Q (outData[30]));
  hi1s1 _______451701(.DIN (_____________________18666), .Q
       (___9____19718));
  hi1s1 _____9_451702(.DIN (_________0_), .Q (outData[20]));
  hi1s1 _____9_451703(.DIN (_____________________18664), .Q
       (________21976));
  hi1s1 _______451704(.DIN (____0_________________18656), .Q
       (_____0__20382));
  hi1s1 _____451705(.DIN (_____________________18668), .Q
       (_____0__22063));
  hi1s1 ______451706(.DIN (______________18870), .Q (_________28939));
  hi1s1 ______451707(.DIN (______________18871), .Q (____9____29052));
  hi1s1 _____451708(.DIN (_____________________18665), .Q
       (_____9__21513));
  hi1s1 _____9_451709(.DIN (_______________18880), .Q (_________31388));
  hi1s1 _______451710(.DIN
       (______________________________________0_____________18889), .Q
       (_________31281));
  ib1s1 _______451711(.DIN (_________________0___18597), .Q
       (_________32644));
  hi1s1 _____9_451712(.DIN (___________0___18877), .Q (_________33835));
  hi1s1 _____451713(.DIN (_________________0___18660), .Q
       (_________34365));
  hi1s1 _______451714(.DIN (_________34465), .Q (______18918));
  hi1s1 _____451715(.DIN (_________________18746), .Q (______18917));
  hi1s1 _______451716(.DIN (_________34448), .Q (______18916));
  hi1s1 _______451717(.DIN (______0__34461), .Q (___0__18915));
  hi1s1 _______451718(.DIN (_________34486), .Q (___9));
  hi1s1 ______451719(.DIN (_________34493), .Q (______18914));
  hi1s1 _______451720(.DIN (______0__18865), .Q (______18913));
  hi1s1 _______451721(.DIN (inData[7]), .Q (______18912));
  hi1s1 _____9_451722(.DIN (_________9_______18811), .Q (____));
  hi1s1 _____9_451723(.DIN (_________34488), .Q (___0));
  hi1s1 _____9_451724(.DIN (_____0___34427), .Q (__9));
  hi1s1 _____0_451725(.DIN (__________________0___18643), .Q
       (_____18911));
  hi1s1 _______451726(.DIN (_________34433), .Q (_____18910));
  hi1s1 ______451727(.DIN (inData[23]), .Q (_____18909));
  hi1s1 _______451728(.DIN (______9__34470), .Q (_____18908));
  hi1s1 ______451729(.DIN (inData[9]), .Q (_____18907));
  hi1s1 _______451730(.DIN (________________18788), .Q (_____18906));
  hi1s1 ______451731(.DIN (_________________9___18642), .Q (___));
  hi1s1 _____0_451732(.DIN (_________34472), .Q (__0));
  hi1s1 _______451733(.DIN (_________18861), .Q (_____9__19186));
  hi1s1 ______451734(.DIN (________18841), .Q (_________28586));
  hi1s1 _____0_451735(.DIN (_____________________18610), .Q
       (_______18969));
  hi1s1 _______451736(.DIN (___________________________________), .Q
       (________19065));
  hi1s1 _______451737(.DIN (_______________0____________________18829),
       .Q (____00__21260));
  hi1s1 ______451738(.DIN (____________9___18758), .Q (____9__19036));
  hi1s1 ______451739(.DIN (_________________18742), .Q
       (___0_____27683));
  hi1s1 _______451740(.DIN (______0__34441), .Q (________19221));
  hi1s1 _______451741(.DIN (_________34464), .Q (___9___18979));
  hi1s1 _______451742(.DIN (_____________________18603), .Q
       (___9___18976));
  hi1s1 _____9_451743(.DIN (_________________18795), .Q
       (_____9__19224));
  hi1s1 ______451744(.DIN (_________18846), .Q (________19191));
  hi1s1 _____0_451745(.DIN (____0____________0___18645), .Q
       (___9___18980));
  hi1s1 _______451746(.DIN (__________________0_), .Q (____0___19058));
  hi1s1 _______451747(.DIN (_________34436), .Q (_______19039));
  hi1s1 _______451748(.DIN (________________18724), .Q
       (_________30491));
  hi1s1 _____0_451749(.DIN (_________________18698), .Q
       (____09__21084));
  hi1s1 _______451750(.DIN (_________18850), .Q (_________32074));
  hi1s1 _____0_451751(.DIN (_____________________18638), .Q
       (________19077));
  hi1s1 _______451752(.DIN (_________9___0_), .Q (___00____27191));
  hi1s1 _______451753(.DIN (_____0___34428), .Q (_____9__23665));
  hi1s1 ______451754(.DIN (____0________________18590), .Q
       (____9___19053));
  hi1s1 _______451755(.DIN (_________34469), .Q (____0_0__30942));
  hi1s1 _______451756(.DIN (inData[8]), .Q (________23682));
  hi1s1 _______451757(.DIN (_____________________18626), .Q (_____0));
  hi1s1 _______451758(.DIN (inData[4]), .Q (____00__19114));
  hi1s1 _____0_451759(.DIN (_________________18731), .Q
       (____0___21449));
  hi1s1 _______451760(.DIN (_____________________18624), .Q
       (_______19048));
  hi1s1 _______451761(.DIN (_____________________18600), .Q
       (________19420));
  hi1s1 _____9_451762(.DIN (________________18736), .Q
       (_________28788));
  hi1s1 _____451763(.DIN (____0________________18649), .Q
       (____0___19059));
  hi1s1 _______451764(.DIN (_________________9___18606), .Q
       (____9___19488));
  hi1s1 _______451765(.DIN (inData[24]), .Q (____0___24155));
  hi1s1 _______451766(.DIN (_________34449), .Q (_________31917));
  hi1s1 _______451767(.DIN (______________________18629), .Q (_____9));
  hi1s1 ______451768(.DIN (outData[13]), .Q (__99____27109));
  hi1s1 _______451769(.DIN (____________________), .Q (___0____19780));
  hi1s1 ______451770(.DIN (____0________________18647), .Q
       (________19580));
  hi1s1 _______451771(.DIN (______________________18630), .Q
       (________19098));
  hi1s1 _____9_451772(.DIN (_____________________18637), .Q
       (________19061));
  hi1s1 _______451773(.DIN (_____________________18620), .Q
       (________19278));
  hi1s1 ______451774(.DIN (outData[9]), .Q (__909___26328));
  hi1s1 _____451775(.DIN (______________________18617), .Q
       (_____0__19068));
  hi1s1 _______451776(.DIN (_________________18711), .Q
       (____0____28155));
  hi1s1 _______451777(.DIN (_____________________18613), .Q
       (___0____19807));
  hi1s1 ______451778(.DIN (____0________________18595), .Q
       (________19518));
  hi1s1 _____0_451779(.DIN
       (______________________________________0__________0), .Q
       (______18932));
  hi1s1 _______451780(.DIN (_____________________18599), .Q
       (________19463));
  hi1s1 _______451781(.DIN (outData[5]), .Q (___9____25205));
  hi1s1 _______451782(.DIN (_____________18895), .Q (outData[14]));
  hi1s1 _______451783(.DIN (outData[10]), .Q (____99__19113));
  hi1s1 ______451784(.DIN (____0_________________18658), .Q
       (________19353));
  hi1s1 _______451785(.DIN (____0________________18652), .Q
       (_____9__20011));
  hi1s1 _______451786(.DIN (_____________________18641), .Q
       (________19139));
  hi1s1 _______451787(.DIN (_____________18894), .Q (outData[12]));
  hi1s1 ______451788(.DIN (____________18893), .Q (outData[7]));
  hi1s1 _____451789(.DIN (_______________18873), .Q (______9__28578));
  hi1s1 _______451790(.DIN (_________9___18903), .Q (outData[29]));
  hi1s1 _______451791(.DIN (inData[20]), .Q (_____0___31003));
  hi1s1 _______451792(.DIN (____0________________18593), .Q
       (________19665));
  hi1s1 _______451793(.DIN (_________________9___18627), .Q
       (___9_0__19727));
  hi1s1 _____9_451794(.DIN (______________18869), .Q (_________28866));
  hi1s1 _______451795(.DIN (___________), .Q (outData[11]));
  hi1s1 _______451796(.DIN (_____________________18635), .Q
       (________20091));
  hi1s1 _______451797(.DIN
       (______________0______________________18824), .Q
       (_________32114));
  hi1s1 ______451798(.DIN (_____________________18623), .Q
       (________20194));
  hi1s1 ______451799(.DIN (______________18868), .Q (_________28603));
  hi1s1 _______451800(.DIN (outData[2]), .Q (___9____24300));
  ib1s1 _______451801(.DIN (_____________________18662), .Q
       (__99____27118));
  hi1s1 _______451802(.DIN (_____________18901), .Q (outData[26]));
  hi1s1 _______451803(.DIN (_____________________18625), .Q
       (___9____19729));
  nb1s1 _____9_451804(.DIN (_________________0___18660), .Q
       (_________34187));
  ib1s1 _______451805(.DIN (____0____________0_), .Q (______18933));
  hi1s1 _______451806(.DIN (_____________________18634), .Q
       (________19996));
  hi1s1 _______451807(.DIN (____0________________18648), .Q
       (_____9__20491));
  hi1s1 _____9_451808(.DIN (_____________________18663), .Q
       (____9___22253));
  hi1s1 _____9_451809(.DIN (__________________0___18670), .Q
       (____0___21991));
  hi1s1 _______451810(.DIN (____0________________18653), .Q
       (________19617));
  hi1s1 _______451811(.DIN
       (______________________________________0_____________18891), .Q
       (______9__30537));
  hi1s1 _______451812(.DIN (_____________________18667), .Q
       (___0____20730));
  hi1s1 _______451813(.DIN
       (______________________________________0__________0__18892), .Q
       (_________29585));
  ib1s1 ______451814(.DIN (_________________0___18607), .Q
       (_____0___33866));
  hi1s1 _____0_451815(.DIN
       (______________________________________0_____________18890), .Q
       (_________30104));
  hi1s1 _______451816(.DIN
       (______________________________________0_____________18887), .Q
       (_________31926));
  hi1s1 _______451817(.DIN (____0________________18591), .Q
       (________22050));
  hi1s1 _______451818(.DIN (_____________18905), .Q (outData[31]));
  hi1s1 _______451819(.DIN (__________________0___18628), .Q
       (_____0__20392));
  hi1s1 _____451820(.DIN (_________________0___18660), .Q
       (_________34393));
  ib1s1 _______451821(.DIN (_______________18882), .Q (____0____31818));
  or2s1 __(.DIN1 (_________34506), .DIN2 (_____9___32470), .Q
       (______9__34507));
  xnr2s1 __451822(.DIN1 (_________32644), .DIN2 (_________32466), .Q
       (_________34506));
  and2s1 _______451823(.DIN1 (_____90__34508), .DIN2 (_________31198),
       .Q (_____9___34509));
  xor2s1 _______451824(.DIN1 (_________31164), .DIN2 (_________31173),
       .Q (_____90__34508));
  and2s1 _______451825(.DIN1 (_____9___34510), .DIN2 (_________29205),
       .Q (_____9___34511));
  xnr2s1 _______451826(.DIN1 (_________33384), .DIN2 (____0____29154),
       .Q (_____9___34510));
  nnd2s1 ______451827(.DIN1 (_____9___34512), .DIN2 (___09____28127),
       .Q (_____9___34513));
  xor2s1 ______451828(.DIN1 (____000__32751), .DIN2 (____0_0__28177),
       .Q (_____9___34512));
  and2s1 _______451829(.DIN1 (_____9___34514), .DIN2 (________20336),
       .Q (_____9___34515));
  xor2s1 _______451830(.DIN1 (_________28661), .DIN2 (____90__25071),
       .Q (_____9___34514));
  or2s1 _______451831(.DIN1 (_____9___34516), .DIN2 (___9____21595), .Q
       (_____99__34517));
  xnr2s1 _______451832(.DIN1 (____00___33677), .DIN2 (________21039),
       .Q (_____9___34516));
  ib1s1 ______________(.DIN (_________34473), .Q (______9__32183));
  nb1s1 ______________451833(.DIN (__9__0__26429), .Q (____9____34518));
  ib1s1 ______________451834(.DIN (____9_9__34520), .Q
       (____9____34519));
  ib1s1 ______________451835(.DIN (_________31230), .Q
       (____9_9__34520));
  and2s1 _______451836(.DIN1 (___9____19756), .DIN2
       (____0________________18649), .Q (____990__34521));
  or2s1 _______451837(.DIN1 (_________34185), .DIN2 (_____0___34422),
       .Q (____99___34522));
  xnr2s1 _______451838(.DIN1 (_________34022), .DIN2 (______0__33107),
       .Q (____99___34523));
  or2s1 _______451839(.DIN1 (_____0___32202), .DIN2 (_____0___33956),
       .Q (____99___34524));
  or2s1 _______451840(.DIN1 (_________33499), .DIN2 (_________33476),
       .Q (____99___34525));
  and2s1 ______451841(.DIN1 (_________________18775), .DIN2
       (_____00__33310), .Q (____99___34526));
  xnr2s1 ______451842(.DIN1 (_____0___33223), .DIN2 (______9__33463),
       .Q (____99___34527));
  xnr2s1 _______451843(.DIN1 (____________9___18791), .DIN2
       (________________18789), .Q (____99___34528));
  xnr2s1 _______451844(.DIN1 (_________18843), .DIN2 (______0__34988),
       .Q (____99___34529));
  and2s1 _______451845(.DIN1 (_________32862), .DIN2 (_________32886),
       .Q (____999__34530));
  xnr2s1 _______451846(.DIN1 (____9_9__31766), .DIN2 (______9__34450),
       .Q (____000__34531));
  or2s1 _______451847(.DIN1 (_________30709), .DIN2 (_____9___32568),
       .Q (____00___34532));
  or2s1 _______451848(.DIN1 (_________32376), .DIN2 (_________32306),
       .Q (____00___34533));
  xnr2s1 _______451849(.DIN1 (_________18866), .DIN2 (________24538),
       .Q (____00___34534));
  xnr2s1 _______451850(.DIN1 (_____________0___18729), .DIN2
       (____0____30978), .Q (____00___34535));
  and2s1 ______451851(.DIN1 (_________31912), .DIN2 (_________30575),
       .Q (____00___34536));
  xnr2s1 ______451852(.DIN1 (_________18863), .DIN2
       (_________________18695), .Q (____00___34537));
  xnr2s1 _______451853(.DIN1 (______0__31201), .DIN2 (_________30341),
       .Q (____00___34538));
  and2s1 _______451854(.DIN1 (_________31038), .DIN2 (_________31144),
       .Q (____00___34539));
  or2s1 _______451855(.DIN1 (_________31010), .DIN2 (_________30615),
       .Q (____009__34540));
  or2s1 _______451856(.DIN1 (_________30790), .DIN2 (_________30602),
       .Q (____0_0__34541));
  or2s1 _______451857(.DIN1 (_________30688), .DIN2 (_________30498),
       .Q (____0____34542));
  or2s1 _______451858(.DIN1 (_________30674), .DIN2 (_____0___30633),
       .Q (____0____34543));
  or2s1 _______451859(.DIN1 (___0_____27729), .DIN2
       (_____________0___18708), .Q (____0____34544));
  xnr2s1 ______451860(.DIN1 (_________30141), .DIN2 (______0__30309),
       .Q (____0____34545));
  xnr2s1 ______451861(.DIN1 (____0_0__30064), .DIN2 (_________30126),
       .Q (____0____34546));
  and2s1 _______451862(.DIN1 (____909__29910), .DIN2 (____0_9__34549),
       .Q (____0____34547));
  xnr2s1 _______451863(.DIN1 (_________29489), .DIN2 (______0__34708),
       .Q (____0____34548));
  xnr2s1 _______451864(.DIN1 (____0____29161), .DIN2 (_____09__29185),
       .Q (____0_9__34549));
  xnr2s1 _______451865(.DIN1 (____00___30907), .DIN2 (____00___30909),
       .Q (____0_0__34550));
  xnr2s1 _______451866(.DIN1 (__9_0___26991), .DIN2 (_________31567),
       .Q (____0____34551));
  or2s1 _______451867(.DIN1 (__9_9___26890), .DIN2 (__9_____26728), .Q
       (____0____34552));
  and2s1 _______451868(.DIN1 (___009__22544), .DIN2 (________22852), .Q
       (____0____34553));
  and2s1 _______451869(.DIN1 (________21378), .DIN2 (________21332), .Q
       (____0____34554));
  xnr2s1 ______451870(.DIN1 (____9___19495), .DIN2 (_____0___34244), .Q
       (____0____34555));
  xnr2s1 ______451871(.DIN1 (_________________18681), .DIN2
       (____9____34519), .Q (____0____34556));
  and2s1 _______451872(.DIN1 (____0____34557), .DIN2 (_________34354),
       .Q (____0____34558));
  nnd2s1 _______451873(.DIN1 (_________34385), .DIN2 (______0__34370),
       .Q (____0____34557));
  or2s1 _______451874(.DIN1 (____0_9__34559), .DIN2
       (_____________0___18798), .Q (____0_0__34560));
  nnd2s1 _______451875(.DIN1 (_____00__34421), .DIN2 (_________34216),
       .Q (____0_9__34559));
  or2s1 _______451876(.DIN1 (____0____34561), .DIN2 (_____9___31993),
       .Q (____0____34562));
  xnr2s1 _______451877(.DIN1 (______0__33983), .DIN2 (_________33984),
       .Q (____0____34561));
  or2s1 _______451878(.DIN1 (____0____34563), .DIN2 (_________33922),
       .Q (____0____34564));
  nnd2s1 _______451879(.DIN1 (______9__33882), .DIN2 (_________29762),
       .Q (____0____34563));
  or2s1 ______451880(.DIN1 (____0____34565), .DIN2 (______0__33883), .Q
       (____0____34566));
  nnd2s1 ______451881(.DIN1 (_________33894), .DIN2 (_________33898),
       .Q (____0____34565));
  and2s1 _______451882(.DIN1 (____0____34567), .DIN2 (_____0___33867),
       .Q (____0____34568));
  xor2s1 _______451883(.DIN1 (_________33894), .DIN2 (______0__33893),
       .Q (____0____34567));
  or2s1 _______451884(.DIN1 (____0_9__34569), .DIN2 (_________31603),
       .Q (____0_0__34570));
  xnr2s1 _______451885(.DIN1 (______9__33856), .DIN2 (_________33855),
       .Q (____0_9__34569));
  or2s1 _______451886(.DIN1 (____0____34571), .DIN2 (________19188), .Q
       (____0____34572));
  nor2s1 _______451887(.DIN1 (_____9__19438), .DIN2 (____0____33734),
       .Q (____0____34571));
  and2s1 _______451888(.DIN1 (____0____34573), .DIN2 (____0____33689),
       .Q (____0____34574));
  xor2s1 _______451889(.DIN1 (____0_9__30961), .DIN2 (_________29840),
       .Q (____0____34573));
  and2s1 ______451890(.DIN1 (____0____34575), .DIN2 (____9_0__30872),
       .Q (____0____34576));
  xor2s1 ______451891(.DIN1 (_________33564), .DIN2 (_________33563),
       .Q (____0____34575));
  or2s1 _______451892(.DIN1 (____0____34577), .DIN2 (______0__30335),
       .Q (____0____34578));
  xnr2s1 _______451893(.DIN1 (_________35106), .DIN2 (_________33559),
       .Q (____0____34577));
  and2s1 _______451894(.DIN1 (____0_9__34579), .DIN2 (_________33201),
       .Q (____0_0__34580));
  xor2s1 _______451895(.DIN1 (_________________0___18607), .DIN2
       (_________33478), .Q (____0_9__34579));
  xnr2s1 _______451896(.DIN1 (____0____34581), .DIN2 (_________33410),
       .Q (____0____34582));
  xor2s1 _______451897(.DIN1 (____99__22260), .DIN2 (_________30439),
       .Q (____0____34581));
  or2s1 ______451898(.DIN1 (____0____34583), .DIN2 (_________33293), .Q
       (____0____34584));
  xnr2s1 ______451899(.DIN1 (_________33385), .DIN2 (______0__33383),
       .Q (____0____34583));
  or2s1 _______451900(.DIN1 (____0____34585), .DIN2 (_________30504),
       .Q (____0____34586));
  xnr2s1 _______451901(.DIN1 (_________33325), .DIN2 (_________33324),
       .Q (____0____34585));
  and2s1 _______451902(.DIN1 (____0_9__34587), .DIN2 (_________30490),
       .Q (____0_0__34588));
  xor2s1 _______451903(.DIN1 (_________33278), .DIN2 (_________33277),
       .Q (____0_9__34587));
  and2s1 _______451904(.DIN1 (____0____34589), .DIN2 (_________33231),
       .Q (____0____34590));
  xor2s1 _______451905(.DIN1 (_________33264), .DIN2 (_________33263),
       .Q (____0____34589));
  and2s1 _______451906(.DIN1 (____0____34591), .DIN2 (_____9___33021),
       .Q (____0____34592));
  xor2s1 _______451907(.DIN1 (_________33174), .DIN2 (_________33173),
       .Q (____0____34591));
  and2s1 ______451908(.DIN1 (____0____34593), .DIN2 (_________32967),
       .Q (____0____34594));
  xor2s1 _____451909(.DIN1 (________21041), .DIN2 (_________32985), .Q
       (____0____34593));
  and2s1 _____9_451910(.DIN1 (____0____34595), .DIN2 (____9____30853),
       .Q (____0____34596));
  xor2s1 _____9_451911(.DIN1 (_____9___32930), .DIN2 (_____9___32929),
       .Q (____0____34595));
  and2s1 _____9_451912(.DIN1 (____0_9__34597), .DIN2 (____0____32813),
       .Q (____0_0__34598));
  xor2s1 _____9_451913(.DIN1 (_____0___32851), .DIN2 (_____0___32850),
       .Q (____0_9__34597));
  or2s1 _____9_451914(.DIN1 (____0____34599), .DIN2 (_____00__32849),
       .Q (____0____34600));
  xnr2s1 _____9_451915(.DIN1 (____00___31810), .DIN2 (____9_9__31801),
       .Q (____0____34599));
  and2s1 _____9_451916(.DIN1 (____0____34601), .DIN2 (______9__32495),
       .Q (____0____34602));
  xor2s1 _____9_451917(.DIN1 (_________33174), .DIN2 (____9_9__32734),
       .Q (____0____34601));
  and2s1 _____451918(.DIN1 (____0____34603), .DIN2 (______9__32444), .Q
       (____0____34604));
  xor2s1 _____451919(.DIN1 (_________32624), .DIN2 (_________32623), .Q
       (____0____34603));
  and2s1 _____0_451920(.DIN1 (____0____34605), .DIN2 (_________32578),
       .Q (____0____34606));
  xor2s1 _____0_451921(.DIN1 (______0__32594), .DIN2 (______9__32593),
       .Q (____0____34605));
  and2s1 _____0_451922(.DIN1 (____0_9__34607), .DIN2 (_________30687),
       .Q (____0_0__34608));
  xor2s1 _____0_451923(.DIN1 (_____0___32570), .DIN2 (_____00__32569),
       .Q (____0_9__34607));
  or2s1 _____0_451924(.DIN1 (____0____34609), .DIN2 (_________32525),
       .Q (____0____34610));
  nnd2s1 _____0_451925(.DIN1 (_________35106), .DIN2 (_________32508),
       .Q (____0____34609));
  or2s1 _____0_451926(.DIN1 (____0____34611), .DIN2 (______0__30152),
       .Q (____0____34612));
  xnr2s1 _____0_451927(.DIN1 (_________35076), .DIN2 (_________32452),
       .Q (____0____34611));
  and2s1 _____451928(.DIN1 (____0____34613), .DIN2 (_________30511), .Q
       (____0____34614));
  xor2s1 ______451929(.DIN1 (____99___31805), .DIN2 (____99___31806),
       .Q (____0____34613));
  or2s1 _______451930(.DIN1 (____0____34615), .DIN2 (_________31920),
       .Q (____0____34616));
  and2s1 _______451931(.DIN1 (____9____31794), .DIN2 (inData[18]), .Q
       (____0____34615));
  or2s1 _______451932(.DIN1 (____0_9__34617), .DIN2 (_____0__24465), .Q
       (____090__34618));
  nor2s1 _______451933(.DIN1 (________24820), .DIN2 (____9____31779),
       .Q (____0_9__34617));
  or2s1 _______451934(.DIN1 (____09___34619), .DIN2 (_________30779),
       .Q (____09___34620));
  xnr2s1 _______451935(.DIN1 (____9____31752), .DIN2 (____9____31753),
       .Q (____09___34619));
  nor2s1 _______451936(.DIN1 (____09___34621), .DIN2 (____9___19682),
       .Q (____09___34622));
  xnr2s1 _______451937(.DIN1 (_________________18683), .DIN2
       (____9____31744), .Q (____09___34621));
  or2s1 ______451938(.DIN1 (____09___34623), .DIN2 (_________31699), .Q
       (____09___34624));
  xnr2s1 ______451939(.DIN1 (_________35012), .DIN2 (_________30125),
       .Q (____09___34623));
  and2s1 _______451940(.DIN1 (____09___34625), .DIN2 (_____9___31626),
       .Q (____09___34626));
  xor2s1 _______451941(.DIN1 (_________34077), .DIN2 (_________31681),
       .Q (____09___34625));
  and2s1 _______451942(.DIN1 (____099__34627), .DIN2 (_________31559),
       .Q (_____00__34628));
  nor2s1 _______451943(.DIN1 (______0__31641), .DIN2 (______0__31491),
       .Q (____099__34627));
  and2s1 _______451944(.DIN1 (_____0___34629), .DIN2 (_________31365),
       .Q (_____0___34630));
  xor2s1 _______451945(.DIN1 (________21041), .DIN2 (_________31517),
       .Q (_____0___34629));
  and2s1 _______451946(.DIN1 (_____0___34631), .DIN2 (_________28371),
       .Q (_____0___34632));
  xor2s1 _______451947(.DIN1 (_________31478), .DIN2 (_________31477),
       .Q (_____0___34631));
  nnd2s1 ______451948(.DIN1 (_____0___34633), .DIN2 (______0__31278),
       .Q (_____0___34634));
  xor2s1 ______451949(.DIN1 (______0__31325), .DIN2 (_________31323),
       .Q (_____0___34633));
  or2s1 _______451950(.DIN1 (_____0___34635), .DIN2 (________20051), .Q
       (_____0___34636));
  xnr2s1 _______451951(.DIN1 (_________________18695), .DIN2
       (_________31289), .Q (_____0___34635));
  and2s1 _______451952(.DIN1 (_____09__34637), .DIN2 (____99___29994),
       .Q (______0__34638));
  xor2s1 _______451953(.DIN1 (_________31295), .DIN2 (_________31287),
       .Q (_____09__34637));
  and2s1 _______451954(.DIN1 (_________34639), .DIN2 (____9____30849),
       .Q (_________34640));
  xor2s1 _______451955(.DIN1 (________21041), .DIN2 (_____9___31266),
       .Q (_________34639));
  or2s1 _______451956(.DIN1 (_________34641), .DIN2 (_________31040),
       .Q (_________34642));
  xnr2s1 _______451957(.DIN1 (_________34023), .DIN2 (_________31163),
       .Q (_________34641));
  and2s1 ______451958(.DIN1 (_________34643), .DIN2 (_________29555),
       .Q (_________34644));
  nnd2s1 ______451959(.DIN1 (______0__31167), .DIN2 (_________29604),
       .Q (_________34643));
  and2s1 _______451960(.DIN1 (_________34645), .DIN2 (_________31055),
       .Q (_________34646));
  xor2s1 _______451961(.DIN1 (____00___31812), .DIN2 (____0____29105),
       .Q (_________34645));
  and2s1 _______451962(.DIN1 (______9__34647), .DIN2 (____00___30910),
       .Q (______0__34648));
  xor2s1 _______451963(.DIN1 (____0____30977), .DIN2 (____0____30976),
       .Q (______9__34647));
  or2s1 _______451964(.DIN1 (_________34649), .DIN2 (_________30749),
       .Q (_________34650));
  xnr2s1 _______451965(.DIN1 (____9____30882), .DIN2 (____9_0__30881),
       .Q (_________34649));
  or2s1 _______451966(.DIN1 (_________34651), .DIN2 (_________30803),
       .Q (_________34652));
  xnr2s1 _______451967(.DIN1 (____9____30874), .DIN2 (____9_9__30863),
       .Q (_________34651));
  or2s1 ______451968(.DIN1 (_________34653), .DIN2 (_________30742), .Q
       (_________34654));
  nor2s1 ______451969(.DIN1 (_________30781), .DIN2 (____9_9__30897),
       .Q (_________34653));
  or2s1 _______451970(.DIN1 (_________34655), .DIN2 (_________29665),
       .Q (_________34656));
  xnr2s1 _______451971(.DIN1 (____9_9__31781), .DIN2 (____9____30839),
       .Q (_________34655));
  or2s1 _______451972(.DIN1 (______9__34657), .DIN2 (_________30788),
       .Q (______0__34658));
  xnr2s1 _______451973(.DIN1 (_________33925), .DIN2 (_________30789),
       .Q (______9__34657));
  and2s1 _______451974(.DIN1 (_________34659), .DIN2 (_________30562),
       .Q (_________34660));
  xor2s1 _______451975(.DIN1 (___0____21656), .DIN2 (____0____29142),
       .Q (_________34659));
  and2s1 _______451976(.DIN1 (_________34661), .DIN2 (_________30252),
       .Q (_________34662));
  xor2s1 _______451977(.DIN1 (_________________0___18633), .DIN2
       (_____9___30541), .Q (_________34661));
  and2s1 ______451978(.DIN1 (_________34663), .DIN2 (_________30499),
       .Q (_________34664));
  nnd2s1 ______451979(.DIN1 (_________30563), .DIN2 (_________30516),
       .Q (_________34663));
  xnr2s1 _______451980(.DIN1 (_________34665), .DIN2 (_________30587),
       .Q (_________34666));
  xor2s1 _______451981(.DIN1 (________________18721), .DIN2
       (_________________0___18633), .Q (_________34665));
  and2s1 _______451982(.DIN1 (______9__34667), .DIN2 (_________30441),
       .Q (______0__34668));
  xor2s1 _______451983(.DIN1 (____9____31746), .DIN2 (____9_0__29012),
       .Q (______9__34667));
  and2s1 _______451984(.DIN1 (_________34669), .DIN2 (_________30214),
       .Q (_________34670));
  xor2s1 _______451985(.DIN1 (_________32901), .DIN2 (______0__30327),
       .Q (_________34669));
  or2s1 _______451986(.DIN1 (_________34671), .DIN2 (____0____30079),
       .Q (_________34672));
  xnr2s1 _______451987(.DIN1 (________19986), .DIN2 (_________30289),
       .Q (_________34671));
  or2s1 ______451988(.DIN1 (_________34673), .DIN2 (_____0___30278), .Q
       (_________34674));
  nor2s1 ______451989(.DIN1 (________________18691), .DIN2
       (_________30293), .Q (_________34673));
  or2s1 _______451990(.DIN1 (_________34675), .DIN2 (__9__0__26459), .Q
       (_________34676));
  nor2s1 _______451991(.DIN1 (__9_0___26516), .DIN2 (_____9___30176),
       .Q (_________34675));
  or2s1 _______451992(.DIN1 (______9__34677), .DIN2 (____99___29997),
       .Q (______0__34678));
  xnr2s1 _______451993(.DIN1 (_________30693), .DIN2 (_________30139),
       .Q (______9__34677));
  or2s1 _______451994(.DIN1 (_________34679), .DIN2 (______9__30127),
       .Q (_________34680));
  xnr2s1 _______451995(.DIN1 (_________30693), .DIN2 (_________30120),
       .Q (_________34679));
  and2s1 _______451996(.DIN1 (_________34681), .DIN2 (____9____29005),
       .Q (_________34682));
  xor2s1 _______451997(.DIN1 (_________30496), .DIN2 (____0____30058),
       .Q (_________34681));
  and2s1 ______451998(.DIN1 (_________34683), .DIN2 (________20094), .Q
       (_________34684));
  nnd2s1 ______451999(.DIN1 (____0____30013), .DIN2 (_____0__22319), .Q
       (_________34683));
  and2s1 _______452000(.DIN1 (_________34685), .DIN2 (_________29730),
       .Q (_________34686));
  xor2s1 _______452001(.DIN1 (____00___31812), .DIN2 (_________29783),
       .Q (_________34685));
  or2s1 _______452002(.DIN1 (______9__34687), .DIN2 (___0_____27348),
       .Q (______0__34688));
  xnr2s1 _______452003(.DIN1 (_________29598), .DIN2 (_________32644),
       .Q (______9__34687));
  or2s1 _______452004(.DIN1 (_________34689), .DIN2 (__9_____26342), .Q
       (_________34690));
  nor2s1 _______452005(.DIN1 (__9_0___26421), .DIN2 (_________29602),
       .Q (_________34689));
  and2s1 _______452006(.DIN1 (_________34691), .DIN2 (_________29574),
       .Q (_________34692));
  xor2s1 _______452007(.DIN1 (_________28737), .DIN2 (______0__28925),
       .Q (_________34691));
  or2s1 ______452008(.DIN1 (_________34693), .DIN2 (_________34704), .Q
       (_________34694));
  xnr2s1 _____452009(.DIN1 (____9_9__31781), .DIN2 (_____0___29534), .Q
       (_________34693));
  or2s1 _____9_452010(.DIN1 (_________34695), .DIN2 (_________29517),
       .Q (_________34696));
  nnd2s1 _____9_452011(.DIN1 (_________35110), .DIN2 (____9__19035), .Q
       (_________34695));
  or2s1 _____9_452012(.DIN1 (______9__34697), .DIN2 (_________29322),
       .Q (______0__34698));
  xnr2s1 _____9_452013(.DIN1 (_________29496), .DIN2 (_________29497),
       .Q (______9__34697));
  and2s1 _____9_452014(.DIN1 (_________34699), .DIN2 (_________29436),
       .Q (_________34700));
  xor2s1 _____9_452015(.DIN1 (_____0___32851), .DIN2 (_________34710),
       .Q (_________34699));
  or2s1 _____9_452016(.DIN1 (_________34701), .DIN2 (_________29371),
       .Q (_________34702));
  xnr2s1 _____9_452017(.DIN1 (____9____32728), .DIN2 (_________34712),
       .Q (_________34701));
  and2s1 _____452018(.DIN1 (_________34703), .DIN2 (______0__34708), .Q
       (_________34704));
  or2s1 _____452019(.DIN1 (_________29495), .DIN2 (_________29489), .Q
       (_________34703));
  or2s1 _____0_452020(.DIN1 (_________34705), .DIN2 (_________29483),
       .Q (_________34706));
  nor2s1 _____0_452021(.DIN1 (________________18754), .DIN2
       (______9__29491), .Q (_________34705));
  or2s1 _____0_452022(.DIN1 (______9__34707), .DIN2 (_____9___29257),
       .Q (______0__34708));
  xnr2s1 _____0_452023(.DIN1 (____0_0__31851), .DIN2 (_________29410),
       .Q (______9__34707));
  and2s1 _____0_452024(.DIN1 (_________34709), .DIN2 (_____09__29365),
       .Q (_________34710));
  or2s1 _____0_452025(.DIN1 (________________18688), .DIN2
       (_________31252), .Q (_________34709));
  or2s1 _____0_452026(.DIN1 (_________34711), .DIN2 (_________28601),
       .Q (_________34712));
  xnr2s1 _____0_452027(.DIN1 (_________29369), .DIN2 (_________32644),
       .Q (_________34711));
  and2s1 _____452028(.DIN1 (_________34713), .DIN2 (_________29251), .Q
       (_________34714));
  xor2s1 ______452029(.DIN1 (_____0__19985), .DIN2 (_____9___29352), .Q
       (_________34713));
  or2s1 _______452030(.DIN1 (_________34715), .DIN2 (_____0___28808),
       .Q (_________34716));
  xnr2s1 _______452031(.DIN1 (______0__31325), .DIN2 (_________29295),
       .Q (_________34715));
  or2s1 _______452032(.DIN1 (______9__34717), .DIN2 (_________29226),
       .Q (_____90__34718));
  xnr2s1 _______452033(.DIN1 (_________29280), .DIN2 (_________29279),
       .Q (______9__34717));
  and2s1 _______452034(.DIN1 (_____9___34719), .DIN2 (_______18994), .Q
       (_____9___34720));
  nnd2s1 _______452035(.DIN1 (_________29207), .DIN2 (____0___19306),
       .Q (_____9___34719));
  and2s1 _______452036(.DIN1 (_____9___34721), .DIN2 (_________28956),
       .Q (_____9___34722));
  xor2s1 _______452037(.DIN1 (_________31951), .DIN2 (____9____29049),
       .Q (_____9___34721));
  and2s1 ______452038(.DIN1 (_____9___34723), .DIN2 (_________28958),
       .Q (_____9___34724));
  nor2s1 ______452039(.DIN1 (____09__22365), .DIN2 (__9__0__26485), .Q
       (_____9___34723));
  and2s1 _______452040(.DIN1 (_____9___34725), .DIN2 (_________28652),
       .Q (_____9___34726));
  nnd2s1 _______452041(.DIN1 (_________28978), .DIN2 (_____9___28700),
       .Q (_____9___34725));
  or2s1 _______452042(.DIN1 (_____99__34727), .DIN2 (_________34966),
       .Q (_____00__34728));
  and2s1 _______452043(.DIN1 (_________28879), .DIN2 (inData[8]), .Q
       (_____99__34727));
  or2s1 _______452044(.DIN1 (_____0___34729), .DIN2 (__9_____26642), .Q
       (_____0___34730));
  xnr2s1 _______452045(.DIN1 (_________28863), .DIN2 (_____00__30545),
       .Q (_____0___34729));
  and2s1 _______452046(.DIN1 (_____0___34731), .DIN2 (________19165),
       .Q (_____0___34732));
  nnd2s1 _______452047(.DIN1 (_________28873), .DIN2 (________19267),
       .Q (_____0___34731));
  or2s1 ______452048(.DIN1 (_____0___34733), .DIN2 (_____9___28699), .Q
       (_____0___34734));
  nor2s1 ______452049(.DIN1 (_________28726), .DIN2 (_____90__28791),
       .Q (_____0___34733));
  or2s1 _______452050(.DIN1 (_____0___34735), .DIN2 (____0____28176),
       .Q (_____0___34736));
  xnr2s1 _______452051(.DIN1 (_________28593), .DIN2 (_________28592),
       .Q (_____0___34735));
  or2s1 _______452052(.DIN1 (_____09__34737), .DIN2 (__9_____26881), .Q
       (______0__34738));
  nnd2s1 _______452053(.DIN1 (__9_0___26992), .DIN2 (_________28673),
       .Q (_____09__34737));
  or2s1 _______452054(.DIN1 (_________34739), .DIN2 (_________28443),
       .Q (_________34740));
  xnr2s1 _______452055(.DIN1 (______9__28560), .DIN2 (_________28559),
       .Q (_________34739));
  or2s1 _______452056(.DIN1 (_________34741), .DIN2 (_________28555),
       .Q (_________34742));
  nnd2s1 _______452057(.DIN1 (________24859), .DIN2 (____9___21802), .Q
       (_________34741));
  and2s1 ______452058(.DIN1 (_________34743), .DIN2 (_________28364),
       .Q (_________34744));
  xor2s1 ______452059(.DIN1 (_________28492), .DIN2 (____00___31810),
       .Q (_________34743));
  and2s1 _______452060(.DIN1 (_________34745), .DIN2 (____00___28139),
       .Q (_________34746));
  xor2s1 _______452061(.DIN1 (_________28365), .DIN2 (_________28366),
       .Q (_________34745));
  or2s1 _______452062(.DIN1 (______9__34747), .DIN2 (_________28287),
       .Q (______0__34748));
  nnd2s1 _______452063(.DIN1 (_________35094), .DIN2 (________25697),
       .Q (______9__34747));
  or2s1 _______452064(.DIN1 (_________34749), .DIN2 (___099___28130),
       .Q (_________34750));
  nnd2s1 _______452065(.DIN1 (__9_____26734), .DIN2 (________24743), .Q
       (_________34749));
  or2s1 _______452066(.DIN1 (_________34751), .DIN2 (___0_____27785),
       .Q (_________34752));
  xnr2s1 _______452067(.DIN1 (______0__33983), .DIN2 (___0_0___27949),
       .Q (_________34751));
  and2s1 ______452068(.DIN1 (_________34753), .DIN2 (___0_____28001),
       .Q (_________34754));
  or2s1 ______452069(.DIN1 (____________0___18704), .DIN2
       (___0_____27933), .Q (_________34753));
  and2s1 _______452070(.DIN1 (_________34755), .DIN2 (___0_0___27853),
       .Q (_________34756));
  nor2s1 _______452071(.DIN1 (________23842), .DIN2 (_____0__25712), .Q
       (_________34755));
  or2s1 _______452072(.DIN1 (______9__34757), .DIN2 (_________31505),
       .Q (______0__34758));
  and2s1 _______452073(.DIN1 (___0_____27597), .DIN2 (___9____26229),
       .Q (______9__34757));
  and2s1 _______452074(.DIN1 (_________34759), .DIN2 (___0__0__27403),
       .Q (_________34760));
  xor2s1 _______452075(.DIN1 (____9____31746), .DIN2 (___0_____27614),
       .Q (_________34759));
  and2s1 _______452076(.DIN1 (_________34761), .DIN2 (___00____27244),
       .Q (_________34762));
  xor2s1 _______452077(.DIN1 (___0_9___27559), .DIN2 (______9__32620),
       .Q (_________34761));
  and2s1 ______452078(.DIN1 (_________34763), .DIN2 (___0_____27914),
       .Q (_________34764));
  nor2s1 ______452079(.DIN1 (____9____29052), .DIN2 (__9_09__26807), .Q
       (_________34763));
  or2s1 _______452080(.DIN1 (_________34765), .DIN2 (__9_____26852), .Q
       (_________34766));
  nnd2s1 _______452081(.DIN1 (________22681), .DIN2 (________23211), .Q
       (_________34765));
  and2s1 _______452082(.DIN1 (______9__34767), .DIN2 (__9_____26362),
       .Q (______0__34768));
  nor2s1 _______452083(.DIN1 (________25020), .DIN2 (__9_____26641), .Q
       (______9__34767));
  and2s1 _______452084(.DIN1 (_________34769), .DIN2 (__9_____26809),
       .Q (_________34770));
  or2s1 _______452085(.DIN1 (___0_____27914), .DIN2 (___0_9___27751),
       .Q (_________34769));
  and2s1 _______452086(.DIN1 (_________34771), .DIN2 (__90____26315),
       .Q (_________34772));
  nor2s1 _______452087(.DIN1 (________22232), .DIN2 (__9_____26480), .Q
       (_________34771));
  and2s1 ______452088(.DIN1 (_________34773), .DIN2 (_____0__25041), .Q
       (_________34774));
  nor2s1 ______452089(.DIN1 (________24075), .DIN2 (__9_9___26418), .Q
       (_________34773));
  nor2s1 _______452090(.DIN1 (_________34775), .DIN2 (________24200),
       .Q (_________34776));
  nnd2s1 _______452091(.DIN1 (__90____26297), .DIN2 (__9_____26631), .Q
       (_________34775));
  nnd2s1 _______452092(.DIN1 (______9__34777), .DIN2 (_____9__26136),
       .Q (______0__34778));
  nor2s1 _______452093(.DIN1 (________24228), .DIN2 (__9_____26535), .Q
       (______9__34777));
  or2s1 _______452094(.DIN1 (_________34779), .DIN2 (________26071), .Q
       (_________34780));
  nnd2s1 _______452095(.DIN1 (________25142), .DIN2 (inData[8]), .Q
       (_________34779));
  nnd2s1 _______452096(.DIN1 (_________34781), .DIN2 (_________34794),
       .Q (_________34782));
  nor2s1 _______452097(.DIN1 (___00___22543), .DIN2 (__90_9), .Q
       (_________34781));
  or2s1 ______452098(.DIN1 (_________34783), .DIN2 (___9____23362), .Q
       (_________34784));
  nnd2s1 ______452099(.DIN1 (______0__34808), .DIN2 (____9___25460), .Q
       (_________34783));
  nor2s1 _______452100(.DIN1 (_________34785), .DIN2 (_____9__25126),
       .Q (_________34786));
  nnd2s1 _______452101(.DIN1 (________25707), .DIN2 (_____0__24809), .Q
       (_________34785));
  and2s1 _______452102(.DIN1 (______9__34787), .DIN2 (________25451),
       .Q (______0__34788));
  and2s1 _______452103(.DIN1 (__9_____26862), .DIN2 (___9____25191), .Q
       (______9__34787));
  or2s1 _______452104(.DIN1 (_________34789), .DIN2 (_____00__34928),
       .Q (_________34790));
  nnd2s1 _______452105(.DIN1 (___00___25277), .DIN2 (___0____24374), .Q
       (_________34789));
  and2s1 _______452106(.DIN1 (_________34791), .DIN2 (________24943),
       .Q (_________34792));
  nor2s1 _______452107(.DIN1 (________24762), .DIN2 (____0___22358), .Q
       (_________34791));
  and2s1 ______452108(.DIN1 (_________34793), .DIN2 (____9___25170), .Q
       (_________34794));
  and2s1 _____452109(.DIN1 (_____9__22971), .DIN2 (________24864), .Q
       (_________34793));
  or2s1 _____9_452110(.DIN1 (_________34795), .DIN2 (________24858), .Q
       (_________34796));
  nnd2s1 _____9_452111(.DIN1 (_____0__24809), .DIN2 (____0___21910), .Q
       (_________34795));
  or2s1 _____9_452112(.DIN1 (______9__34797), .DIN2 (________24811), .Q
       (______0__34798));
  nnd2s1 _____9_452113(.DIN1 (________25139), .DIN2 (_____9__24198), .Q
       (______9__34797));
  or2s1 _____9_452114(.DIN1 (_________34799), .DIN2 (________19236), .Q
       (_________34800));
  nnd2s1 _____9_452115(.DIN1 (_______________18874), .DIN2
       (________23900), .Q (_________34799));
  and2s1 _____9_452116(.DIN1 (_________34801), .DIN2 (___0____24399),
       .Q (_________34802));
  nor2s1 _____9_452117(.DIN1 (________24232), .DIN2 (___9____25198), .Q
       (_________34801));
  and2s1 _____452118(.DIN1 (_________34803), .DIN2 (________24229), .Q
       (_________34804));
  nor2s1 _____452119(.DIN1 (____0___24157), .DIN2 (___0_9__24400), .Q
       (_________34803));
  nnd2s1 _____0_452120(.DIN1 (_________34805), .DIN2 (________23244),
       .Q (_________34806));
  nor2s1 _____0_452121(.DIN1 (________25123), .DIN2 (_________34864),
       .Q (_________34805));
  and2s1 _____0_452122(.DIN1 (______9__34807), .DIN2 (_____0__25790),
       .Q (______0__34808));
  nor2s1 _____0_452123(.DIN1 (________26101), .DIN2 (________24536), .Q
       (______9__34807));
  or2s1 _____0_452124(.DIN1 (_________34809), .DIN2 (________24692), .Q
       (_________34810));
  nor2s1 _____0_452125(.DIN1 (________24459), .DIN2 (________24458), .Q
       (_________34809));
  or2s1 _____0_452126(.DIN1 (_________34811), .DIN2 (________26092), .Q
       (_________34812));
  nnd2s1 _____0_452127(.DIN1 (________24229), .DIN2 (_____0__24956), .Q
       (_________34811));
  or2s1 _____452128(.DIN1 (_________34813), .DIN2 (_____0__24035), .Q
       (_________34814));
  nnd2s1 ______452129(.DIN1 (________24031), .DIN2 (_____9__24838), .Q
       (_________34813));
  and2s1 _______452130(.DIN1 (_________34815), .DIN2 (____00__24063),
       .Q (_________34816));
  nor2s1 _______452131(.DIN1 (________24030), .DIN2 (___0____22592), .Q
       (_________34815));
  and2s1 _______452132(.DIN1 (______9__34817), .DIN2 (________24006),
       .Q (_____90__34818));
  nor2s1 _______452133(.DIN1 (___09___24423), .DIN2 (_____00__34928),
       .Q (______9__34817));
  or2s1 _______452134(.DIN1 (_____9___34819), .DIN2 (_________32219),
       .Q (_____9___34820));
  nnd2s1 _______452135(.DIN1 (inData[16]), .DIN2 (_________34485), .Q
       (_____9___34819));
  nor2s1 _______452136(.DIN1 (_____9___34821), .DIN2 (__90____26262),
       .Q (_____9___34822));
  nnd2s1 _______452137(.DIN1 (________23952), .DIN2 (________24817), .Q
       (_____9___34821));
  and2s1 ______452138(.DIN1 (_____9___34823), .DIN2 (____9___24154), .Q
       (_____9___34824));
  nor2s1 ______452139(.DIN1 (________24762), .DIN2 (______0__34908), .Q
       (_____9___34823));
  and2s1 _______452140(.DIN1 (_____9___34825), .DIN2 (______9__28444),
       .Q (_____9___34826));
  nor2s1 _______452141(.DIN1 (_________28461), .DIN2 (____00__23974),
       .Q (_____9___34825));
  nor2s1 _______452142(.DIN1 (_____99__34827), .DIN2 (____0___23090),
       .Q (_____00__34828));
  nnd2s1 _______452143(.DIN1 (____0___24704), .DIN2 (_________34910),
       .Q (_____99__34827));
  and2s1 _______452144(.DIN1 (_____0___34829), .DIN2 (_____0__23601),
       .Q (_____0___34830));
  nor2s1 _______452145(.DIN1 (________23136), .DIN2 (________24083), .Q
       (_____0___34829));
  nor2s1 _______452146(.DIN1 (_____0___34831), .DIN2 (______0__34898),
       .Q (_____0___34832));
  nnd2s1 _______452147(.DIN1 (________24669), .DIN2 (________22203), .Q
       (_____0___34831));
  and2s1 ______452148(.DIN1 (_____0___34833), .DIN2 (____0___22630), .Q
       (_____0___34834));
  nor2s1 ______452149(.DIN1 (________24475), .DIN2 (_____9__23843), .Q
       (_____0___34833));
  or2s1 _______452150(.DIN1 (_____0___34835), .DIN2 (________24845), .Q
       (_____0___34836));
  nnd2s1 _______452151(.DIN1 (________23788), .DIN2 (________25399), .Q
       (_____0___34835));
  nor2s1 _______452152(.DIN1 (_____09__34837), .DIN2 (________23845),
       .Q (______0__34838));
  nnd2s1 _______452153(.DIN1 (________22931), .DIN2 (___9____22466), .Q
       (_____09__34837));
  nor2s1 _______452154(.DIN1 (_________34839), .DIN2 (________23844),
       .Q (_________34840));
  nnd2s1 _______452155(.DIN1 (___9____24253), .DIN2 (________24939), .Q
       (_________34839));
  or2s1 _______452156(.DIN1 (_________34841), .DIN2 (________23927), .Q
       (_________34842));
  nnd2s1 _______452157(.DIN1 (___9____23426), .DIN2 (_____9___34922),
       .Q (_________34841));
  or2s1 ______452158(.DIN1 (_________34843), .DIN2 (_________34442), .Q
       (_________34844));
  nnd2s1 ______452159(.DIN1 (inData[0]), .DIN2 (_____0___33034), .Q
       (_________34843));
  nor2s1 _______452160(.DIN1 (_________34845), .DIN2 (_____0___34930),
       .Q (_________34846));
  nnd2s1 _______452161(.DIN1 (____0_9__28185), .DIN2 (________24474),
       .Q (_________34845));
  nor2s1 _______452162(.DIN1 (______9__34847), .DIN2 (________23000),
       .Q (______0__34848));
  nnd2s1 _______452163(.DIN1 (___0____23480), .DIN2 (__9_9___26791), .Q
       (______9__34847));
  or2s1 _______452164(.DIN1 (_________34849), .DIN2 (________24111), .Q
       (_________34850));
  nnd2s1 _______452165(.DIN1 (______9__32271), .DIN2
       (____________0___18686), .Q (_________34849));
  nnd2s1 _______452166(.DIN1 (_________34851), .DIN2 (________23871),
       .Q (_________34852));
  nor2s1 _______452167(.DIN1 (___90___24245), .DIN2 (________23593), .Q
       (_________34851));
  and2s1 ______452168(.DIN1 (_________34853), .DIN2 (___09___23525), .Q
       (_________34854));
  nor2s1 ______452169(.DIN1 (________23315), .DIN2 (________23910), .Q
       (_________34853));
  or2s1 _______452170(.DIN1 (_________34855), .DIN2 (________23752), .Q
       (_________34856));
  nnd2s1 _______452171(.DIN1 (________23314), .DIN2 (________24970), .Q
       (_________34855));
  and2s1 _______452172(.DIN1 (______9__34857), .DIN2 (________23316),
       .Q (______0__34858));
  nor2s1 _______452173(.DIN1 (________22412), .DIN2 (________23831), .Q
       (______9__34857));
  nor2s1 _______452174(.DIN1 (_________34859), .DIN2 (________22907),
       .Q (_________34860));
  nnd2s1 _______452175(.DIN1 (_____0__23223), .DIN2 (________25509), .Q
       (_________34859));
  or2s1 _______452176(.DIN1 (_________34861), .DIN2 (________23218), .Q
       (_________34862));
  nnd2s1 _______452177(.DIN1 (________23114), .DIN2 (____9___24154), .Q
       (_________34861));
  or2s1 ______452178(.DIN1 (_________34863), .DIN2 (_____9__23868), .Q
       (_________34864));
  nnd2s1 ______452179(.DIN1 (________23226), .DIN2 (________24726), .Q
       (_________34863));
  nnd2s1 _______452180(.DIN1 (_________34865), .DIN2 (________23652),
       .Q (_________34866));
  nor2s1 _______452181(.DIN1 (___9_0__24316), .DIN2 (________24207), .Q
       (_________34865));
  and2s1 _______452182(.DIN1 (______9__34867), .DIN2 (________24094),
       .Q (______0__34868));
  nor2s1 _______452183(.DIN1 (________22950), .DIN2 (___0_9__22563), .Q
       (______9__34867));
  nnd2s1 _______452184(.DIN1 (_________34869), .DIN2 (_____0__24646),
       .Q (_________34870));
  nor2s1 _______452185(.DIN1 (________24024), .DIN2 (________23872), .Q
       (_________34869));
  or2s1 _______452186(.DIN1 (_________34871), .DIN2 (__9_____26743), .Q
       (_________34872));
  nnd2s1 _______452187(.DIN1 (________23332), .DIN2 (__99____27091), .Q
       (_________34871));
  and2s1 ______452188(.DIN1 (_________34873), .DIN2 (___0__0__27609),
       .Q (_________34874));
  nor2s1 ______452189(.DIN1 (____09__23983), .DIN2 (___9_9__23422), .Q
       (_________34873));
  nnd2s1 _______452190(.DIN1 (_________34875), .DIN2 (____9___24515),
       .Q (_________34876));
  nor2s1 _______452191(.DIN1 (____9___23973), .DIN2 (________22834), .Q
       (_________34875));
  or2s1 _______452192(.DIN1 (______9__34877), .DIN2 (_____0__22833), .Q
       (______0__34878));
  nnd2s1 _______452193(.DIN1 (___0____23469), .DIN2 (________23332), .Q
       (______9__34877));
  or2s1 _______452194(.DIN1 (_________34879), .DIN2 (_________32604),
       .Q (_________34880));
  and2s1 _______452195(.DIN1 (____0___22631), .DIN2 (inData[24]), .Q
       (_________34879));
  and2s1 _______452196(.DIN1 (_________34881), .DIN2 (___0____23508),
       .Q (_________34882));
  nor2s1 _______452197(.DIN1 (________23932), .DIN2 (__9__0__26637), .Q
       (_________34881));
  and2s1 ______452198(.DIN1 (_________34883), .DIN2 (___00___23444), .Q
       (_________34884));
  nor2s1 ______452199(.DIN1 (___90___23347), .DIN2 (________23919), .Q
       (_________34883));
  or2s1 _______452200(.DIN1 (_________34885), .DIN2 (________23204), .Q
       (_________34886));
  nnd2s1 _______452201(.DIN1 (________23840), .DIN2 (________22768), .Q
       (_________34885));
  and2s1 _______452202(.DIN1 (______9__34887), .DIN2 (________23274),
       .Q (______0__34888));
  nor2s1 _______452203(.DIN1 (___9____25186), .DIN2 (_____0__22772), .Q
       (______9__34887));
  nor2s1 _______452204(.DIN1 (_________34889), .DIN2 (________22162),
       .Q (_________34890));
  nnd2s1 _______452205(.DIN1 (__9_____26555), .DIN2 (________24830), .Q
       (_________34889));
  or2s1 _______452206(.DIN1 (_________34891), .DIN2 (________23144), .Q
       (_________34892));
  nnd2s1 _______452207(.DIN1 (________24735), .DIN2 (____0___22361), .Q
       (_________34891));
  and2s1 ______452208(.DIN1 (_________34893), .DIN2 (____9_0__33597),
       .Q (_________34894));
  or2s1 _____452209(.DIN1 (_____0___31003), .DIN2 (_____0___34426), .Q
       (_________34893));
  nor2s1 _____9_452210(.DIN1 (_________34895), .DIN2 (________23139),
       .Q (_________34896));
  nnd2s1 _____9_452211(.DIN1 (____99__23711), .DIN2 (________22661), .Q
       (_________34895));
  or2s1 _____9_452212(.DIN1 (______9__34897), .DIN2 (________23113), .Q
       (______0__34898));
  and2s1 _____9_452213(.DIN1 (_____9__20856), .DIN2 (___00___20703), .Q
       (______9__34897));
  nor2s1 _____9_452214(.DIN1 (_________34899), .DIN2 (________22775),
       .Q (_________34900));
  nnd2s1 _____9_452215(.DIN1 (___00____27182), .DIN2 (________23292),
       .Q (_________34899));
  or2s1 _____9_452216(.DIN1 (_________34901), .DIN2 (____9___23163), .Q
       (_________34902));
  nnd2s1 _____9_452217(.DIN1 (____0___22721), .DIN2 (__9_____26354), .Q
       (_________34901));
  or2s1 _____452218(.DIN1 (_________34903), .DIN2 (___9____24313), .Q
       (_________34904));
  nnd2s1 _____452219(.DIN1 (________23698), .DIN2 (____9___22982), .Q
       (_________34903));
  nor2s1 _____0_452220(.DIN1 (_________34905), .DIN2 (________24644),
       .Q (_________34906));
  nnd2s1 _____0_452221(.DIN1 (________25774), .DIN2 (____9___23795), .Q
       (_________34905));
  or2s1 _____0_452222(.DIN1 (______9__34907), .DIN2 (________23198), .Q
       (______0__34908));
  nnd2s1 _____0_452223(.DIN1 (________22765), .DIN2 (_____0__23695), .Q
       (______9__34907));
  nor2s1 _____0_452224(.DIN1 (_________34909), .DIN2 (________23218),
       .Q (_________34910));
  nnd2s1 _____0_452225(.DIN1 (________22845), .DIN2 (_____0__25090), .Q
       (_________34909));
  nnd2s1 _____0_452226(.DIN1 (_________34911), .DIN2 (________23014),
       .Q (_________34912));
  nor2s1 _____0_452227(.DIN1 (____9___23883), .DIN2 (_____9__24578), .Q
       (_________34911));
  and2s1 _____452228(.DIN1 (_________34913), .DIN2 (_____9__22408), .Q
       (_________34914));
  nor2s1 ______452229(.DIN1 (________22940), .DIN2 (____9___24884), .Q
       (_________34913));
  nor2s1 _______452230(.DIN1 (_________34915), .DIN2 (___99___24331),
       .Q (_________34916));
  nnd2s1 _______452231(.DIN1 (________23539), .DIN2 (___0____22595), .Q
       (_________34915));
  and2s1 _______452232(.DIN1 (______9__34917), .DIN2 (____09__24992),
       .Q (_____90__34918));
  and2s1 _______452233(.DIN1 (______0__28974), .DIN2 (___9____26218),
       .Q (______9__34917));
  or2s1 _______452234(.DIN1 (_____9___34919), .DIN2 (____0___22268), .Q
       (_____9___34920));
  nnd2s1 _______452235(.DIN1 (___009__23445), .DIN2 (____9___24151), .Q
       (_____9___34919));
  nor2s1 _______452236(.DIN1 (_____9___34921), .DIN2 (___9____24263),
       .Q (_____9___34922));
  nnd2s1 _______452237(.DIN1 (____0___25465), .DIN2 (____99__25750), .Q
       (_____9___34921));
  and2s1 ______452238(.DIN1 (_____9___34923), .DIN2 (____0___22180), .Q
       (_____9___34924));
  nor2s1 ______452239(.DIN1 (__9_____26435), .DIN2 (________22371), .Q
       (_____9___34923));
  or2s1 _______452240(.DIN1 (_____9___34925), .DIN2 (_________34976),
       .Q (_____9___34926));
  nnd2s1 _______452241(.DIN1 (________25604), .DIN2 (________22275), .Q
       (_____9___34925));
  nnd2s1 _______452242(.DIN1 (_____99__34927), .DIN2 (________23014),
       .Q (_____00__34928));
  nor2s1 _______452243(.DIN1 (__9__0__26749), .DIN2 (__9_0___26897), .Q
       (_____99__34927));
  and2s1 _______452244(.DIN1 (_____0___34929), .DIN2 (___0____21644),
       .Q (_____0___34930));
  nor2s1 _______452245(.DIN1 (____0___22810), .DIN2 (________21409), .Q
       (_____0___34929));
  and2s1 _______452246(.DIN1 (_____0___34931), .DIN2 (____0___22630),
       .Q (_____0___34932));
  nor2s1 _______452247(.DIN1 (____90__23704), .DIN2 (___099__22625), .Q
       (_____0___34931));
  or2s1 ______452248(.DIN1 (_____0___34933), .DIN2 (________22641), .Q
       (_____0___34934));
  nnd2s1 ______452249(.DIN1 (________22143), .DIN2 (________24571), .Q
       (_____0___34933));
  nnd2s1 _______452250(.DIN1 (_____0___34935), .DIN2 (________25378),
       .Q (_____0___34936));
  nor2s1 _______452251(.DIN1 (________24780), .DIN2 (________23273), .Q
       (_____0___34935));
  nnd2s1 _______452252(.DIN1 (_____09__34937), .DIN2 (________21937),
       .Q (______0__34938));
  nor2s1 _______452253(.DIN1 (____9___22799), .DIN2 (________23248), .Q
       (_____09__34937));
  nor2s1 _______452254(.DIN1 (_________34939), .DIN2 (________24563),
       .Q (_________34940));
  nnd2s1 _______452255(.DIN1 (____9___23885), .DIN2 (________23222), .Q
       (_________34939));
  or2s1 _______452256(.DIN1 (_________34941), .DIN2 (________22398), .Q
       (_________34942));
  nnd2s1 _______452257(.DIN1 (________23207), .DIN2 (________22321), .Q
       (_________34941));
  nnd2s1 ______452258(.DIN1 (_________34943), .DIN2 (________22140), .Q
       (_________34944));
  nor2s1 ______452259(.DIN1 (________23182), .DIN2 (________22204), .Q
       (_________34943));
  or2s1 _______452260(.DIN1 (_________34945), .DIN2 (___0____24389), .Q
       (_________34946));
  nnd2s1 _______452261(.DIN1 (___9____22462), .DIN2 (________22741), .Q
       (_________34945));
  and2s1 _______452262(.DIN1 (______9__34947), .DIN2 (________22054),
       .Q (______0__34948));
  nor2s1 _______452263(.DIN1 (________24183), .DIN2 (________22205), .Q
       (______9__34947));
  nor2s1 _______452264(.DIN1 (_________34949), .DIN2 (_____9__24181),
       .Q (_________34950));
  nnd2s1 _______452265(.DIN1 (________24859), .DIN2 (________24822), .Q
       (_________34949));
  nnd2s1 _______452266(.DIN1 (_________34951), .DIN2 (________24944),
       .Q (_________34952));
  nor2s1 _______452267(.DIN1 (___0____23488), .DIN2 (_____9__25145), .Q
       (_________34951));
  and2s1 ______452268(.DIN1 (_________34953), .DIN2 (___9_0__22500), .Q
       (_________34954));
  nor2s1 ______452269(.DIN1 (___0____22565), .DIN2 (____9___22986), .Q
       (_________34953));
  nor2s1 _______452270(.DIN1 (_________34955), .DIN2 (___0_0___27370),
       .Q (_________34956));
  nnd2s1 _______452271(.DIN1 (________22682), .DIN2 (________22955), .Q
       (_________34955));
  and2s1 _______452272(.DIN1 (______9__34957), .DIN2 (____0___22364),
       .Q (______0__34958));
  nor2s1 _______452273(.DIN1 (____0___22358), .DIN2 (________25980), .Q
       (______9__34957));
  or2s1 _______452274(.DIN1 (_________34959), .DIN2 (____99__24517), .Q
       (_________34960));
  nnd2s1 _______452275(.DIN1 (________22665), .DIN2 (_____9__25596), .Q
       (_________34959));
  or2s1 _______452276(.DIN1 (_________34961), .DIN2 (___9____22469), .Q
       (_________34962));
  nnd2s1 _______452277(.DIN1 (____9___23885), .DIN2 (________25452), .Q
       (_________34961));
  and2s1 ______452278(.DIN1 (_________34963), .DIN2 (____9___23800), .Q
       (_________34964));
  nor2s1 ______452279(.DIN1 (___9____23387), .DIN2 (____0___22359), .Q
       (_________34963));
  and2s1 _______452280(.DIN1 (_________34965), .DIN2 (___900__21543),
       .Q (_________34966));
  nor2s1 _______452281(.DIN1 (____0____29098), .DIN2 (____9___22167),
       .Q (_________34965));
  and2s1 _______452282(.DIN1 (______9__34967), .DIN2 (___0____21708),
       .Q (______0__34968));
  nor2s1 _______452283(.DIN1 (________22730), .DIN2 (________22683), .Q
       (______9__34967));
  nor2s1 _______452284(.DIN1 (_________34969), .DIN2 (____0___21078),
       .Q (_________34970));
  nnd2s1 _______452285(.DIN1 (___090__21711), .DIN2 (_____9__22435), .Q
       (_________34969));
  and2s1 _______452286(.DIN1 (_________34971), .DIN2 (________21105),
       .Q (_________34972));
  nor2s1 _______452287(.DIN1 (________21836), .DIN2 (_____9__22156), .Q
       (_________34971));
  and2s1 ______452288(.DIN1 (_________34973), .DIN2 (____0___21361), .Q
       (_________34974));
  nor2s1 ______452289(.DIN1 (___9____21618), .DIN2 (_____9__21970), .Q
       (_________34973));
  or2s1 _______452290(.DIN1 (_________34975), .DIN2 (__90_0__26281), .Q
       (_________34976));
  nnd2s1 _______452291(.DIN1 (________25380), .DIN2 (________21435), .Q
       (_________34975));
  nor2s1 _______452292(.DIN1 (______9__34977), .DIN2 (___9_0__22472),
       .Q (______0__34978));
  nnd2s1 _______452293(.DIN1 (____00__24792), .DIN2 (__90_0__26271), .Q
       (______9__34977));
  and2s1 _______452294(.DIN1 (_________34979), .DIN2 (________22029),
       .Q (_________34980));
  nor2s1 _______452295(.DIN1 (________22410), .DIN2 (___0____21700), .Q
       (_________34979));
  or2s1 _______452296(.DIN1 (_________34981), .DIN2 (____9___21807), .Q
       (_________34982));
  nnd2s1 _______452297(.DIN1 (________22129), .DIN2 (___9____20684), .Q
       (_________34981));
  or2s1 ______452298(.DIN1 (_________34983), .DIN2 (____9___20413), .Q
       (_________34984));
  nnd2s1 ______452299(.DIN1 (________21150), .DIN2 (________19557), .Q
       (_________34983));
  and2s1 _______452300(.DIN1 (_________34985), .DIN2 (________21525),
       .Q (_________34986));
  nor2s1 _______452301(.DIN1 (____9___21984), .DIN2 (________21862), .Q
       (_________34985));
  or2s1 _______452302(.DIN1 (______9__34987), .DIN2 (_____0__21140), .Q
       (______0__34988));
  nnd2s1 _______452303(.DIN1 (_____9__20078), .DIN2 (_____9__20283), .Q
       (______9__34987));
  and2s1 _______452304(.DIN1 (_________34989), .DIN2 (________22141),
       .Q (_________34990));
  nor2s1 _______452305(.DIN1 (____9___21537), .DIN2 (________22017), .Q
       (_________34989));
  or2s1 _______452306(.DIN1 (_________34991), .DIN2 (_________18856),
       .Q (_________34992));
  or2s1 _______452307(.DIN1 (____99__21810), .DIN2 (____9___21068), .Q
       (_________34991));
  or2s1 ______452308(.DIN1 (_________34993), .DIN2 (___9____21618), .Q
       (_________34994));
  nnd2s1 _____452309(.DIN1 (________21034), .DIN2 (_____0__22118), .Q
       (_________34993));
  and2s1 _____9_452310(.DIN1 (_________34995), .DIN2 (________21122),
       .Q (_________34996));
  nor2s1 _____9_452311(.DIN1 (_____9__20313), .DIN2 (_____9__21038), .Q
       (_________34995));
  or2s1 _____9_452312(.DIN1 (______9__34997), .DIN2 (____9___21898), .Q
       (______0__34998));
  nnd2s1 _____9_452313(.DIN1 (_____0__21056), .DIN2 (________21381), .Q
       (______9__34997));
  and2s1 _____9_452314(.DIN1 (_________34999), .DIN2 (________20497),
       .Q (_________35000));
  nor2s1 _____9_452315(.DIN1 (________21879), .DIN2 (________21089), .Q
       (_________34999));
  and2s1 _____9_452316(.DIN1 (_________35001), .DIN2 (___99___20694),
       .Q (_________35002));
  nor2s1 _____9_452317(.DIN1 (____90__20972), .DIN2 (___0____19840), .Q
       (_________35001));
  and2s1 _____452318(.DIN1 (_________35003), .DIN2 (________22663), .Q
       (_________35004));
  nor2s1 ____452319(.DIN1 (________21893), .DIN2 (________21224), .Q
       (_________35003));
  or2s1 ____90_452320(.DIN1 (_________35005), .DIN2 (___9____21610), .Q
       (_________35006));
  nnd2s1 ____90_452321(.DIN1 (________20941), .DIN2 (____9___19587), .Q
       (_________35005));
  or2s1 ____90_452322(.DIN1 (______9__35007), .DIN2 (________20965), .Q
       (______0__35008));
  nnd2s1 ____90_452323(.DIN1 (___0____20710), .DIN2 (________19456), .Q
       (______9__35007));
  or2s1 ____90_452324(.DIN1 (_________35009), .DIN2 (________21424), .Q
       (_________35010));
  nnd2s1 ____90_452325(.DIN1 (____9___21257), .DIN2 (_____0__21885), .Q
       (_________35009));
  or2s1 ____90_452326(.DIN1 (_________35011), .DIN2 (___0_9__20715), .Q
       (_________35012));
  or2s1 ____90_452327(.DIN1 (___9____20675), .DIN2 (____0___20891), .Q
       (_________35011));
  or2s1 ____452328(.DIN1 (_________35013), .DIN2 (________20853), .Q
       (_________35014));
  nnd2s1 ____9_452329(.DIN1 (_____9__22147), .DIN2 (_____9__19152), .Q
       (_________35013));
  and2s1 ____9__452330(.DIN1 (_________35015), .DIN2 (________21012),
       .Q (_________35016));
  nor2s1 ____9__452331(.DIN1 (____00__21355), .DIN2 (___9____20660), .Q
       (_________35015));
  or2s1 ____9__452332(.DIN1 (______9__35017), .DIN2 (________21114), .Q
       (_____90__35018));
  nnd2s1 ____9__452333(.DIN1 (___9____20685), .DIN2 (________21893), .Q
       (______9__35017));
  or2s1 ____9__452334(.DIN1 (_____9___35019), .DIN2 (_____9__21093), .Q
       (_____9___35020));
  nnd2s1 ____9__452335(.DIN1 (____0___21816), .DIN2 (____9___21441), .Q
       (_____9___35019));
  and2s1 ____9__452336(.DIN1 (_____9___35021), .DIN2 (_____0__21365),
       .Q (_____9___35022));
  nor2s1 ____9__452337(.DIN1 (___0____21692), .DIN2 (________20450), .Q
       (_____9___35021));
  and2s1 ____9_452338(.DIN1 (_____9___35023), .DIN2 (_____0__21504), .Q
       (_____9___35024));
  nor2s1 ____9_452339(.DIN1 (___9____19725), .DIN2 (____0___20425), .Q
       (_____9___35023));
  or2s1 ____9__452340(.DIN1 (_____9___35025), .DIN2 (________20389), .Q
       (_____9___35026));
  or2s1 ____9__452341(.DIN1 (________20057), .DIN2 (________21089), .Q
       (_____9___35025));
  and2s1 ____9__452342(.DIN1 (_____99__35027), .DIN2 (____0____30080),
       .Q (_____00__35028));
  or2s1 ____9__452343(.DIN1 (_______19014), .DIN2
       (______________0___________________0), .Q (_____99__35027));
  and2s1 ____9__452344(.DIN1 (_____0___35029), .DIN2 (____9___21256),
       .Q (_____0___35030));
  nor2s1 ____9__452345(.DIN1 (________21750), .DIN2 (________21014), .Q
       (_____0___35029));
  nor2s1 ____9__452346(.DIN1 (_____0___35031), .DIN2 (________21113),
       .Q (_____0___35032));
  nnd2s1 ____9__452347(.DIN1 (________22141), .DIN2 (___9____20657), .Q
       (_____0___35031));
  and2s1 ____9_452348(.DIN1 (_____0___35033), .DIN2 (___0____21690), .Q
       (_____0___35034));
  nor2s1 ____9_452349(.DIN1 (________21113), .DIN2 (________19613), .Q
       (_____0___35033));
  and2s1 ____9__452350(.DIN1 (_____0___35035), .DIN2 (_____0__20837),
       .Q (_____0___35036));
  nor2s1 ____9__452351(.DIN1 (________21018), .DIN2 (___9____21568), .Q
       (_____0___35035));
  or2s1 ____9__452352(.DIN1 (_____09__35037), .DIN2 (________21407), .Q
       (______0__35038));
  nnd2s1 ____9__452353(.DIN1 (________19257), .DIN2 (________21141), .Q
       (_____09__35037));
  or2s1 ____9__452354(.DIN1 (_________35039), .DIN2 (_____9__21229), .Q
       (_________35040));
  nnd2s1 ____9__452355(.DIN1 (____0___20517), .DIN2 (____9___21441), .Q
       (_________35039));
  or2s1 ____9__452356(.DIN1 (_________35041), .DIN2 (_________34071),
       .Q (_________35042));
  and2s1 ____9__452357(.DIN1 (________20363), .DIN2 (inData[2]), .Q
       (_________35041));
  or2s1 ____9_452358(.DIN1 (_________35043), .DIN2 (________20897), .Q
       (_________35044));
  nnd2s1 ____9_452359(.DIN1 (inData[16]), .DIN2
       (_________________18683), .Q (_________35043));
  or2s1 ____9__452360(.DIN1 (_________35045), .DIN2 (________19613), .Q
       (_________35046));
  or2s1 ____9__452361(.DIN1 (____9___21898), .DIN2 (____0___20887), .Q
       (_________35045));
  or2s1 ____9__452362(.DIN1 (______9__35047), .DIN2 (________20845), .Q
       (______0__35048));
  nnd2s1 ____9__452363(.DIN1 (____0___20983), .DIN2 (________21776), .Q
       (______9__35047));
  or2s1 ____9__452364(.DIN1 (_________35049), .DIN2 (________19667), .Q
       (_________35050));
  nnd2s1 ____9__452365(.DIN1 (________20166), .DIN2 (_____0__21191), .Q
       (_________35049));
  or2s1 ____9__452366(.DIN1 (_________35051), .DIN2 (________20897), .Q
       (_________35052));
  nnd2s1 ____9__452367(.DIN1 (inData[20]), .DIN2 (_________34489), .Q
       (_________35051));
  nnd2s1 ____9_452368(.DIN1 (_________35053), .DIN2 (____0___20511), .Q
       (_________35054));
  nor2s1 ____9_452369(.DIN1 (________21409), .DIN2 (________20821), .Q
       (_________35053));
  or2s1 ____9__452370(.DIN1 (_________35055), .DIN2 (_____9__20172), .Q
       (_________35056));
  nnd2s1 ____9__452371(.DIN1 (___0____21698), .DIN2 (________21369), .Q
       (_________35055));
  and2s1 ____9__452372(.DIN1 (______9__35057), .DIN2 (________21206),
       .Q (______0__35058));
  nor2s1 ____9__452373(.DIN1 (________21197), .DIN2 (___9____20615), .Q
       (______9__35057));
  and2s1 ____9__452374(.DIN1 (_________35059), .DIN2 (________20243),
       .Q (_________35060));
  nor2s1 ____9__452375(.DIN1 (________21505), .DIN2 (_____0__20352), .Q
       (_________35059));
  or2s1 ____9__452376(.DIN1 (_________35061), .DIN2 (________21495), .Q
       (_________35062));
  nnd2s1 ____9__452377(.DIN1 (________20570), .DIN2 (________20569), .Q
       (_________35061));
  or2s1 ____9_452378(.DIN1 (_________35063), .DIN2 (________20868), .Q
       (_________35064));
  nnd2s1 ____9_452379(.DIN1 (________21893), .DIN2 (________20566), .Q
       (_________35063));
  and2s1 ____9__452380(.DIN1 (_________35065), .DIN2 (________20408),
       .Q (_________35066));
  nor2s1 ____9__452381(.DIN1 (________19974), .DIN2 (____90__20972), .Q
       (_________35065));
  or2s1 ____9__452382(.DIN1 (______9__35067), .DIN2 (________21134), .Q
       (______0__35068));
  nnd2s1 ____9__452383(.DIN1 (________20209), .DIN2 (________19907), .Q
       (______9__35067));
  and2s1 ____9__452384(.DIN1 (_________35069), .DIN2 (________20493),
       .Q (_________35070));
  nor2s1 ____9__452385(.DIN1 (________20854), .DIN2 (___0____21699), .Q
       (_________35069));
  or2s1 ____9__452386(.DIN1 (_________35071), .DIN2 (________21479), .Q
       (_________35072));
  nnd2s1 ____9__452387(.DIN1 (________19886), .DIN2 (____90__21066), .Q
       (_________35071));
  or2s1 ____9_452388(.DIN1 (_________35073), .DIN2 (________21502), .Q
       (_________35074));
  nnd2s1 ____9_452389(.DIN1 (____90__21066), .DIN2 (________21023), .Q
       (_________35073));
  or2s1 ____9__452390(.DIN1 (_________35075), .DIN2 (____09__20235), .Q
       (_________35076));
  nnd2s1 ____9__452391(.DIN1 (_____9__19965), .DIN2 (________20829), .Q
       (_________35075));
  or2s1 ____9__452392(.DIN1 (______9__35077), .DIN2 (____0___20328), .Q
       (______0__35078));
  nor2s1 ____9__452393(.DIN1 (_____________________18604), .DIN2
       (_____9__19177), .Q (______9__35077));
  nnd2s1 ____9__452394(.DIN1 (_________35079), .DIN2 (_____0__20254),
       .Q (_________35080));
  nor2s1 ____9__452395(.DIN1 (___9____20651), .DIN2 (___0_0__21696), .Q
       (_________35079));
  or2s1 ____9__452396(.DIN1 (_________35081), .DIN2 (___0____19804), .Q
       (_________35082));
  nnd2s1 ____9__452397(.DIN1 (_________28604), .DIN2 (inData[14]), .Q
       (_________35081));
  and2s1 ____9_452398(.DIN1 (_________35083), .DIN2 (____0___20984), .Q
       (_________35084));
  or2s1 ____9_452399(.DIN1 (________22050), .DIN2 (________20286), .Q
       (_________35083));
  and2s1 ____9__452400(.DIN1 (_________35085), .DIN2 (____0___19502),
       .Q (_________35086));
  nor2s1 ____9__452401(.DIN1 (___9____19701), .DIN2 (___9____19742), .Q
       (_________35085));
  nor2s1 ____9__452402(.DIN1 (______9__35087), .DIN2 (________19462),
       .Q (______0__35088));
  nnd2s1 ____9__452403(.DIN1 (_____9__19458), .DIN2 (_____0__19380), .Q
       (______9__35087));
  and2s1 ____9__452404(.DIN1 (_________35089), .DIN2 (________19645),
       .Q (_________35090));
  nor2s1 ____9__452405(.DIN1 (____09__19601), .DIN2
       (_________________0___18607), .Q (_________35089));
  and2s1 ____9__452406(.DIN1 (_________35091), .DIN2 (________19322),
       .Q (_________35092));
  nor2s1 ____9__452407(.DIN1 (_________________0___18607), .DIN2
       (____09__19408), .Q (_________35091));
  or2s1 ____9_452408(.DIN1 (_________35093), .DIN2 (___0_9__19817), .Q
       (_________35094));
  and2s1 ____452409(.DIN1 (_____9__19543), .DIN2
       (_____________________18641), .Q (_________35093));
  or2s1 ____99_452410(.DIN1 (_________35095), .DIN2
       (_________________18748), .Q (_________35096));
  nnd2s1 ____99_452411(.DIN1 (____0____29098), .DIN2 (inData[12]), .Q
       (_________35095));
  or2s1 ____99_452412(.DIN1 (______9__35097), .DIN2 (________19526), .Q
       (______0__35098));
  and2s1 ____99_452413(.DIN1 (____99__19398), .DIN2
       (_____________________18621), .Q (______9__35097));
  or2s1 ____99_452414(.DIN1 (_________35099), .DIN2 (________19283), .Q
       (_________35100));
  nnd2s1 ____99_452415(.DIN1 (____9___19587), .DIN2 (_________18852),
       .Q (_________35099));
  or2s1 ____99_452416(.DIN1 (_________35101), .DIN2
       (______________0___________________9__18827), .Q
       (_________35102));
  nnd2s1 ____99_452417(.DIN1 (___9____20638), .DIN2 (inData[18]), .Q
       (_________35101));
  or2s1 ____452418(.DIN1 (_________35103), .DIN2 (______9__33390), .Q
       (_________35104));
  xor2s1 ____452419(.DIN1 (_________29500), .DIN2 (______0__33446), .Q
       (_________35103));
endmodule

