
module iir_core_obf ( inData, clk, reset, outData );
  input [31:0] inData;
  output [31:0] outData;
  input clk, reset;
  wire   ___, _____, _______1____2________________1____________________,
         _______26____2________________26____________________,
         _______25____2________________25____________________,
         _______23____2________________23____________________,
         _______22____2________________22____________________,
         _______21____2________________21____________________,
         _______20____2________________20____________________,
         _______17____2________________17____________________,
         _______16____2________________16____________________,
         _______9____2________________9____________________,
         _______8____2________________8____________________,
         _______5____2________________5____________________,
         _______4____2________________4____________________,
         _______2____2________________2____________________,
         _______0____2________________0____________________,
         _______28____2________________28____________________,
         _______27____2________________27____________________,
         _______18____2________________18____________________,
         _______15____2________________15____________________,
         _______13____2________________13____________________,
         _______10____2________________10____________________,
         _______7____2________________7____________________,
         ____3____________9_____, ____0___________0_5_____,
         ____1____________11_____, _________________________________6_________,
         _________________________________________2_________,
         ______________________________70________,
         _______14____2________________14____________________,
         _______24____2________________24____________________,
         _______11____2________________11____________________,
         _________________________________31_________,
         _________________________________27_________,
         _________________________________25_________,
         _________________________________24_________,
         _________________________________17_________,
         _________________________________11_________,
         _________________________________10_________,
         _________________________________9_________,
         _________________________________5_________,
         _________________________________2_________,
         _________________________________1_________,
         _________________________________0_________,
         _____________________________225________,
         _____________________________227________,
         _____________________________236________,
         _____________________________237________,
         _____________________________239________,
         _____________________________243________,
         _____________________________245________,
         _____________________________248________,
         _____________________________249________,
         _____________________________250________,
         _____________________________251________,
         _____________________________254________,
         _____________________________194________,
         _____________________________197________,
         _____________________________198________,
         _____________________________199________,
         _____________________________200________,
         _____________________________202________,
         _____________________________205________,
         _____________________________208________,
         _____________________________210________,
         _____________________________211________,
         _____________________________217________,
         _____________________________220________,
         _____________________________162________,
         _____________________________165________,
         _____________________________167________,
         _____________________________168________,
         _____________________________173________,
         _____________________________176________,
         _____________________________177________,
         _____________________________179________,
         _____________________________181________,
         _____________________________183________,
         _____________________________184________,
         _____________________________132________,
         _____________________________133________,
         _____________________________135________,
         _____________________________140________,
         _____________________________141________,
         _____________________________142________,
         _____________________________145________,
         _____________________________146________,
         _____________________________150________,
         _____________________________153________,
         _____________________________154________,
         _____________________________98________,
         _____________________________99________,
         _____________________________101________,
         _____________________________109________,
         _____________________________111________,
         _____________________________115________,
         _____________________________116________,
         _____________________________119________,
         _____________________________122________,
         _____________________________125________,
         _____________________________126________,
         _____________________________71________,
         _____________________________74________,
         _____________________________78________,
         _____________________________79________,
         _____________________________86________,
         _____________________________90________,
         _____________________________91________,
         _____________________________93________,
         _____________________________35________,
         _____________________________37________,
         _____________________________41________,
         _____________________________44________,
         _____________________________48________,
         _____________________________52________,
         _____________________________5________,
         _____________________________8________,
         _____________________________9________,
         _____________________________12________,
         _____________________________13________,
         _____________________________16________,
         _____________________________17________,
         _____________________________19________,
         _____________________________20________,
         _____________________________22________,
         _____________________________24________,
         _____________________________29________,
         _________________________________________3_________,
         _________________________________________18_________,
         _________________________________________22_________,
         _________________________________________23_________,
         _________________________________________0_________,
         _________________________________________0________1____________,
         _________________________________________0________3____________,
         ______________________________129________,
         ______________________________130________,
         ______________________________131________,
         ______________________________132________,
         ______________________________137________,
         ______________________________140________,
         ______________________________143________,
         ______________________________146________,
         ______________________________148________,
         ______________________________150________,
         ______________________________152________,
         ______________________________154________,
         ______________________________155________,
         ______________________________158________,
         ______________________________68________,
         ______________________________74________,
         ______________________________78________,
         ______________________________82________,
         ______________________________83________,
         ______________________________84________,
         ______________________________87________,
         ______________________________96________,
         ______________________________2________,
         ______________________________6________,
         ______________________________7________,
         ______________________________10________,
         ______________________________11________,
         ______________________________16________,
         ______________________________22________,
         ______________________________23________,
         ______________________________24________,
         ______________________________26________,
         ______________________________27________,
         ______________________________28________,
         ______________________________30________,
         ______________________________32________,
         __________________________________19_________,
         __________________________________7_________,
         _______29____2________________29____________________,
         _____________________________258________,
         _____________________________259________,
         _____________________________261________,
         _____________________________262________,
         _____________________________267________,
         _____________________________272________,
         _____________________________277________,
         _____________________________281________,
         _____________________________284________,
         _____________________________287________,
         ______________________________162________,
         ______________________________98________,
         ______________________________62________,
         ______________________________161________,
         ______________________________164________,
         ______________________________165________,
         ______________________________166________,
         ______________________________168________,
         ______________________________172________,
         ______________________________173________,
         ______________________________179________,
         ______________________________181________,
         ______________________________185________,
         ______________________________188________,
         ______________________________97________,
         ______________________________99________,
         ______________________________100________,
         ______________________________101________,
         ______________________________116________,
         ______________________________117________,
         ______________________________118________,
         ______________________________119________,
         ______________________________122________,
         ______________________________123________,
         ______________________________124________,
         ______________________________126________,
         ______________________________33________,
         ______________________________36________,
         ______________________________38________,
         ______________________________39________,
         ______________________________41________,
         ______________________________43________,
         ______________________________44________,
         ______________________________47________,
         ______________________________50________,
         ______________________________54________,
         ______________________________56________,
         ______________________________57________,
         ______________________________61________,
         __________________________________________2_________,
         __________________________________________3_________,
         __________________________________________6_________,
         __________________________________________7_________,
         __________________________________________11_________,
         __________________________________________14_________,
         __________________________________________15_________,
         __________________________________________17_________,
         __________________________________________19_________,
         __________________________________________23_________,
         __________________________________________4_________,
         __________________________________________8_________,
         __________________________________________25________0____________,
         ____3____________1_____, ____3____________2_____,
         ____1____________4_____, ____0___________0_12_____,
         ____0___________0_9_____, ____0___________0_8_____,
         ____0____________0_____, ____0____________11_____,
         ____0____________6_____, ____0____________4_____,
         ____0____________7_____, ____0____________1_____,
         ____0____________8_____, ____0____________3_____,
         ____0____________5_____, ____0____________9_____,
         ____0____________2_____, ____1____________9_____,
         ____1____________8_____, ____1____________2_____,
         ____1____________5_____, ____1____________7_____,
         ____1____________10_____, ____1____________1_____,
         ____1____________3_____, ____2____________10_____,
         ____2____________7_____, ____2____________11_____,
         ____2____________8_____, ____2____________6_____,
         ____2____________13_____, ____2____________9_____,
         ____2____________12_____, _____________________________216________,
         _____________________________190________,
         _____________________________120________,
         _____________________________127________,
         _____________________________92________,
         _____________________________49________,
         _____________________________7________,
         ______________________________77________,
         ______________________________8________,
         __________________________________18_________,
         __________________________________12_________,
         _____________________________191________,
         _________________________________26_________,
         _____________________________30________,
         _________________________________23_________,
         _____________________________255________,
         _____________________________222________,
         _____________________________39________,
         ______________________________90________,
         ______________________________18________,
         _____________________________201________,
         _____________________________213________,
         _____________________________224________,
         ______________________________141________,
         ______________________________17________,
         ______________________________20________,
         _________________________________30_________,
         _________________________________20_________,
         _________________________________19_________,
         _____________________________131________,
         _____________________________139________,
         _____________________________155________,
         _____________________________72________,
         _____________________________73________,
         _____________________________76________,
         _____________________________77________,
         _____________________________50________,
         _____________________________6________,
         _____________________________11________,
         _________________________________________16_________,
         _________________________________________24_________,
         ______________________________85________,
         _____________________________209________,
         _____________________________174________,
         _____________________________54________,
         ______________________________157________,
         ______________________________21________,
         __________________________________24_________,
         ______________________________182________,
         __________________________________1_________,
         ______________________________105________,
         _____________________________180________,
         ______________________________14________,
         _____________________________192________,
         ______________________________92________,
         __________________________________30_________,
         ______________________________171________,
         _________________________________29_________,
         _____________________________43________,
         ______________________________159________,
         _____________________________128________,
         ______________________________89________,
         _____________________________64________,
         _____________________________223________,
         _____________________________97________,
         _________________________________13_________,
         _____________________________31________,
         _____________________________256________,
         ______________________________71________,
         _____________________________226________,
         _____________________________241________,
         _________________________________________0________4____________,
         _________________________________________1_________,
         _________________________________________10_________,
         _____________________________67________,
         __________________________________9_________,
         _____________________________232________,
         _________________________________________0________0____________,
         _____________________________95________,
         _____________________________188________,
         _________________________________22_________,
         _____________________________160________,
         _____________________________195________,
         _______30____2________________30____________________,
         _____________________________242________,
         _________________________________________21_________,
         __________________________________20_________,
         __________________________________17_________,
         __________________________________16_________,
         ______________________________153________,
         _____________________________286________,
         _____________________________285________,
         ______________________________63________,
         ______________________________106________,
         __________________________________________5_________,
         ______________________________58________,
         ______________________________180________,
         ______________________________46________,
         _____________________________271________,
         _____________________________62________,
         ______________________________156________,
         __________________________________11_________,
         __________________________________8_________,
         __________________________________3_________,
         ______________________________133________,
         ______________________________139________,
         ______________________________149________,
         ______________________________151________,
         ______________________________79________,
         ______________________________134________,
         _____________________________275________,
         _____________________________279________,
         _____________________________264________,
         ______________________________163________,
         __________________________________________22_________,
         _____________________________268________,
         _____________________________151________,
         ______________________________76________,
         _____________________________152________,
         _____________________________117________,
         _____________________________118________,
         _____________________________121________,
         _____________________________10________,
         _________________________________________15_________,
         ______________________________138________,
         ______________________________49________,
         ______________________________80________,
         ______________________________183________,
         _________________________________14_________,
         __________________________________5_________,
         __________________________________________18_________,
         __________________________________10_________,
         _____________________________263________,
         ______________________________102________,
         ______________________________110________,
         ______________________________114________,
         __________________________________________25________5____________,
         ______________________________37________,
         ______________________________187________,
         _____________________________229________,
         _____________________________113________,
         _____________________________114________,
         __________________________________________24_________,
         _____________________________112________,
         ______________________________73________,
         ______________________________127________,
         ______________________________175________,
         __________________________________________13_________,
         _____________________________189________,
         ______________________________170________, ____3____________8_____,
         ______________________________103________,
         _____________________________66________,
         _____________________________129________,
         ______________________________167________,
         ______________________________190________,
         __________________________________________25________1____________,
         _____________________________193________,
         ______________________________184________,
         ______________________________112________,
         _________________________________21_________,
         _____________________________273________,
         _____________________________47________,
         ______________________________66________,
         __________________________________22_________,
         _____________________________84________,
         ______________________________145________,
         _____________________________82________,
         _____________________________25________,
         __________________________________31_________,
         __________________________________________20_________,
         ______________________________51________,
         ______________________________192________,
         ______________________________69________,
         ______________________________94________,
         _____________________________61________,
         ______________________________135________,
         ______________________________45________,
         _____________________________157________,
         _____________________________68________,
         _____________________________228________,
         _____________________________123________,
         ______________________________186________,
         ______________________________109________,
         ______________________________42________,
         __________________________________________10_________,
         ____3____________0_____, _____________________________196________,
         _____________________________178________,
         _____________________________147________,
         _____________________________104________,
         _____________________________89________,
         _____________________________42________,
         _____________________________45________,
         _____________________________46________,
         _____________________________23________,
         _________________________________________4_________,
         ______________________________93________,
         ______________________________29________,
         _____________________________53________,
         _____________________________244________,
         _____________________________149________,
         _____________________________124________,
         _____________________________36________,
         _____________________________56________,
         ______________________________142________,
         ______________________________160________,
         _________________________________________0________5____________,
         ______________________________67________,
         ______________________________34________, ____0____________12_____,
         ______________________________108________,
         ______________________________177________,
         ______________________________64________,
         _____________________________269________,
         _____________________________235________,
         _____________________________231________,
         ______________________________48________,
         _____________________________130________,
         ______________________________40________,
         _____________________________257________,
         ______________________________125________,
         __________________________________________25________3____________,
         _____________________________260________, ____2____________5_____,
         ____2____________4_____, ______________________________52________,
         _________________________________8_________,
         _____________________________100________,
         _____________________________69________,
         _____________________________134________,
         _____________________________158________,
         _________________________________________20_________,
         _________________________________28_________,
         _____________________________204________,
         _____________________________221________,
         _________________________________________0________2____________,
         __________________________________27_________,
         _____________________________182________,
         _____________________________15________,
         _____________________________252________,
         ______________________________88________, ____2____________3_____,
         ____3____________7_____, _____________________________103________,
         _____________________________88________,
         _____________________________212________,
         _____________________________57________,
         ______________________________35________,
         __________________________________________25_________,
         _____________________________28________,
         ______________________________111________,
         __________________________________________1_________,
         _____________________________288________,
         _____________________________169________,
         _________________________________7_________,
         ______________________________144________,
         _____________________________246________,
         _____________________________4________,
         _____________________________14________,
         ______________________________178________,
         _____________________________186________,
         _____________________________240________,
         __________________________________28_________,
         _____________________________33________,
         _____________________________65________,
         ______________________________9________,
         ______________________________13________,
         _________________________________4_________,
         ______________________________4________,
         _________________________________________25_________,
         __________________________________________25________4____________,
         _____________________________144________,
         _____________________________219________,
         _____________________________207________,
         _________________________________________8_________,
         ____0___________0_1_____, _____________________________107________,
         _____________________________80________,
         _____________________________26________,
         _________________________________________11_________,
         _____________________________148________,
         _____________________________55________,
         ______________________________19________,
         ______________________________147________,
         _____________________________27________,
         ______________________________91________,
         _____________________________282________,
         _____________________________214________,
         ______________________________72________,
         ______________________________12________,
         _____________________________233________,
         ______________________________176________,
         __________________________________________25________2____________,
         _____________________________266________,
         _____________________________2________,
         _________________________________________5_________,
         _____________________________171________, ____2____________0_____,
         _____________________________21________,
         _____________________________32________,
         _____________________________203________,
         __________________________________13_________,
         __________________________________6_________, ____2____________1_____,
         _____________________________276________,
         _____________________________234________, ____0____________15_____,
         _____________________________63________,
         _____________________________175________,
         _____________________________59________,
         _____________________________161________,
         _____________________________85________,
         _____________________________143________,
         _____________________________156________,
         _____________________________108________,
         _____________________________58________,
         _____________________________253________,
         ______________________________1________,
         _____________________________187________,
         ______________________________60________, ____1____________6_____,
         ______________________________53________, ____0____________10_____,
         ______________________________107________,
         _____________________________34________,
         __________________________________25_________,
         _________________________________________6_________,
         __________________________________________12_________,
         _____________________________280________,
         _____________________________283________,
         __________________________________________0_________,
         _____________________________83________,
         _____________________________215________,
         __________________________________________9_________,
         _____________________________70________,
         _____________________________137________,
         __________________________________15_________,
         ______________________________121________,
         _____________________________106________,
         ______________________________113________,
         _____________________________278________,
         _____________________________102________,
         _____________________________185________,
         _____________________________18________,
         _____________________________274________,
         _____________________________75________,
         _____________________________38________,
         ______________________________189________,
         _____________________________138________,
         ______________________________115________,
         _____________________________166________,
         _____________________________170________,
         __________________________________4_________,
         ____0____________14_____, _____________________________230________,
         __________________________________2_________,
         _____________________________159________,
         _________________________________3_________,
         _________________________________15_________,
         _____________________________164________,
         ______________________________136________,
         ______________________________81________,
         _________________________________16_________, ____3____________4_____,
         _____________________________1________,
         _____________________________110________,
         _____________________________3________,
         ______________________________5________,
         ______________________________25________,
         __________________________________________16_________,
         ____2____________2_____, ____3____________10_____,
         _____________________________60________, ____0___________0_2_____,
         ____0___________0_4_____,
         _________________________________18_________,
         ____0____________13_____, ______________________________174________,
         ______________________________75________,
         __________________________________23_________,
         ______________________________104________,
         __________________________________14_________,
         _________________________________________9_________,
         _____________________________163________,
         _____________________________105________,
         _____________________________81________,
         ______________________________120________,
         ______________________________169________,
         __________________________________29_________,
         _____________________________247________,
         _____________________________172________,
         ______________________________95________,
         _____________________________96________,
         _________________________________12_________,
         ____0___________0_6_____, ____0___________0_7_____,
         __________________________________________21_________,
         _____________________________270________,
         _____________________________265________, ____3____________5_____,
         _____________________________94________,
         ______________________________191________,
         __________________________________26_________,
         ____0___________0_3_____, ______________________________128________,
         ______________________________55________,
         ______________________________59________, ____0___________0_0_____,
         _____________________________206________,
         __________________________________0_________,
         _______6____2________________6____________________,
         _____________________________87________,
         _____________________________136________, ____0___________0_11_____,
         _____________________________238________, ____3____________3_____,
         ______________________________65________,
         _____________________________218________,
         _____________________________51________, ____1____________0_____,
         ____0___________0_10_____, ______________________________15________,
         ______________________________86________,
         __________________________________21_________, _14172, _15544, _15546,
         _15547, _15550, _15551, _15553, _15555, _15560, _922,
         _______12____2________________12____________________,
         _______31____2________________31____________________,
         _____________________________40________, ____3____________6_____,
         _______19____2________________19____________________,
         _______3____2________________3____________________,
         ____0___________0_13_____, ______________________________3________,
         ______________________________31________,
         _________________________________________7_________,
         _________________________________________12_________,
         _________________________________________19_________,
         _________________________________________13_________,
         _________________________________________14_________,
         _________________________________________17_________, _15563, _15561,
         _353, _355, _356, _359, _382, _398, _408, _414, _420, _424, _433,
         _438, _441, _640, _648, _652, _654, _1824, _1825, _1826, _1827, _1851,
         _1852, _1853, _1860, _1863, _1876, _1877, _1986, _2006, _2015, _2022,
         _2023, _2025, _2026, _2027, _2030, _2031, _2056, _2057, _2061, _2062,
         _2063, _2064, _2175, _2179, _2180, _2181, _2182, _2203, _2214, _2216,
         _2217, _2238, _2251, _2252, _2253, _2273, _2274, _2320, _2395, _2429,
         _2432, _2439, _2440, _2472, _2473, _2474, _2571, _2575, _2576, _2590,
         _2598, _2599, _2624, _2625, _2627, _2628, _2637, _2642, _2643, _2684,
         _2697, _2698, _2699, _2711, _2718, _2722, _2724, _2730, _2731, _26204,
         _26205, _26206, _26207, _26208, _26209, _26210, _26211, _26212,
         _26213, _26214, _26215, _26216, _26217, _26218, _26219, _26220,
         _26221, _26222, _26223, _26224, _26225, _26226, _26227, _26228,
         _26229, _26230, _26231, _26232, _26233, _26234, _26235, _26236,
         _26237, _26238, _26239, _26240, _26241, _26242, _26243, _26244,
         _26245, _26246, _26247, _26248, _26249, _26250, _26251, _26252,
         _26253, _26254, _26255, _26256, _26257, _26258, _26259, _26260,
         _26261, _26262, _26263, _26264, _26265, _26266, _26267, _26268,
         _26269, _26270, _26271, _26272, _26273, _26274, _26275, _26276,
         _26277, _26278, _26279, _26280, _26281, _26282, _26283, _26284,
         _26285, _26286, _26287, _26288, _26289, _26290, _26291, _26292,
         _26293, _26294, _26295, _26296, _26297, _26298, _26299, _26300,
         _26301, _26302, _26303, _26304, _26305, _26306, _26307, _26308,
         _26309, _26310, _26311, _26312, _26313, _26314, _26315, _26316,
         _26317, _26318, _26319, _26320, _26321, _26322, _26323, _26324,
         _26325, _26326, _26327, _26328, _26329, _26330, _26331, _26332,
         _26333, _26334, _26335, _26336, _26337, _26338, _26339, _26340,
         _26341, _26342, _26343, _26344, _26345, _26346, _26347, _26348,
         _26349, _26350, _26351, _26352, _26353, _26354, _26355, _26356,
         _26357, _26358, _26359, _26360, _26361, _26362, _26363, _26364,
         _26365, _26366, _26367, _26368, _26369, _26370, _26371, _26372,
         _26373, _26374, _26375, _26376, _26377, _26378, _26379, _26380,
         _26381, _26382, _26383, _26384, _26385, _26386, _26387, _26388,
         _26389, _26390, _26391, _26392, _26393, _26394, _26395, _26396,
         _26397, _26398, _26399, _26400, _26401, _26402, _26403, _26404,
         _26405, _26406, _26407, _26408, _26409, _26410, _26411, _26412,
         _26413, _26414, _26415, _26416, _26417, _26418, _26419, _26420,
         _26421, _26422, _26423, _26424, _26425, _26426, _26427, _26428,
         _26429, _26430, _26431, _26432, _26433, _26434, _26435, _26436,
         _26437, _26438, _26439, _26440, _26441, _26442, _26443, _26444,
         _26445, _26446, _26447, _26448, _26449, _26450, _26451, _26452,
         _26453, _26454, _26455, _26456, _26457, _26458, _26459, _26460,
         _26461, _26462, _26463, _26464, _26465, _26466, _26467, _26468,
         _26469, _26470, _26471, _26472, _26473, _26474, _26475, _26476,
         _26477, _26478, _26479, _26480, _26481, _26482, _26483, _26484,
         _26485, _26486, _26487, _26488, _26489, _26490, _26491, _26492,
         _26493, _26494, _26495, _26496, _26497, _26498, _26499, _26500,
         _26501, _26502, _26503, _26504, _26505, _26506, _26507, _26508,
         _26509, _26510, _26511, _26512, _26513, _26514, _26515, _26516,
         _26517, _26518, _26519, _26520, _26521, _26522, _26523, _26524,
         _26525, _26526, _26527, _26528, _26529, _26530, _26531, _26532,
         _26533, _26534, _26535, _26536, _26537, _26538, _26539, _26540,
         _26541, _26542, _26543, _26544, _26545, _26546, _26547, _26548,
         _26549, _26550, _26551, _26552, _26553, _26554, _26555, _26556,
         _26557, _26558, _26559, _26560, _26561, _26562, _26563, _26564,
         _26565, _26566, _26567, _26568, _26569, _26570, _26571, _26572,
         _26573, _26574, _26575, _26576, _26577, _26578, _26579, _26580,
         _26581, _26582, _26583, _26584, _26585, _26586, _26587, _26588,
         _26589, _26590, _26591, _26592, _26593, _26594, _26595, _26596,
         _26597, _26598, _26599, _26600, _26601, _26602, _26603, _26604,
         _26605, _26606, _26607, _26608, _26609, _26610, _26611, _26612,
         _26613, _26614, _26615, _26616, _26617, _26618, _26619, _26620,
         _26621, _26622, _26623, _26624, _26625, _26626, _26627, _26628,
         _26629, _26630, _26631, _26632, _26633, _26634, _26635, _26636,
         _26637, _26638, _26639, _26640, _26641, _26642, _26643, _26644,
         _26645, _26646, _26647, _26648, _26649, _26650, _26651, _26652,
         _26653, _26654, _26655, _26656, _26657, _26658, _26659, _26660,
         _26661, _26662, _26663, _26664, _26665, _26666, _26667, _26668,
         _26669, _26670, _26671, _26672, _26673, _26674, _26675, _26676,
         _26677, _26678, _26679, _26680, _26681, _26682, _26683, _26684,
         _26685, _26686, _26687, _26688, _26689, _26690, _26691, _26692,
         _26693, _26694, _26695, _26696, _26697, _26698, _26699, _26700,
         _26701, _26702, _26703, _26704, _26705, _26706, _26707, _26708,
         _26709, _26710, _26711, _26712, _26713, _26714, _26715, _26716,
         _26717, _26718, _26719, _26720, _26721, _26722, _26723, _26724,
         _26725, _26726, _26727, _26728, _26729, _26730, _26731, _26732,
         _26733, _26734, _26735, _26736, _26737, _26738, _26739, _26740,
         _26741, _26742, _26743, _26744, _26745, _26746, _26747, _26748,
         _26749, _26750, _26751, _26752, _26753, _26754, _26755, _26756,
         _26757, _26758, _26759, _26760, _26761, _26762, _26763, _26764,
         _26765, _26766, _26767, _26768, _26769, _26770, _26771, _26772,
         _26773, _26774, _26775, _26776, _26777, _26778, _26779, _26780,
         _26781, _26782, _26783, _26784, _26785, _26786, _26787, _26788,
         _26789, _26790, _26791, _26792, _26793, _26794, _26795, _26796,
         _26797, _26798, _26799, _26800, _26801, _26802, _26803, _26804,
         _26805, _26806, _26807, _26808, _26809, _26810, _26811, _26812,
         _26813, _26814, _26815, _26816, _26817, _26818, _26819, _26820,
         _26821, _26822, _26823, _26824, _26825, _26826, _26827, _26828,
         _26829, _26830, _26831, _26832, _26833, _26834, _26835, _26836,
         _26837, _26838, _26839, _26840, _26841, _26842, _26843, _26844,
         _26845, _26846, _26847, _26848, _26849, _26850, _26851, _26852,
         _26853, _26854, _26855, _26856, _26857, _26858, _26859, _26860,
         _26861, _26862, _26863, _26864, _26865, _26866, _26867, _26868,
         _26869, _26870, _26871, _26872, _26873, _26874, _26875, _26876,
         _26877, _26878, _26879, _26880, _26881, _26882, _26883, _26884,
         _26885, _26886, _26887, _26888, _26889, _26890, _26891, _26892,
         _26893, _26894, _26895, _26896, _26897, _26898, _26899, _26900,
         _26901, _26902, _26903, _26904, _26905, _26906, _26907, _26908,
         _26909, _26910, _26911, _26912, _26913, _26914, _26915, _26916,
         _26917, _26918, _26919, _26920, _26921, _26922, _26923, _26924,
         _26925, _26926, _26927, _26928, _26929, _26930, _26931, _26932,
         _26933, _26934, _26935, _26936, _26937, _26938, _26939, _26940,
         _26941, _26942, _26943, _26944, _26945, _26946, _26947, _26948,
         _26949, _26950, _26951, _26952, _26953, _26954, _26955, _26956,
         _26957, _26958, _26959, _26960, _26961, _26962, _26963, _26964,
         _26965, _26966, _26967, _26968, _26969, _26970, _26971, _26972,
         _26973, _26974, _26975, _26976, _26977, _26978, _26979, _26980,
         _26981, _26982, _26983, _26984, _26985, _26986, _26987, _26988,
         _26989, _26990, _26991, _26992, _26993, _26994, _26995, _26996,
         _26997, _26998, _26999, _27000, _27001, _27002, _27003, _27004,
         _27005, _27006, _27007, _27008, _27009, _27010, _27011, _27012,
         _27013, _27014, _27015, _27016, _27017, _27018, _27019, _27020,
         _27021, _27022, _27023, _27024, _27025, _27026, _27027, _27028,
         _27029, _27030, _27031, _27032, _27033, _27034, _27035, _27036,
         _27037, _27038, _27039, _27040, _27041, _27042, _27043, _27044,
         _27045, _27046, _27047, _27048, _27049, _27050, _27051, _27052,
         _27053, _27054, _27055, _27056, _27057, _27058, _27059, _27060,
         _27061, _27062, _27063, _27064, _27065, _27066, _27067, _27068,
         _27069, _27070, _27071, _27072, _27073, _27074, _27075, _27076,
         _27077, _27078, _27079, _27080, _27081, _27082, _27083, _27084,
         _27085, _27086, _27087, _27088, _27089, _27090, _27091, _27092,
         _27093, _27094, _27095, _27096, _27097, _27098, _27099, _27100,
         _27101, _27102, _27103, _27104, _27105, _27106, _27107, _27108,
         _27109, _27110, _27111, _27112, _27113, _27114, _27115, _27116,
         _27117, _27118, _27119, _27120, _27121, _27122, _27123, _27124,
         _27125, _27126, _27127, _27128, _27129, _27130, _27131, _27132,
         _27133, _27134, _27135, _27136, _27137, _27138, _27139, _27140,
         _27141, _27142, _27143, _27144, _27145, _27146, _27147, _27148,
         _27149, _27150, _27151, _27152, _27153, _27154, _27155, _27156,
         _27157, _27158, _27159, _27160, _27161, _27162, _27163, _27164,
         _27165, _27166, _27167, _27168, _27169, _27170, _27171, _27172,
         _27173, _27174, _27175, _27176, _27177, _27178, _27179, _27180,
         _27181, _27182, _27183, _27184, _27185, _27186, _27187, _27188,
         _27189, _27190, _27191, _27192, _27193, _27194, _27195, _27196,
         _27197, _27198, _27199, _27200, _27201, _27202, _27203, _27204,
         _27205, _27206, _27207, _27208, _27209, _27210, _27211, _27212,
         _27213, _27214, _27215, _27216, _27217, _27218, _27219, _27220,
         _27221, _27222, _27223, _27224, _27225, _27226, _27227, _27228,
         _27229, _27230, _27231, _27232, _27233, _27234, _27235, _27236,
         _27237, _27238, _27239, _27240, _27241, _27242, _27243, _27244,
         _27245, _27246, _27247, _27248, _27249, _27250, _27251, _27252,
         _27253, _27254, _27255, _27256, _27257, _27258, _27259, _27260,
         _27261, _27262, _27263, _27264, _27265, _27266, _27267, _27268,
         _27269, _27270, _27271, _27272, _27273, _27274, _27275, _27276,
         _27277, _27278, _27279, _27280, _27281, _27282, _27283, _27284,
         _27285, _27286, _27287, _27288, _27289, _27290, _27291, _27292,
         _27293, _27294, _27295, _27296, _27297, _27298, _27299, _27300,
         _27301, _27302, _27303, _27304, _27305, _27306, _27307, _27308,
         _27309, _27310, _27311, _27312, _27313, _27314, _27315, _27316,
         _27317, _27318, _27319, _27320, _27321, _27322, _27323, _27324,
         _27325, _27326, _27327, _27328, _27329, _27330, _27331, _27332,
         _27333, _27334, _27335, _27336, _27337, _27338, _27339, _27340,
         _27341, _27342, _27343, _27344, _27345, _27346, _27347, _27348,
         _27349, _27350, _27351, _27352, _27353, _27354, _27355, _27356,
         _27357, _27358, _27359, _27360, _27361, _27362, _27363, _27364,
         _27365, _27366, _27367, _27368, _27369, _27370, _27371, _27372,
         _27373, _27374, _27375, _27376, _27377, _27378, _27379, _27380,
         _27381, _27382, _27383, _27384, _27385, _27386, _27387, _27388,
         _27389, _27390, _27391, _27392, _27393, _27394, _27395, _27396,
         _27397, _27398, _27399, _27400, _27401, _27402, _27403, _27404,
         _27405, _27406, _27407, _27408, _27409, _27410, _27411, _27412,
         _27413, _27414, _27415, _27416, _27417, _27418, _27419, _27420,
         _27421, _27422, _27423, _27424, _27425, _27426, _27427, _27428,
         _27429, _27430, _27431, _27432, _27433, _27434, _27435, _27436,
         _27437, _27438, _27439, _27440, _27441, _27442, _27443, _27444,
         _27445, _27446, _27447, _27448, _27449, _27450, _27451, _27452,
         _27453, _27454, _27455, _27456, _27457, _27458, _27459, _27460,
         _27461, _27462, _27463, _27464, _27465, _27466, _27467, _27468,
         _27469, _27470, _27471, _27472, _27473, _27474, _27475, _27476,
         _27477, _27478, _27479, _27480, _27481, _27482, _27483, _27484,
         _27485, _27486, _27487, _27488, _27489, _27490, _27491, _27492,
         _27493, _27494, _27495, _27496, _27497, _27498, _27499, _27500,
         _27501, _27502, _27503, _27504, _27505, _27506, _27507, _27508,
         _27509, _27510, _27511, _27512, _27513, _27514, _27515, _27516,
         _27517, _27518, _27519, _27520, _27521, _27522, _27523, _27524,
         _27525, _27526, _27527, _27528, _27529, _27530, _27531, _27532,
         _27533, _27534, _27535, _27536, _27537, _27538, _27539, _27540,
         _27541, _27542, _27543, _27544, _27545, _27546, _27547, _27548,
         _27549, _27550, _27551, _27552, _27553, _27554, _27555, _27556,
         _27557, _27558, _27559, _27560, _27561, _27562, _27563, _27564,
         _27565, _27566, _27567, _27568, _27569, _27570, _27571, _27572,
         _27573, _27574, _27575, _27576, _27577, _27578, _27579, _27580,
         _27581, _27582, _27583, _27584, _27585, _27586, _27587, _27588,
         _27589, _27590, _27591, _27592, _27593, _27594, _27595, _27596,
         _27597, _27598, _27599, _27600, _27601, _27602, _27603, _27604,
         _27605, _27606, _27607, _27608, _27609, _27610, _27611, _27612,
         _27613, _27614, _27615, _27616, _27617, _27618, _27619, _27620,
         _27621, _27622, _27623, _27624, _27625, _27626, _27627, _27628,
         _27629, _27630, _27631, _27632, _27633, _27634, _27635, _27636,
         _27637, _27638, _27639, _27640, _27641, _27642, _27643, _27644,
         _27645, _27646, _27647, _27648, _27649, _27650, _27651, _27652,
         _27653, _27654, _27655, _27656, _27657, _27658, _27659, _27660,
         _27661, _27662, _27663, _27664, _27665, _27666, _27667, _27668,
         _27669, _27670, _27671, _27672, _27673, _27674, _27675, _27676,
         _27677, _27678, _27679, _27680, _27681, _27682, _27683, _27684,
         _27685, _27686, _27687, _27688, _27689, _27690, _27691, _27692,
         _27693, _27694, _27695, _27696, _27697, _27698, _27699, _27700,
         _27701, _27702, _27703, _27704, _27705, _27706, _27707, _27708,
         _27709, _27710, _27711, _27712, _27713, _27714, _27715, _27716,
         _27717, _27718, _27719, _27720, _27721, _27722, _27723, _27724,
         _27725, _27726, _27727, _27728, _27729, _27730, _27731, _27732,
         _27733, _27734, _27735, _27736, _27737, _27738, _27739, _27740,
         _27741, _27742, _27743, _27744, _27745, _27746, _27747, _27748,
         _27749, _27750, _27751, _27752, _27753, _27754, _27755, _27756,
         _27757, _27758, _27759, _27760, _27761, _27762, _27763, _27764,
         _27765, _27766, _27767, _27768, _27769, _27770, _27771, _27772,
         _27773, _27774, _27775, _27776, _27777, _27778, _27779, _27780,
         _27781, _27782, _27783, _27784, _27785, _27786, _27787, _27788,
         _27789, _27790, _27791, _27792, _27793, _27794, _27795, _27796,
         _27797, _27798, _27799, _27800, _27801, _27802, _27803, _27804,
         _27805, _27806, _27807, _27808, _27809, _27810, _27811, _27812,
         _27813, _27814, _27815, _27816, _27817, _27818, _27819, _27820,
         _27821, _27822, _27823, _27824, _27825, _27826, _27827, _27828,
         _27829, _27830, _27831, _27832, _27833, _27834, _27835, _27836,
         _27837, _27838, _27839, _27840, _27841, _27842, _27843, _27844,
         _27845, _27846, _27847, _27848, _27849, _27850, _27851, _27852,
         _27853, _27854, _27855, _27856, _27857, _27858, _27859, _27860,
         _27861, _27862, _27863, _27864, _27865, _27866, _27867, _27868,
         _27869, _27870, _27871, _27872, _27873, _27874, _27875, _27876,
         _27877, _27878, _27879, _27880, _27881, _27882, _27883, _27884,
         _27885, _27886, _27887, _27888, _27889, _27890, _27891, _27892,
         _27893, _27894, _27895, _27896, _27897, _27898, _27899, _27900,
         _27901, _27902, _27903, _27904, _27905, _27906, _27907, _27908,
         _27909, _27910, _27911, _27912, _27913, _27914, _27915, _27916,
         _27917, _27918, _27919, _27920, _27921, _27922, _27923, _27924,
         _27925, _27926, _27927, _27928, _27929, _27930, _27931, _27932,
         _27933, _27934, _27935, _27936, _27937, _27938, _27939, _27940,
         _27941, _27942, _27943, _27944, _27945, _27946, _27947, _27948,
         _27949, _27950, _27951, _27952, _27953, _27954, _27955, _27956,
         _27957, _27958, _27959, _27960, _27961, _27962, _27963, _27964,
         _27965, _27966, _27967, _27968, _27969, _27970, _27971, _27972,
         _27973, _27974, _27975, _27976, _27977, _27978, _27979, _27980,
         _27981, _27982, _27983, _27984, _27985, _27986, _27987, _27988,
         _27989, _27990, _27991, _27992, _27993, _27994, _27995, _27996,
         _27997, _27998, _27999, _28000, _28001, _28002, _28003, _28004,
         _28005, _28006, _28007, _28008, _28009, _28010, _28011, _28012,
         _28013, _28014, _28015, _28016, _28017, _28018, _28019, _28020,
         _28021, _28022, _28023, _28024, _28025, _28026, _28027, _28028,
         _28029, _28030, _28031, _28032, _28033, _28034, _28035, _28036,
         _28037, _28038, _28039, _28040, _28041, _28042, _28043, _28044,
         _28045, _28046, _28047, _28048, _28049, _28050, _28051, _28052,
         _28053, _28054, _28055, _28056, _28057, _28058, _28059, _28060,
         _28061, _28062, _28063, _28064, _28065, _28066, _28067, _28068,
         _28069, _28070, _28071, _28072, _28073, _28074, _28075, _28076,
         _28077, _28078, _28079, _28080, _28081, _28082, _28083, _28084,
         _28085, _28086, _28087, _28088, _28089, _28090, _28091, _28092,
         _28093, _28094, _28095, _28096, _28097, _28098, _28099, _28100,
         _28101, _28102, _28103, _28104, _28105, _28106, _28107, _28108,
         _28109, _28110, _28111, _28112, _28113, _28114, _28115, _28116,
         _28117, _28118, _28119, _28120, _28121, _28122, _28123, _28124,
         _28125, _28126, _28127, _28128, _28129, _28130, _28131, _28132,
         _28133, _28134, _28135, _28136, _28137, _28138, _28139, _28140,
         _28141, _28142, _28143, _28144, _28145, _28146, _28147, _28148,
         _28149, _28150, _28151, _28152, _28153, _28154, _28155, _28156,
         _28157, _28158, _28159, _28160, _28161, _28162, _28163, _28164,
         _28165, _28166, _28167, _28168, _28169, _28170, _28171, _28172,
         _28173, _28174, _28175, _28176, _28177, _28178, _28179, _28180,
         _28181, _28182, _28183, _28184, _28185, _28186, _28187, _28188,
         _28189, _28190, _28191, _28192, _28193, _28194, _28195, _28196,
         _28197, _28198, _28199, _28200, _28201, _28202, _28203, _28204,
         _28205, _28206, _28207, _28208, _28209, _28210, _28211, _28212,
         _28213, _28214, _28215, _28216, _28217, _28218, _28219, _28220,
         _28221, _28222, _28223, _28224, _28225, _28226, _28227, _28228,
         _28229, _28230, _28231, _28232, _28233, _28234, _28235, _28236,
         _28237, _28238, _28239, _28240, _28241, _28242, _28243, _28244,
         _28245, _28246, _28247, _28248, _28249, _28250, _28251, _28252,
         _28253, _28254, _28255, _28256, _28257, _28258, _28259, _28260,
         _28261, _28262, _28263, _28264, _28265, _28266, _28267, _28268,
         _28269, _28270, _28271, _28272, _28273, _28274, _28275, _28276,
         _28277, _28278, _28279, _28280, _28281, _28282, _28283, _28284,
         _28285, _28286, _28287, _28288, _28289, _28290, _28291, _28292,
         _28293, _28294, _28295, _28296, _28297, _28298, _28299, _28300,
         _28301, _28302, _28303, _28304, _28305, _28306, _28307, _28308,
         _28309, _28310, _28311, _28312, _28313, _28314, _28315, _28316,
         _28317, _28318, _28319, _28320, _28321, _28322, _28323, _28324,
         _28325, _28326, _28327, _28328, _28329, _28330, _28331, _28332,
         _28333, _28334, _28335, _28336, _28337, _28338, _28339, _28340,
         _28341, _28342, _28343, _28344, _28345, _28346, _28347, _28348,
         _28349, _28350, _28351, _28352, _28353, _28354, _28355, _28356,
         _28357, _28358, _28359, _28360, _28361, _28362, _28363, _28364,
         _28365, _28366, _28367, _28368, _28369, _28370, _28371, _28372,
         _28373, _28374, _28375, _28376, _28377, _28378, _28379, _28380,
         _28381, _28382, _28383, _28384, _28385, _28386, _28387, _28388,
         _28389, _28390, _28391, _28392, _28393, _28394, _28395, _28396,
         _28397, _28398, _28399, _28400, _28401, _28402, _28403, _28404,
         _28405, _28406, _28407, _28408, _28409, _28410, _28411, _28412,
         _28413, _28414, _28415, _28416, _28417, _28418, _28419, _28420,
         _28421, _28422, _28423, _28424, _28425, _28426, _28427, _28428,
         _28429, _28430, _28431, _28432, _28433, _28434, _28435, _28436,
         _28437, _28438, _28439, _28440, _28441, _28442, _28443, _28444,
         _28445, _28446, _28447, _28448, _28449, _28450, _28451, _28452,
         _28453, _28454, _28455, _28456, _28457, _28458, _28459, _28460,
         _28461, _28462, _28463, _28464, _28465, _28466, _28467, _28468,
         _28469, _28470, _28471, _28472, _28473, _28474, _28475, _28476,
         _28477, _28478, _28479, _28480, _28481, _28482, _28483, _28484,
         _28485, _28486, _28487, _28488, _28489, _28490, _28491, _28492,
         _28493, _28494, _28495, _28496, _28497, _28498, _28499, _28500,
         _28501, _28502, _28503, _28504, _28505, _28506, _28507, _28508,
         _28509, _28510, _28511, _28512, _28513, _28514, _28515, _28516,
         _28517, _28518, _28519, _28520, _28521, _28522, _28523, _28524,
         _28525, _28526, _28527, _28528, _28529, _28530, _28531, _28532,
         _28533, _28534, _28535, _28536, _28537, _28538, _28539, _28540,
         _28541, _28542, _28543, _28544, _28545, _28546, _28547, _28548,
         _28549, _28550, _28551, _28552, _28553, _28554, _28555, _28556,
         _28557, _28558, _28559, _28560, _28561, _28562, _28563, _28564,
         _28565, _28566, _28567, _28568, _28569, _28570, _28571, _28572,
         _28573, _28574, _28575, _28576, _28577, _28578, _28579, _28580,
         _28581, _28582, _28583, _28584, _28585, _28586, _28587, _28588,
         _28589, _28590, _28591, _28592, _28593, _28594, _28595, _28596,
         _28597, _28598, _28599, _28600, _28601, _28602, _28603, _28604,
         _28605, _28606, _28607, _28608, _28609, _28610, _28611, _28612,
         _28613, _28614, _28615, _28616, _28617, _28618, _28619, _28620,
         _28621, _28622, _28623, _28624, _28625, _28626, _28627, _28628,
         _28629, _28630, _28631, _28632, _28633, _28634, _28635, _28636,
         _28637, _28638, _28639, _28640, _28641, _28642, _28643, _28644,
         _28645, _28646, _28647, _28648, _28649, _28650, _28651, _28652,
         _28653, _28654, _28655, _28656, _28657, _28658, _28659, _28660,
         _28661, _28662, _28663, _28664, _28665, _28666, _28667, _28668,
         _28669, _28670, _28671, _28672, _28673, _28674, _28675, _28676,
         _28677, _28678, _28679, _28680, _28681, _28682, _28683, _28684,
         _28685, _28686, _28687, _28688, _28689, _28690, _28691, _28692,
         _28693, _28694, _28695, _28696, _28697, _28698, _28699, _28700,
         _28701, _28702, _28703, _28704, _28705, _28706, _28707, _28708,
         _28709, _28710, _28711, _28712, _28713, _28714, _28715, _28716,
         _28717, _28718, _28719, _28720, _28721, _28722, _28723, _28724,
         _28725, _28726, _28727, _28728, _28729, _28730, _28731, _28732,
         _28733, _28734, _28735, _28736, _28737, _28738, _28739, _28740,
         _28741, _28742, _28743, _28744, _28745, _28746, _28747, _28748,
         _28749, _28750, _28751, _28752, _28753, _28754, _28755, _28756,
         _28757, _28758, _28759, _28760, _28761, _28762, _28763, _28764,
         _28765, _28766, _28767, _28768, _28769, _28770, _28771, _28772,
         _28773, _28774, _28775, _28776, _28777, _28778, _28779, _28780,
         _28781, _28782, _28783, _28784, _28785, _28786, _28787, _28788,
         _28789, _28790, _28791, _28792, _28793, _28794, _28795, _28796,
         _28797, _28798, _28799, _28800, _28801, _28802, _28803, _28804,
         _28805, _28806, _28807, _28808, _28809, _28810, _28811, _28812,
         _28813, _28814, _28815, _28816, _28817, _28818, _28819, _28820,
         _28821, _28822, _28823, _28824, _28825, _28826, _28827, _28828,
         _28829, _28830, _28831, _28832, _28833, _28834, _28835, _28836,
         _28837, _28838, _28839, _28840, _28841, _28842, _28843, _28844,
         _28845, _28846, _28847, _28848, _28849, _28850, _28851, _28852,
         _28853, _28854, _28855, _28856, _28857, _28858, _28859, _28860,
         _28861, _28862, _28863, _28864, _28865, _28866, _28867, _28868,
         _28869, _28870, _28871, _28872, _28873, _28874, _28875, _28876,
         _28877, _28878, _28879, _28880, _28881, _28882, _28883, _28884,
         _28885, _28886, _28887, _28888, _28889, _28890, _28891, _28892,
         _28893, _28894, _28895, _28896, _28897, _28898, _28899, _28900,
         _28901, _28902, _28903, _28904, _28905, _28906, _28907, _28908,
         _28909, _28910, _28911, _28912, _28913, _28914, _28915, _28916,
         _28917, _28918, _28919, _28920, _28921, _28922, _28923, _28924,
         _28925, _28926, _28927, _28928, _28929, _28930, _28931, _28932,
         _28933, _28934, _28935, _28936, _28937, _28938, _28939, _28940,
         _28941, _28942, _28943, _28944, _28945, _28946, _28947, _28948,
         _28949, _28950, _28951, _28952, _28953, _28954, _28955, _28956,
         _28957, _28958, _28959, _28960, _28961, _28962, _28963, _28964,
         _28965, _28966, _28967, _28968, _28969, _28970, _28971, _28972,
         _28973, _28974, _28975, _28976, _28977, _28978, _28979, _28980,
         _28981, _28982, _28983, _28984, _28985, _28986, _28987, _28988,
         _28989, _28990, _28991, _28992, _28993, _28994, _28995, _28996,
         _28997, _28998, _28999, _29000, _29001, _29002, _29003, _29004,
         _29005, _29006, _29007, _29008, _29009, _29010, _29011, _29012,
         _29013, _29014, _29015, _29016, _29017, _29018, _29019, _29020,
         _29021, _29022, _29023, _29024, _29025, _29026, _29027, _29028,
         _29029, _29030, _29031, _29032, _29033, _29034, _29035, _29036,
         _29037, _29038, _29039, _29040, _29041, _29042, _29043, _29044,
         _29045, _29046, _29047, _29048, _29049, _29050, _29051, _29052,
         _29053, _29054, _29055, _29056, _29057, _29058, _29059, _29060,
         _29061, _29062, _29063, _29064, _29065, _29066, _29067, _29068,
         _29069, _29070, _29071, _29072, _29073, _29074, _29075, _29076,
         _29077, _29078, _29079, _29080, _29081, _29082, _29083, _29084,
         _29085, _29086, _29087, _29088, _29089, _29090, _29091, _29092,
         _29093, _29094, _29095, _29096, _29097, _29098, _29099, _29100,
         _29101, _29102, _29103, _29104, _29105, _29106, _29107, _29108,
         _29109, _29110, _29111, _29112, _29113, _29114, _29115, _29116,
         _29117, _29118, _29119, _29120, _29121, _29122, _29123, _29124,
         _29125, _29126, _29127, _29128, _29129, _29130, _29131, _29132,
         _29133, _29134, _29135, _29136, _29137, _29138, _29139, _29140,
         _29141, _29142, _29143, _29144, _29145, _29146, _29147, _29148,
         _29149, _29150, _29151, _29152, _29153, _29154, _29155, _29156,
         _29157, _29158, _29159, _29160, _29161, _29162, _29163, _29164,
         _29165, _29166, _29167, _29168, _29169, _29170, _29171, _29172,
         _29173, _29174, _29175, _29176, _29177, _29178, _29179, _29180,
         _29181, _29182, _29183, _29184, _29185, _29186, _29187, _29188,
         _29189, _29190, _29191, _29192, _29193, _29194, _29195, _29196,
         _29197, _29198, _29199, _29200, _29201, _29202, _29203, _29204,
         _29205, _29206, _29207, _29208, _29209, _29210, _29211, _29212,
         _29213, _29214, _29215, _29216, _29217, _29218, _29219, _29220,
         _29221, _29222, _29223, _29224, _29225, _29226, _29227, _29228,
         _29229, _29230, _29231, _29232, _29233, _29234, _29235, _29236,
         _29237, _29238, _29239, _29240, _29241, _29242, _29243, _29244,
         _29245, _29246, _29247, _29248, _29249, _29250, _29251, _29252,
         _29253, _29254, _29255, _29256, _29257, _29258, _29259, _29260,
         _29261, _29262, _29263, _29264, _29265, _29266, _29267, _29268,
         _29269, _29270, _29271, _29272, _29273, _29274, _29275, _29276,
         _29277, _29278, _29279, _29280, _29281, _29282, _29283, _29284,
         _29285, _29286, _29287, _29288, _29289, _29290, _29291, _29292,
         _29293, _29294, _29295, _29296, _29297, _29298, _29299, _29300,
         _29301, _29302, _29303, _29304, _29305, _29306, _29307, _29308,
         _29309, _29310, _29311, _29312, _29313, _29314, _29315, _29316,
         _29317, _29318, _29319, _29320, _29321, _29322, _29323, _29324,
         _29325, _29326, _29327, _29328, _29329, _29330, _29331, _29332,
         _29333, _29334, _29335, _29336, _29337, _29338, _29339, _29340,
         _29341, _29342, _29343, _29344, _29345, _29346, _29347, _29348,
         _29349, _29350, _29351, _29352, _29353, _29354, _29355, _29356,
         _29357, _29358, _29359, _29360, _29361, _29362, _29363, _29364,
         _29365, _29366, _29367, _29368, _29369, _29370, _29371, _29372,
         _29373, _29374, _29375, _29376, _29377, _29378, _29379, _29380,
         _29381, _29382, _29383, _29384, _29385, _29386, _29387, _29388,
         _29389, _29390, _29391, _29392, _29393, _29394, _29395, _29396,
         _29397, _29398, _29399, _29400, _29401, _29402, _29403, _29404,
         _29405, _29406, _29407, _29408, _29409, _29410, _29411, _29412,
         _29413, _29414, _29415, _29416, _29417, _29418, _29419, _29420,
         _29421, _29422, _29423, _29424, _29425, _29426, _29427, _29428,
         _29429, _29430, _29431, _29432, _29433, _29434, _29435, _29436,
         _29437, _29438, _29439, _29440, _29441, _29442, _29443, _29444,
         _29445, _29446, _29447, _29448, _29449, _29450, _29451, _29452,
         _29453, _29454, _29455, _29456, _29457, _29458, _29459, _29460,
         _29461, _29462, _29463, _29464, _29465, _29466, _29467, _29468,
         _29469, _29470, _29471, _29472, _29473, _29474, _29475, _29476,
         _29477, _29478, _29479, _29480, _29481, _29482, _29483, _29484,
         _29485, _29486, _29487, _29488, _29489, _29490, _29491, _29492,
         _29493, _29494, _29495, _29496, _29497, _29498, _29499, _29500,
         _29501, _29502, _29503, _29504, _29505, _29506, _29507, _29508,
         _29509, _29510, _29511, _29512, _29513, _29514, _29515, _29516,
         _29517, _29518, _29519, _29520, _29521, _29522, _29523, _29524,
         _29525, _29526, _29527, _29528, _29529, _29530, _29531, _29532,
         _29533, _29534, _29535, _29536, _29537, _29538, _29539, _29540,
         _29541, _29542, _29543, _29544, _29545, _29546, _29547, _29548,
         _29549, _29550, _29551, _29552, _29553, _29554, _29555, _29556,
         _29557, _29558, _29559, _29560, _29561, _29562, _29563, _29564,
         _29565, _29566, _29567, _29568, _29569, _29570, _29571, _29572,
         _29573, _29574, _29575, _29576, _29577, _29578, _29579, _29580,
         _29581, _29582, _29583, _29584, _29585, _29586, _29587, _29588,
         _29589, _29590, _29591, _29592, _29593, _29594, _29595, _29596,
         _29597, _29598, _29599, _29600, _29601, _29602, _29603, _29604,
         _29605, _29606, _29607, _29608, _29609, _29610, _29611, _29612,
         _29613, _29614, _29615, _29616, _29617, _29618, _29619, _29620,
         _29621, _29622, _29623, _29624, _29625, _29626, _29627, _29628,
         _29629, _29630, _29631, _29632, _29633, _29634, _29635, _29636,
         _29637, _29638, _29639, _29640, _29641, _29642, _29643, _29644,
         _29645, _29646, _29647, _29648, _29649, _29650, _29651, _29652,
         _29653, _29654, _29655, _29656, _29657, _29658, _29659, _29660,
         _29661, _29662, _29663, _29664, _29665, _29666, _29667, _29668,
         _29669, _29670, _29671, _29672, _29673, _29674, _29675, _29676,
         _29677, _29678, _29679, _29680, _29681, _29682, _29683, _29684,
         _29685, _29686, _29687, _29688, _29689, _29690, _29691, _29692,
         _29693, _29694, _29695, _29696, _29697, _29698, _29699, _29700,
         _29701, _29702, _29703, _29704, _29705, _29706, _29707, _29708,
         _29709, _29710, _29711, _29712, _29713, _29714, _29715, _29716,
         _29717, _29718, _29719, _29720, _29721, _29722, _29723, _29724,
         _29725, _29726, _29727, _29728, _29729, _29730, _29731, _29732,
         _29733, _29734, _29735, _29736, _29737, _29738, _29739, _29740,
         _29741, _29742, _29743, _29744, _29745, _29746, _29747, _29748,
         _29749, _29750, _29751, _29752, _29753, _29754, _29755, _29756,
         _29757, _29758, _29759, _29760, _29761, _29762, _29763, _29764,
         _29765, _29766, _29767, _29768, _29769, _29770, _29771, _29772,
         _29773, _29774, _29775, _29776, _29777, _29778, _29779, _29780,
         _29781, _29782, _29783, _29784, _29785, _29786, _29787, _29788,
         _29789, _29790, _29791, _29792, _29793, _29794, _29795, _29796,
         _29797, _29798, _29799, _29800, _29801, _29802, _29803, _29804,
         _29805, _29806, _29807, _29808, _29809, _29810, _29811, _29812,
         _29813, _29814, _29815, _29816, _29817, _29818, _29819, _29820,
         _29821, _29822, _29823, _29824, _29825, _29826, _29827, _29828,
         _29829, _29830, _29831, _29832, _29833, _29834, _29835, _29836,
         _29837, _29838, _29839, _29840, _29841, _29842, _29843, _29844,
         _29845, _29846, _29847, _29848, _29849, _29850, _29851, _29852,
         _29853, _29854, _29855, _29856, _29857, _29858, _29859, _29860,
         _29861, _29862, _29863, _29864, _29865, _29866, _29867, _29868,
         _29869, _29870, _29871, _29872, _29873, _29874, _29875, _29876,
         _29877, _29878, _29879, _29880, _29881, _29882, _29883, _29884,
         _29885, _29886, _29887, _29888, _29889, _29890, _29891, _29892,
         _29893, _29894, _29895, _29896, _29897, _29898, _29899, _29900,
         _29901, _29902, _29903, _29904, _29905, _29906, _29907, _29908,
         _29909, _29910, _29911, _29912, _29913, _29914, _29915, _29916,
         _29917, _29918, _29919, _29920, _29921, _29922, _29923, _29924,
         _29925, _29926, _29927, _29928, _29929, _29930, _29931, _29932,
         _29933, _29934, _29935, _29936, _29937, _29938, _29939, _29940,
         _29941, _29942, _29943, _29944, _29945, _29946, _29947, _29948,
         _29949, _29950, _29951, _29952, _29953, _29954, _29955, _29956,
         _29957, _29958, _29959, _29960, _29961, _29962, _29963, _29964,
         _29965, _29966, _29967, _29968, _29969, _29970, _29971, _29972,
         _29973, _29974, _29975, _29976, _29977, _29978, _29979, _29980,
         _29981, _29982, _29983, _29984, _29985, _29986, _29987, _29988,
         _29989, _29990, _29991, _29992, _29993, _29994, _29995, _29996,
         _29997, _29998, _29999, _30000, _30001, _30002, _30003, _30004,
         _30005, _30006, _30007, _30008, _30009, _30010, _30011, _30012,
         _30013, _30014, _30015, _30016, _30017, _30018, _30019, _30020,
         _30021, _30022, _30023, _30024, _30025, _30026, _30027, _30028,
         _30029, _30030, _30031, _30032, _30033, _30034, _30035, _30036,
         _30037, _30038, _30039, _30040, _30041, _30042, _30043, _30044,
         _30045, _30046, _30047, _30048, _30049, _30050, _30051, _30052,
         _30053, _30054, _30055, _30056, _30057, _30058, _30059, _30060,
         _30061, _30062, _30063, _30064, _30065, _30066, _30067, _30068,
         _30069, _30070, _30071, _30072, _30073, _30074, _30075, _30076,
         _30077, _30078, _30079, _30080, _30081, _30082, _30083, _30084,
         _30085, _30086, _30087, _30088, _30089, _30090, _30091, _30092,
         _30093, _30094, _30095, _30096, _30097, _30098, _30099, _30100,
         _30101, _30102, _30103, _30104, _30105, _30106, _30107, _30108,
         _30109, _30110, _30111, _30112, _30113, _30114, _30115, _30116,
         _30117, _30118, _30119, _30120, _30121, _30122, _30123, _30124,
         _30125, _30126, _30127, _30128, _30129, _30130, _30131, _30132,
         _30133, _30134, _30135, _30136, _30137, _30138, _30139, _30140,
         _30141, _30142, _30143, _30144, _30145, _30146, _30147, _30148,
         _30149, _30150, _30151, _30152, _30153, _30154, _30155, _30156,
         _30157, _30158, _30159, _30160, _30161, _30162, _30163, _30164,
         _30165, _30166, _30167, _30168, _30169, _30170, _30171, _30172,
         _30173, _30174, _30175, _30176, _30177, _30178, _30179, _30180,
         _30181, _30182, _30183, _30184, _30185, _30186, _30187, _30188,
         _30189, _30190, _30191, _30192, _30193, _30194, _30195, _30196,
         _30197, _30198, _30199, _30200, _30201, _30202, _30203, _30204,
         _30205, _30206, _30207, _30208, _30209, _30210, _30211, _30212,
         _30213, _30214, _30215, _30216, _30217, _30218, _30219, _30220,
         _30221, _30222, _30223, _30224, _30225, _30226, _30227, _30228,
         _30229, _30230, _30231, _30232, _30233, _30234, _30235, _30236,
         _30237, _30238, _30239, _30240, _30241, _30242, _30243, _30244,
         _30245, _30246, _30247, _30248, _30249, _30250, _30251, _30252,
         _30253, _30254, _30255, _30256, _30257, _30258, _30259, _30260,
         _30261, _30262, _30263, _30264, _30265, _30266, _30267, _30268,
         _30269, _30270, _30271, _30272, _30273, _30274, _30275, _30276,
         _30277, _30278, _30279, _30280, _30281, _30282, _30283, _30284,
         _30285, _30286, _30287, _30288, _30289, _30290, _30291, _30292,
         _30293, _30294, _30295, _30296, _30297, _30298, _30299, _30300,
         _30301, _30302, _30303, _30304, _30305, _30306, _30307, _30308,
         _30309, _30310, _30311, _30312, _30313, _30314, _30315, _30316,
         _30317, _30318, _30319, _30320, _30321, _30322, _30323, _30324,
         _30325, _30326, _30327, _30328, _30329, _30330, _30331, _30332,
         _30333, _30334, _30335, _30336, _30337, _30338, _30339, _30340,
         _30341, _30342, _30343, _30344, _30345, _30346, _30347, _30348,
         _30349, _30350, _30351, _30352, _30353, _30354, _30355, _30356,
         _30357, _30358, _30359, _30360, _30361, _30362, _30363, _30364,
         _30365, _30366, _30367, _30368, _30369, _30370, _30371, _30372,
         _30373, _30374, _30375, _30376, _30377, _30378, _30379, _30380,
         _30381, _30382, _30383, _30384, _30385, _30386, _30387, _30388,
         _30389, _30390, _30391, _30392, _30393, _30394, _30395, _30396,
         _30397, _30398, _30399, _30400, _30401, _30402, _30403, _30404,
         _30405, _30406, _30407, _30408, _30409, _30410, _30411, _30412,
         _30413, _30414, _30415, _30416, _30417, _30418, _30419, _30420,
         _30421, _30422, _30423, _30424, _30425, _30426, _30427, _30428,
         _30429, _30430, _30431, _30432, _30433, _30434, _30435, _30436,
         _30437, _30438, _30439, _30440, _30441, _30442, _30443, _30444,
         _30445, _30446, _30447, _30448, _30449, _30450, _30451, _30452,
         _30453, _30454, _30455, _30456, _30457, _30458, _30459, _30460,
         _30461, _30462, _30463, _30464, _30465, _30466, _30467, _30468,
         _30469, _30470, _30471, _30472, _30473, _30474, _30475, _30476,
         _30477, _30478, _30479, _30480, _30481, _30482, _30483, _30484,
         _30485, _30486, _30487, _30488, _30489, _30490, _30491, _30492,
         _30493, _30494, _30495, _30496, _30497, _30498, _30499, _30500,
         _30501, _30502, _30503, _30504, _30505, _30506, _30507, _30508,
         _30509, _30510, _30511, _30512, _30513, _30514, _30515, _30516,
         _30517, _30518, _30519, _30520, _30521, _30522, _30523, _30524,
         _30525, _30526, _30527, _30528, _30529, _30530, _30531, _30532,
         _30533, _30534, _30535, _30536, _30537, _30538, _30539, _30540,
         _30541, _30542, _30543, _30544, _30545, _30546, _30547, _30548,
         _30549, _30550, _30551, _30552, _30553, _30554, _30555, _30556,
         _30557, _30558, _30559, _30560, _30561, _30562, _30563, _30564,
         _30565, _30566, _30567, _30568, _30569, _30570, _30571, _30572,
         _30573, _30574, _30575, _30576, _30577, _30578, _30579, _30580,
         _30581, _30582, _30583, _30584, _30585, _30586, _30587, _30588,
         _30589, _30590, _30591, _30592, _30593, _30594, _30595, _30596,
         _30597, _30598, _30599, _30600, _30601, _30602, _30603, _30604,
         _30605, _30606, _30607, _30608, _30609, _30610, _30611, _30612,
         _30613, _30614, _30615, _30616, _30617, _30618, _30619, _30620,
         _30621, _30622, _30623, _30624, _30625, _30626, _30627, _30628,
         _30629, _30630, _30631, _30632, _30633, _30634, _30635, _30636,
         _30637, _30638, _30639, _30640, _30641, _30642, _30643, _30644,
         _30645, _30646, _30647, _30648, _30649, _30650, _30651, _30652,
         _30653, _30654, _30655, _30656, _30657, _30658, _30659, _30660,
         _30661, _30662, _30663, _30664, _30665, _30666, _30667, _30668,
         _30669, _30670, _30671, _30672, _30673, _30674, _30675, _30676,
         _30677, _30678, _30679, _30680, _30681, _30682, _30683, _30684,
         _30685, _30686, _30687, _30688, _30689, _30690, _30691, _30692,
         _30693, _30694, _30695, _30696, _30697, _30698, _30699, _30700,
         _30701, _30702, _30703, _30704, _30705, _30706, _30707, _30708,
         _30709, _30710, _30711, _30712, _30713, _30714, _30715, _30716,
         _30717, _30718, _30719, _30720, _30721, _30722, _30723, _30724,
         _30725, _30726, _30727, _30728, _30729, _30730, _30731, _30732,
         _30733, _30734, _30735, _30736, _30737, _30738, _30739, _30740,
         _30741, _30742, _30743, _30744, _30745, _30746, _30747, _30748,
         _30749, _30750, _30751, _30752, _30753, _30754, _30755, _30756,
         _30757, _30758, _30759, _30760, _30761, _30762, _30763, _30764,
         _30765, _30766, _30767, _30768, _30769, _30770, _30771, _30772,
         _30773, _30774, _30775, _30776, _30777, _30778, _30779, _30780,
         _30781, _30782, _30783, _30784, _30785, _30786, _30787, _30788,
         _30789, _30790, _30791, _30792, _30793, _30794, _30795, _30796,
         _30797, _30798, _30799, _30800, _30801, _30802, _30803, _30804,
         _30805, _30806, _30807, _30808, _30809, _30810, _30811, _30812,
         _30813, _30814, _30815, _30816, _30817, _30818, _30819, _30820,
         _30821, _30822, _30823, _30824, _30825, _30826, _30827, _30828,
         _30829, _30830, _30831, _30832, _30833, _30834, _30835, _30836,
         _30837, _30838, _30839, _30840, _30841, _30842, _30843, _30844,
         _30845, _30846, _30847, _30848, _30849, _30850, _30851, _30852,
         _30853, _30854, _30855, _30856, _30857, _30858, _30859, _30860,
         _30861, _30862, _30863, _30864, _30865, _30866, _30867, _30868,
         _30869, _30870, _30871, _30872, _30873, _30874, _30875, _30876,
         _30877, _30878, _30879, _30880, _30881, _30882, _30883, _30884,
         _30885, _30886, _30887, _30888, _30889, _30890, _30891, _30892,
         _30893, _30894, _30895, _30896, _30897, _30898, _30899, _30900,
         _30901, _30902, _30903, _30904, _30905, _30906, _30907, _30908,
         _30909, _30910, _30911, _30912, _30913, _30914, _30915, _30916,
         _30917, _30918, _30919, _30920, _30921, _30922, _30923, _30924,
         _30925, _30926, _30927, _30928, _30929, _30930, _30931, _30932,
         _30933, _30934, _30935, _30936, _30937, _30938, _30939, _30940,
         _30941, _30942, _30943, _30944, _30945, _30946, _30947, _30948,
         _30949, _30950, _30951, _30952, _30953, _30954, _30955, _30956,
         _30957, _30958, _30959, _30960, _30961, _30962, _30963, _30964,
         _30965, _30966, _30967, _30968, _30969, _30970, _30971, _30972,
         _30973, _30974, _30975, _30976, _30977, _30978, _30979, _30980,
         _30981, _30982, _30983, _30984, _30985, _30986, _30987, _30988,
         _30989, _30990, _30991, _30992, _30993, _30994, _30995, _30996,
         _30997, _30998, _30999, _31000, _31001, _31002, _31003, _31004,
         _31005, _31006, _31007, _31008, _31009, _31010, _31011, _31012,
         _31013, _31014, _31015, _31016, _31017, _31018, _31019, _31020,
         _31021, _31022, _31023, _31024, _31025, _31026, _31027, _31028,
         _31029, _31030, _31031, _31032, _31033, _31034, _31035, _31036,
         _31037, _31038, _31039, _31040, _31041, _31042, _31043, _31044,
         _31045, _31046, _31047, _31048, _31049, _31050, _31051, _31052,
         _31053, _31054, _31055, _31056, _31057, _31058, _31059, _31060,
         _31061, _31062, _31063, _31064, _31065, _31066, _31067, _31068,
         _31069, _31070, _31071, _31072, _31073, _31074, _31075, _31076,
         _31077, _31078, _31079, _31080, _31081, _31082, _31083, _31084,
         _31085, _31086, _31087, _31088, _31089, _31090, _31091, _31092,
         _31093, _31094, _31095, _31096, _31097, _31098, _31099, _31100,
         _31101, _31102, _31103, _31104, _31105, _31106, _31107, _31108,
         _31109, _31110, _31111, _31112, _31113, _31114, _31115, _31116,
         _31117, _31118, _31119, _31120, _31121, _31122, _31123, _31124,
         _31125, _31126, _31127, _31128, _31129, _31130, _31131, _31132,
         _31133, _31134, _31135, _31136, _31137, _31138, _31139, _31140,
         _31141, _31142, _31143, _31144, _31145, _31146, _31147, _31148,
         _31149, _31150, _31151, _31152, _31153, _31154, _31155, _31156,
         _31157, _31158, _31159, _31160, _31161, _31162, _31163, _31164,
         _31165, _31166, _31167, _31168, _31169, _31170, _31171, _31172,
         _31173, _31174, _31175, _31176, _31177, _31178, _31179, _31180,
         _31181, _31182, _31183, _31184, _31185, _31186, _31187, _31188,
         _31189, _31190, _31191, _31192, _31193, _31194, _31195, _31196,
         _31197, _31198, _31199, _31200, _31201, _31202, _31203, _31204,
         _31205, _31206, _31207, _31208, _31209, _31210, _31211, _31212,
         _31213, _31214, _31215, _31216, _31217, _31218, _31219, _31220,
         _31221, _31222, _31223, _31224, _31225, _31226, _31227, _31228,
         _31229, _31230, _31231, _31232, _31233, _31234, _31235, _31236,
         _31237, _31238, _31239, _31240, _31241, _31242, _31243, _31244,
         _31245, _31246, _31247, _31248, _31249, _31250, _31251, _31252,
         _31253, _31254, _31255, _31256, _31257, _31258, _31259, _31260,
         _31261, _31262, _31263, _31264, _31265, _31266, _31267, _31268,
         _31269, _31270, _31271, _31272, _31273, _31274, _31275, _31276,
         _31277, _31278, _31279, _31280, _31281, _31282, _31283, _31284,
         _31285, _31286, _31287, _31288, _31289, _31290, _31291, _31292,
         _31293, _31294, _31295, _31296, _31297, _31298, _31299, _31300,
         _31301, _31302, _31303, _31304, _31305, _31306, _31307, _31308,
         _31309, _31310, _31311, _31312, _31313, _31314, _31315, _31316,
         _31317, _31318, _31319, _31320, _31321, _31322, _31323, _31324,
         _31325, _31326, _31327, _31328, _31329, _31330, _31331, _31332,
         _31333, _31334, _31335, _31336, _31337, _31338, _31339, _31340,
         _31341, _31342, _31343, _31344, _31345, _31346, _31347, _31348,
         _31349, _31350, _31351, _31352, _31353, _31354, _31355, _31356,
         _31357, _31358, _31359, _31360, _31361, _31362, _31363, _31364,
         _31365, _31366, _31367, _31368, _31369, _31370, _31371, _31372,
         _31373, _31374, _31375, _31376, _31377, _31378, _31379, _31380,
         _31381, _31382, _31383, _31384, _31385, _31386, _31387, _31388,
         _31389, _31390, _31391, _31392, _31393, _31394, _31395, _31396,
         _31397, _31398, _31399, _31400, _31401, _31402, _31403, _31404,
         _31405, _31406, _31407, _31408, _31409, _31410, _31411, _31412,
         _31413, _31414, _31415, _31416, _31417, _31418, _31419, _31420,
         _31421, _31422, _31423, _31424, _31425, _31426, _31427, _31428,
         _31429, _31430, _31431, _31432, _31433, _31434, _31435, _31436,
         _31437, _31438, _31439, _31440, _31441, _31442, _31443, _31444,
         _31445, _31446, _31447, _31448, _31449, _31450, _31451, _31452,
         _31453, _31454, _31455, _31456, _31457, _31458, _31459, _31460,
         _31461, _31462, _31463, _31464, _31465, _31466, _31467, _31468,
         _31469, _31470, _31471, _31472, _31473, _31474, _31475, _31476,
         _31477, _31478, _31479, _31480, _31481, _31482, _31483, _31484,
         _31485, _31486, _31487, _31488, _31489, _31490, _31491, _31492,
         _31493, _31494, _31495, _31496, _31497, _31498, _31499, _31500,
         _31501, _31502, _31503, _31504, _31505, _31506, _31507, _31508,
         _31509, _31510, _31511, _31512, _31513, _31514, _31515, _31516,
         _31517, _31518, _31519, _31520, _31521, _31522, _31523, _31524,
         _31525, _31526, _31527, _31528, _31529, _31530, _31531, _31532,
         _31533, _31534, _31535, _31536, _31537, _31538, _31539, _31540,
         _31541, _31542, _31543, _31544, _31545, _31546, _31547, _31548,
         _31549, _31550, _31551, _31552, _31553, _31554, _31555, _31556,
         _31557, _31558, _31559, _31560, _31561, _31562, _31563, _31564,
         _31565, _31566, _31567, _31568, _31569, _31570, _31571, _31572,
         _31573, _31574, _31575, _31576, _31577, _31578, _31579, _31580,
         _31581, _31582, _31583, _31584, _31585, _31586, _31587, _31588,
         _31589, _31590, _31591, _31592, _31593, _31594, _31595, _31596,
         _31597, _31598, _31599, _31600, _31601, _31602, _31603, _31604,
         _31605, _31606, _31607, _31608, _31609, _31610, _31611, _31612,
         _31613, _31614, _31615, _31616, _31617, _31618, _31619, _31620,
         _31621, _31622, _31623, _31624, _31625, _31626, _31627, _31628,
         _31629, _31630, _31631, _31632, _31633, _31634, _31635, _31636,
         _31637, _31638, _31639, _31640, _31641, _31642, _31643, _31644,
         _31645, _31646, _31647, _31648, _31649, _31650, _31651, _31652,
         _31653, _31654, _31655, _31656, _31657, _31658, _31659, _31660,
         _31661, _31662, _31663, _31664, _31665, _31666, _31667, _31668,
         _31669, _31670, _31671, _31672, _31673, _31674, _31675, _31676,
         _31677, _31678, _31679, _31680, _31681, _31682, _31683, _31684,
         _31685, _31686, _31687, _31688, _31689, _31690, _31691, _31692,
         _31693, _31694, _31695, _31696, _31697, _31698, _31699, _31700,
         _31701, _31702, _31703, _31704, _31705, _31706, _31707, _31708,
         _31709, _31710, _31711, _31712, _31713, _31714, _31715, _31716,
         _31717, _31718, _31719, _31720, _31721, _31722, _31723, _31724,
         _31725, _31726, _31727, _31728, _31729, _31730, _31731, _31732,
         _31733, _31734, _31735, _31736, _31737, _31738, _31739, _31740,
         _31741, _31742, _31743, _31744, _31745, _31746, _31747, _31748,
         _31749, _31750, _31751, _31752, _31753, _31754, _31755, _31756,
         _31757, _31758, _31759, _31760, _31761, _31762, _31763, _31764,
         _31765, _31766, _31767, _31768, _31769, _31770, _31771, _31772,
         _31773, _31774, _31775, _31776, _31777, _31778, _31779, _31780,
         _31781, _31782, _31783, _31784, _31785, _31786, _31787, _31788,
         _31789, _31790, _31791, _31792, _31793, _31794, _31795, _31796,
         _31797, _31798, _31799, _31800, _31801, _31802, _31803, _31804,
         _31805, _31806, _31807, _31808, _31809, _31810, _31811, _31812,
         _31813, _31814, _31815, _31816, _31817, _31818, _31819, _31820,
         _31821, _31822, _31823, _31824, _31825, _31826, _31827, _31828,
         _31829, _31830, _31831, _31832, _31833, _31834, _31835, _31836,
         _31837, _31838, _31839, _31840, _31841, _31842, _31843, _31844,
         _31845, _31846, _31847, _31848, _31849, _31850, _31851, _31852,
         _31853, _31854, _31855, _31856, _31857, _31858, _31859, _31860,
         _31861, _31862, _31863, _31864, _31865, _31866, _31867, _31868,
         _31869, _31870, _31871, _31872, _31873, _31874, _31875, _31876,
         _31877, _31878, _31879, _31880, _31881, _31882, _31883, _31884,
         _31885, _31886, _31887, _31888, _31889, _31890, _31891, _31892,
         _31893, _31894, _31895, _31896, _31897, _31898, _31899, _31900,
         _31901, _31902, _31903, _31904, _31905, _31906, _31907, _31908,
         _31909, _31910, _31911, _31912, _31913, _31914, _31915, _31916,
         _31917, _31918, _31919, _31920, _31921, _31922, _31923, _31924,
         _31925, _31926, _31927, _31928, _31929, _31930, _31931, _31932,
         _31933, _31934, _31935, _31936, _31937, _31938, _31939, _31940,
         _31941, _31942, _31943, _31944, _31945, _31946, _31947, _31948,
         _31949, _31950, _31951, _31952, _31953, _31954, _31955, _31956,
         _31957, _31958, _31959, _31960, _31961, _31962, _31963, _31964,
         _31965, _31966, _31967, _31968, _31969, _31970, _31971, _31972,
         _31973, _31974, _31975, _31976, _31977, _31978, _31979, _31980,
         _31981, _31982, _31983, _31984, _31985, _31986, _31987, _31988,
         _31989, _31990, _31991, _31992, _31993, _31994, _31995, _31996,
         _31997, _31998, _31999, _32000, _32001, _32002, _32003, _32004,
         _32005, _32006, _32007, _32008, _32009, _32010, _32011, _32012,
         _32013, _32014, _32015, _32016, _32017, _32018, _32019, _32020,
         _32021, _32022, _32023, _32024, _32025, _32026, _32027, _32028,
         _32029, _32030, _32031, _32032, _32033, _32034, _32035, _32036,
         _32037, _32038, _32039, _32040, _32041, _32042, _32043, _32044,
         _32045, _32046, _32047, _32048, _32049, _32050, _32051, _32052,
         _32053, _32054, _32055, _32056, _32057, _32058, _32059, _32060,
         _32061, _32062, _32063, _32064, _32065, _32066, _32067, _32068,
         _32069, _32070, _32071, _32072, _32073, _32074, _32075, _32076,
         _32077, _32078, _32079, _32080, _32081, _32082, _32083, _32084,
         _32085, _32086, _32087, _32088, _32089, _32090, _32091, _32092,
         _32093, _32094, _32095, _32096, _32097, _32098, _32099, _32100,
         _32101, _32102, _32103, _32104, _32105, _32106, _32107, _32108,
         _32109, _32110, _32111, _32112, _32113, _32114, _32115, _32116,
         _32117, _32118, _32119, _32120, _32121, _32122, _32123, _32124,
         _32125, _32126, _32127, _32128, _32129, _32130, _32131, _32132,
         _32133, _32134, _32135, _32136, _32137, _32138, _32139, _32140,
         _32141, _32142, _32143, _32144, _32145, _32146, _32147, _32148,
         _32149, _32150, _32151, _32152, _32153, _32154, _32155, _32156,
         _32157, _32158, _32159, _32160, _32161, _32162, _32163, _32164,
         _32165, _32166, _32167, _32168, _32169, _32170, _32171, _32172,
         _32173, _32174, _32175, _32176, _32177, _32178, _32179, _32180,
         _32181, _32182, _32183, _32184, _32185, _32186, _32187, _32188,
         _32189, _32190, _32191, _32192, _32193, _32194, _32195, _32196,
         _32197, _32198, _32199, _32200, _32201, _32202, _32203, _32204,
         _32205, _32206, _32207, _32208, _32209, _32210, _32211, _32212,
         _32213, _32214, _32215, _32216, _32217, _32218, _32219, _32220,
         _32221, _32222, _32223, _32224, _32225, _32226, _32227, _32228,
         _32229, _32230, _32231, _32232, _32233, _32234, _32235, _32236,
         _32237, _32238, _32239, _32240, _32241, _32242, _32243, _32244,
         _32245, _32246, _32247, _32248, _32249, _32250, _32251, _32252,
         _32253, _32254, _32255, _32256, _32257, _32258, _32259, _32260,
         _32261, _32262, _32263, _32264, _32265, _32266, _32267, _32268,
         _32269, _32270, _32271, _32272, _32273, _32274, _32275, _32276,
         _32277, _32278, _32279, _32280, _32281, _32282, _32283, _32284,
         _32285, _32286, _32287, _32288, _32289, _32290, _32291, _32292,
         _32293, _32294, _32295, _32296, _32297, _32298, _32299, _32300,
         _32301, _32302, _32303, _32304, _32305, _32306, _32307, _32308,
         _32309, _32310, _32311, _32312, _32313, _32314, _32315, _32316,
         _32317, _32318, _32319, _32320, _32321, _32322, _32323, _32324,
         _32325, _32326, _32327, _32328, _32329, _32330, _32331, _32332,
         _32333, _32334, _32335, _32336, _32337, _32338, _32339, _32340,
         _32341, _32342, _32343, _32344, _32345, _32346, _32347, _32348,
         _32349, _32350, _32351, _32352, _32353, _32354, _32355, _32356,
         _32357, _32358, _32359, _32360, _32361, _32362, _32363, _32364,
         _32365, _32366, _32367, _32368, _32369, _32370, _32371, _32372,
         _32373, _32374, _32375, _32376, _32377, _32378, _32379, _32380,
         _32381, _32382, _32383, _32384, _32385, _32386, _32387, _32388,
         _32389, _32390, _32391, _32392, _32393, _32394, _32395, _32396,
         _32397, _32398, _32399, _32400, _32401, _32402, _32403, _32404,
         _32405, _32406, _32407, _32408, _32409, _32410, _32411, _32412,
         _32413, _32414, _32415, _32416, _32417, _32418, _32419, _32420,
         _32421, _32422, _32423, _32424, _32425, _32426, _32427, _32428,
         _32429, _32430, _32431, _32432, _32433, _32434, _32435, _32436,
         _32437, _32438, _32439, _32440, _32441, _32442, _32443, _32444,
         _32445, _32446, _32447, _32448, _32449, _32450, _32451, _32452,
         _32453, _32454, _32455, _32456, _32457, _32458, _32459, _32460,
         _32461, _32462, _32463, _32464, _32465, _32466, _32467, _32468,
         _32469, _32470, _32471, _32472, _32473, _32474, _32475, _32476,
         _32477, _32478, _32479, _32480, _32481, _32482, _32483, _32484,
         _32485, _32486, _32487, _32488, _32489, _32490, _32491, _32492,
         _32493, _32494, _32495, _32496, _32497, _32498, _32499, _32500,
         _32501, _32502, _32503, _32504, _32505, _32506, _32507, _32508,
         _32509, _32510, _32511, _32512, _32513, _32514, _32515, _32516,
         _32517, _32518, _32519, _32520, _32521, _32522, _32523, _32524,
         _32525, _32526, _32527, _32528, _32529, _32530, _32531, _32532,
         _32533, _32534, _32535, _32536, _32537, _32538, _32539, _32540,
         _32541, _32542, _32543, _32544, _32545, _32546, _32547, _32548,
         _32549, _32550, _32551, _32552, _32553, _32554, _32555, _32556,
         _32557, _32558, _32559, _32560, _32561, _32562, _32563, _32564,
         _32565, _32566, _32567, _32568, _32569, _32570, _32571, _32572,
         _32573, _32574, _32575, _32576, _32577, _32578, _32579, _32580,
         _32581, _32582, _32583, _32584, _32585, _32586, _32587, _32588,
         _32589, _32590, _32591, _32592, _32593, _32594, _32595, _32596,
         _32597, _32598, _32599, _32600, _32601, _32602, _32603, _32604,
         _32605, _32606, _32607, _32608, _32609, _32610, _32611, _32612,
         _32613, _32614, _32615, _32616, _32617, _32618, _32619, _32620,
         _32621, _32622, _32623, _32624, _32625, _32626, _32627, _32628,
         _32629, _32630, _32631, _32632, _32633, _32634, _32635, _32636,
         _32637, _32638, _32639, _32640, _32641, _32642, _32643, _32644,
         _32645, _32646, _32647, _32648, _32649, _32650, _32651, _32652,
         _32653, _32654, _32655, _32656, _32657, _32658, _32659, _32660,
         _32661, _32662, _32663, _32664, _32665, _32666, _32667, _32668,
         _32669, _32670, _32671, _32672, _32673, _32674, _32675, _32676,
         _32677, _32678, _32679, _32680, _32681, _32682, _32683, _32684,
         _32685, _32686, _32687, _32688, _32689, _32690, _32691, _32692,
         _32693, _32694, _32695, _32696, _32697, _32698, _32699, _32700,
         _32701, _32702, _32703, _32704, _32705, _32706, _32707, _32708,
         _32709, _32710, _32711, _32712, _32713, _32714, _32715, _32716,
         _32717, _32718, _32719, _32720, _32721, _32722, _32723, _32724,
         _32725, _32726, _32727, _32728, _32729, _32730, _32731, _32732,
         _32733, _32734, _32735, _32736, _32737, _32738, _32739, _32740,
         _32741, _32742, _32743, _32744, _32745, _32746, _32747, _32748,
         _32749, _32750, _32751, _32752, _32753, _32754, _32755, _32756,
         _32757, _32758, _32759, _32760, _32761, _32762, _32763, _32764,
         _32765, _32766, _32767, _32768, _32769, _32770, _32771, _32772,
         _32773, _32774, _32775, _32776, _32777, _32778, _32779, _32780,
         _32781, _32782, _32783, _32784, _32785, _32786, _32787, _32788,
         _32789, _32790, _32791, _32792, _32793, _32794, _32795, _32796,
         _32797, _32798, _32799, _32800, _32801, _32802, _32803, _32804,
         _32805, _32806, _32807, _32808, _32809, _32810, _32811, _32812,
         _32813, _32814, _32815, _32816, _32817, _32818, _32819, _32820,
         _32821, _32822, _32823, _32824, _32825, _32826, _32827, _32828,
         _32829, _32830, _32831, _32832, _32833, _32834, _32835, _32836,
         _32837, _32838, _32839, _32840, _32841, _32842, _32843, _32844,
         _32845, _32846, _32847, _32848, _32849, _32850, _32851, _32852,
         _32853, _32854, _32855, _32856, _32857, _32858, _32859, _32860,
         _32861, _32862, _32863, _32864, _32865, _32866, _32867, _32868,
         _32869, _32870, _32871, _32872, _32873, _32874, _32875, _32876,
         _32877, _32878, _32879, _32880, _32881, _32882, _32883, _32884,
         _32885, _32886, _32887, _32888, _32889, _32890, _32891, _32892,
         _32893, _32894, _32895, _32896, _32897, _32898, _32899, _32900,
         _32901, _32902, _32903, _32904, _32905, _32906, _32907, _32908,
         _32909, _32910, _32911, _32912, _32913, _32914, _32915, _32916,
         _32917, _32918, _32919, _32920, _32921, _32922, _32923, _32924,
         _32925, _32926, _32927, _32928, _32929, _32930, _32931, _32932,
         _32933, _32934, _32935, _32936, _32937, _32938, _32939, _32940,
         _32941, _32942, _32943, _32944, _32945, _32946, _32947, _32948,
         _32949, _32950, _32951, _32952, _32953, _32954, _32955, _32956,
         _32957, _32958, _32959, _32960, _32961, _32962, _32963, _32964,
         _32965, _32966, _32967, _32968, _32969, _32970, _32971, _32972,
         _32973, _32974, _32975, _32976, _32977, _32978, _32979, _32980,
         _32981, _32982, _32983, _32984, _32985, _32986, _32987, _32988,
         _32989, _32990, _32991, _32992, _32993, _32994, _32995, _32996,
         _32997, _32998, _32999, _33000, _33001, _33002, _33003, _33004,
         _33005, _33006, _33007, _33008, _33009, _33010, _33011, _33012,
         _33013, _33014, _33015, _33016, _33017, _33018, _33019, _33020,
         _33021, _33022, _33023, _33024, _33025, _33026, _33027, _33028,
         _33029, _33030, _33031, _33032, _33033, _33034, _33035, _33036,
         _33037, _33038, _33039, _33040, _33041, _33042, _33043, _33044,
         _33045, _33046, _33047, _33048, _33049, _33050, _33051, _33052,
         _33053, _33054, _33055, _33056, _33057, _33058, _33059, _33060,
         _33061, _33062, _33063, _33064, _33065, _33066, _33067, _33068,
         _33069, _33070, _33071, _33072, _33073, _33074, _33075, _33076,
         _33077, _33078, _33079, _33080, _33081, _33082, _33083, _33084,
         _33085, _33086, _33087, _33088, _33089, _33090, _33091, _33092,
         _33093, _33094, _33095, _33096, _33097, _33098, _33099, _33100,
         _33101, _33102, _33103, _33104, _33105, _33106, _33107, _33108,
         _33109, _33110, _33111, _33112, _33113, _33114, _33115, _33116,
         _33117, _33118, _33119, _33120, _33121, _33122, _33123, _33124,
         _33125, _33126, _33127, _33128, _33129, _33130, _33131, _33132,
         _33133, _33134, _33135, _33136, _33137, _33138, _33139, _33140,
         _33141, _33142, _33143, _33144, _33145, _33146, _33147, _33148,
         _33149, _33150, _33151, _33152, _33153, _33154, _33155, _33156,
         _33157, _33158, _33159, _33160, _33161, _33162, _33163, _33164,
         _33165, _33166, _33167, _33168, _33169, _33170, _33171, _33172,
         _33173, _33174, _33175, _33176, _33177, _33178, _33179, _33180,
         _33181, _33182, _33183, _33184, _33185, _33186, _33187, _33188,
         _33189, _33190, _33191, _33192, _33193, _33194, _33195, _33196,
         _33197, _33198, _33199, _33200, _33201, _33202, _33203, _33204,
         _33205, _33206, _33207, _33208, _33209, _33210, _33211, _33212,
         _33213, _33214, _33215, _33216, _33217, _33218, _33219, _33220,
         _33221, _33222, _33223, _33224, _33225, _33226, _33227, _33228,
         _33229, _33230, _33231, _33232, _33233, _33234, _33235, _33236,
         _33237, _33238, _33239, _33240, _33241, _33242, _33243, _33244,
         _33245, _33246, _33247, _33248, _33249, _33250, _33251, _33252,
         _33253, _33254, _33255, _33256, _33257, _33258, _33259, _33260,
         _33261, _33262, _33263, _33264, _33265, _33266, _33267, _33268,
         _33269, _33270, _33271, _33272, _33273, _33274, _33275, _33276,
         _33277, _33278, _33279, _33280, _33281, _33282, _33283, _33284,
         _33285, _33286, _33287, _33288, _33289, _33290, _33291, _33292,
         _33293, _33294, _33295, _33296, _33297, _33298, _33299, _33300,
         _33301, _33302, _33303, _33304, _33305, _33306, _33307, _33308,
         _33309, _33310, _33311, _33312, _33313, _33314, _33315, _33316,
         _33317, _33318, _33319, _33320, _33321, _33322, _33323, _33324,
         _33325, _33326, _33327, _33328, _33329, _33330, _33331, _33332,
         _33333, _33334, _33335, _33336, _33337, _33338, _33339, _33340,
         _33341, _33342, _33343, _33344, _33345, _33346, _33347, _33348,
         _33349, _33350, _33351, _33352, _33353, _33354, _33355, _33356,
         _33357, _33358, _33359, _33360, _33361, _33362, _33363, _33364,
         _33365, _33366, _33367, _33368, _33369, _33370, _33371, _33372,
         _33373, _33374, _33375, _33376, _33377, _33378, _33379, _33380,
         _33381, _33382, _33383, _33384, _33385, _33386, _33387, _33388,
         _33389, _33390, _33391, _33392, _33393, _33394, _33395, _33396,
         _33397, _33398, _33399, _33400, _33401, _33402, _33403, _33404,
         _33405, _33406, _33407, _33408, _33409, _33410, _33411, _33412,
         _33413, _33414, _33415, _33416, _33417, _33418, _33419, _33420,
         _33421, _33422, _33423, _33424, _33425, _33426, _33427, _33428,
         _33429, _33430, _33431, _33432, _33433, _33434, _33435, _33436,
         _33437, _33438, _33439, _33440, _33441, _33442, _33443, _33444,
         _33445, _33446, _33447, _33448, _33449, _33450, _33451, _33452,
         _33453, _33454, _33455, _33456, _33457, _33458, _33459, _33460,
         _33461, _33462, _33463, _33464, _33465, _33466, _33467, _33468,
         _33469, _33470, _33471, _33472, _33473, _33474, _33475, _33476,
         _33477, _33478, _33479, _33480, _33481, _33482, _33483, _33484,
         _33485, _33486, _33487, _33488, _33489, _33490, _33491, _33492,
         _33493, _33494, _33495, _33496, _33497, _33498, _33499, _33500,
         _33501, _33502, _33503, _33504, _33505, _33506, _33507, _33508,
         _33509, _33510, _33511, _33512, _33513, _33514, _33515, _33516,
         _33517, _33518, _33519, _33520, _33521, _33522, _33523, _33524,
         _33525, _33526, _33527, _33528, _33529, _33530, _33531, _33532,
         _33533, _33534, _33535, _33536, _33537, _33538, _33539, _33540,
         _33541, _33542, _33543, _33544, _33545, _33546, _33547, _33548,
         _33549, _33550, _33551, _33552, _33553, _33554, _33555, _33556,
         _33557, _33558, _33559, _33560, _33561, _33562, _33563, _33564,
         _33565, _33566, _33567, _33568, _33569, _33570, _33571, _33572,
         _33573, _33574, _33575, _33576, _33577, _33578, _33579, _33580,
         _33581, _33582, _33583, _33584, _33585, _33586, _33587, _33588,
         _33589, _33590, _33591, _33592, _33593, _33594, _33595, _33596,
         _33597, _33598, _33599, _33600, _33601, _33602, _33603, _33604,
         _33605, _33606, _33607, _33608, _33609, _33610, _33611, _33612,
         _33613, _33614, _33615, _33616, _33617, _33618, _33619, _33620,
         _33621, _33622, _33623, _33624, _33625, _33626, _33627, _33628,
         _33629, _33630, _33631, _33632, _33633, _33634, _33635, _33636,
         _33637, _33638, _33639, _33640, _33641, _33642, _33643, _33644,
         _33645, _33646, _33647, _33648, _33649, _33650, _33651, _33652,
         _33653, _33654, _33655, _33656, _33657, _33658, _33659, _33660,
         _33661, _33662, _33663, _33664, _33665, _33666, _33667, _33668,
         _33669, _33670, _33671, _33672, _33673, _33674, _33675, _33676,
         _33677, _33678, _33679, _33680, _33681, _33682, _33683, _33684,
         _33685, _33686, _33687, _33688, _33689, _33690, _33691, _33692,
         _33693, _33694, _33695, _33696, _33697, _33698, _33699, _33700,
         _33701, _33702, _33703, _33704, _33705, _33706, _33707, _33708,
         _33709, _33710, _33711, _33712, _33713, _33714, _33715, _33716,
         _33717, _33718, _33719, _33720, _33721, _33722, _33723, _33724,
         _33725, _33726, _33727, _33728, _33729, _33730, _33731, _33732,
         _33733, _33734, _33735, _33736, _33737, _33738, _33739, _33740,
         _33741, _33742, _33743, _33744, _33745, _33746, _33747, _33748,
         _33749, _33750, _33751, _33752, _33753, _33754, _33755, _33756,
         _33757, _33758, _33759, _33760, _33761, _33762, _33763, _33764,
         _33765, _33766, _33767, _33768, _33769, _33770, _33771, _33772,
         _33773, _33774, _33775, _33776, _33777, _33778, _33779, _33780,
         _33781, _33782, _33783, _33784, _33785, _33786, _33787, _33788,
         _33789, _33790, _33791, _33792, _33793, _33794, _33795, _33796,
         _33797, _33798, _33799, _33800, _33801, _33802, _33803, _33804,
         _33805, _33806, _33807, _33808, _33809, _33810, _33811, _33812,
         _33813, _33814, _33815, _33816, _33817, _33818, _33819, _33820,
         _33821, _33822, _33823, _33824, _33825, _33826, _33827, _33828,
         _33829, _33830, _33831, _33832, _33833, _33834, _33835, _33836,
         _33837, _33838, _33839, _33840, _33841, _33842, _33843, _33844,
         _33845, _33846, _33847, _33848, _33849, _33850, _33851, _33852,
         _33853, _33854, _33855, _33856, _33857, _33858, _33859, _33860,
         _33861, _33862, _33863, _33864, _33865, _33866, _33867, _33868,
         _33869, _33870, _33871, _33872, _33873, _33874, _33875, _33876,
         _33877, _33878, _33879, _33880, _33881, _33882, _33883, _33884,
         _33885, _33886, _33887, _33888, _33889, _33890, _33891, _33892,
         _33893, _33894, _33895, _33896, _33897, _33898, _33899, _33900,
         _33901, _33902, _33903, _33904, _33905, _33906, _33907, _33908,
         _33909, _33910, _33911, _33912, _33913, _33914, _33915, _33916,
         _33917, _33918, _33919, _33920, _33921, _33922, _33923, _33924,
         _33925, _33926, _33927, _33928, _33929, _33930, _33931, _33932,
         _33933, _33934, _33935, _33936, _33937, _33938, _33939, _33940,
         _33941, _33942, _33943, _33944, _33945, _33946, _33947, _33948,
         _33949, _33950, _33951, _33952, _33953, _33954, _33955, _33956,
         _33957, _33958, _33959, _33960, _33961, _33962, _33963, _33964,
         _33965, _33966, _33967, _33968, _33969, _33970, _33971, _33972,
         _33973, _33974, _33975, _33976, _33977, _33978, _33979, _33980,
         _33981, _33982, _33983, _33984, _33985, _33986, _33987, _33988,
         _33989, _33990, _33991, _33992, _33993, _33994, _33995, _33996,
         _33997, _33998, _33999, _34000, _34001, _34002, _34003, _34004,
         _34005, _34006, _34007, _34008, _34009, _34010, _34011, _34012,
         _34013, _34014, _34015, _34016, _34017, _34018, _34019, _34020,
         _34021, _34022, _34023, _34024, _34025, _34026, _34027, _34028,
         _34029, _34030, _34031, _34032, _34033, _34034, _34035, _34036,
         _34037, _34038, _34039, _34040, _34041, _34042, _34043, _34044,
         _34045, _34046, _34047, _34048, _34049, _34050, _34051, _34052,
         _34053, _34054, _34055, _34056, _34057, _34058, _34059, _34060,
         _34061, _34062, _34063, _34064, _34065, _34066, _34067, _34068,
         _34069, _34070, _34071, _34072, _34073, _34074, _34075, _34076,
         _34077, _34078, _34079, _34080, _34081, _34082, _34083, _34084,
         _34085, _34086, _34087, _34088, _34089, _34090, _34091, _34092,
         _34093, _34094, _34095, _34096, _34097, _34098, _34099, _34100,
         _34101, _34102, _34103, _34104, _34105, _34106, _34107, _34108,
         _34109, _34110, _34111, _34112, _34113, _34114, _34115, _34116,
         _34117, _34118, _34119, _34120, _34121, _34122, _34123, _34124,
         _34125, _34126, _34127, _34128, _34129, _34130, _34131, _34132,
         _34133, _34134, _34135, _34136, _34137, _34138, _34139, _34140,
         _34141, _34142, _34143, _34144, _34145, _34146, _34147, _34148,
         _34149, _34150, _34151, _34152, _34153, _34154, _34155, _34156,
         _34157, _34158, _34159, _34160, _34161, _34162, _34163, _34164,
         _34165, _34166, _34167, _34168, _34169, _34170, _34171, _34172,
         _34173, _34174, _34175, _34176, _34177, _34178, _34179, _34180,
         _34181, _34182, _34183, _34184, _34185, _34186, _34187, _34188,
         _34189, _34190, _34191, _34192, _34193, _34194, _34195, _34196,
         _34197, _34198, _34199, _34200, _34201, _34202, _34203, _34204,
         _34205, _34206, _34207, _34208, _34209, _34210, _34211, _34212,
         _34213, _34214, _34215, _34216, _34217, _34218, _34219, _34220,
         _34221, _34222, _34223, _34224, _34225, _34226, _34227, _34228,
         _34229, _34230, _34231, _34232, _34233, _34234, _34235, _34236,
         _34237, _34238, _34239, _34240, _34241, _34242, _34243, _34244,
         _34245, _34246, _34247, _34248, _34249, _34250, _34251, _34252,
         _34253, _34254, _34255, _34256, _34257, _34258, _34259, _34260,
         _34261, _34262, _34263, _34264, _34265, _34266, _34267, _34268,
         _34269, _34270, _34271, _34272, _34273, _34274, _34275, _34276,
         _34277, _34278, _34279, _34280, _34281, _34282, _34283, _34284,
         _34285, _34286, _34287, _34288, _34289, _34290, _34291, _34292,
         _34293, _34294, _34295, _34296, _34297, _34298, _34299, _34300,
         _34301, _34302, _34303, _34304, _34305, _34306, _34307, _34308,
         _34309, _34310, _34311, _34312, _34313, _34314, _34315, _34316,
         _34317, _34318, _34319, _34320, _34321, _34322, _34323, _34324,
         _34325, _34326, _34327, _34328, _34329, _34330, _34331, _34332,
         _34333, _34334, _34335, _34336, _34337, _34338, _34339, _34340,
         _34341, _34342, _34343, _34344, _34345, _34346, _34347, _34348,
         _34349, _34350, _34351, _34352, _34353, _34354, _34355, _34356,
         _34357, _34358, _34359, _34360, _34361, _34362, _34363, _34364,
         _34365, _34366, _34367, _34368, _34369, _34370, _34371, _34372,
         _34373, _34374, _34375, _34376, _34377, _34378, _34379, _34380,
         _34381, _34382, _34383, _34384, _34385, _34386, _34387, _34388,
         _34389, _34390, _34391, _34392, _34393, _34394, _34395, _34396,
         _34397, _34398, _34399, _34400, _34401, _34402, _34403, _34404,
         _34405, _34406, _34407, _34408, _34409, _34410, _34411, _34412,
         _34413, _34414, _34415, _34416, _34417, _34418, _34419, _34420,
         _34421, _34422, _34423, _34424, _34425, _34426, _34427, _34428,
         _34429, _34430, _34431, _34432, _34433, _34434, _34435, _34436,
         _34437, _34438, _34439, _34440, _34441, _34442, _34443, _34444,
         _34445, _34446, _34447, _34448, _34449, _34450, _34451, _34452,
         _34453, _34454, _34455, _34456, _34457, _34458, _34459, _34460,
         _34461, _34462, _34463, _34464, _34465, _34466, _34467, _34468,
         _34469, _34470, _34471, _34472, _34473, _34474, _34475, _34476,
         _34477, _34478, _34479, _34480, _34481, _34482, _34483, _34484,
         _34485, _34486, _34487, _34488, _34489, _34490, _34491, _34492,
         _34493, _34494, _34495, _34496, _34497, _34498, _34499, _34500,
         _34501, _34502, _34503, _34504, _34505, _34506, _34507, _34508,
         _34509, _34510, _34511, _34512, _34513, _34514, _34515, _34516,
         _34517, _34518, _34519, _34520, _34521, _34522, _34523, _34524,
         _34525, _34526, _34527, _34528, _34529, _34530, _34531, _34532,
         _34533, _34534, _34535, _34536, _34537, _34538, _34539, _34540,
         _34541, _34542, _34543, _34544, _34545, _34546, _34547, _34548,
         _34549, _34550, _34551, _34552, _34553, _34554, _34555, _34556,
         _34557, _34558, _34559, _34560, _34561, _34562, _34563, _34564,
         _34565, _34566, _34567, _34568, _34569, _34570, _34571, _34572,
         _34573, _34574, _34575, _34576, _34577, _34578, _34579, _34580,
         _34581, _34582, _34583, _34584, _34585, _34586, _34587, _34588,
         _34589, _34590, _34591, _34592, _34593, _34594, _34595, _34596,
         _34597, _34598, _34599, _34600, _34601, _34602, _34603, _34604,
         _34605, _34606, _34607, _34608, _34609, _34610, _34611, _34612,
         _34613, _34614, _34615, _34616, _34617, _34618, _34619, _34620,
         _34621, _34622, _34623, _34624, _34625, _34626, _34627, _34628,
         _34629, _34630, _34631, _34632, _34633, _34634, _34635, _34636,
         _34637, _34638, _34639, _34640, _34641, _34642, _34643, _34644,
         _34645, _34646, _34647, _34648, _34649, _34650, _34651, _34652,
         _34653, _34654, _34655, _34656, _34657, _34658, _34659, _34660,
         _34661, _34662, _34663, _34664, _34665, _34666, _34667, _34668,
         _34669, _34670, _34671, _34672, _34673, _34674, _34675, _34676,
         _34677, _34678, _34679, _34680, _34681, _34682, _34683, _34684,
         _34685, _34686, _34687, _34688, _34689, _34690, _34691, _34692,
         _34693, _34694, _34695, _34696, _34697, _34698, _34699, _34700,
         _34701, _34702, _34703, _34704, _34705, _34706, _34707, _34708,
         _34709, _34710, _34711, _34712, _34713, _34714, _34715, _34716,
         _34717, _34718, _34719, _34720, _34721, _34722, _34723, _34724,
         _34725, _34726, _34727, _34728, _34729, _34730, _34731, _34732,
         _34733, _34734, _34735, _34736, _34737, _34738, _34739, _34740,
         _34741, _34742, _34743, _34744, _34745, _34746, _34747, _34748,
         _34749, _34750, _34751, _34752, _34753, _34754, _34755, _34756,
         _34757, _34758, _34759, _34760, _34761, _34762, _34763, _34764,
         _34765, _34766, _34767, _34768, _34769, _34770, _34771, _34772,
         _34773, _34774, _34775, _34776, _34777, _34778, _34779, _34780,
         _34781, _34782, _34783, _34784, _34785, _34786, _34787, _34788,
         _34789, _34790, _34791, _34792, _34793, _34794, _34795, _34796,
         _34797, _34798, _34799, _34800, _34801, _34802, _34803, _34804,
         _34805, _34806, _34807, _34808, _34809, _34810, _34811, _34812,
         _34813, _34814, _34815, _34816, _34817, _34818, _34819, _34820,
         _34821, _34822, _34823, _34824, _34825, _34826, _34827, _34828,
         _34829, _34830, _34831, _34832, _34833, _34834, _34835, _34836,
         _34837, _34838, _34839, _34840, _34841, _34842, _34843, _34844,
         _34845, _34846, _34847, _34848, _34849, _34850, _34851, _34852,
         _34853, _34854, _34855, _34856, _34857, _34858, _34859, _34860,
         _34861, _34862, _34863, _34864, _34865, _34866, _34867, _34868,
         _34869, _34870, _34871, _34872, _34873, _34874, _34875, _34876,
         _34877, _34878, _34879, _34880, _34881, _34882, _34883, _34884,
         _34885, _34886, _34887, _34888, _34889, _34890, _34891, _34892,
         _34893, _34894, _34895, _34896, _34897, _34898, _34899, _34900,
         _34901, _34902, _34903, _34904, _34905, _34906, _34907, _34908,
         _34909, _34910, _34911, _34912, _34913, _34914, _34915, _34916,
         _34917, _34918, _34919, _34920, _34921, _34922, _34923, _34924,
         _34925, _34926, _34927, _34928, _34929, _34930, _34931, _34932,
         _34933, _34934, _34935, _34936, _34937, _34938, _34939, _34940,
         _34941, _34942, _34943, _34944, _34945, _34946, _34947, _34948,
         _34949, _34950, _34951, _34952, _34953, _34954, _34955, _34956,
         _34957, _34958, _34959, _34960, _34961, _34962, _34963, _34964,
         _34965, _34966, _34967, _34968, _34969, _34970, _34971, _34972,
         _34973, _34974, _34975, _34976, _34977, _34978, _34979, _34980,
         _34981, _34982, _34983, _34984, _34985, _34986, _34987, _34988,
         _34989, _34990, _34991, _34992, _34993, _34994, _34995, _34996,
         _34997, _34998, _34999, _35000, _35001, _35002, _35003, _35004,
         _35005, _35006, _35007, _35008, _35009, _35010, _35011, _35012,
         _35013, _35014, _35015, _35016, _35017, _35018, _35019, _35020,
         _35021, _35022, _35023, _35024, _35025, _35026, _35027, _35028,
         _35029, _35030, _35031, _35032, _35033, _35034, _35035, _35036,
         _35037, _35038, _35039, _35040, _35041, _35042, _35043, _35044,
         _35045, _35046, _35047, _35048, _35049, _35050, _35051, _35052,
         _35053, _35054, _35055, _35056, _35057, _35058, _35059, _35060,
         _35061, _35062, _35063, _35064, _35065, _35066, _35067, _35068,
         _35069, _35070, _35071, _35072, _35073, _35074, _35075, _35076,
         _35077, _35078, _35079, _35080, _35081, _35082, _35083, _35084,
         _35085, _35086, _35087, _35088, _35089, _35090, _35091, _35092,
         _35093, _35094, _35095, _35096, _35097, _35098, _35099, _35100,
         _35101, _35102, _35103, _35104, _35105, _35106, _35107, _35108,
         _35109, _35110, _35111, _35112, _35113, _35114, _35115, _35116,
         _35117, _35118, _35119, _35120, _35121, _35122, _35123, _35124,
         _35125, _35126, _35127, _35128, _35129, _35130, _35131, _35132,
         _35133, _35134, _35135, _35136, _35137, _35138, _35139, _35140,
         _35141, _35142, _35143, _35144, _35145, _35146, _35147, _35148,
         _35149, _35150, _35151, _35152, _35153, _35154, _35155, _35156,
         _35157, _35158, _35159, _35160, _35161, _35162, _35163, _35164,
         _35165, _35166, _35167, _35168, _35169, _35170, _35171, _35172,
         _35173, _35174, _35175, _35176, _35177, _35178, _35179, _35180,
         _35181, _35182, _35183, _35184, _35185, _35186, _35187, _35188,
         _35189, _35190, _35191, _35192, _35193, _35194, _35195, _35196,
         _35197, _35198, _35199, _35200, _35201, _35202, _35203, _35204,
         _35205, _35206, _35207, _35208, _35209, _35210, _35211, _35212,
         _35213, _35214, _35215, _35216, _35217, _35218, _35219, _35220,
         _35221, _35222, _35223, _35224, _35225, _35226, _35227, _35228,
         _35229, _35230, _35231, _35232, _35233, _35234, _35235, _35236,
         _35237, _35238, _35239, _35240, _35241, _35242, _35243, _35244,
         _35245, _35246, _35247, _35248, _35249, _35250, _35251, _35252,
         _35253, _35254, _35255, _35256, _35257, _35258, _35259, _35260,
         _35261, _35262, _35263, _35264, _35265, _35266, _35267, _35268,
         _35269, _35270, _35271, _35272, _35273, _35274, _35275, _35276,
         _35277, _35278, _35279, _35280, _35281, _35282, _35283, _35284,
         _35285, _35286, _35287, _35288, _35289, _35290, _35291, _35292,
         _35293, _35294, _35295, _35296, _35297, _35298, _35299, _35300,
         _35301, _35302, _35303, _35304, _35305, _35306, _35307, _35308,
         _35309, _35310, _35311, _35312, _35313, _35314, _35315, _35316,
         _35317, _35318, _35319, _35320, _35321, _35322, _35323, _35324,
         _35325, _35326, _35327, _35328, _35329, _35330, _35331, _35332,
         _35333, _35334, _35335, _35336, _35337, _35338, _35339, _35340,
         _35341, _35342, _35343, _35344, _35345, _35346, _35347, _35348,
         _35349, _35350, _35351, _35352, _35353, _35354, _35355, _35356,
         _35357, _35358, _35359, _35360, _35361, _35362, _35363, _35364,
         _35365, _35366, _35367, _35368, _35369, _35370, _35371, _35372,
         _35373, _35374, _35375, _35376, _35377, _35378, _35379, _35380,
         _35381, _35382, _35383, _35384, _35385, _35386, _35387, _35388,
         _35389, _35390, _35391, _35392, _35393, _35394, _35395, _35396,
         _35397, _35398, _35399, _35400, _35401, _35402, _35403, _35404,
         _35405, _35406, _35407, _35408, _35409, _35410, _35411, _35412,
         _35413, _35414, _35415, _35416, _35417, _35418, _35419, _35420,
         _35421, _35422, _35423, _35424, _35425, _35426, _35427, _35428,
         _35429, _35430, _35431, _35432, _35433, _35434, _35435, _35436,
         _35437, _35438, _35439, _35440, _35441, _35442, _35443, _35444,
         _35445, _35446, _35447, _35448, _35449, _35450, _35451, _35452,
         _35453, _35454, _35455, _35456, _35457, _35458, _35459, _35460,
         _35461, _35462, _35463, _35464, _35465, _35466, _35467, _35468,
         _35469, _35470, _35471, _35472, _35473, _35474, _35475, _35476,
         _35477, _35478, _35479, _35480, _35481, _35482, _35483, _35484,
         _35485, _35486, _35487, _35488, _35489, _35490, _35491, _35492,
         _35493, _35494, _35495, _35496, _35497, _35498, _35499, _35500,
         _35501, _35502, _35503, _35504, _35505, _35506, _35507, _35508,
         _35509, _35510, _35511, _35512, _35513, _35514, _35515, _35516,
         _35517, _35518, _35519, _35520, _35521, _35522, _35523, _35524,
         _35525, _35526, _35527, _35528, _35529, _35530, _35531, _35532,
         _35533, _35534, _35535, _35536, _35537, _35538, _35539, _35540,
         _35541, _35542, _35543, _35544, _35545, _35546, _35547, _35548,
         _35549, _35550, _35551, _35552, _35553, _35554, _35555, _35556,
         _35557, _35558, _35559, _35560, _35561, _35562, _35563, _35564,
         _35565, _35566, _35567, _35568, _35569, _35570, _35571, _35572,
         _35573, _35574, _35575, _35576, _35577, _35578, _35579, _35580,
         _35581, _35582, _35583, _35584, _35585, _35586, _35587, _35588,
         _35589, _35590, _35591, _35592, _35593, _35594, _35595, _35596,
         _35597, _35598, _35599, _35600, _35601, _35602, _35603, _35604,
         _35605, _35606, _35607, _35608, _35609, _35610, _35611, _35612,
         _35613, _35614, _35615, _35616, _35617, _35618, _35619, _35620,
         _35621, _35622, _35623, _35624, _35625, _35626, _35627, _35628,
         _35629, _35630, _35631, _35632, _35633, _35634, _35635, _35636,
         _35637, _35638, _35639, _35640, _35641, _35642, _35643, _35644,
         _35645, _35646, _35647, _35648, _35649, _35650, _35651, _35652,
         _35653, _35654, _35655, _35656, _35657, _35658, _35659, _35660,
         _35661, _35662, _35663, _35664, _35665, _35666, _35667, _35668,
         _35669, _35670, _35671, _35672, _35673, _35674, _35675, _35676,
         _35677, _35678, _35679, _35680, _35681, _35682, _35683, _35684,
         _35685, _35686, _35687, _35688, _35689, _35690, _35691, _35692,
         _35693, _35694, _35695, _35696, _35697, _35698, _35699, _35700,
         _35701, _35702, _35703, _35704, _35705, _35706, _35707, _35708,
         _35709, _35710, _35711, _35712, _35713, _35714, _35715, _35716,
         _35717, _35718, _35719, _35720, _35721, _35722, _35723, _35724,
         _35725, _35726, _35727, _35728, _35729, _35730, _35731, _35732,
         _35733, _35734, _35735, _35736, _35737, _35738, _35739, _35740,
         _35741, _35742, _35743, _35744, _35745, _35746, _35747, _35748,
         _35749, _35750, _35751, _35752, _35753, _35754, _35755, _35756,
         _35757, _35758, _35759, _35760, _35761, _35762, _35763, _35764,
         _35765, _35766, _35767, _35768, _35769, _35770, _35771, _35772,
         _35773, _35774, _35775, _35776, _35777, _35778, _35779, _35780,
         _35781, _35782, _35783, _35784, _35785, _35786, _35787, _35788,
         _35789, _35790, _35791, _35792, _35793, _35794, _35795, _35796,
         _35797, _35798, _35799, _35800, _35801, _35802, _35803, _35804,
         _35805, _35806, _35807, _35808, _35809, _35810, _35811, _35812,
         _35813, _35814, _35815, _35816, _35817, _35818, _35819, _35820,
         _35821, _35822, _35823, _35824, _35825, _35826, _35827, _35828,
         _35829, _35830, _35831, _35832, _35833, _35834, _35835, _35836,
         _35837, _35838, _35839, _35840, _35841, _35842, _35843, _35844,
         _35845, _35846, _35847, _35848, _35849, _35850, _35851, _35852,
         _35853, _35854, _35855, _35856, _35857, _35858, _35859, _35860,
         _35861, _35862, _35863, _35864, _35865, _35866, _35867, _35868,
         _35869, _35870, _35871, _35872, _35873, _35874, _35875, _35876,
         _35877, _35878, _35879, _35880, _35881, _35882, _35883, _35884,
         _35885, _35886, _35887, _35888, _35889, _35890, _35891, _35892,
         _35893, _35894, _35895, _35896, _35897, _35898, _35899, _35900,
         _35901, _35902, _35903, _35904, _35905, _35906, _35907, _35908,
         _35909, _35910, _35911, _35912, _35913, _35914, _35915, _35916,
         _35917, _35918, _35919, _35920, _35921, _35922, _35923, _35924,
         _35925, _35926, _35927, _35928, _35929, _35930, _35931, _35932,
         _35933, _35934, _35935, _35936, _35937, _35938, _35939, _35940,
         _35941, _35942, _35943, _35944, _35945, _35946, _35947, _35948,
         _35949, _35950, _35951, _35952, _35953, _35954, _35955, _35956,
         _35957, _35958, _35959, _35960, _35961, _35962, _35963, _35964,
         _35965, _35966, _35967, _35968, _35969, _35970, _35971, _35972,
         _35973, _35974, _35975, _35976, _35977, _35978, _35979, _35980,
         _35981, _35982, _35983, _35984, _35985, _35986, _35987, _35988,
         _35989, _35990, _35991, _35992, _35993, _35994, _35995, _35996,
         _35997, _35998, _35999, _36000, _36001, _36002, _36003, _36004,
         _36005, _36006, _36007, _36008, _36009, _36010, _36011, _36012,
         _36013, _36014, _36015, _36016, _36017, _36018, _36019, _36020,
         _36021, _36022, _36023, _36024, _36025, _36026, _36027, _36028,
         _36029, _36030, _36031, _36032, _36033, _36034, _36035, _36036,
         _36037, _36038, _36039, _36040, _36041, _36042, _36043, _36044,
         _36045, _36046, _36047, _36048, _36049, _36050, _36051, _36052,
         _36053, _36054, _36055, _36056, _36057, _36058, _36059, _36060,
         _36061, _36062, _36063, _36064, _36065, _36066, _36067, _36068,
         _36069, _36070, _36071, _36072, _36073, _36074, _36075, _36076,
         _36077, _36078, _36079, _36080, _36081, _36082, _36083, _36084,
         _36085, _36086, _36087, _36088, _36089, _36090, _36091, _36092,
         _36093, _36094, _36095, _36096, _36097, _36098, _36099, _36100,
         _36101, _36102, _36103, _36104, _36105, _36106, _36107, _36108,
         _36109, _36110, _36111, _36112, _36113, _36114, _36115, _36116,
         _36117, _36118, _36119, _36120, _36121, _36122, _36123, _36124,
         _36125, _36126, _36127, _36128, _36129, _36130, _36131, _36132,
         _36133, _36134, _36135, _36136, _36137, _36138, _36139, _36140,
         _36141, _36142, _36143, _36144, _36145, _36146, _36147, _36148,
         _36149, _36150, _36151, _36152, _36153, _36154, _36155, _36156,
         _36157, _36158, _36159, _36160, _36161, _36162, _36163, _36164,
         _36165, _36166, _36167, _36168, _36169, _36170, _36171, _36172,
         _36173, _36174, _36175, _36176, _36177, _36178, _36179, _36180,
         _36181, _36182, _36183, _36184, _36185, _36186, _36187, _36188,
         _36189, _36190, _36191, _36192, _36193, _36194, _36195, _36196,
         _36197, _36198, _36199, _36200, _36201, _36202, _36203, _36204,
         _36205, _36206, _36207, _36208, _36209, _36210, _36211, _36212,
         _36213, _36214, _36215, _36216, _36217, _36218, _36219, _36220,
         _36221, _36222, _36223, _36224, _36225, _36226, _36227, _36228,
         _36229, _36230, _36231, _36232, _36233, _36234, _36235, _36236,
         _36237, _36238, _36239, _36240, _36241, _36242, _36243, _36244,
         _36245, _36246, _36247, _36248, _36249, _36250, _36251, _36252,
         _36253, _36254, _36255, _36256, _36257, _36258, _36259, _36260,
         _36261, _36262, _36263, _36264, _36265, _36266, _36267, _36268,
         _36269, _36270, _36271, _36272, _36273, _36274, _36275, _36276,
         _36277, _36278, _36279, _36280, _36281, _36282, _36283, _36284,
         _36285, _36286, _36287, _36288, _36289, _36290, _36291, _36292,
         _36293, _36294, _36295, _36296, _36297, _36298, _36299, _36300,
         _36301, _36302, _36303, _36304, _36305, _36306, _36307, _36308,
         _36309, _36310, _36311, _36312, _36313, _36314, _36315, _36316,
         _36317, _36318, _36319, _36320, _36321, _36322, _36323, _36324,
         _36325, _36326, _36327, _36328, _36329, _36330, _36331, _36332,
         _36333, _36334, _36335, _36336, _36337, _36338, _36339, _36340,
         _36341, _36342, _36343, _36344, _36345, _36346, _36347, _36348,
         _36349, _36350, _36351, _36352, _36353, _36354, _36355, _36356,
         _36357, _36358, _36359, _36360, _36361, _36362, _36363, _36364,
         _36365, _36366, _36367, _36368, _36369, _36370, _36371, _36372,
         _36373, _36374, _36375, _36376, _36377, _36378, _36379, _36380,
         _36381, _36382, _36383, _36384, _36385, _36386, _36387, _36388,
         _36389, _36390, _36391, _36392, _36393, _36394, _36395, _36396,
         _36397, _36398, _36399, _36400, _36401, _36402, _36403, _36404,
         _36405, _36406, _36407, _36408, _36409, _36410, _36411, _36412,
         _36413, _36414, _36415, _36416, _36417, _36418, _36419, _36420,
         _36421, _36422, _36423, _36424, _36425, _36426, _36427, _36428,
         _36429, _36430, _36431, _36432, _36433, _36434, _36435, _36436,
         _36437, _36438, _36439, _36440, _36441, _36442, _36443, _36444,
         _36445, _36446, _36447, _36448, _36449, _36450, _36451, _36452,
         _36453, _36454, _36455, _36456, _36457, _36458, _36459, _36460,
         _36461, _36462, _36463, _36464, _36465, _36466, _36467, _36468,
         _36469, _36470, _36471, _36472, _36473, _36474, _36475, _36476,
         _36477, _36478, _36479, _36480, _36481, _36482, _36483, _36484,
         _36485, _36486, _36487, _36488, _36489, _36490, _36491, _36492,
         _36493, _36494, _36495, _36496, _36497, _36498, _36499, _36500,
         _36501, _36502, _36503, _36504, _36505, _36506, _36507, _36508,
         _36509, _36510, _36511, _36512, _36513, _36514, _36515, _36516,
         _36517, _36518, _36519, _36520, _36521, _36522, _36523, _36524,
         _36525, _36526, _36527, _36528, _36529, _36530, _36531, _36532,
         _36533, _36534, _36535, _36536, _36537, _36538, _36539, _36540,
         _36541, _36542, _36543, _36544, _36545, _36546, _36547, _36548,
         _36549, _36550, _36551, _36552, _36553, _36554, _36555, _36556,
         _36557, _36558, _36559, _36560, _36561, _36562, _36563, _36564,
         _36565, _36566, _36567, _36568, _36569, _36570, _36571, _36572,
         _36573, _36574, _36575, _36576, _36577, _36578, _36579, _36580,
         _36581, _36582, _36583, _36584, _36585, _36586, _36587, _36588,
         _36589, _36590, _36591, _36592, _36593, _36594, _36595, _36596,
         _36597, _36598, _36599, _36600, _36601, _36602, _36603, _36604,
         _36605, _36606, _36607, _36608, _36609, _36610, _36611, _36612,
         _36613, _36614, _36615, _36616, _36617, _36618, _36619, _36620,
         _36621, _36622, _36623, _36624, _36625, _36626, _36627, _36628,
         _36629, _36630, _36631, _36632, _36633, _36634, _36635, _36636,
         _36637, _36638, _36639, _36640, _36641, _36642, _36643, _36644,
         _36645, _36646, _36647, _36648, _36649, _36650, _36651, _36652,
         _36653, _36654, _36655, _36656, _36657, _36658, _36659, _36660,
         _36661, _36662, _36663, _36664, _36665, _36666, _36667, _36668,
         _36669, _36670, _36671, _36672, _36673, _36674, _36675, _36676,
         _36677, _36678, _36679, _36680, _36681, _36682, _36683, _36684,
         _36685, _36686, _36687, _36688, _36689, _36690, _36691, _36692,
         _36693, _36694, _36695, _36696, _36697, _36698, _36699, _36700,
         _36701, _36702, _36703, _36704, _36705, _36706, _36707, _36708,
         _36709, _36710, _36711, _36712, _36713, _36714, _36715, _36716,
         _36717, _36718, _36719, _36720, _36721, _36722, _36723, _36724,
         _36725, _36726, _36727, _36728, _36729, _36730, _36731, _36732,
         _36733, _36734, _36735, _36736, _36737, _36738, _36739, _36740,
         _36741, _36742, _36743, _36744, _36745, _36746, _36747, _36748,
         _36749, _36750, _36751, _36752, _36753, _36754, _36755, _36756,
         _36757, _36758, _36759, _36760, _36761, _36762, _36763, _36764,
         _36765, _36766, _36767, _36768, _36769, _36770, _36771, _36772,
         _36773, _36774, _36775, _36776, _36777, _36778, _36779, _36780,
         _36781, _36782, _36783, _36784, _36785, _36786, _36787, _36788,
         _36789, _36790, _36791, _36792, _36793, _36794, _36795, _36796,
         _36797, _36798, _36799, _36800, _36801, _36802, _36803, _36804,
         _36805, _36806, _36807, _36808, _36809, _36810, _36811, _36812,
         _36813, _36814, _36815, _36816, _36817, _36818, _36819, _36820,
         _36821, _36822, _36823, _36824, _36825, _36826, _36827, _36828,
         _36829, _36830, _36831, _36832, _36833, _36834, _36835, _36836,
         _36837, _36838, _36839, _36840, _36841, _36842, _36843, _36844,
         _36845, _36846, _36847, _36848, _36849, _36850, _36851, _36852,
         _36853, _36854, _36855, _36856, _36857, _36858, _36859, _36860,
         _36861, _36862, _36863, _36864, _36865, _36866, _36867, _36868,
         _36869, _36870, _36871, _36872, _36873, _36874, _36875, _36876,
         _36877, _36878, _36879, _36880, _36881, _36882, _36883, _36884,
         _36885, _36886, _36887, _36888, _36889, _36890, _36891, _36892,
         _36893, _36894, _36895, _36896, _36897, _36898, _36899, _36900,
         _36901, _36902, _36903, _36904, _36905, _36906, _36907, _36908,
         _36909, _36910, _36911, _36912, _36913, _36914, _36915, _36916,
         _36917, _36918, _36919, _36920, _36921, _36922, _36923, _36924,
         _36925, _36926, _36927, _36928, _36929, _36930, _36931, _36932,
         _36933, _36934, _36935, _36936, _36937, _36938, _36939, _36940,
         _36941, _36942, _36943, _36944, _36945, _36946, _36947, _36948,
         _36949, _36950, _36951, _36952, _36953, _36954, _36955, _36956,
         _36957, _36958, _36959, _36960, _36961, _36962, _36963, _36964,
         _36965, _36966, _36967, _36968, _36969, _36970, _36971, _36972,
         _36973, _36974, _36975, _36976, _36977, _36978, _36979, _36980,
         _36981, _36982, _36983, _36984, _36985, _36986, _36987, _36988,
         _36989, _36990, _36991, _36992, _36993, _36994, _36995, _36996,
         _36997, _36998, _36999, _37000, _37001, _37002, _37003, _37004,
         _37005, _37006, _37007, _37008, _37009, _37010, _37011, _37012,
         _37013, _37014, _37015, _37016, _37017, _37018, _37019, _37020,
         _37021, _37022, _37023, _37024, _37025, _37026, _37027, _37028,
         _37029, _37030, _37031, _37032, _37033, _37034, _37035, _37036,
         _37037, _37038, _37039, _37040, _37041, _37042, _37043, _37044,
         _37045, _37046, _37047, _37048, _37049, _37050, _37051, _37052,
         _37053, _37054, _37055, _37056, _37057, _37058, _37059, _37060,
         _37061, _37062, _37063, _37064, _37065, _37066, _37067, _37068,
         _37069, _37070, _37071, _37072, _37073, _37074, _37075, _37076,
         _37077, _37078, _37079, _37080, _37081, _37082, _37083, _37084,
         _37085, _37086, _37087, _37088, _37089, _37090, _37091, _37092,
         _37093, _37094, _37095, _37096, _37097, _37098, _37099, _37100,
         _37101, _37102, _37103, _37104, _37105, _37106, _37107, _37108,
         _37109, _37110, _37111, _37112, _37113, _37114, _37115, _37116,
         _37117, _37118, _37119, _37120, _37121, _37122, _37123, _37124,
         _37125, _37126, _37127, _37128, _37129, _37130, _37131, _37132,
         _37133, _37134, _37135, _37136, _37137, _37138, _37139, _37140,
         _37141, _37142, _37143, _37144, _37145, _37146, _37147, _37148,
         _37149, _37150, _37151, _37152, _37153, _37154, _37155, _37156,
         _37157, _37158, _37159, _37160, _37161, _37162, _37163, _37164,
         _37165, _37166, _37167, _37168, _37169, _37170, _37171, _37172,
         _37173, _37174, _37175, _37176, _37177, _37178, _37179, _37180,
         _37181, _37182, _37183, _37184, _37185, _37186, _37187, _37188,
         _37189, _37190, _37191, _37192, _37193, _37194, _37195, _37196,
         _37197, _37198, _37199, _37200, _37201, _37202, _37203, _37204,
         _37205, _37206, _37207, _37208, _37209, _37210, _37211, _37212,
         _37213, _37214, _37215, _37216, _37217, _37218, _37219, _37220,
         _37221, _37222, _37223, _37224, _37225, _37226, _37227, _37228,
         _37229, _37230, _37231, _37232, _37233, _37234, _37235, _37236,
         _37237, _37238, _37239, _37240, _37241, _37242, _37243, _37244,
         _37245, _37246, _37247, _37248, _37249, _37250, _37251, _37252,
         _37253, _37254, _37255, _37256, _37257, _37258, _37259, _37260,
         _37261, _37262, _37263, _37264, _37265, _37266, _37267, _37268,
         _37269, _37270, _37271, _37272, _37273, _37274, _37275, _37276,
         _37277, _37278, _37279, _37280, _37281, _37282, _37283, _37284,
         _37285, _37286, _37287, _37288, _37289, _37290, _37291, _37292,
         _37293, _37294, _37295, _37296, _37297, _37298, _37299, _37300,
         _37301, _37302, _37303, _37304, _37305, _37306, _37307, _37308,
         _37309, _37310, _37311, _37312, _37313, _37314, _37315, _37316,
         _37317, _37318, _37319, _37320, _37321, _37322, _37323, _37324,
         _37325, _37326, _37327, _37328, _37329, _37330, _37331, _37332,
         _37333, _37334, _37335, _37336, _37337, _37338, _37339, _37340,
         _37341, _37342, _37343, _37344, _37345, _37346, _37347, _37348,
         _37349, _37350, _37351, _37352, _37353, _37354, _37355, _37356,
         _37357, _37358, _37359, _37360, _37361, _37362, _37363, _37364,
         _37365, _37366, _37367, _37368, _37369, _37370, _37371, _37372,
         _37373, _37374, _37375, _37376, _37377, _37378, _37379, _37380,
         _37381, _37382, _37383, _37384, _37385, _37386, _37387, _37388,
         _37389, _37390, _37391, _37392, _37393, _37394, _37395, _37396,
         _37397, _37398, _37399, _37400, _37401, _37402, _37403, _37404,
         _37405, _37406, _37407, _37408, _37409, _37410, _37411, _37412,
         _37413, _37414, _37415, _37416, _37417, _37418, _37419, _37420,
         _37421, _37422, _37423, _37424, _37425, _37426, _37427, _37428,
         _37429, _37430, _37431, _37432, _37433, _37434, _37435, _37436,
         _37437, _37438, _37439, _37440, _37441, _37442, _37443, _37444,
         _37445, _37446, _37447, _37448, _37449, _37450, _37451, _37452,
         _37453, _37454, _37455, _37456, _37457, _37458, _37459, _37460,
         _37461, _37462, _37463, _37464, _37465, _37466, _37467, _37468,
         _37469, _37470, _37471, _37472, _37473, _37474, _37475, _37476,
         _37477, _37478, _37479, _37480, _37481, _37482, _37483, _37484,
         _37485, _37486, _37487, _37488, _37489, _37490, _37491, _37492,
         _37493, _37494, _37495, _37496, _37497, _37498, _37499, _37500,
         _37501, _37502, _37503, _37504, _37505, _37506, _37507, _37508,
         _37509, _37510, _37511, _37512, _37513, _37514, _37515, _37516,
         _37517, _37518, _37519, _37520, _37521, _37522, _37523, _37524,
         _37525, _37526, _37527, _37528, _37529, _37530, _37531, _37532,
         _37533, _37534, _37535, _37536, _37537, _37538, _37539, _37540,
         _37541, _37542, _37543, _37544, _37545, _37546, _37547, _37548,
         _37549, _37550, _37551, _37552, _37553, _37554, _37555, _37556,
         _37557, _37558, _37559, _37560, _37561, _37562, _37563, _37564,
         _37565, _37566, _37567, _37568, _37569, _37570, _37571, _37572,
         _37573, _37574, _37575, _37576, _37577, _37578, _37579, _37580,
         _37581, _37582, _37583, _37584, _37585, _37586, _37587, _37588,
         _37589, _37590, _37591, _37592, _37593, _37594, _37595, _37596,
         _37597, _37598, _37599, _37600, _37601, _37602, _37603, _37604,
         _37605, _37606, _37607, _37608, _37609, _37610, _37611, _37612,
         _37613, _37614, _37615, _37616, _37617, _37618, _37619, _37620,
         _37621, _37622, _37623, _37624, _37625, _37626, _37627, _37628,
         _37629, _37630, _37631, _37632, _37633, _37634, _37635, _37636,
         _37637, _37638, _37639, _37640, _37641, _37642, _37643, _37644,
         _37645, _37646, _37647, _37648, _37649, _37650, _37651, _37652,
         _37653, _37654, _37655, _37656, _37657, _37658, _37659, _37660,
         _37661, _37662, _37663, _37664, _37665, _37666, _37667, _37668,
         _37669, _37670, _37671, _37672, _37673, _37674, _37675, _37676,
         _37677, _37678, _37679, _37680, _37681, _37682, _37683, _37684,
         _37685, _37686, _37687, _37688, _37689, _37690, _37691, _37692,
         _37693, _37694, _37695, _37696, _37697, _37698, _37699, _37700,
         _37701, _37702, _37703, _37704, _37705, _37706, _37707, _37708,
         _37709, _37710, _37711, _37712, _37713, _37714, _37715, _37716,
         _37717, _37718, _37719, _37720, _37721, _37722, _37723, _37724,
         _37725, _37726, _37727, _37728, _37729, _37730, _37731, _37732,
         _37733, _37734, _37735, _37736, _37737, _37738, _37739, _37740,
         _37741, _37742, _37743, _37744, _37745, _37746, _37747, _37748,
         _37749, _37750, _37751, _37752, _37753, _37754, _37755, _37756,
         _37757, _37758, _37759, _37760, _37761, _37762, _37763, _37764,
         _37765, _37766, _37767, _37768, _37769, _37770, _37771, _37772,
         _37773, _37774, _37775, _37776, _37777, _37778, _37779, _37780,
         _37781, _37782, _37783, _37784, _37785, _37786, _37787, _37788,
         _37789, _37790, _37791, _37792, _37793, _37794, _37795, _37796,
         _37797, _37798, _37799, _37800, _37801, _37802, _37803, _37804,
         _37805, _37806, _37807, _37808, _37809, _37810, _37811, _37812,
         _37813, _37814, _37815, _37816, _37817, _37818, _37819, _37820,
         _37821, _37822, _37823, _37824, _37825, _37826, _37827, _37828,
         _37829, _37830, _37831, _37832, _37833, _37834, _37835, _37836,
         _37837, _37838, _37839, _37840, _37841, _37842, _37843, _37844,
         _37845, _37846, _37847, _37848, _37849, _37850, _37851, _37852,
         _37853, _37854, _37855, _37856, _37857, _37858, _37859, _37860,
         _37861, _37862, _37863, _37864, _37865, _37866, _37867, _37868,
         _37869, _37870, _37871, _37872, _37873, _37874, _37875, _37876,
         _37877, _37878, _37879, _37880, _37881, _37882, _37883, _37884,
         _37885, _37886, _37887, _37888, _37889, _37890, _37891, _37892,
         _37893, _37894, _37895, _37896, _37897, _37898, _37899, _37900,
         _37901, _37902, _37903, _37904, _37905, _37906, _37907, _37908,
         _37909, _37910, _37911, _37912, _37913, _37914, _37915, _37916,
         _37917, _37918, _37919, _37920, _37921, _37922, _37923, _37924,
         _37925, _37926, _37927, _37928, _37929, _37930, _37931, _37932,
         _37933, _37934, _37935, _37936, _37937, _37938, _37939, _37940,
         _37941, _37942, _37943, _37944, _37945, _37946, _37947, _37948,
         _37949, _37950, _37951, _37952, _37953, _37954, _37955, _37956,
         _37957, _37958, _37959, _37960, _37961, _37962, _37963, _37964,
         _37965, _37966, _37967, _37968, _37969, _37970, _37971, _37972,
         _37973, _37974, _37975, _37976, _37977, _37978, _37979, _37980,
         _37981, _37982, _37983, _37984, _37985, _37986, _37987, _37988,
         _37989, _37990, _37991, _37992, _37993, _37994, _37995, _37996,
         _37997, _37998, _37999, _38000, _38001, _38002, _38003, _38004,
         _38005, _38006, _38007, _38008, _38009, _38010, _38011, _38012,
         _38013, _38014, _38015, _38016, _38017, _38018, _38019, _38020,
         _38021, _38022, _38023, _38024, _38025, _38026, _38027, _38028,
         _38029, _38030, _38031, _38032, _38033, _38034, _38035, _38036,
         _38037, _38038, _38039, _38040, _38041, _38042, _38043, _38044,
         _38045, _38046, _38047, _38048, _38049, _38050, _38051, _38052,
         _38053, _38054, _38055, _38056, _38057, _38058, _38059, _38060,
         _38061, _38062, _38063, _38064, _38065, _38066, _38067, _38068,
         _38069, _38070, _38071, _38072, _38073, _38074, _38075, _38076,
         _38077, _38078, _38079, _38080, _38081, _38082, _38083, _38084,
         _38085, _38086, _38087, _38088, _38089, _38090, _38091, _38092,
         _38093, _38094, _38095, _38096, _38097, _38098, _38099, _38100,
         _38101, _38102, _38103, _38104, _38105, _38106, _38107, _38108,
         _38109, _38110, _38111, _38112, _38113, _38114, _38115, _38116,
         _38117, _38118, _38119, _38120, _38121, _38122, _38123, _38124,
         _38125, _38126, _38127, _38128, _38129, _38130, _38131, _38132,
         _38133, _38134, _38135, _38136, _38137, _38138, _38139, _38140,
         _38141, _38142, _38143, _38144, _38145, _38146, _38147, _38148,
         _38149, _38150, _38151, _38152, _38153, _38154, _38155, _38156,
         _38157, _38158, _38159, _38160, _38161, _38162, _38163, _38164,
         _38165, _38166, _38167, _38168, _38169, _38170, _38171, _38172,
         _38173, _38174, _38175, _38176, _38177, _38178, _38179, _38180,
         _38181, _38182, _38183, _38184, _38185, _38186, _38187, _38188,
         _38189, _38190, _38191, _38192, _38193, _38194, _38195, _38196,
         _38197, _38198, _38199, _38200, _38201, _38202, _38203, _38204,
         _38205, _38206, _38207, _38208, _38209, _38210, _38211, _38212,
         _38213, _38214, _38215, _38216, _38217, _38218, _38219, _38220,
         _38221, _38222, _38223, _38224, _38225, _38226, _38227, _38228,
         _38229, _38230, _38231, _38232, _38233, _38234, _38235, _38236,
         _38237, _38238, _38239, _38240, _38241, _38242, _38243, _38244,
         _38245, _38246, _38247, _38248, _38249, _38250, _38251, _38252,
         _38253, _38254, _38255, _38256, _38257, _38258, _38259, _38260,
         _38261, _38262, _38263, _38264, _38265, _38266, _38267, _38268,
         _38269, _38270, _38271, _38272, _38273, _38274, _38275, _38276,
         _38277, _38278, _38279, _38280, _38281, _38282, _38283, _38284,
         _38285, _38286, _38287, _38288, _38289, _38290, _38291, _38292,
         _38293, _38294, _38295, _38296, _38297, _38298, _38299, _38300,
         _38301, _38302, _38303, _38304, _38305, _38306, _38307, _38308,
         _38309, _38310, _38311, _38312, _38313, _38314, _38315, _38316,
         _38317, _38318, _38319, _38320, _38321, _38322, _38323, _38324,
         _38325, _38326, _38327, _38328, _38329, _38330, _38331, _38332,
         _38333, _38334, _38335, _38336, _38337, _38338, _38339, _38340,
         _38341, _38342, _38343, _38344, _38345, _38346, _38347, _38348,
         _38349, _38350, _38351, _38352, _38353, _38354, _38355, _38356,
         _38357, _38358, _38359, _38360, _38361, _38362, _38363, _38364,
         _38365, _38366, _38367, _38368, _38369, _38370, _38371, _38372,
         _38373, _38374, _38375, _38376, _38377, _38378, _38379, _38380,
         _38381, _38382, _38383, _38384, _38385, _38386, _38387, _38388,
         _38389, _38390, _38391, _38392, _38393, _38394, _38395, _38396,
         _38397, _38398, _38399, _38400, _38401, _38402, _38403, _38404,
         _38405, _38406, _38407, _38408, _38409, _38410, _38411, _38412,
         _38413, _38414, _38415, _38416, _38417, _38418, _38419, _38420,
         _38421, _38422, _38423, _38424, _38425, _38426, _38427, _38428,
         _38429, _38430, _38431, _38432, _38433, _38434, _38435, _38436,
         _38437, _38438, _38439, _38440, _38441, _38442, _38443, _38444,
         _38445, _38446, _38447, _38448, _38449, _38450, _38451, _38452,
         _38453, _38454, _38455, _38456, _38457, _38458, _38459, _38460,
         _38461, _38462, _38463, _38464, _38465, _38466, _38467, _38468,
         _38469, _38470, _38471, _38472, _38473, _38474, _38475, _38476,
         _38477, _38478, _38479, _38480, _38481, _38482, _38483, _38484,
         _38485, _38486, _38487, _38488, _38489, _38490, _38491, _38492,
         _38493, _38494, _38495, _38496, _38497, _38498, _38499, _38500,
         _38501, _38502, _38503, _38504, _38505, _38506, _38507, _38508,
         _38509, _38510, _38511, _38512, _38513, _38514, _38515, _38516,
         _38517, _38518, _38519, _38520, _38521, _38522, _38523, _38524,
         _38525, _38526, _38527, _38528, _38529, _38530, _38531, _38532,
         _38533, _38534, _38535, _38536, _38537, _38538, _38539, _38540,
         _38541, _38542, _38543, _38544, _38545, _38546, _38547, _38548,
         _38549, _38550, _38551, _38552, _38553, _38554, _38555, _38556,
         _38557, _38558, _38559, _38560, _38561, _38562, _38563, _38564,
         _38565, _38566, _38567, _38568, _38569, _38570, _38571, _38572,
         _38573, _38574, _38575, _38576, _38577, _38578, _38579, _38580,
         _38581, _38582, _38583, _38584, _38585, _38586, _38587, _38588,
         _38589, _38590, _38591, _38592, _38593, _38594, _38595, _38596,
         _38597, _38598, _38599, _38600, _38601, _38602, _38603, _38604,
         _38605, _38606, _38607, _38608, _38609, _38610, _38611, _38612,
         _38613, _38614, _38615, _38616, _38617, _38618, _38619, _38620,
         _38621, _38622, _38623, _38624, _38625, _38626, _38627, _38628,
         _38629, _38630, _38631, _38632, _38633, _38634, _38635, _38636,
         _38637, _38638, _38639, _38640, _38641, _38642, _38643, _38644,
         _38645, _38646, _38647, _38648, _38649, _38650, _38651, _38652,
         _38653, _38654, _38655, _38656, _38657, _38658, _38659, _38660,
         _38661, _38662, _38663, _38664, _38665, _38666, _38667, _38668,
         _38669, _38670, _38671, _38672, _38673, _38674, _38675, _38676,
         _38677, _38678, _38679, _38680, _38681, _38682, _38683, _38684,
         _38685, _38686, _38687, _38688, _38689, _38690, _38691, _38692,
         _38693, _38694, _38695, _38696, _38697, _38698, _38699, _38700,
         _38701, _38702, _38703, _38704, _38705, _38706, _38707, _38708,
         _38709, _38710, _38711, _38712, _38713, _38714, _38715, _38716,
         _38717, _38718, _38719, _38720, _38721, _38722, _38723, _38724,
         _38725, _38726, _38727, _38728, _38729, _38730, _38731, _38732,
         _38733, _38734, _38735, _38736, _38737, _38738, _38739, _38740,
         _38741, _38742, _38743, _38744, _38745, _38746, _38747, _38748,
         _38749, _38750, _38751, _38752, _38753, _38754, _38755, _38756,
         _38757, _38758, _38759, _38760, _38761, _38762, _38763, _38764,
         _38765, _38766, _38767, _38768, _38769, _38770, _38771, _38772,
         _38773, _38774, _38775, _38776, _38777, _38778, _38779, _38780,
         _38781, _38782, _38783, _38784, _38785, _38786, _38787, _38788,
         _38789, _38790, _38791, _38792, _38793, _38794, _38795, _38796,
         _38797, _38798, _38799, _38800, _38801, _38802, _38803, _38804,
         _38805, _38806, _38807, _38808, _38809, _38810, _38811, _38812,
         _38813, _38814, _38815, _38816, _38817, _38818, _38819, _38820,
         _38821, _38822, _38823, _38824, _38825, _38826, _38827, _38828,
         _38829, _38830, _38831, _38832, _38833, _38834, _38835, _38836,
         _38837, _38838, _38839, _38840, _38841, _38842, _38843, _38844,
         _38845, _38846, _38847, _38848, _38849, _38850, _38851, _38852,
         _38853, _38854, _38855, _38856, _38857, _38858, _38859, _38860,
         _38861, _38862, _38863, _38864, _38865, _38866, _38867, _38868,
         _38869, _38870, _38871, _38872, _38873, _38874, _38875, _38876,
         _38877, _38878, _38879, _38880, _38881, _38882, _38883, _38884,
         _38885, _38886, _38887, _38888, _38889, _38890, _38891, _38892,
         _38893, _38894, _38895, _38896, _38897, _38898, _38899, _38900,
         _38901, _38902, _38903, _38904, _38905, _38906, _38907, _38908,
         _38909, _38910, _38911, _38912, _38913, _38914, _38915, _38916,
         _38917, _38918, _38919, _38920, _38921, _38922, _38923, _38924,
         _38925, _38926, _38927, _38928, _38929, _38930, _38931, _38932,
         _38933, _38934, _38935, _38936, _38937, _38938, _38939, _38940,
         _38941, _38942, _38943, _38944, _38945, _38946, _38947, _38948,
         _38949, _38950, _38951, _38952, _38953, _38954, _38955, _38956,
         _38957, _38958, _38959, _38960, _38961, _38962, _38963, _38964,
         _38965, _38966, _38967, _38968, _38969, _38970, _38971, _38972,
         _38973, _38974, _38975, _38976, _38977, _38978, _38979, _38980,
         _38981, _38982, _38983, _38984, _38985, _38986, _38987, _38988,
         _38989, _38990, _38991, _38992, _38993, _38994, _38995, _38996,
         _38997, _38998, _38999, _39000, _39001, _39002, _39003, _39004,
         _39005, _39006, _39007, _39008, _39009, _39010, _39011, _39012,
         _39013, _39014, _39015, _39016, _39017, _39018, _39019, _39020,
         _39021, _39022, _39023, _39024, _39025, _39026, _39027, _39028,
         _39029, _39030, _39031, _39032, _39033, _39034, _39035, _39036,
         _39037, _39038, _39039, _39040, _39041, _39042, _39043, _39044,
         _39045, _39046, _39047, _39048, _39049, _39050, _39051, _39052,
         _39053, _39054, _39055, _39056, _39057, _39058, _39059, _39060,
         _39061, _39062, _39063, _39064, _39065, _39066, _39067, _39068,
         _39069, _39070, _39071, _39072, _39073, _39074, _39075, _39076,
         _39077, _39078, _39079, _39080, _39081, _39082, _39083, _39084,
         _39085, _39086, _39087, _39088, _39089, _39090, _39091, _39092,
         _39093, _39094, _39095, _39096, _39097, _39098, _39099, _39100,
         _39101, _39102, _39103, _39104, _39105, _39106, _39107, _39108,
         _39109, _39110, _39111, _39112, _39113, _39114, _39115, _39116,
         _39117, _39118, _39119, _39120, _39121, _39122, _39123, _39124,
         _39125, _39126, _39127, _39128, _39129, _39130, _39131, _39132,
         _39133, _39134, _39135, _39136, _39137, _39138, _39139, _39140,
         _39141, _39142, _39143, _39144, _39145, _39146, _39147, _39148,
         _39149, _39150, _39151, _39152, _39153, _39154, _39155, _39156,
         _39157, _39158, _39159, _39160, _39161, _39162, _39163, _39164,
         _39165, _39166, _39167, _39168, _39169, _39170, _39171, _39172,
         _39173, _39174, _39175, _39176, _39177, _39178, _39179, _39180,
         _39181, _39182, _39183, _39184, _39185, _39186, _39187, _39188,
         _39189, _39190, _39191, _39192, _39193, _39194, _39195, _39196,
         _39197, _39198, _39199, _39200, _39201, _39202, _39203, _39204,
         _39205, _39206, _39207, _39208, _39209, _39210, _39211, _39212,
         _39213, _39214, _39215, _39216, _39217, _39218, _39219, _39220,
         _39221, _39222, _39223, _39224, _39225, _39226, _39227, _39228,
         _39229, _39230, _39231, _39232, _39233, _39234, _39235, _39236,
         _39237, _39238, _39239, _39240, _39241, _39242, _39243, _39244,
         _39245, _39246, _39247, _39248, _39249, _39250, _39251, _39252,
         _39253, _39254, _39255, _39256, _39257, _39258, _39259, _39260,
         _39261, _39262, _39263, _39264, _39265, _39266, _39267, _39268,
         _39269, _39270, _39271, _39272, _39273, _39274, _39275, _39276,
         _39277, _39278, _39279, _39280, _39281, _39282, _39283, _39284,
         _39285, _39286, _39287, _39288, _39289, _39290, _39291, _39292,
         _39293, _39294, _39295, _39296, _39297, _39298, _39299, _39300,
         _39301, _39302, _39303, _39304, _39305, _39306, _39307, _39308,
         _39309, _39310, _39311, _39312, _39313, _39314, _39315, _39316,
         _39317, _39318, _39319, _39320, _39321, _39322, _39323, _39324,
         _39325, _39326, _39327, _39328, _39329, _39330, _39331, _39332,
         _39333, _39334, _39335, _39336, _39337, _39338, _39339, _39340,
         _39341, _39342, _39343, _39344, _39345, _39346, _39347, _39348,
         _39349, _39350, _39351, _39352, _39353, _39354, _39355, _39356,
         _39357, _39358, _39359, _39360, _39361, _39362, _39363, _39364,
         _39365, _39366, _39367, _39368, _39369, _39370, _39371, _39372,
         _39373, _39374, _39375, _39376, _39377, _39378, _39379, _39380,
         _39381, _39382, _39383, _39384, _39385, _39386, _39387, _39388,
         _39389, _39390, _39391, _39392, _39393, _39394, _39395, _39396,
         _39397, _39398, _39399, _39400, _39401, _39402, _39403, _39404,
         _39405, _39406, _39407, _39408, _39409, _39410, _39411, _39412,
         _39413, _39414, _39415, _39416, _39417, _39418, _39419, _39420,
         _39421, _39422, _39423, _39424, _39425, _39426, _39427, _39428,
         _39429, _39430, _39431, _39432, _39433, _39434, _39435, _39436,
         _39437, _39438, _39439, _39440, _39441, _39442, _39443, _39444,
         _39445, _39446, _39447, _39448, _39449, _39450, _39451, _39452,
         _39453, _39454, _39455, _39456, _39457, _39458, _39459, _39460,
         _39461, _39462, _39463, _39464, _39465, _39466, _39467, _39468,
         _39469, _39470, _39471, _39472, _39473, _39474, _39475, _39476,
         _39477, _39478, _39479, _39480, _39481, _39482, _39483, _39484,
         _39485, _39486, _39487, _39488, _39489, _39490, _39491, _39492,
         _39493, _39494, _39495, _39496, _39497, _39498, _39499, _39500,
         _39501, _39502, _39503, _39504, _39505, _39506, _39507, _39508,
         _39509, _39510, _39511, _39512, _39513, _39514, _39515, _39516,
         _39517, _39518, _39519, _39520, _39521, _39522, _39523, _39524,
         _39525, _39526, _39527, _39528, _39529, _39530, _39531, _39532,
         _39533, _39534, _39535, _39536, _39537, _39538, _39539, _39540,
         _39541, _39542, _39543, _39544, _39545, _39546, _39547, _39548,
         _39549, _39550, _39551, _39552, _39553, _39554, _39555, _39556,
         _39557, _39558, _39559, _39560, _39561, _39562, _39563, _39564,
         _39565, _39566, _39567, _39568, _39569, _39570, _39571, _39572,
         _39573, _39574, _39575, _39576, _39577, _39578, _39579, _39580,
         _39581, _39582, _39583, _39584, _39585, _39586, _39587, _39588,
         _39589, _39590, _39591, _39592, _39593, _39594, _39595, _39596,
         _39597, _39598, _39599, _39600, _39601, _39602, _39603, _39604,
         _39605, _39606, _39607, _39608, _39609, _39610, _39611, _39612,
         _39613, _39614, _39615, _39616, _39617, _39618, _39619, _39620,
         _39621, _39622, _39623, _39624, _39625, _39626, _39627, _39628,
         _39629, _39630, _39631, _39632, _39633, _39634, _39635, _39636,
         _39637, _39638, _39639, _39640, _39641, _39642, _39643, _39644,
         _39645, _39646, _39647, _39648, _39649, _39650, _39651, _39652,
         _39653, _39654, _39655, _39656, _39657, _39658, _39659, _39660,
         _39661, _39662, _39663, _39664, _39665, _39666, _39667, _39668,
         _39669, _39670, _39671, _39672, _39673, _39674, _39675, _39676,
         _39677, _39678, _39679, _39680, _39681, _39682, _39683, _39684,
         _39685, _39686, _39687, _39688, _39689, _39690, _39691, _39692,
         _39693, _39694, _39695, _39696, _39697, _39698, _39699, _39700,
         _39701, _39702, _39703, _39704, _39705, _39706, _39707, _39708,
         _39709, _39710, _39711, _39712, _39713, _39714, _39715, _39716,
         _39717, _39718, _39719, _39720, _39721, _39722, _39723, _39724,
         _39725, _39726, _39727, _39728, _39729, _39730, _39731, _39732,
         _39733, _39734, _39735, _39736, _39737, _39738, _39739, _39740,
         _39741, _39742, _39743, _39744, _39745, _39746, _39747, _39748,
         _39749, _39750, _39751, _39752, _39753, _39754, _39755, _39756,
         _39757, _39758, _39759, _39760, _39761, _39762, _39763, _39764,
         _39765, _39766, _39767, _39768, _39769, _39770, _39771, _39772,
         _39773, _39774, _39775, _39776, _39777, _39778, _39779, _39780,
         _39781, _39782, _39783, _39784, _39785, _39786, _39787, _39788,
         _39789, _39790, _39791, _39792, _39793, _39794, _39795, _39796,
         _39797, _39798, _39799, _39800, _39801, _39802, _39803, _39804,
         _39805, _39806, _39807, _39808, _39809, _39810, _39811, _39812,
         _39813, _39814, _39815, _39816, _39817, _39818, _39819, _39820,
         _39821, _39822, _39823, _39824, _39825, _39826, _39827, _39828,
         _39829, _39830, _39831, _39832, _39833, _39834, _39835, _39836,
         _39837, _39838, _39839, _39840, _39841, _39842, _39843, _39844,
         _39845, _39846, _39847, _39848, _39849, _39850, _39851, _39852,
         _39853, _39854, _39855, _39856, _39857, _39858, _39859, _39860,
         _39861, _39862, _39863, _39864, _39865, _39866, _39867, _39868,
         _39869, _39870, _39871, _39872, _39873, _39874, _39875, _39876,
         _39877, _39878, _39879, _39880, _39881, _39882, _39883, _39884,
         _39885, _39886, _39887, _39888, _39889, _39890, _39891, _39892,
         _39893, _39894, _39895, _39896, _39897, _39898, _39899, _39900,
         _39901, _39902, _39903, _39904, _39905, _39906, _39907, _39908,
         _39909, _39910, _39911, _39912, _39913, _39914, _39915, _39916,
         _39917, _39918, _39919, _39920, _39921, _39922, _39923, _39924,
         _39925, _39926, _39927, _39928, _39929, _39930, _39931, _39932,
         _39933, _39934, _39935, _39936, _39937, _39938, _39939, _39940,
         _39941, _39942, _39943, _39944, _39945, _39946, _39947, _39948,
         _39949, _39950, _39951, _39952, _39953, _39954, _39955, _39956,
         _39957, _39958, _39959, _39960, _39961, _39962, _39963, _39964,
         _39965, _39966, _39967, _39968, _39969, _39970, _39971, _39972,
         _39973, _39974, _39975, _39976, _39977, _39978, _39979, _39980,
         _39981, _39982, _39983, _39984, _39985, _39986, _39987, _39988,
         _39989, _39990, _39991, _39992, _39993, _39994, _39995, _39996,
         _39997, _39998, _39999, _40000, _40001, _40002, _40003, _40004,
         _40005, _40006, _40007, _40008, _40009, _40010, _40011, _40012,
         _40013, _40014, _40015, _40016, _40017, _40018, _40019, _40020,
         _40021, _40022, _40023, _40024, _40025, _40026, _40027, _40028,
         _40029, _40030, _40031, _40032, _40033, _40034, _40035, _40036,
         _40037, _40038, _40039, _40040, _40041, _40042, _40043, _40044,
         _40045, _40046, _40047, _40048, _40049, _40050, _40051, _40052,
         _40053, _40054, _40055, _40056, _40057, _40058, _40059, _40060,
         _40061, _40062, _40063, _40064, _40065, _40066, _40067, _40068,
         _40069, _40070, _40071, _40072, _40073, _40074, _40075, _40076,
         _40077, _40078, _40079, _40080, _40081, _40082, _40083, _40084,
         _40085, _40086, _40087, _40088, _40089, _40090, _40091, _40092,
         _40093, _40094, _40095, _40096, _40097, _40098, _40099, _40100,
         _40101, _40102, _40103, _40104, _40105, _40106, _40107, _40108,
         _40109, _40110, _40111, _40112, _40113, _40114, _40115, _40116,
         _40117, _40118, _40119, _40120, _40121, _40122, _40123, _40124,
         _40125, _40126, _40127, _40128, _40129, _40130, _40131, _40132,
         _40133, _40134, _40135, _40136, _40137, _40138, _40139, _40140,
         _40141, _40142, _40143, _40144, _40145, _40146, _40147, _40148,
         _40149, _40150, _40151, _40152, _40153, _40154, _40155, _40156,
         _40157, _40158, _40159, _40160, _40161, _40162, _40163, _40164,
         _40165, _40166, _40167, _40168, _40169, _40170, _40171, _40172,
         _40173, _40174, _40175, _40176, _40177, _40178, _40179, _40180,
         _40181, _40182, _40183, _40184, _40185, _40186, _40187, _40188,
         _40189, _40190, _40191, _40192, _40193, _40194, _40195, _40196,
         _40197, _40198, _40199, _40200, _40201, _40202, _40203, _40204,
         _40205, _40206, _40207, _40208, _40209, _40210, _40211, _40212,
         _40213, _40214, _40215, _40216, _40217, _40218, _40219, _40220,
         _40221, _40222, _40223, _40224, _40225, _40226, _40227, _40228,
         _40229, _40230, _40231, _40232, _40233, _40234, _40235, _40236,
         _40237, _40238, _40239, _40240, _40241, _40242, _40243, _40244,
         _40245, _40246, _40247, _40248, _40249, _40250, _40251, _40252,
         _40253, _40254, _40255, _40256, _40257, _40258, _40259, _40260,
         _40261, _40262, _40263, _40264, _40265, _40266, _40267, _40268,
         _40269, _40270, _40271, _40272, _40273, _40274, _40275, _40276,
         _40277, _40278, _40279, _40280, _40281, _40282, _40283, _40284,
         _40285, _40286, _40287, _40288, _40289, _40290, _40291, _40292,
         _40293, _40294, _40295, _40296, _40297, _40298, _40299, _40300,
         _40301, _40302, _40303, _40304, _40305, _40306, _40307, _40308,
         _40309, _40310, _40311, _40312, _40313, _40314, _40315, _40316,
         _40317, _40318, _40319, _40320, _40321, _40322, _40323, _40324,
         _40325, _40326, _40327, _40328, _40329, _40330, _40331, _40332,
         _40333, _40334, _40335, _40336, _40337, _40338, _40339, _40340,
         _40341, _40342, _40343, _40344, _40345, _40346, _40347, _40348,
         _40349, _40350, _40351, _40352, _40353, _40354, _40355, _40356,
         _40357, _40358, _40359, _40360, _40361, _40362, _40363, _40364,
         _40365, _40366, _40367, _40368, _40369, _40370, _40371, _40372,
         _40373, _40374, _40375, _40376, _40377, _40378, _40379, _40380,
         _40381, _40382, _40383, _40384, _40385, _40386, _40387, _40388,
         _40389, _40390, _40391, _40392, _40393, _40394, _40395, _40396,
         _40397, _40398, _40399, _40400, _40401, _40402, _40403, _40404,
         _40405, _40406, _40407, _40408, _40409, _40410, _40411, _40412,
         _40413, _40414, _40415, _40416, _40417, _40418, _40419, _40420,
         _40421, _40422, _40423, _40424, _40425, _40426, _40427, _40428,
         _40429, _40430, _40431, _40432, _40433, _40434, _40435, _40436,
         _40437, _40438, _40439, _40440, _40441, _40442, _40443, _40444,
         _40445, _40446, _40447, _40448, _40449, _40450, _40451, _40452,
         _40453, _40454, _40455, _40456, _40457, _40458, _40459, _40460,
         _40461, _40462, _40463, _40464, _40465, _40466, _40467, _40468,
         _40469, _40470, _40471, _40472, _40473, _40474, _40475, _40476,
         _40477, _40478, _40479, _40480, _40481, _40482, _40483, _40484,
         _40485, _40486, _40487, _40488, _40489, _40490, _40491, _40492,
         _40493, _40494, _40495, _40496, _40497, _40498, _40499, _40500,
         _40501, _40502, _40503, _40504, _40505, _40506, _40507, _40508,
         _40509, _40510, _40511, _40512, _40513, _40514, _40515, _40516,
         _40517, _40518, _40519, _40520, _40521, _40522, _40523, _40524,
         _40525, _40526, _40527, _40528, _40529, _40530, _40531, _40532,
         _40533, _40534, _40535, _40536, _40537, _40538, _40539, _40540,
         _40541, _40542, _40543, _40544, _40545, _40546, _40547, _40548,
         _40549, _40550, _40551, _40552, _40553, _40554, _40555, _40556,
         _40557, _40558, _40559, _40560, _40561, _40562, _40563, _40564,
         _40565, _40566, _40567, _40568, _40569, _40570, _40571, _40572,
         _40573, _40574, _40575, _40576, _40577, _40578, _40579, _40580,
         _40581, _40582, _40583, _40584, _40585, _40586, _40587, _40588,
         _40589, _40590, _40591, _40592, _40593, _40594, _40595, _40596,
         _40597, _40598, _40599, _40600, _40601, _40602, _40603, _40604,
         _40605, _40606, _40607, _40608, _40609, _40610, _40611, _40612,
         _40613, _40614, _40615, _40616, _40617, _40618, _40619, _40620,
         _40621, _40622, _40623, _40624, _40625, _40626, _40627, _40628,
         _40629, _40630, _40631, _40632, _40633, _40634, _40635, _40636,
         _40637, _40638, _40639, _40640, _40641, _40642, _40643, _40644,
         _40645, _40646, _40647, _40648, _40649, _40650, _40651, _40652,
         _40653, _40654, _40655, _40656, _40657, _40658, _40659, _40660,
         _40661, _40662, _40663, _40664, _40665, _40666, _40667, _40668,
         _40669, _40670, _40671, _40672, _40673, _40674, _40675, _40676,
         _40677, _40678, _40679, _40680, _40681, _40682, _40683, _40684,
         _40685, _40686, _40687, _40688, _40689, _40690, _40691, _40692,
         _40693, _40694, _40695, _40696, _40697, _40698, _40699, _40700,
         _40701, _40702, _40703, _40704, _40705, _40706, _40707, _40708,
         _40709, _40710, _40711, _40712, _40713, _40714, _40715, _40716,
         _40717, _40718, _40719, _40720, _40721, _40722, _40723, _40724,
         _40725, _40726, _40727, _40728, _40729, _40730, _40731, _40732,
         _40733, _40734, _40735, _40736, _40737, _40738, _40739, _40740,
         _40741, _40742, _40743, _40744, _40745, _40746, _40747, _40748,
         _40749, _40750, _40751, _40752, _40753, _40754, _40755, _40756,
         _40757, _40758, _40759, _40760, _40761, _40762, _40763, _40764,
         _40765, _40766, _40767, _40768, _40769, _40770, _40771, _40772,
         _40773, _40774, _40775, _40776, _40777, _40778, _40779, _40780,
         _40781, _40782, _40783, _40784, _40785, _40786, _40787, _40788,
         _40789, _40790, _40791, _40792, _40793, _40794, _40795, _40796,
         _40797, _40798, _40799, _40800, _40801, _40802, _40803, _40804,
         _40805, _40806, _40807, _40808, _40809, _40810, _40811, _40812,
         _40813, _40814, _40815, _40816, _40817, _40818, _40819, _40820,
         _40821, _40822, _40823, _40824, _40825, _40826, _40827, _40828,
         _40829, _40830, _40831, _40832, _40833, _40834, _40835, _40836,
         _40837, _40838, _40839, _40840, _40841, _40842, _40843, _40844,
         _40845, _40846, _40847, _40848, _40849, _40850, _40851, _40852,
         _40853, _40854, _40855, _40856, _40857, _40858, _40859, _40860,
         _40861, _40862, _40863, _40864, _40865, _40866, _40867, _40868,
         _40869, _40870, _40871, _40872, _40873, _40874, _40875, _40876,
         _40877, _40878, _40879, _40880, _40881, _40882, _40883, _40884,
         _40885, _40886, _40887, _40888, _40889, _40890, _40891, _40892,
         _40893, _40894, _40895, _40896, _40897, _40898, _40899, _40900,
         _40901, _40902, _40903, _40904, _40905, _40906, _40907, _40908,
         _40909, _40910, _40911, _40912, _40913, _40914, _40915, _40916,
         _40917, _40918, _40919, _40920, _40921, _40922, _40923, _40924,
         _40925, _40926, _40927, _40928, _40929, _40930, _40931, _40932,
         _40933, _40934, _40935, _40936, _40937, _40938, _40939, _40940,
         _40941, _40942, _40943, _40944, _40945, _40946, _40947, _40948,
         _40949, _40950, _40951, _40952, _40953, _40954, _40955, _40956,
         _40957, _40958, _40959, _40960, _40961, _40962, _40963, _40964,
         _40965, _40966, _40967, _40968, _40969, _40970, _40971, _40972,
         _40973, _40974, _40975, _40976, _40977, _40978, _40979, _40980,
         _40981, _40982, _40983, _40984, _40985, _40986, _40987, _40988,
         _40989, _40990, _40991, _40992, _40993, _40994, _40995, _40996,
         _40997, _40998, _40999, _41000, _41001, _41002, _41003, _41004,
         _41005, _41006, _41007, _41008, _41009, _41010, _41011, _41012,
         _41013, _41014, _41015, _41016, _41017, _41018, _41019, _41020,
         _41021, _41022, _41023, _41024, _41025, _41026, _41027, _41028,
         _41029, _41030, _41031, _41032, _41033, _41034, _41035, _41036,
         _41037, _41038, _41039, _41040, _41041, _41042, _41043, _41044,
         _41045, _41046, _41047, _41048, _41049, _41050, _41051, _41052,
         _41053, _41054, _41055, _41056, _41057, _41058, _41059, _41060,
         _41061, _41062, _41063, _41064, _41065, _41066, _41067, _41068,
         _41069, _41070, _41071, _41072, _41073, _41074, _41075, _41076,
         _41077, _41078, _41079, _41080, _41081, _41082, _41083, _41084,
         _41085, _41086, _41087, _41088, _41089, _41090, _41091, _41092,
         _41093, _41094, _41095, _41096, _41097, _41098, _41099, _41100,
         _41101, _41102, _41103, _41104, _41105, _41106, _41107, _41108,
         _41109, _41110, _41111, _41112, _41113, _41114, _41115, _41116,
         _41117, _41118, _41119, _41120, _41121, _41122, _41123, _41124,
         _41125, _41126, _41127, _41128, _41129, _41130, _41131, _41132,
         _41133, _41134, _41135, _41136, _41137, _41138, _41139, _41140,
         _41141, _41142, _41143, _41144, _41145, _41146, _41147, _41148,
         _41149, _41150, _41151, _41152, _41153, _41154, _41155, _41156,
         _41157, _41158, _41159, _41160, _41161, _41162, _41163, _41164,
         _41165, _41166, _41167, _41168, _41169, _41170, _41171, _41172,
         _41173, _41174, _41175, _41176, _41177, _41178, _41179, _41180,
         _41181, _41182, _41183, _41184, _41185, _41186, _41187, _41188,
         _41189, _41190, _41191, _41192, _41193, _41194, _41195, _41196,
         _41197, _41198, _41199, _41200, _41201, _41202, _41203, _41204,
         _41205, _41206, _41207, _41208, _41209, _41210, _41211, _41212,
         _41213, _41214, _41215, _41216, _41217, _41218, _41219, _41220,
         _41221, _41222, _41223, _41224, _41225, _41226, _41227, _41228,
         _41229, _41230, _41231, _41232, _41233, _41234, _41235, _41236,
         _41237, _41238, _41239, _41240, _41241, _41242, _41243, _41244,
         _41245, _41246, _41247, _41248, _41249, _41250, _41251, _41252,
         _41253, _41254, _41255, _41256, _41257, _41258, _41259, _41260,
         _41261, _41262, _41263, _41264, _41265, _41266, _41267, _41268,
         _41269, _41270, _41271, _41272, _41273, _41274, _41275, _41276,
         _41277, _41278, _41279, _41280, _41281, _41282, _41283, _41284,
         _41285, _41286, _41287, _41288, _41289, _41290, _41291, _41292,
         _41293, _41294, _41295, _41296, _41297, _41298, _41299, _41300,
         _41301, _41302, _41303, _41304, _41305, _41306, _41307, _41308,
         _41309, _41310, _41311, _41312, _41313, _41314, _41315, _41316,
         _41317, _41318, _41319, _41320, _41321, _41322, _41323, _41324,
         _41325, _41326, _41327, _41328, _41329, _41330, _41331, _41332,
         _41333, _41334, _41335, _41336, _41337, _41338, _41339, _41340,
         _41341, _41342, _41343, _41344, _41345, _41346, _41347, _41348,
         _41349, _41350, _41351, _41352, _41353, _41354, _41355, _41356,
         _41357, _41358, _41359, _41360, _41361, _41362, _41363, _41364,
         _41365, _41366, _41367, _41368, _41369, _41370, _41371, _41372,
         _41373, _41374, _41375, _41376, _41377, _41378, _41379, _41380,
         _41381, _41382, _41383, _41384, _41385, _41386, _41387, _41388,
         _41389, _41390, _41391, _41392, _41393, _41394, _41395, _41396,
         _41397, _41398, _41399, _41400, _41401, _41402, _41403, _41404,
         _41405, _41406, _41407, _41408, _41409, _41410, _41411, _41412,
         _41413, _41414, _41415, _41416, _41417, _41418, _41419, _41420,
         _41421, _41422, _41423, _41424, _41425, _41426, _41427, _41428,
         _41429, _41430, _41431, _41432, _41433, _41434, _41435, _41436,
         _41437, _41438, _41439, _41440, _41441, _41442, _41443, _41444,
         _41445, _41446, _41447, _41448, _41449, _41450, _41451, _41452,
         _41453, _41454, _41455, _41456, _41457, _41458, _41459, _41460,
         _41461, _41462, _41463, _41464, _41465, _41466, _41467, _41468,
         _41469, _41470, _41471, _41472, _41473, _41474, _41475, _41476,
         _41477, _41478, _41479, _41480, _41481, _41482, _41483, _41484,
         _41485, _41486, _41487, _41488, _41489, _41490, _41491, _41492,
         _41493, _41494, _41495, _41496, _41497, _41498, _41499, _41500,
         _41501, _41502, _41503, _41504, _41505, _41506, _41507, _41508,
         _41509, _41510, _41511, _41512, _41513, _41514, _41515, _41516,
         _41517, _41518, _41519, _41520, _41521, _41522, _41523, _41524,
         _41525, _41526, _41527, _41528, _41529, _41530, _41531, _41532,
         _41533, _41534, _41535, _41536, _41537, _41538, _41539, _41540,
         _41541, _41542, _41543, _41544, _41545, _41546, _41547, _41548,
         _41549, _41550, _41551, _41552, _41553, _41554, _41555, _41556,
         _41557, _41558, _41559, _41560, _41561, _41562, _41563, _41564,
         _41565, _41566, _41567, _41568, _41569, _41570, _41571, _41572,
         _41573, _41574, _41575, _41576, _41577, _41578, _41579, _41580,
         _41581, _41582, _41583, _41584, _41585, _41586, _41587, _41588,
         _41589, _41590, _41591, _41592, _41593, _41594, _41595, _41596,
         _41597, _41598, _41599, _41600, _41601, _41602, _41603, _41604,
         _41605, _41606, _41607, _41608, _41609, _41610, _41611, _41612,
         _41613, _41614, _41615, _41616, _41617, _41618, _41619, _41620,
         _41621, _41622, _41623, _41624, _41625, _41626, _41627, _41628,
         _41629, _41630, _41631, _41632, _41633, _41634, _41635, _41636,
         _41637, _41638, _41639, _41640, _41641, _41642, _41643, _41644,
         _41645, _41646, _41647, _41648, _41649, _41650, _41651, _41652,
         _41653, _41654, _41655, _41656, _41657, _41658, _41659, _41660,
         _41661, _41662, _41663, _41664, _41665, _41666, _41667, _41668,
         _41669, _41670, _41671, _41672, _41673, _41674, _41675, _41676,
         _41677, _41678, _41679, _41680, _41681, _41682, _41683, _41684,
         _41685, _41686, _41687, _41688, _41689, _41690, _41691, _41692,
         _41693, _41694, _41695, _41696, _41697, _41698, _41699, _41700,
         _41701, _41702, _41703, _41704, _41705, _41706, _41707, _41708,
         _41709, _41710, _41711, _41712, _41713, _41714, _41715, _41716,
         _41717, _41718, _41719, _41720, _41721, _41722, _41723, _41724,
         _41725, _41726, _41727, _41728, _41729, _41730, _41731, _41732,
         _41733, _41734, _41735, _41736, _41737, _41738, _41739, _41740,
         _41741, _41742, _41743, _41744, _41745, _41746, _41747, _41748,
         _41749, _41750, _41751, _41752, _41753, _41754, _41755, _41756,
         _41757, _41758, _41759, _41760, _41761, _41762, _41763, _41764,
         _41765, _41766, _41767, _41768, _41769, _41770, _41771, _41772,
         _41773, _41774, _41775, _41776, _41777, _41778, _41779, _41780,
         _41781, _41782, _41783, _41784, _41785, _41786, _41787, _41788,
         _41789, _41790, _41791, _41792, _41793, _41794, _41795, _41796,
         _41797, _41798, _41799, _41800, _41801, _41802, _41803, _41804,
         _41805, _41806, _41807, _41808, _41809, _41810, _41811, _41812,
         _41813, _41814, _41815, _41816, _41817, _41818, _41819, _41820,
         _41821, _41822, _41823, _41824, _41825, _41826, _41827, _41828,
         _41829, _41830, _41831, _41832, _41833, _41834, _41835, _41836,
         _41837, _41838, _41839, _41840, _41841, _41842, _41843, _41844,
         _41845, _41846, _41847, _41848, _41849, _41850, _41851, _41852,
         _41853, _41854, _41855, _41856, _41857, _41858, _41859, _41860,
         _41861, _41862, _41863, _41864, _41865, _41866, _41867, _41868,
         _41869, _41870, _41871, _41872, _41873, _41874, _41875, _41876,
         _41877, _41878, _41879, _41880, _41881, _41882, _41883, _41884,
         _41885, _41886, _41887, _41888, _41889, _41890, _41891, _41892,
         _41893, _41894, _41895, _41896, _41897, _41898, _41899, _41900,
         _41901, _41902, _41903, _41904, _41905, _41906, _41907, _41908,
         _41909, _41910, _41911, _41912, _41913, _41914, _41915, _41916,
         _41917, _41918, _41919, _41920, _41921, _41922, _41923, _41924,
         _41925, _41926, _41927, _41928, _41929, _41930, _41931, _41932,
         _41933, _41934, _41935, _41936, _41937, _41938, _41939, _41940,
         _41941, _41942, _41943, _41944, _41945, _41946, _41947, _41948,
         _41949, _41950, _41951, _41952, _41953, _41954, _41955, _41956,
         _41957, _41958, _41959, _41960, _41961, _41962, _41963, _41964,
         _41965, _41966, _41967, _41968, _41969, _41970, _41971, _41972,
         _41973, _41974, _41975, _41976, _41977, _41978, _41979, _41980,
         _41981, _41982, _41983, _41984, _41985, _41986, _41987, _41988,
         _41989, _41990, _41991, _41992, _41993, _41994, _41995, _41996,
         _41997, _41998, _41999, _42000, _42001, _42002, _42003, _42004,
         _42005, _42006, _42007, _42008, _42009, _42010, _42011, _42012,
         _42013, _42014, _42015, _42016, _42017, _42018, _42019, _42020,
         _42021, _42022, _42023, _42024, _42025, _42026, _42027, _42028,
         _42029, _42030, _42031, _42032, _42033, _42034, _42035, _42036,
         _42037, _42038, _42039, _42040, _42041, _42042, _42043, _42044,
         _42045, _42046, _42047, _42048, _42049, _42050, _42051, _42052,
         _42053, _42054, _42055, _42056, _42057, _42058, _42059, _42060,
         _42061, _42062, _42063, _42064, _42065, _42066, _42067, _42068,
         _42069, _42070, _42071, _42072, _42073, _42074, _42075, _42076,
         _42077, _42078, _42079, _42080, _42081, _42082, _42083, _42084,
         _42085, _42086, _42087, _42088, _42089, _42090, _42091, _42092,
         _42093, _42094, _42095, _42096, _42097, _42098, _42099, _42100,
         _42101, _42102, _42103, _42104, _42105, _42106, _42107, _42108,
         _42109, _42110, _42111, _42112, _42113, _42114, _42115, _42116,
         _42117, _42118, _42119, _42120, _42121, _42122, _42123, _42124,
         _42125, _42126, _42127, _42128, _42129, _42130, _42131, _42132,
         _42133, _42134, _42135, _42136, _42137, _42138, _42139, _42140,
         _42141, _42142, _42143, _42144, _42145, _42146, _42147, _42148,
         _42149, _42150, _42151, _42152, _42153, _42154, _42155, _42156,
         _42157, _42158, _42159, _42160, _42161, _42162, _42163, _42164,
         _42165, _42166, _42167, _42168, _42169, _42170, _42171, _42172,
         _42173, _42174, _42175, _42176, _42177, _42178, _42179, _42180,
         _42181, _42182, _42183, _42184, _42185, _42186, _42187, _42188,
         _42189, _42190, _42191, _42192, _42193, _42194, _42195, _42196,
         _42197, _42198, _42199, _42200, _42201, _42202, _42203, _42204,
         _42205, _42206, _42207, _42208, _42209, _42210, _42211, _42212,
         _42213, _42214, _42215, _42216, _42217, _42218, _42219, _42220,
         _42221, _42222, _42223, _42224, _42225, _42226, _42227, _42228,
         _42229, _42230, _42231, _42232, _42233, _42234, _42235, _42236,
         _42237, _42238, _42239, _42240, _42241, _42242, _42243, _42244,
         _42245, _42246, _42247, _42248, _42249, _42250, _42251, _42252,
         _42253, _42254, _42255, _42256, _42257, _42258, _42259, _42260,
         _42261, _42262, _42263, _42264, _42265, _42266, _42267, _42268,
         _42269, _42270, _42271, _42272, _42273, _42274, _42275, _42276,
         _42277, _42278, _42279, _42280, _42281, _42282, _42283, _42284,
         _42285, _42286, _42287, _42288, _42289, _42290, _42291, _42292,
         _42293, _42294, _42295, _42296, _42297, _42298, _42299, _42300,
         _42301, _42302, _42303, _42304, _42305, _42306, _42307, _42308,
         _42309, _42310, _42311, _42312, _42313, _42314, _42315, _42316,
         _42317, _42318, _42319, _42320, _42321, _42322, _42323, _42324,
         _42325, _42326, _42327, _42328, _42329, _42330, _42331, _42332,
         _42333, _42334, _42335, _42336, _42337, _42338, _42339, _42340,
         _42341, _42342, _42343, _42344, _42345, _42346, _42347, _42348,
         _42349, _42350, _42351, _42352, _42353, _42354, _42355, _42356,
         _42357, _42358, _42359, _42360, _42361, _42362, _42363, _42364,
         _42365, _42366, _42367, _42368, _42369, _42370, _42371, _42372,
         _42373, _42374, _42375, _42376, _42377, _42378, _42379, _42380,
         _42381, _42382, _42383, _42384, _42385, _42386, _42387, _42388,
         _42389, _42390, _42391, _42392, _42393, _42394, _42395, _42396,
         _42397, _42398, _42399, _42400, _42401, _42402, _42403, _42404,
         _42405, _42406, _42407, _42408, _42409, _42410, _42411, _42412,
         _42413, _42414, _42415, _42416, _42417, _42418, _42419, _42420,
         _42421, _42422, _42423, _42424, _42425, _42426, _42427, _42428,
         _42429, _42430, _42431, _42432, _42433, _42434, _42435, _42436,
         _42437, _42438, _42439, _42440, _42441, _42442, _42443, _42444,
         _42445, _42446, _42447, _42448, _42449, _42450, _42451, _42452,
         _42453, _42454, _42455, _42456, _42457, _42458, _42459, _42460,
         _42461, _42462, _42463, _42464, _42465, _42466, _42467, _42468,
         _42469, _42470, _42471, _42472, _42473, _42474, _42475, _42476,
         _42477, _42478, _42479, _42480, _42481, _42482, _42483, _42484,
         _42485, _42486, _42487, _42488, _42489, _42490, _42491, _42492,
         _42493, _42494, _42495, _42496, _42497, _42498, _42499, _42500,
         _42501, _42502, _42503, _42504, _42505, _42506, _42507, _42508,
         _42509, _42510, _42511, _42512, _42513, _42514, _42515, _42516,
         _42517, _42518, _42519, _42520, _42521, _42522, _42523, _42524,
         _42525, _42526, _42527, _42528, _42529, _42530, _42531, _42532,
         _42533, _42534, _42535, _42536, _42537, _42538, _42539, _42540,
         _42541, _42542, _42543, _42544, _42545, _42546, _42547, _42548,
         _42549, _42550, _42551, _42552, _42553, _42554, _42555, _42556,
         _42557, _42558, _42559, _42560, _42561, _42562, _42563, _42564,
         _42565, _42566, _42567, _42568, _42569, _42570, _42571, _42572,
         _42573, _42574, _42575, _42576, _42577, _42578, _42579, _42580,
         _42581, _42582, _42583, _42584, _42585, _42586, _42587, _42588,
         _42589, _42590, _42591, _42592, _42593, _42594, _42595, _42596,
         _42597, _42598, _42599, _42600, _42601, _42602, _42603, _42604,
         _42605, _42606, _42607, _42608, _42609, _42610, _42611, _42612,
         _42613, _42614, _42615, _42616, _42617, _42618, _42619, _42620,
         _42621, _42622, _42623, _42624, _42625, _42626, _42627, _42628,
         _42629, _42630, _42631, _42632, _42633, _42634, _42635, _42636,
         _42637, _42638, _42639, _42640, _42641, _42642, _42643, _42644,
         _42645, _42646, _42647, _42648, _42649, _42650, _42651, _42652,
         _42653, _42654, _42655, _42656, _42657, _42658, _42659, _42660,
         _42661, _42662, _42663, _42664, _42665, _42666, _42667, _42668,
         _42669, _42670, _42671, _42672, _42673, _42674, _42675, _42676,
         _42677, _42678, _42679, _42680, _42681, _42682, _42683, _42684,
         _42685, _42686, _42687, _42688, _42689, _42690, _42691, _42692,
         _42693, _42694, _42695, _42696, _42697, _42698, _42699, _42700,
         _42701, _42702, _42703, _42704, _42705, _42706, _42707, _42708,
         _42709, _42710, _42711, _42712, _42713, _42714, _42715, _42716,
         _42717, _42718, _42719, _42720, _42721, _42722, _42723, _42724,
         _42725, _42726, _42727, _42728, _42729, _42730, _42731, _42732,
         _42733, _42734, _42735, _42736, _42737, _42738, _42739, _42740,
         _42741, _42742, _42743, _42744, _42745, _42746, _42747, _42748,
         _42749, _42750, _42751, _42752, _42753, _42754, _42755, _42756,
         _42757, _42758, _42759, _42760, _42761, _42762, _42763, _42764,
         _42765, _42766, _42767, _42768, _42769, _42770, _42771, _42772,
         _42773, _42774, _42775, _42776, _42777, _42778, _42779, _42780,
         _42781, _42782, _42783, _42784, _42785, _42786, _42787, _42788,
         _42789, _42790, _42791, _42792, _42793, _42794, _42795, _42796,
         _42797, _42798, _42799, _42800, _42801, _42802, _42803, _42804,
         _42805, _42806, _42807, _42808, _42809, _42810, _42811, _42812,
         _42813, _42814, _42815, _42816, _42817, _42818, _42819, _42820,
         _42821, _42822, _42823, _42824, _42825, _42826, _42827, _42828,
         _42829, _42830, _42831, _42832, _42833, _42834, _42835, _42836,
         _42837, _42838, _42839, _42840, _42841, _42842, _42843, _42844,
         _42845, _42846, _42847, _42848, _42849, _42850, _42851, _42852,
         _42853, _42854, _42855, _42856, _42857, _42858, _42859, _42860,
         _42861, _42862, _42863, _42864, _42865, _42866, _42867, _42868,
         _42869, _42870, _42871, _42872, _42873, _42874, _42875, _42876,
         _42877, _42878, _42879, _42880, _42881, _42882, _42883, _42884,
         _42885, _42886, _42887, _42888, _42889, _42890, _42891, _42892,
         _42893, _42894, _42895, _42896, _42897, _42898, _42899, _42900,
         _42901, _42902, _42903, _42904, _42905, _42906, _42907, _42908,
         _42909, _42910, _42911, _42912, _42913, _42914, _42915, _42916,
         _42917, _42918, _42919, _42920, _42921, _42922, _42923, _42924,
         _42925, _42926, _42927, _42928, _42929, _42930, _42931, _42932,
         _42933, _42934, _42935, _42936, _42937, _42938, _42939, _42940,
         _42941, _42942, _42943, _42944, _42945, _42946, _42947, _42948,
         _42949, _42950, _42951, _42952, _42953, _42954, _42955, _42956,
         _42957, _42958, _42959, _42960, _42961, _42962, _42963, _42964,
         _42965, _42966, _42967, _42968, _42969, _42970, _42971, _42972,
         _42973, _42974, _42975, _42976, _42977, _42978, _42979, _42980,
         _42981, _42982, _42983, _42984, _42985, _42986, _42987, _42988,
         _42989, _42990, _42991, _42992, _42993, _42994, _42995, _42996,
         _42997, _42998, _42999, _43000, _43001, _43002, _43003, _43004,
         _43005, _43006, _43007, _43008, _43009, _43010, _43011, _43012,
         _43013, _43014, _43015, _43016, _43017, _43018, _43019, _43020,
         _43021, _43022, _43023, _43024, _43025, _43026, _43027, _43028,
         _43029, _43030, _43031, _43032, _43033, _43034, _43035, _43036,
         _43037, _43038, _43039, _43040, _43041, _43042, _43043, _43044,
         _43045, _43046, _43047, _43048, _43049, _43050, _43051, _43052,
         _43053, _43054, _43055, _43056, _43057, _43058, _43059, _43060,
         _43061, _43062, _43063, _43064, _43065, _43066, _43067, _43068,
         _43069, _43070, _43071, _43072, _43073, _43074, _43075, _43076,
         _43077, _43078, _43079, _43080, _43081, _43082, _43083, _43084,
         _43085, _43086, _43087, _43088, _43089, _43090, _43091, _43092,
         _43093, _43094, _43095, _43096, _43097, _43098, _43099, _43100,
         _43101, _43102, _43103, _43104, _43105, _43106, _43107, _43108,
         _43109, _43110, _43111, _43112, _43113, _43114, _43115, _43116,
         _43117, _43118, _43119, _43120, _43121, _43122, _43123, _43124,
         _43125, _43126, _43127, _43128, _43129, _43130, _43131, _43132,
         _43133, _43134, _43135, _43136, _43137, _43138, _43139, _43140,
         _43141, _43142, _43143, _43144, _43145, _43146, _43147, _43148,
         _43149, _43150, _43151, _43152, _43153, _43154, _43155, _43156,
         _43157, _43158, _43159, _43160, _43161, _43162, _43163, _43164,
         _43165, _43166, _43167, _43168, _43169, _43170, _43171, _43172,
         _43173, _43174, _43175, _43176, _43177, _43178, _43179, _43180,
         _43181, _43182, _43183, _43184, _43185, _43186, _43187, _43188,
         _43189, _43190, _43191, _43192, _43193, _43194, _43195, _43196,
         _43197, _43198, _43199, _43200, _43201, _43202, _43203, _43204,
         _43205, _43206, _43207, _43208, _43209, _43210, _43211, _43212,
         _43213, _43214, _43215, _43216, _43217, _43218, _43219, _43220,
         _43221, _43222, _43223, _43224, _43225, _43226, _43227, _43228,
         _43229, _43230, _43231, _43232, _43233, _43234, _43235, _43236,
         _43237, _43238, _43239, _43240, _43241, _43242, _43243, _43244,
         _43245, _43246, _43247, _43248, _43249, _43250, _43251, _43252,
         _43253, _43254, _43255, _43256, _43257, _43258, _43259, _43260,
         _43261, _43262, _43263, _43264, _43265, _43266, _43267, _43268,
         _43269, _43270, _43271, _43272, _43273, _43274, _43275, _43276,
         _43277, _43278, _43279, _43280, _43281, _43282, _43283, _43284,
         _43285, _43286, _43287, _43288, _43289, _43290, _43291, _43292,
         _43293, _43294, _43295, _43296, _43297, _43298, _43299, _43300,
         _43301, _43302, _43303, _43304, _43305, _43306, _43307, _43308,
         _43309, _43310, _43311, _43312, _43313, _43314, _43315, _43316,
         _43317, _43318, _43319, _43320, _43321, _43322, _43323, _43324,
         _43325, _43326, _43327, _43328, _43329, _43330, _43331, _43332,
         _43333, _43334, _43335, _43336, _43337, _43338, _43339, _43340,
         _43341, _43342, _43343, _43344, _43345, _43346, _43347, _43348,
         _43349, _43350, _43351, _43352, _43353, _43354, _43355, _43356,
         _43357, _43358, _43359, _43360, _43361, _43362, _43363, _43364,
         _43365, _43366, _43367, _43368, _43369, _43370, _43371, _43372,
         _43373, _43374, _43375, _43376, _43377, _43378, _43379, _43380,
         _43381, _43382, _43383, _43384, _43385, _43386, _43387, _43388,
         _43389, _43390, _43391, _43392, _43393, _43394, _43395, _43396,
         _43397, _43398, _43399, _43400, _43401, _43402, _43403, _43404,
         _43405, _43406, _43407, _43408, _43409, _43410, _43411, _43412,
         _43413, _43414, _43415, _43416, _43417, _43418, _43419, _43420,
         _43421, _43422, _43423, _43424, _43425, _43426, _43427, _43428,
         _43429, _43430, _43431, _43432, _43433, _43434, _43435, _43436,
         _43437, _43438, _43439, _43440, _43441, _43442, _43443, _43444,
         _43445, _43446, _43447, _43448, _43449, _43450, _43451, _43452,
         _43453, _43454, _43455, _43456, _43457, _43458, _43459, _43460,
         _43461, _43462, _43463, _43464, _43465, _43466, _43467, _43468,
         _43469, _43470, _43471, _43472, _43473, _43474, _43475, _43476,
         _43477, _43478, _43479, _43480, _43481, _43482, _43483, _43484,
         _43485, _43486, _43487, _43488, _43489, _43490, _43491, _43492,
         _43493, _43494, _43495, _43496, _43497, _43498, _43499, _43500,
         _43501, _43502, _43503, _43504, _43505, _43506, _43507, _43508,
         _43509, _43510, _43511, _43512, _43513, _43514, _43515, _43516,
         _43517, _43518, _43519, _43520, _43521, _43522, _43523, _43524,
         _43525, _43526, _43527, _43528, _43529, _43530, _43531, _43532,
         _43533, _43534, _43535, _43536, _43537, _43538, _43539, _43540,
         _43541, _43542, _43543, _43544, _43545, _43546, _43547, _43548,
         _43549, _43550, _43551, _43552, _43553, _43554, _43555, _43556,
         _43557, _43558, _43559, _43560, _43561, _43562, _43563, _43564,
         _43565, _43566, _43567, _43568, _43569, _43570, _43571, _43572,
         _43573, _43574, _43575, _43576, _43577, _43578, _43579, _43580,
         _43581, _43582, _43583, _43584, _43585, _43586, _43587, _43588,
         _43589, _43590, _43591, _43592, _43593, _43594, _43595, _43596,
         _43597, _43598, _43599, _43600, _43601, _43602, _43603, _43604,
         _43605, _43606, _43607, _43608, _43609, _43610, _43611, _43612,
         _43613, _43614, _43615, _43616, _43617, _43618, _43619, _43620,
         _43621, _43622, _43623, _43624, _43625, _43626, _43627, _43628,
         _43629, _43630, _43631, _43632, _43633, _43634, _43635, _43636,
         _43637, _43638, _43639, _43640, _43641, _43642, _43643, _43644,
         _43645, _43646, _43647, _43648, _43649, _43650, _43651, _43652,
         _43653, _43654, _43655, _43656, _43657, _43658, _43659, _43660,
         _43661, _43662, _43663, _43664, _43665, _43666, _43667, _43668,
         _43669, _43670, _43671, _43672, _43673, _43674, _43675, _43676,
         _43677, _43678, _43679, _43680, _43681, _43682, _43683, _43684,
         _43685, _43686, _43687, _43688, _43689, _43690, _43691, _43692,
         _43693, _43694, _43695, _43696, _43697, _43698, _43699, _43700,
         _43701, _43702, _43703, _43704, _43705, _43706, _43707, _43708,
         _43709, _43710, _43711, _43712, _43713, _43714, _43715, _43716,
         _43717, _43718, _43719, _43720, _43721, _43722, _43723, _43724,
         _43725, _43726, _43727, _43728, _43729, _43730, _43731, _43732,
         _43733, _43734, _43735, _43736, _43737, _43738, _43739, _43740,
         _43741, _43742, _43743, _43744, _43745, _43746, _43747, _43748,
         _43749, _43750, _43751, _43752, _43753, _43754, _43755, _43756,
         _43757, _43758, _43759, _43760, _43761, _43762, _43763, _43764,
         _43765, _43766, _43767, _43768, _43769, _43770, _43771, _43772,
         _43773, _43774, _43775, _43776, _43777, _43778, _43779, _43780,
         _43781, _43782, _43783, _43784, _43785, _43786, _43787, _43788,
         _43789, _43790, _43791, _43792, _43793, _43794, _43795, _43796,
         _43797, _43798, _43799, _43800, _43801, _43802, _43803, _43804,
         _43805, _43806, _43807, _43808, _43809, _43810, _43811, _43812,
         _43813, _43814, _43815, _43816, _43817, _43818, _43819, _43820,
         _43821, _43822, _43823, _43824, _43825, _43826, _43827, _43828,
         _43829, _43830, _43831, _43832, _43833, _43834, _43835, _43836,
         _43837, _43838, _43839, _43840, _43841, _43842, _43843, _43844,
         _43845, _43846, _43847, _43848, _43849, _43850, _43851, _43852,
         _43853, _43854, _43855, _43856, _43857, _43858, _43859, _43860,
         _43861, _43862, _43863, _43864, _43865, _43866, _43867, _43868,
         _43869, _43870, _43871, _43872, _43873, _43874, _43875, _43876,
         _43877, _43878, _43879, _43880, _43881, _43882, _43883, _43884,
         _43885, _43886, _43887, _43888, _43889, _43890, _43891, _43892,
         _43893, _43894, _43895, _43896, _43897, _43898, _43899, _43900,
         _43901, _43902, _43903, _43904, _43905, _43906, _43907, _43908,
         _43909, _43910, _43911, _43912, _43913, _43914, _43915, _43916,
         _43917, _43918, _43919, _43920, _43921, _43922, _43923, _43924,
         _43925, _43926, _43927, _43928, _43929, _43930, _43931, _43932,
         _43933, _43934, _43935, _43936, _43937, _43938, _43939, _43940,
         _43941, _43942, _43943, _43944, _43945, _43946, _43947, _43948,
         _43949, _43950, _43951, _43952, _43953, _43954, _43955, _43956,
         _43957, _43958, _43959, _43960, _43961, _43962, _43963, _43964,
         _43965, _43966, _43967, _43968, _43969, _43970, _43971, _43972,
         _43973, _43974, _43975, _43976, _43977, _43978, _43979, _43980,
         _43981, _43982, _43983, _43984, _43985, _43986, _43987, _43988,
         _43989, _43990, _43991, _43992, _43993, _43994, _43995, _43996,
         _43997, _43998, _43999, _44000, _44001, _44002, _44003, _44004,
         _44005, _44006, _44007, _44008, _44009, _44010, _44011, _44012,
         _44013, _44014, _44015, _44016, _44017, _44018, _44019, _44020,
         _44021, _44022, _44023, _44024, _44025, _44026, _44027, _44028,
         _44029, _44030, _44031, _44032, _44033, _44034, _44035, _44036,
         _44037, _44038, _44039, _44040, _44041, _44042, _44043, _44044,
         _44045, _44046, _44047, _44048, _44049, _44050, _44051, _44052,
         _44053, _44054, _44055, _44056, _44057, _44058, _44059, _44060,
         _44061, _44062, _44063, _44064, _44065, _44066, _44067, _44068,
         _44069, _44070, _44071, _44072, _44073, _44074, _44075, _44076,
         _44077, _44078, _44079, _44080, _44081, _44082, _44083, _44084,
         _44085, _44086, _44087, _44088, _44089, _44090, _44091, _44092,
         _44093, _44094, _44095, _44096, _44097, _44098, _44099, _44100,
         _44101, _44102, _44103, _44104, _44105, _44106, _44107, _44108,
         _44109, _44110, _44111, _44112, _44113, _44114, _44115, _44116,
         _44117, _44118, _44119, _44120, _44121, _44122, _44123, _44124,
         _44125, _44126, _44127, _44128, _44129, _44130, _44131, _44132,
         _44133, _44134, _44135, _44136, _44137, _44138, _44139, _44140,
         _44141, _44142, _44143, _44144, _44145, _44146, _44147, _44148,
         _44149, _44150, _44151, _44152, _44153, _44154, _44155, _44156,
         _44157, _44158, _44159, _44160, _44161, _44162, _44163, _44164,
         _44165, _44166, _44167, _44168, _44169, _44170, _44171, _44172,
         _44173, _44174, _44175, _44176, _44177, _44178, _44179, _44180,
         _44181, _44182, _44183, _44184, _44185, _44186, _44187, _44188,
         _44189, _44190, _44191, _44192, _44193, _44194, _44195, _44196,
         _44197, _44198, _44199, _44200, _44201, _44202, _44203, _44204,
         _44205, _44206, _44207, _44208, _44209, _44210, _44211, _44212,
         _44213, _44214, _44215, _44216, _44217, _44218, _44219, _44220,
         _44221, _44222, _44223, _44224, _44225, _44226, _44227, _44228,
         _44229, _44230, _44231, _44232, _44233, _44234, _44235, _44236,
         _44237, _44238, _44239, _44240, _44241, _44242, _44243, _44244,
         _44245, _44246, _44247, _44248, _44249, _44250, _44251, _44252,
         _44253, _44254, _44255, _44256, _44257, _44258, _44259, _44260,
         _44261, _44262, _44263, _44264, _44265, _44266, _44267, _44268,
         _44269, _44270, _44271, _44272, _44273, _44274, _44275, _44276,
         _44277, _44278, _44279, _44280, _44281, _44282, _44283, _44284,
         _44285, _44286, _44287, _44288, _44289, _44290, _44291, _44292,
         _44293, _44294, _44295, _44296, _44297, _44298, _44299, _44300,
         _44301, _44302, _44303, _44304, _44305, _44306, _44307, _44308,
         _44309, _44310, _44311, _44312, _44313, _44314, _44315, _44316,
         _44317, _44318, _44319, _44320, _44321, _44322, _44323, _44324,
         _44325, _44326, _44327, _44328, _44329, _44330, _44331, _44332,
         _44333, _44334, _44335, _44336, _44337, _44338, _44339, _44340,
         _44341, _44342, _44343, _44344, _44345, _44346, _44347, _44348,
         _44349, _44350, _44351, _44352, _44353, _44354, _44355, _44356,
         _44357, _44358, _44359, _44360, _44361, _44362, _44363, _44364,
         _44365, _44366, _44367, _44368, _44369, _44370, _44371, _44372,
         _44373, _44374, _44375, _44376, _44377, _44378, _44379, _44380,
         _44381, _44382, _44383, _44384, _44385, _44386, _44387, _44388,
         _44389, _44390, _44391, _44392, _44393, _44394, _44395, _44396,
         _44397, _44398, _44399, _44400, _44401, _44402, _44403, _44404,
         _44405, _44406, _44407, _44408, _44409, _44410, _44411, _44412,
         _44413, _44414, _44415, _44416, _44417, _44418, _44419, _44420,
         _44421, _44422, _44423, _44424, _44425, _44426, _44427, _44428,
         _44429, _44430, _44431, _44432, _44433, _44434, _44435, _44436,
         _44437, _44438, _44439, _44440, _44441, _44442, _44443, _44444,
         _44445, _44446, _44447, _44448, _44449, _44450, _44451, _44452,
         _44453, _44454, _44455, _44456, _44457, _44458, _44459, _44460,
         _44461, _44462, _44463, _44464, _44465, _44466, _44467, _44468,
         _44469, _44470, _44471, _44472, _44473, _44474, _44475, _44476,
         _44477, _44478, _44479, _44480, _44481, _44482, _44483, _44484,
         _44485, _44486, _44487, _44488, _44489, _44490, _44491, _44492,
         _44493, _44494, _44495, _44496, _44497, _44498, _44499, _44500,
         _44501, _44502, _44503, _44504, _44505, _44506, _44507, _44508,
         _44509, _44510, _44511, _44512, _44513, _44514, _44515, _44516,
         _44517, _44518, _44519, _44520, _44521, _44522, _44523, _44524,
         _44525, _44526, _44527, _44528, _44529, _44530, _44531, _44532,
         _44533, _44534, _44535, _44536, _44537, _44538, _44539, _44540,
         _44541, _44542, _44543, _44544, _44545, _44546, _44547, _44548,
         _44549, _44550, _44551, _44552, _44553, _44554, _44555, _44556,
         _44557, _44558, _44559, _44560, _44561, _44562, _44563, _44564,
         _44565, _44566, _44567, _44568, _44569, _44570, _44571, _44572,
         _44573, _44574, _44575, _44576, _44577, _44578, _44579, _44580,
         _44581, _44582, _44583, _44584, _44585, _44586, _44587, _44588,
         _44589, _44590, _44591, _44592, _44593, _44594, _44595, _44596,
         _44597, _44598, _44599, _44600, _44601, _44602, _44603, _44604,
         _44605, _44606, _44607, _44608, _44609, _44610, _44611, _44612,
         _44613, _44614, _44615, _44616, _44617, _44618, _44619, _44620,
         _44621, _44622, _44623, _44624, _44625, _44626, _44627, _44628,
         _44629, _44630, _44631, _44632, _44633, _44634, _44635, _44636,
         _44637, _44638, _44639, _44640, _44641, _44642, _44643, _44644,
         _44645, _44646, _44647, _44648, _44649, _44650, _44651, _44652,
         _44653, _44654, _44655, _44656, _44657, _44658, _44659, _44660,
         _44661, _44662, _44663, _44664, _44665, _44666, _44667, _44668,
         _44669, _44670, _44671, _44672, _44673, _44674, _44675, _44676,
         _44677, _44678, _44679, _44680, _44681, _44682, _44683, _44684,
         _44685, _44686, _44687, _44688, _44689, _44690, _44691, _44692,
         _44693, _44694, _44695, _44696, _44697, _44698, _44699, _44700,
         _44701, _44702, _44703, _44704, _44705, _44706, _44707, _44708,
         _44709, _44710, _44711, _44712, _44713, _44714, _44715, _44716,
         _44717, _44718, _44719, _44720, _44721, _44722, _44723, _44724,
         _44725, _44726, _44727, _44728, _44729, _44730, _44731, _44732,
         _44733, _44734, _44735, _44736, _44737, _44738, _44739, _44740,
         _44741, _44742, _44743, _44744, _44745, _44746, _44747, _44748,
         _44749, _44750, _44751, _44752, _44753, _44754, _44755, _44756,
         _44757, _44758, _44759, _44760, _44761, _44762, _44763, _44764,
         _44765, _44766, _44767, _44768, _44769, _44770, _44771, _44772,
         _44773, _44774, _44775, _44776, _44777, _44778, _44779, _44780,
         _44781, _44782, _44783, _44784, _44785, _44786, _44787, _44788,
         _44789, _44790, _44791, _44792, _44793, _44794, _44795, _44796,
         _44797, _44798, _44799, _44800, _44801, _44802, _44803, _44804,
         _44805, _44806, _44807, _44808, _44809, _44810, _44811, _44812,
         _44813, _44814, _44815, _44816, _44817, _44818, _44819, _44820,
         _44821, _44822, _44823, _44824, _44825, _44826, _44827, _44828,
         _44829, _44830, _44831, _44832, _44833, _44834, _44835, _44836,
         _44837, _44838, _44839, _44840, _44841, _44842, _44843, _44844,
         _44845, _44846, _44847, _44848, _44849, _44850, _44851, _44852,
         _44853, _44854, _44855, _44856, _44857, _44858, _44859, _44860,
         _44861, _44862, _44863, _44864, _44865, _44866, _44867, _44868,
         _44869, _44870, _44871, _44872, _44873, _44874, _44875, _44876,
         _44877, _44878, _44879, _44880, _44881, _44882, _44883, _44884,
         _44885, _44886, _44887, _44888, _44889, _44890, _44891, _44892,
         _44893, _44894, _44895, _44896, _44897, _44898, _44899, _44900,
         _44901, _44902, _44903, _44904, _44905, _44906, _44907, _44908,
         _44909, _44910, _44911, _44912, _44913, _44914, _44915, _44916,
         _44917, _44918, _44919, _44920, _44921, _44922, _44923, _44924,
         _44925, _44926, _44927, _44928, _44929, _44930, _44931, _44932,
         _44933, _44934, _44935, _44936, _44937, _44938, _44939, _44940,
         _44941, _44942, _44943, _44944, _44945, _44946, _44947, _44948,
         _44949, _44950, _44951, _44952, _44953, _44954, _44955, _44956,
         _44957, _44958, _44959, _44960, _44961, _44962, _44963, _44964,
         _44965, _44966, _44967, _44968, _44969, _44970, _44971, _44972,
         _44973, _44974, _44975, _44976, _44977, _44978, _44979, _44980,
         _44981, _44982, _44983, _44984, _44985, _44986, _44987, _44988,
         _44989, _44990, _44991, _44992, _44993, _44994, _44995, _44996,
         _44997, _44998, _44999, _45000, _45001, _45002, _45003, _45004,
         _45005, _45006, _45007, _45008, _45009, _45010, _45011, _45012,
         _45013, _45014, _45015, _45016, _45017, _45018, _45019, _45020,
         _45021, _45022, _45023, _45024, _45025, _45026, _45027, _45028,
         _45029, _45030, _45031, _45032, _45033, _45034, _45035, _45036,
         _45037, _45038, _45039, _45040, _45041, _45042, _45043, _45044,
         _45045, _45046, _45047, _45048, _45049, _45050, _45051, _45052,
         _45053, _45054, _45055, _45056, _45057, _45058, _45059, _45060,
         _45061, _45062, _45063, _45064, _45065, _45066, _45067, _45068,
         _45069, _45070, _45071, _45072, _45073, _45074, _45075, _45076,
         _45077, _45078, _45079, _45080, _45081, _45082, _45083, _45084,
         _45085, _45086, _45087, _45088, _45089, _45090, _45091, _45092,
         _45093, _45094, _45095, _45096, _45097, _45098, _45099, _45100,
         _45101, _45102, _45103, _45104, _45105, _45106, _45107, _45108,
         _45109, _45110, _45111, _45112, _45113, _45114, _45115, _45116,
         _45117, _45118, _45119, _45120, _45121, _45122, _45123, _45124,
         _45125, _45126, _45127, _45128, _45129, _45130, _45131, _45132,
         _45133, _45134, _45135, _45136, _45137, _45138, _45139, _45140,
         _45141, _45142, _45143, _45144, _45145, _45146, _45147, _45148,
         _45149, _45150, _45151, _45152, _45153, _45154, _45155, _45156,
         _45157, _45158, _45159, _45160, _45161, _45162, _45163, _45164,
         _45165, _45166, _45167, _45168, _45169, _45170, _45171, _45172,
         _45173, _45174, _45175, _45176, _45177, _45178, _45179, _45180,
         _45181, _45182, _45183, _45184, _45185, _45186, _45187, _45188,
         _45189, _45190, _45191, _45192, _45193, _45194, _45195, _45196,
         _45197, _45198, _45199, _45200, _45201, _45202, _45203, _45204,
         _45205, _45206, _45207, _45208, _45209, _45210, _45211, _45212,
         _45213, _45214, _45215, _45216, _45217, _45218, _45219, _45220,
         _45221, _45222, _45223, _45224, _45225, _45226, _45227, _45228,
         _45229, _45230, _45231, _45232, _45233, _45234, _45235, _45236,
         _45237, _45238, _45239, _45240, _45241, _45242, _45243, _45244,
         _45245, _45246, _45247, _45248, _45249, _45250, _45251, _45252,
         _45253, _45254, _45255, _45256, _45257, _45258, _45259, _45260,
         _45261, _45262, _45263, _45264, _45265, _45266, _45267, _45268,
         _45269, _45270, _45271, _45272, _45273, _45274, _45275, _45276,
         _45277, _45278, _45279, _45280, _45281, _45282, _45283, _45284,
         _45285, _45286, _45287, _45288, _45289, _45290, _45291, _45292,
         _45293, _45294, _45295, _45296, _45297, _45298, _45299, _45300,
         _45301, _45302, _45303, _45304, _45305, _45306, _45307, _45308,
         _45309, _45310, _45311, _45312, _45313, _45314, _45315, _45316,
         _45317, _45318, _45319, _45320, _45321, _45322, _45323, _45324,
         _45325, _45326, _45327, _45328, _45329, _45330, _45331, _45332,
         _45333, _45334, _45335, _45336, _45337, _45338, _45339, _45340,
         _45341, _45342, _45343, _45344, _45345, _45346, _45347, _45348,
         _45349, _45350, _45351, _45352, _45353, _45354, _45355, _45356,
         _45357, _45358, _45359, _45360, _45361, _45362, _45363, _45364,
         _45365, _45366, _45367, _45368, _45369, _45370, _45371, _45372,
         _45373, _45374, _45375, _45376, _45377, _45378, _45379, _45380,
         _45381, _45382, _45383, _45384, _45385, _45386, _45387, _45388,
         _45389, _45390, _45391, _45392, _45393, _45394, _45395, _45396,
         _45397, _45398, _45399, _45400, _45401, _45402, _45403, _45404,
         _45405, _45406, _45407, _45408, _45409, _45410, _45411, _45412,
         _45413, _45414, _45415, _45416, _45417, _45418, _45419, _45420,
         _45421, _45422, _45423, _45424, _45425, _45426, _45427, _45428,
         _45429, _45430, _45431, _45432, _45433, _45434, _45435, _45436,
         _45437, _45438, _45439, _45440, _45441, _45442, _45443, _45444,
         _45445, _45446, _45447, _45448, _45449, _45450, _45451, _45452,
         _45453, _45454, _45455, _45456, _45457, _45458, _45459, _45460,
         _45461, _45462, _45463, _45464, _45465, _45466, _45467, _45468,
         _45469, _45470, _45471, _45472, _45473, _45474, _45475, _45476,
         _45477, _45478, _45479, _45480, _45481, _45482, _45483, _45484,
         _45485, _45486, _45487, _45488, _45489, _45490, _45491, _45492,
         _45493, _45494, _45495, _45496, _45497, _45498, _45499, _45500,
         _45501, _45502, _45503, _45504, _45505, _45506, _45507, _45508,
         _45509, _45510, _45511, _45512, _45513, _45514, _45515, _45516,
         _45517, _45518, _45519, _45520, _45521, _45522, _45523, _45524,
         _45525, _45526, _45527, _45528, _45529, _45530, _45531, _45532,
         _45533, _45534, _45535, _45536, _45537, _45538, _45539, _45540,
         _45541, _45542, _45543, _45544, _45545, _45546, _45547, _45548,
         _45549, _45550, _45551, _45552, _45553, _45554, _45555, _45556,
         _45557, _45558, _45559, _45560, _45561, _45562, _45563, _45564,
         _45565, _45566, _45567, _45568, _45569, _45570, _45571, _45572,
         _45573, _45574, _45575, _45576, _45577, _45578, _45579, _45580,
         _45581, _45582, _45583, _45584, _45585, _45586, _45587, _45588,
         _45589, _45590, _45591, _45592, _45593, _45594, _45595, _45596,
         _45597, _45598, _45599, _45600, _45601, _45602, _45603, _45604,
         _45605, _45606, _45607, _45608, _45609, _45610, _45611, _45612,
         _45613, _45614, _45615, _45616, _45617, _45618, _45619, _45620,
         _45621, _45622, _45623, _45624, _45625, _45626, _45627, _45628,
         _45629, _45630, _45631, _45632, _45633, _45634, _45635, _45636,
         _45637, _45638, _45639, _45640, _45641, _45642, _45643, _45644,
         _45645, _45646, _45647, _45648, _45649, _45650, _45651, _45652,
         _45653, _45654, _45655, _45656, _45657, _45658, _45659, _45660,
         _45661, _45662, _45663, _45664, _45665, _45666, _45667, _45668,
         _45669, _45670, _45671, _45672, _45673, _45674, _45675, _45676,
         _45677, _45678, _45679, _45680, _45681, _45682, _45683, _45684,
         _45685, _45686, _45687, _45688, _45689, _45690, _45691, _45692,
         _45693, _45694, _45695, _45696, _45697, _45698, _45699, _45700,
         _45701, _45702, _45703, _45704, _45705, _45706, _45707, _45708,
         _45709, _45710, _45711, _45712, _45713, _45714, _45715, _45716,
         _45717, _45718, _45719, _45720, _45721, _45722, _45723, _45724,
         _45725, _45726, _45727, _45728, _45729, _45730, _45731, _45732,
         _45733, _45734, _45735, _45736, _45737, _45738, _45739, _45740,
         _45741, _45742, _45743, _45744, _45745, _45746, _45747, _45748,
         _45749, _45750, _45751, _45752, _45753, _45754, _45755, _45756,
         _45757, _45758, _45759, _45760, _45761, _45762, _45763, _45764,
         _45765, _45766, _45767, _45768, _45769, _45770, _45771, _45772,
         _45773, _45774, _45775, _45776, _45777, _45778, _45779, _45780,
         _45781, _45782, _45783, _45784, _45785, _45786, _45787, _45788,
         _45789, _45790, _45791, _45792, _45793, _45794, _45795, _45796,
         _45797, _45798, _45799, _45800, _45801, _45802, _45803, _45804,
         _45805, _45806, _45807, _45808, _45809, _45810, _45811, _45812,
         _45813, _45814, _45815, _45816, _45817, _45818, _45819, _45820,
         _45821, _45822, _45823, _45824, _45825, _45826, _45827, _45828,
         _45829, _45830, _45831, _45832, _45833, _45834, _45835, _45836,
         _45837, _45838, _45839, _45840, _45841, _45842, _45843, _45844,
         _45845, _45846, _45847, _45848, _45849, _45850, _45851, _45852,
         _45853, _45854, _45855, _45856, _45857, _45858, _45859, _45860,
         _45861, _45862, _45863, _45864, _45865, _45866, _45867, _45868,
         _45869, _45870, _45871, _45872, _45873, _45874, _45875, _45876,
         _45877, _45878, _45879, _45880, _45881, _45882, _45883, _45884,
         _45885, _45886, _45887, _45888, _45889, _45890, _45891, _45892,
         _45893, _45894, _45895, _45896, _45897, _45898, _45899, _45900,
         _45901, _45902, _45903, _45904, _45905, _45906, _45907, _45908,
         _45909, _45910, _45911, _45912, _45913, _45914, _45915, _45916,
         _45917, _45918, _45919, _45920, _45921, _45922, _45923, _45924,
         _45925, _45926, _45927, _45928, _45929, _45930, _45931, _45932,
         _45933, _45934, _45935, _45936, _45937, _45938, _45939, _45940,
         _45941, _45942, _45943, _45944, _45945, _45946, _45947, _45948,
         _45949, _45950, _45951, _45952, _45953, _45954, _45955, _45956,
         _45957, _45958, _45959, _45960, _45961, _45962, _45963, _45964,
         _45965, _45966, _45967, _45968, _45969, _45970, _45971, _45972,
         _45973, _45974, _45975, _45976, _45977, _45978, _45979, _45980,
         _45981, _45982, _45983, _45984, _45985, _45986, _45987, _45988,
         _45989, _45990, _45991, _45992, _45993, _45994, _45995, _45996,
         _45997, _45998, _45999, _46000, _46001, _46002, _46003, _46004,
         _46005, _46006, _46007, _46008, _46009, _46010, _46011, _46012,
         _46013, _46014, _46015, _46016, _46017, _46018, _46019, _46020,
         _46021, _46022, _46023, _46024, _46025, _46026, _46027, _46028,
         _46029, _46030, _46031, _46032, _46033, _46034, _46035, _46036,
         _46037, _46038, _46039, _46040, _46041, _46042, _46043, _46044,
         _46045, _46046, _46047, _46048, _46049, _46050, _46051, _46052,
         _46053, _46054, _46055, _46056, _46057, _46058, _46059, _46060,
         _46061, _46062, _46063, _46064, _46065, _46066, _46067, _46068,
         _46069, _46070, _46071, _46072, _46073, _46074, _46075, _46076,
         _46077, _46078, _46079, _46080, _46081, _46082, _46083, _46084,
         _46085, _46086, _46087, _46088, _46089, _46090, _46091, _46092,
         _46093, _46094, _46095, _46096, _46097, _46098, _46099, _46100,
         _46101, _46102, _46103, _46104, _46105, _46106, _46107, _46108,
         _46109, _46110, _46111, _46112, _46113, _46114, _46115, _46116,
         _46117, _46118, _46119, _46120, _46121, _46122, _46123, _46124,
         _46125, _46126, _46127, _46128, _46129, _46130, _46131, _46132,
         _46133, _46134, _46135, _46136, _46137, _46138, _46139, _46140,
         _46141, _46142, _46143, _46144, _46145, _46146, _46147, _46148,
         _46149, _46150, _46151, _46152, _46153, _46154, _46155, _46156,
         _46157, _46158, _46159, _46160, _46161, _46162, _46163, _46164,
         _46165, _46166, _46167, _46168, _46169, _46170, _46171, _46172,
         _46173, _46174, _46175, _46176, _46177, _46178, _46179, _46180,
         _46181, _46182, _46183, _46184, _46185, _46186, _46187, _46188,
         _46189, _46190, _46191, _46192, _46193, _46194, _46195, _46196,
         _46197, _46198, _46199, _46200, _46201, _46202, _46203, _46204,
         _46205, _46206, _46207, _46208, _46209, _46210, _46211, _46212,
         _46213, _46214, _46215, _46216, _46217, _46218, _46219, _46220,
         _46221, _46222, _46223, _46224, _46225, _46226, _46227, _46228,
         _46229, _46230, _46231, _46232, _46233, _46234, _46235, _46236,
         _46237, _46238, _46239, _46240, _46241, _46242, _46243, _46244,
         _46245, _46246, _46247, _46248, _46249, _46250, _46251, _46252,
         _46253, _46254, _46255, _46256, _46257, _46258, _46259, _46260,
         _46261, _46262, _46263, _46264, _46265, _46266, _46267, _46268,
         _46269, _46270, _46271, _46272, _46273, _46274, _46275, _46276,
         _46277, _46278, _46279, _46280, _46281, _46282, _46283, _46284,
         _46285, _46286, _46287, _46288, _46289, _46290, _46291, _46292,
         _46293, _46294, _46295, _46296, _46297, _46298, _46299, _46300,
         _46301, _46302, _46303, _46304, _46305, _46306, _46307, _46308,
         _46309, _46310, _46311, _46312, _46313, _46314, _46315, _46316,
         _46317, _46318, _46319, _46320, _46321, _46322, _46323, _46324,
         _46325, _46326, _46327, _46328, _46329, _46330, _46331, _46332,
         _46333, _46334, _46335, _46336, _46337, _46338, _46339, _46340,
         _46341, _46342, _46343, _46344, _46345, _46346, _46347, _46348,
         _46349, _46350, _46351, _46352, _46353, _46354, _46355, _46356,
         _46357, _46358, _46359, _46360, _46361, _46362, _46363, _46364,
         _46365, _46366, _46367, _46368, _46369, _46370, _46371, _46372,
         _46373, _46374, _46375, _46376, _46377, _46378, _46379, _46380,
         _46381, _46382, _46383, _46384, _46385, _46386, _46387, _46388,
         _46389, _46390, _46391, _46392, _46393, _46394, _46395, _46396,
         _46397, _46398, _46399, _46400, _46401, _46402, _46403, _46404,
         _46405, _46406, _46407, _46408, _46409, _46410, _46411, _46412,
         _46413, _46414, _46415, _46416, _46417, _46418, _46419, _46420,
         _46421, _46422, _46423, _46424, _46425, _46426, _46427, _46428,
         _46429, _46430, _46431, _46432, _46433, _46434, _46435, _46436,
         _46437, _46438, _46439, _46440, _46441, _46442, _46443, _46444,
         _46445, _46446, _46447, _46448, _46449, _46450, _46451, _46452,
         _46453, _46454, _46455, _46456, _46457, _46458, _46459, _46460,
         _46461, _46462, _46463, _46464, _46465, _46466, _46467, _46468,
         _46469, _46470, _46471, _46472, _46473, _46474, _46475, _46476,
         _46477, _46478, _46479, _46480, _46481, _46482, _46483, _46484,
         _46485, _46486, _46487, _46488, _46489, _46490, _46491, _46492,
         _46493, _46494, _46495, _46496, _46497, _46498, _46499, _46500,
         _46501, _46502, _46503, _46504, _46505, _46506, _46507, _46508,
         _46509, _46510, _46511, _46512, _46513, _46514, _46515, _46516,
         _46517, _46518, _46519, _46520, _46521, _46522, _46523, _46524,
         _46525, _46526, _46527, _46528, _46529, _46530, _46531, _46532,
         _46533, _46534, _46535, _46536, _46537, _46538, _46539, _46540,
         _46541, _46542, _46543, _46544, _46545, _46546, _46547, _46548,
         _46549, _46550, _46551, _46552, _46553, _46554, _46555, _46556,
         _46557, _46558, _46559, _46560, _46561, _46562, _46563, _46564,
         _46565, _46566, _46567, _46568, _46569, _46570, _46571, _46572,
         _46573, _46574, _46575, _46576, _46577, _46578, _46579, _46580,
         _46581, _46582, _46583, _46584, _46585, _46586, _46587, _46588,
         _46589, _46590, _46591, _46592, _46593, _46594, _46595, _46596,
         _46597, _46598, _46599, _46600, _46601, _46602, _46603, _46604,
         _46605, _46606, _46607, _46608, _46609, _46610, _46611, _46612,
         _46613, _46614, _46615, _46616, _46617, _46618, _46619, _46620,
         _46621, _46622, _46623, _46624, _46625, _46626, _46627, _46628,
         _46629, _46630, _46631, _46632, _46633, _46634, _46635, _46636,
         _46637, _46638, _46639, _46640, _46641, _46642, _46643, _46644,
         _46645, _46646, _46647, _46648, _46649, _46650, _46651, _46652,
         _46653, _46654, _46655, _46656, _46657, _46658, _46659, _46660,
         _46661, _46662, _46663, _46664, _46665, _46666, _46667, _46668,
         _46669, _46670, _46671, _46672, _46673, _46674, _46675, _46676,
         _46677, _46678, _46679, _46680, _46681, _46682, _46683, _46684,
         _46685, _46686, _46687, _46688, _46689, _46690, _46691, _46692,
         _46693, _46694, _46695, _46696, _46697, _46698, _46699, _46700,
         _46701, _46702, _46703, _46704, _46705, _46706, _46707, _46708,
         _46709, _46710, _46711, _46712, _46713, _46714, _46715, _46716,
         _46717, _46718, _46719, _46720, _46721, _46722, _46723, _46724,
         _46725, _46726, _46727, _46728, _46729, _46730, _46731, _46732,
         _46733, _46734, _46735, _46736, _46737, _46738, _46739, _46740,
         _46741, _46742, _46743, _46744, _46745, _46746, _46747, _46748,
         _46749, _46750, _46751, _46752, _46753, _46754, _46755, _46756,
         _46757, _46758, _46759, _46760, _46761, _46762, _46763, _46764,
         _46765, _46766, _46767, _46768, _46769, _46770, _46771, _46772,
         _46773, _46774, _46775, _46776, _46777, _46778, _46779, _46780,
         _46781, _46782, _46783, _46784, _46785, _46786, _46787, _46788,
         _46789, _46790, _46791, _46792, _46793, _46794, _46795, _46796,
         _46797, _46798, _46799, _46800, _46801, _46802, _46803, _46804,
         _46805, _46806, _46807, _46808, _46809, _46810, _46811, _46812,
         _46813, _46814, _46815, _46816, _46817, _46818, _46819, _46820,
         _46821, _46822, _46823, _46824, _46825, _46826, _46827, _46828,
         _46829, _46830, _46831, _46832, _46833, _46834, _46835, _46836,
         _46837, _46838, _46839, _46840, _46841, _46842, _46843, _46844,
         _46845, _46846, _46847, _46848, _46849, _46850, _46851, _46852,
         _46853, _46854, _46855, _46856, _46857, _46858, _46859, _46860,
         _46861, _46862, _46863, _46864, _46865, _46866, _46867, _46868,
         _46869, _46870, _46871, _46872, _46873, _46874, _46875, _46876,
         _46877, _46878, _46879, _46880, _46881, _46882, _46883, _46884,
         _46885, _46886, _46887, _46888, _46889, _46890, _46891, _46892,
         _46893, _46894, _46895, _46896, _46897, _46898, _46899, _46900,
         _46901, _46902, _46903, _46904, _46905, _46906, _46907, _46908,
         _46909, _46910, _46911, _46912, _46913, _46914, _46915, _46916,
         _46917, _46918, _46919, _46920, _46921, _46922, _46923, _46924,
         _46925, _46926, _46927, _46928, _46929, _46930, _46931, _46932,
         _46933, _46934, _46935, _46936, _46937, _46938, _46939, _46940,
         _46941, _46942, _46943, _46944, _46945, _46946, _46947, _46948,
         _46949, _46950, _46951, _46952, _46953, _46954, _46955, _46956,
         _46957, _46958, _46959, _46960, _46961, _46962, _46963, _46964,
         _46965, _46966, _46967, _46968, _46969, _46970, _46971, _46972,
         _46973, _46974, _46975, _46976, _46977, _46978, _46979, _46980,
         _46981, _46982, _46983, _46984, _46985, _46986, _46987, _46988,
         _46989, _46990, _46991, _46992, _46993, _46994, _46995, _46996,
         _46997, _46998, _46999, _47000, _47001, _47002, _47003, _47004,
         _47005, _47006, _47007, _47008, _47009, _47010, _47011, _47012,
         _47013, _47014, _47015, _47016, _47017, _47018, _47019, _47020,
         _47021, _47022, _47023, _47024, _47025, _47026, _47027, _47028,
         _47029, _47030, _47031, _47032, _47033, _47034, _47035, _47036,
         _47037, _47038, _47039, _47040, _47041, _47042, _47043, _47044,
         _47045, _47046, _47047, _47048, _47049, _47050, _47051, _47052,
         _47053, _47054, _47055, _47056, _47057, _47058, _47059, _47060,
         _47061, _47062, _47063, _47064, _47065, _47066, _47067, _47068,
         _47069, _47070, _47071, _47072, _47073, _47074, _47075, _47076,
         _47077, _47078, _47079, _47080, _47081, _47082, _47083, _47084,
         _47085, _47086, _47087, _47088, _47089, _47090, _47091, _47092,
         _47093, _47094, _47095, _47096, _47097, _47098, _47099, _47100,
         _47101, _47102, _47103, _47104, _47105, _47106, _47107, _47108,
         _47109, _47110, _47111, _47112, _47113, _47114, _47115, _47116,
         _47117, _47118, _47119, _47120, _47121, _47122, _47123, _47124,
         _47125, _47126, _47127, _47128, _47129, _47130, _47131, _47132,
         _47133, _47134, _47135, _47136, _47137, _47138, _47139, _47140,
         _47141, _47142, _47143, _47144, _47145, _47146, _47147, _47148,
         _47149, _47150, _47151, _47152, _47153, _47154, _47155, _47156,
         _47157, _47158, _47159, _47160, _47161, _47162, _47163, _47164,
         _47165, _47166, _47167, _47168, _47169, _47170, _47171, _47172,
         _47173, _47174, _47175, _47176, _47177, _47178, _47179, _47180,
         _47181, _47182, _47183, _47184, _47185, _47186, _47187, _47188,
         _47189, _47190, _47191, _47192, _47193, _47194, _47195, _47196,
         _47197, _47198, _47199, _47200, _47201, _47202, _47203, _47204,
         _47205, _47206, _47207, _47208, _47209, _47210, _47211, _47212,
         _47213, _47214, _47215, _47216, _47217, _47218, _47219, _47220,
         _47221, _47222, _47223, _47224, _47225, _47226, _47227, _47228,
         _47229, _47230, _47231, _47232, _47233, _47234, _47235, _47236,
         _47237, _47238, _47239, _47240, _47241, _47242, _47243, _47244,
         _47245, _47246, _47247, _47248, _47249, _47250, _47251, _47252,
         _47253, _47254, _47255, _47256, _47257, _47258, _47259, _47260,
         _47261, _47262, _47263, _47264, _47265, _47266, _47267, _47268,
         _47269, _47270, _47271, _47272, _47273, _47274, _47275, _47276,
         _47277, _47278, _47279, _47280, _47281, _47282, _47283, _47284,
         _47285, _47286, _47287, _47288, _47289, _47290, _47291, _47292,
         _47293, _47294, _47295, _47296, _47297, _47298, _47299, _47300,
         _47301, _47302, _47303, _47304, _47305, _47306, _47307, _47308,
         _47309, _47310, _47311, _47312, _47313, _47314, _47315, _47316,
         _47317, _47318, _47319, _47320, _47321, _47322, _47323, _47324,
         _47325, _47326, _47327, _47328, _47329, _47330, _47331, _47332,
         _47333, _47334, _47335, _47336, _47337, _47338, _47339, _47340,
         _47341, _47342, _47343, _47344, _47345, _47346, _47347, _47348,
         _47349, _47350, _47351, _47352, _47353, _47354, _47355, _47356,
         _47357, _47358, _47359, _47360, _47361, _47362, _47363, _47364,
         _47365, _47366, _47367, _47368, _47369, _47370, _47371, _47372,
         _47373, _47374, _47375, _47376, _47377, _47378, _47379, _47380,
         _47381, _47382, _47383, _47384, _47385, _47386, _47387, _47388,
         _47389, _47390, _47391, _47392, _47393, _47394, _47395, _47396,
         _47397, _47398, _47399, _47400, _47401, _47402, _47403, _47404,
         _47405, _47406, _47407, _47408, _47409, _47410, _47411, _47412,
         _47413, _47414, _47415, _47416, _47417, _47418, _47419, _47420,
         _47421, _47422, _47423, _47424, _47425, _47426, _47427, _47428,
         _47429, _47430, _47431, _47432, _47433, _47434, _47435, _47436,
         _47437, _47438, _47439, _47440, _47441, _47442, _47443, _47444,
         _47445, _47446, _47447, _47448, _47449, _47450, _47451, _47452,
         _47453, _47454, _47455, _47456, _47457, _47458, _47459, _47460,
         _47461, _47462, _47463, _47464, _47465, _47466, _47467, _47468,
         _47469, _47470, _47471, _47472, _47473, _47474, _47475, _47476,
         _47477, _47478, _47479, _47480, _47481, _47482, _47483, _47484,
         _47485, _47486, _47487, _47488, _47489, _47490, _47491, _47492,
         _47493, _47494, _47495, _47496, _47497, _47498, _47499, _47500,
         _47501, _47502, _47503, _47504, _47505, _47506, _47507, _47508,
         _47509, _47510, _47511, _47512, _47513, _47514, _47515, _47516,
         _47517, _47518, _47519, _47520, _47521, _47522, _47523, _47524,
         _47525, _47526, _47527, _47528, _47529, _47530, _47531, _47532,
         _47533, _47534, _47535, _47536, _47537, _47538, _47539, _47540,
         _47541, _47542, _47543, _47544, _47545, _47546, _47547, _47548,
         _47549, _47550, _47551, _47552, _47553, _47554, _47555, _47556,
         _47557, _47558, _47559, _47560, _47561, _47562, _47563, _47564,
         _47565, _47566, _47567, _47568, _47569, _47570, _47571, _47572,
         _47573, _47574, _47575, _47576, _47577, _47578, _47579, _47580,
         _47581, _47582, _47583, _47584, _47585, _47586, _47587, _47588,
         _47589, _47590, _47591, _47592, _47593, _47594, _47595, _47596,
         _47597, _47598, _47599, _47600, _47601, _47602, _47603, _47604,
         _47605, _47606, _47607, _47608, _47609, _47610, _47611, _47612,
         _47613, _47614, _47615, _47616, _47617, _47618, _47619, _47620,
         _47621, _47622, _47623, _47624, _47625, _47626, _47627, _47628,
         _47629, _47630, _47631, _47632, _47633, _47634, _47635, _47636,
         _47637, _47638, _47639, _47640, _47641, _47642, _47643, _47644,
         _47645, _47646, _47647, _47648, _47649, _47650, _47651, _47652,
         _47653, _47654, _47655, _47656, _47657, _47658, _47659, _47660,
         _47661, _47662, _47663, _47664, _47665, _47666, _47667, _47668,
         _47669, _47670, _47671, _47672, _47673, _47674, _47675, _47676,
         _47677, _47678, _47679, _47680, _47681, _47682, _47683, _47684,
         _47685, _47686, _47687, _47688, _47689, _47690, _47691, _47692,
         _47693, _47694, _47695, _47696, _47697, _47698, _47699, _47700,
         _47701, _47702, _47703, _47704, _47705, _47706, _47707, _47708,
         _47709, _47710, _47711, _47712, _47713, _47714, _47715, _47716,
         _47717, _47718, _47719, _47720, _47721, _47722, _47723, _47724,
         _47725, _47726, _47727, _47728, _47729, _47730, _47731, _47732,
         _47733, _47734, _47735, _47736, _47737, _47738, _47739, _47740,
         _47741, _47742, _47743, _47744, _47745, _47746, _47747, _47748,
         _47749, _47750, _47751, _47752, _47753, _47754, _47755, _47756,
         _47757, _47758, _47759, _47760, _47761, _47762, _47763, _47764,
         _47765, _47766, _47767, _47768, _47769, _47770, _47771, _47772,
         _47773, _47774, _47775, _47776, _47777, _47778, _47779, _47780,
         _47781, _47782, _47783, _47784, _47785, _47786, _47787, _47788,
         _47789, _47790, _47791, _47792, _47793, _47794, _47795, _47796,
         _47797, _47798, _47799, _47800, _47801, _47802, _47803, _47804,
         _47805, _47806, _47807, _47808, _47809, _47810, _47811, _47812,
         _47813, _47814, _47815, _47816, _47817, _47818, _47819, _47820,
         _47821, _47822, _47823, _47824, _47825, _47826, _47827, _47828,
         _47829, _47830, _47831, _47832, _47833, _47834, _47835, _47836,
         _47837, _47838, _47839, _47840, _47841, _47842, _47843, _47844,
         _47845, _47846, _47847, _47848, _47849, _47850, _47851, _47852,
         _47853, _47854, _47855, _47856, _47857, _47858, _47859, _47860,
         _47861, _47862, _47863, _47864, _47865, _47866, _47867, _47868,
         _47869, _47870, _47871, _47872, _47873, _47874, _47875, _47876,
         _47877, _47878, _47879, _47880, _47881, _47882, _47883, _47884,
         _47885, _47886, _47887, _47888, _47889, _47890, _47891, _47892,
         _47893, _47894, _47895, _47896, _47897, _47898, _47899, _47900,
         _47901, _47902, _47903, _47904, _47905, _47906, _47907, _47908,
         _47909, _47910, _47911, _47912, _47913, _47914, _47915, _47916,
         _47917, _47918, _47919, _47920, _47921, _47922, _47923, _47924,
         _47925, _47926, _47927, _47928, _47929, _47930, _47931, _47932,
         _47933, _47934, _47935, _47936, _47937, _47938, _47939, _47940,
         _47941, _47942, _47943, _47944, _47945, _47946, _47947, _47948,
         _47949, _47950, _47951, _47952, _47953, _47954, _47955, _47956,
         _47957, _47958, _47959, _47960, _47961, _47962, _47963, _47964,
         _47965, _47966, _47967, _47968, _47969, _47970, _47971, _47972,
         _47973, _47974, _47975, _47976, _47977, _47978, _47979, _47980,
         _47981, _47982, _47983, _47984, _47985, _47986, _47987, _47988,
         _47989, _47990, _47991, _47992, _47993, _47994, _47995, _47996,
         _47997, _47998, _47999, _48000, _48001, _48002, _48003, _48004,
         _48005, _48006, _48007, _48008, _48009, _48010, _48011, _48012,
         _48013, _48014, _48015, _48016, _48017, _48018, _48019, _48020,
         _48021, _48022, _48023, _48024, _48025, _48026, _48027, _48028,
         _48029, _48030, _48031, _48032, _48033, _48034, _48035, _48036,
         _48037, _48038, _48039, _48040, _48041, _48042, _48043, _48044,
         _48045, _48046, _48047, _48048, _48049, _48050, _48051, _48052,
         _48053, _48054, _48055, _48056, _48057, _48058, _48059, _48060,
         _48061, _48062, _48063, _48064, _48065, _48066, _48067, _48068,
         _48069, _48070, _48071, _48072, _48073, _48074, _48075, _48076,
         _48077, _48078, _48079, _48080, _48081, _48082, _48083, _48084,
         _48085, _48086, _48087, _48088, _48089, _48090, _48091, _48092,
         _48093, _48094, _48095, _48096, _48097, _48098, _48099, _48100,
         _48101, _48102, _48103, _48104, _48105, _48106, _48107, _48108,
         _48109, _48110, _48111, _48112, _48113, _48114, _48115, _48116,
         _48117, _48118, _48119, _48120, _48121, _48122, _48123, _48124,
         _48125, _48126, _48127, _48128, _48129, _48130, _48131, _48132,
         _48133, _48134, _48135, _48136, _48137, _48138, _48139, _48140,
         _48141, _48142, _48143, _48144, _48145, _48146, _48147, _48148,
         _48149, _48150, _48151, _48152, _48153, _48154, _48155, _48156,
         _48157, _48158, _48159, _48160, _48161, _48162, _48163, _48164,
         _48165, _48166, _48167, _48168, _48169, _48170, _48171, _48172,
         _48173, _48174, _48175, _48176, _48177, _48178, _48179, _48180,
         _48181, _48182, _48183, _48184, _48185, _48186, _48187, _48188,
         _48189, _48190, _48191, _48192, _48193, _48194, _48195, _48196,
         _48197, _48198, _48199, _48200, _48201, _48202, _48203, _48204,
         _48205, _48206, _48207, _48208, _48209, _48210, _48211, _48212,
         _48213, _48214, _48215, _48216, _48217, _48218, _48219, _48220,
         _48221, _48222, _48223, _48224, _48225, _48226, _48227, _48228,
         _48229, _48230, _48231, _48232, _48233, _48234, _48235, _48236,
         _48237, _48238, _48239, _48240, _48241, _48242, _48243, _48244,
         _48245, _48246, _48247, _48248, _48249, _48250, _48251, _48252,
         _48253, _48254, _48255, _48256, _48257, _48258, _48259, _48260,
         _48261, _48262, _48263, _48264, _48265, _48266, _48267, _48268,
         _48269, _48270, _48271, _48272, _48273, _48274, _48275, _48276,
         _48277, _48278, _48279, _48280, _48281, _48282, _48283, _48284,
         _48285, _48286, _48287, _48288, _48289, _48290, _48291, _48292,
         _48293, _48294, _48295, _48296, _48297, _48298, _48299, _48300,
         _48301, _48302, _48303, _48304, _48305, _48306, _48307, _48308,
         _48309, _48310, _48311, _48312, _48313, _48314, _48315, _48316,
         _48317, _48318, _48319, _48320, _48321, _48322, _48323, _48324,
         _48325, _48326, _48327, _48328, _48329, _48330, _48331, _48332,
         _48333, _48334, _48335, _48336, _48337, _48338, _48339, _48340,
         _48341, _48342, _48343, _48344, _48345, _48346, _48347, _48348,
         _48349, _48350, _48351, _48352, _48353, _48354, _48355, _48356,
         _48357, _48358, _48359, _48360, _48361, _48362, _48363, _48364,
         _48365, _48366, _48367, _48368, _48369, _48370, _48371, _48372,
         _48373, _48374, _48375, _48376, _48377, _48378, _48379, _48380,
         _48381, _48382, _48383, _48384, _48385, _48386, _48387, _48388,
         _48389, _48390, _48391, _48392, _48393, _48394, _48395, _48396,
         _48397, _48398, _48399, _48400, _48401, _48402, _48403, _48404,
         _48405, _48406, _48407, _48408, _48409, _48410, _48411, _48412,
         _48413, _48414, _48415, _48416, _48417, _48418, _48419, _48420,
         _48421, _48422, _48423, _48424, _48425, _48426, _48427, _48428,
         _48429, _48430, _48431, _48432, _48433, _48434, _48435, _48436,
         _48437, _48438, _48439, _48440, _48441, _48442, _48443, _48444,
         _48445, _48446, _48447, _48448, _48449, _48450, _48451, _48452,
         _48453, _48454, _48455, _48456, _48457, _48458, _48459, _48460,
         _48461, _48462, _48463, _48464, _48465, _48466, _48467, _48468,
         _48469, _48470, _48471, _48472, _48473, _48474, _48475, _48476,
         _48477, _48478, _48479, _48480, _48481, _48482, _48483, _48484,
         _48485, _48486, _48487, _48488, _48489, _48490, _48491, _48492,
         _48493, _48494, _48495, _48496, _48497, _48498, _48499, _48500,
         _48501, _48502, _48503, _48504, _48505, _48506, _48507, _48508,
         _48509, _48510, _48511, _48512, _48513, _48514, _48515, _48516,
         _48517, _48518, _48519, _48520, _48521, _48522, _48523, _48524,
         _48525, _48526, _48527, _48528, _48529, _48530, _48531, _48532,
         _48533, _48534, _48535, _48536, _48537, _48538, _48539, _48540,
         _48541, _48542, _48543, _48544, _48545, _48546, _48547, _48548,
         _48549, _48550, _48551, _48552, _48553, _48554, _48555, _48556,
         _48557, _48558, _48559, _48560, _48561, _48562, _48563, _48564,
         _48565, _48566, _48567, _48568, _48569, _48570, _48571, _48572,
         _48573, _48574, _48575, _48576, _48577, _48578, _48579, _48580,
         _48581, _48582, _48583, _48584, _48585, _48586, _48587, _48588,
         _48589, _48590, _48591, _48592, _48593, _48594, _48595, _48596,
         _48597, _48598, _48599, _48600, _48601, _48602, _48603, _48604,
         _48605, _48606, _48607, _48608, _48609, _48610, _48611, _48612,
         _48613, _48614, _48615, _48616, _48617, _48618, _48619, _48620,
         _48621, _48622, _48623, _48624, _48625, _48626, _48627, _48628,
         _48629, _48630, _48631, _48632, _48633, _48634, _48635, _48636,
         _48637, _48638, _48639, _48640, _48641, _48642, _48643, _48644,
         _48645, _48646, _48647, _48648, _48649, _48650, _48651, _48652,
         _48653, _48654, _48655, _48656, _48657, _48658, _48659, _48660,
         _48661, _48662, _48663, _48664, _48665, _48666, _48667, _48668,
         _48669, _48670, _48671, _48672, _48673, _48674, _48675, _48676,
         _48677, _48678, _48679, _48680, _48681, _48682, _48683, _48684,
         _48685, _48686, _48687, _48688, _48689, _48690, _48691, _48692,
         _48693, _48694, _48695, _48696, _48697, _48698, _48699, _48700,
         _48701, _48702, _48703, _48704, _48705, _48706, _48707, _48708,
         _48709, _48710, _48711, _48712, _48713, _48714, _48715, _48716,
         _48717, _48718, _48719, _48720, _48721, _48722, _48723, _48724,
         _48725, _48726, _48727, _48728, _48729, _48730, _48731, _48732,
         _48733, _48734, _48735, _48736, _48737, _48738, _48739, _48740,
         _48741, _48742, _48743, _48744, _48745, _48746, _48747, _48748,
         _48749, _48750, _48751, _48752, _48753, _48754, _48755, _48756,
         _48757, _48758, _48759, _48760, _48761, _48762, _48763, _48764,
         _48765, _48766, _48767, _48768, _48769, _48770, _48771, _48772,
         _48773, _48774, _48775, _48776, _48777, _48778, _48779, _48780,
         _48781, _48782, _48783, _48784, _48785, _48786, _48787, _48788,
         _48789, _48790, _48791, _48792, _48793, _48794, _48795, _48796,
         _48797, _48798, _48799, _48800, _48801, _48802, _48803, _48804,
         _48805, _48806, _48807, _48808, _48809, _48810, _48811, _48812,
         _48813, _48814, _48815, _48816, _48817, _48818, _48819, _48820,
         _48821, _48822, _48823, _48824, _48825, _48826, _48827, _48828,
         _48829, _48830, _48831, _48832, _48833, _48834, _48835, _48836,
         _48837, _48838, _48839, _48840, _48841, _48842, _48843, _48844,
         _48845, _48846, _48847, _48848, _48849, _48850, _48851, _48852,
         _48853, _48854, _48855, _48856, _48857, _48858, _48859, _48860,
         _48861, _48862, _48863, _48864, _48865, _48866, _48867, _48868,
         _48869, _48870, _48871, _48872, _48873, _48874, _48875, _48876,
         _48877, _48878, _48879, _48880, _48881, _48882, _48883, _48884,
         _48885, _48886, _48887, _48888, _48889, _48890, _48891, _48892,
         _48893, _48894, _48895, _48896, _48897, _48898, _48899, _48900,
         _48901, _48902, _48903, _48904, _48905, _48906, _48907, _48908,
         _48909, _48910, _48911, _48912, _48913, _48914, _48915, _48916,
         _48917, _48918, _48919, _48920, _48921, _48922, _48923, _48924,
         _48925, _48926, _48927, _48928, _48929, _48930, _48931, _48932,
         _48933, _48934, _48935, _48936, _48937, _48938, _48939, _48940,
         _48941, _48942, _48943, _48944, _48945, _48946, _48947, _48948,
         _48949, _48950, _48951, _48952, _48953, _48954, _48955, _48956,
         _48957, _48958, _48959, _48960, _48961, _48962, _48963, _48964,
         _48965, _48966, _48967, _48968, _48969, _48970, _48971, _48972,
         _48973, _48974, _48975, _48976, _48977, _48978, _48979, _48980,
         _48981, _48982, _48983, _48984, _48985, _48986, _48987, _48988,
         _48989, _48990, _48991, _48992, _48993, _48994, _48995, _48996,
         _48997, _48998, _48999, _49000, _49001, _49002, _49003, _49004,
         _49005, _49006, _49007, _49008, _49009, _49010, _49011, _49012,
         _49013, _49014, _49015, _49016, _49017, _49018, _49019, _49020,
         _49021, _49022, _49023, _49024, _49025, _49026, _49027, _49028,
         _49029, _49030, _49031, _49032, _49033, _49034, _49035, _49036,
         _49037, _49038, _49039, _49040, _49041, _49042, _49043, _49044,
         _49045, _49046, _49047, _49048, _49049, _49050, _49051, _49052,
         _49053, _49054, _49055, _49056, _49057, _49058, _49059, _49060,
         _49061, _49062, _49063, _49064, _49065, _49066, _49067, _49068,
         _49069, _49070, _49071, _49072, _49073, _49074, _49075, _49076,
         _49077, _49078, _49079, _49080, _49081, _49082, _49083, _49084,
         _49085, _49086, _49087, _49088, _49089, _49090, _49091, _49092,
         _49093, _49094, _49095, _49096, _49097, _49098, _49099, _49100,
         _49101, _49102, _49103, _49104, _49105, _49106, _49107, _49108,
         _49109, _49110, _49111, _49112, _49113, _49114, _49115, _49116,
         _49117, _49118, _49119, _49120, _49121, _49122, _49123, _49124,
         _49125, _49126, _49127, _49128, _49129, _49130, _49131, _49132,
         _49133, _49134, _49135, _49136, _49137, _49138, _49139, _49140,
         _49141, _49142, _49143, _49144, _49145, _49146, _49147, _49148,
         _49149, _49150, _49151, _49152, _49153, _49154, _49155, _49156,
         _49157, _49158, _49159, _49160, _49161, _49162, _49163, _49164,
         _49165, _49166, _49167, _49168, _49169, _49170, _49171, _49172,
         _49173, _49174, _49175, _49176, _49177, _49178, _49179, _49180,
         _49181, _49182, _49183, _49184, _49185, _49186, _49187, _49188,
         _49189, _49190, _49191, _49192, _49193, _49194, _49195, _49196,
         _49197, _49198, _49199, _49200, _49201, _49202, _49203, _49204,
         _49205, _49206, _49207, _49208, _49209, _49210, _49211, _49212,
         _49213, _49214, _49215, _49216, _49217, _49218, _49219, _49220,
         _49221, _49222, _49223, _49224, _49225, _49226, _49227, _49228,
         _49229, _49230, _49231, _49232, _49233, _49234, _49235, _49236,
         _49237, _49238, _49239, _49240, _49241, _49242, _49243, _49244,
         _49245, _49246, _49247, _49248, _49249, _49250, _49251, _49252,
         _49253, _49254, _49255, _49256, _49257, _49258, _49259, _49260,
         _49261, _49262, _49263, _49264, _49265, _49266, _49267, _49268,
         _49269, _49270, _49271, _49272, _49273, _49274, _49275, _49276,
         _49277, _49278, _49279, _49280, _49281, _49282, _49283, _49284,
         _49285, _49286, _49287, _49288, _49289, _49290, _49291, _49292,
         _49293, _49294, _49295, _49296, _49297, _49298, _49299, _49300,
         _49301, _49302, _49303, _49304, _49305, _49306, _49307, _49308,
         _49309, _49310, _49311, _49312, _49313, _49314, _49315, _49316,
         _49317, _49318, _49319, _49320, _49321, _49322, _49323, _49324,
         _49325, _49326, _49327, _49328, _49329, _49330, _49331, _49332,
         _49333, _49334, _49335, _49336, _49337, _49338, _49339, _49340,
         _49341, _49342, _49343, _49344, _49345, _49346, _49347, _49348,
         _49349, _49350, _49351, _49352, _49353, _49354, _49355, _49356,
         _49357, _49358, _49359, _49360, _49361, _49362, _49363, _49364,
         _49365, _49366, _49367, _49368, _49369, _49370, _49371, _49372,
         _49373, _49374, _49375, _49376, _49377, _49378, _49379, _49380,
         _49381, _49382, _49383, _49384, _49385, _49386, _49387, _49388,
         _49389, _49390, _49391, _49392, _49393, _49394, _49395, _49396,
         _49397, _49398, _49399, _49400, _49401, _49402, _49403, _49404,
         _49405, _49406, _49407, _49408, _49409, _49410, _49411, _49412,
         _49413, _49414, _49415, _49416, _49417, _49418, _49419, _49420,
         _49421, _49422, _49423, _49424, _49425, _49426, _49427, _49428,
         _49429, _49430, _49431, _49432, _49433, _49434, _49435, _49436,
         _49437, _49438, _49439, _49440, _49441, _49442, _49443, _49444,
         _49445, _49446, _49447, _49448, _49449, _49450, _49451, _49452,
         _49453, _49454, _49455, _49456, _49457, _49458, _49459, _49460,
         _49461, _49462, _49463, _49464, _49465, _49466, _49467, _49468,
         _49469, _49470, _49471, _49472, _49473, _49474, _49475, _49476,
         _49477, _49478, _49479, _49480, _49481, _49482, _49483, _49484,
         _49485, _49486, _49487, _49488, _49489, _49490, _49491, _49492,
         _49493, _49494, _49495, _49496, _49497, _49498, _49499, _49500,
         _49501, _49502, _49503, _49504, _49505, _49506, _49507, _49508,
         _49509, _49510, _49511, _49512, _49513, _49514, _49515, _49516,
         _49517, _49518, _49519, _49520, _49521, _49522, _49523, _49524,
         _49525, _49526, _49527, _49528, _49529, _49530, _49531, _49532,
         _49533, _49534, _49535, _49536, _49537, _49538, _49539, _49540,
         _49541, _49542, _49543, _49544, _49545, _49546, _49547, _49548,
         _49549, _49550, _49551, _49552, _49553, _49554, _49555, _49556,
         _49557, _49558, _49559, _49560, _49561, _49562, _49563, _49564,
         _49565, _49566, _49567, _49568, _49569, _49570, _49571, _49572,
         _49573, _49574, _49575, _49576, _49577, _49578, _49579, _49580,
         _49581, _49582, _49583, _49584, _49585, _49586, _49587, _49588,
         _49589, _49590, _49591, _49592, _49593, _49594, _49595, _49596,
         _49597, _49598, _49599, _49600, _49601, _49602, _49603, _49604,
         _49605, _49606, _49607, _49608, _49609, _49610, _49611, _49612,
         _49613, _49614, _49615, _49616, _49617, _49618, _49619, _49620,
         _49621, _49622, _49623, _49624, _49625, _49626, _49627, _49628,
         _49629, _49630, _49631, _49632, _49633, _49634, _49635, _49636,
         _49637, _49638, _49639, _49640, _49641, _49642, _49643, _49644,
         _49645, _49646, _49647, _49648, _49649, _49650, _49651, _49652,
         _49653, _49654, _49655, _49656, _49657, _49658, _49659, _49660,
         _49661, _49662, _49663, _49664, _49665, _49666, _49667, _49668,
         _49669, _49670, _49671, _49672, _49673, _49674, _49675, _49676,
         _49677, _49678, _49679, _49680, _49681, _49682, _49683, _49684,
         _49685, _49686, _49687, _49688, _49689, _49690, _49691, _49692,
         _49693, _49694, _49695, _49696, _49697, _49698, _49699, _49700,
         _49701, _49702, _49703, _49704, _49705, _49706, _49707, _49708,
         _49709, _49710, _49711, _49712, _49713, _49714, _49715, _49716,
         _49717, _49718, _49719, _49720, _49721, _49722, _49723, _49724,
         _49725, _49726, _49727, _49728, _49729, _49730, _49731, _49732,
         _49733, _49734, _49735, _49736, _49737, _49738, _49739, _49740,
         _49741, _49742, _49743, _49744, _49745, _49746, _49747, _49748,
         _49749, _49750, _49751, _49752, _49753, _49754, _49755, _49756,
         _49757, _49758, _49759, _49760, _49761, _49762, _49763, _49764,
         _49765, _49766, _49767, _49768, _49769, _49770, _49771, _49772,
         _49773, _49774, _49775, _49776, _49777, _49778, _49779, _49780,
         _49781, _49782, _49783, _49784, _49785, _49786, _49787, _49788,
         _49789, _49790, _49791, _49792, _49793, _49794, _49795, _49796,
         _49797, _49798, _49799, _49800, _49801, _49802, _49803, _49804,
         _49805, _49806, _49807, _49808, _49809, _49810, _49811, _49812,
         _49813, _49814, _49815, _49816, _49817, _49818, _49819, _49820,
         _49821, _49822, _49823, _49824, _49825, _49826, _49827, _49828,
         _49829, _49830, _49831, _49832, _49833, _49834, _49835, _49836,
         _49837, _49838, _49839, _49840, _49841, _49842, _49843, _49844,
         _49845, _49846, _49847, _49848, _49849, _49850, _49851, _49852,
         _49853, _49854, _49855, _49856, _49857, _49858, _49859, _49860,
         _49861, _49862, _49863, _49864, _49865, _49866, _49867, _49868,
         _49869, _49870, _49871, _49872, _49873, _49874, _49875, _49876,
         _49877, _49878, _49879, _49880, _49881, _49882, _49883, _49884,
         _49885, _49886, _49887, _49888, _49889, _49890, _49891, _49892,
         _49893, _49894, _49895, _49896, _49897, _49898, _49899, _49900,
         _49901, _49902, _49903, _49904, _49905, _49906, _49907, _49908,
         _49909, _49910, _49911, _49912, _49913, _49914, _49915, _49916,
         _49917, _49918, _49919, _49920, _49921, _49922, _49923, _49924,
         _49925, _49926, _49927, _49928, _49929, _49930, _49931, _49932,
         _49933, _49934, _49935, _49936, _49937, _49938, _49939, _49940,
         _49941, _49942, _49943, _49944, _49945, _49946, _49947, _49948,
         _49949, _49950, _49951, _49952, _49953, _49954, _49955, _49956,
         _49957, _49958, _49959, _49960, _49961, _49962, _49963, _49964,
         _49965, _49966, _49967, _49968, _49969, _49970, _49971, _49972,
         _49973, _49974, _49975, _49976, _49977, _49978, _49979, _49980,
         _49981, _49982, _49983, _49984, _49985, _49986, _49987, _49988,
         _49989, _49990, _49991, _49992, _49993, _49994, _49995, _49996,
         _49997, _49998, _49999, _50000, _50001, _50002, _50003, _50004,
         _50005, _50006, _50007, _50008, _50009, _50010, _50011, _50012,
         _50013, _50014, _50015, _50016, _50017, _50018, _50019, _50020,
         _50021, _50022, _50023, _50024, _50025, _50026, _50027, _50028,
         _50029, _50030, _50031, _50032, _50033, _50034, _50035, _50036,
         _50037, _50038, _50039, _50040, _50041, _50042, _50043, _50044,
         _50045, _50046, _50047, _50048, _50049, _50050, _50051, _50052,
         _50053, _50054, _50055, _50056, _50057, _50058, _50059, _50060,
         _50061, _50062, _50063, _50064, _50065, _50066, _50067, _50068,
         _50069, _50070, _50071, _50072, _50073, _50074, _50075, _50076,
         _50077, _50078, _50079, _50080, _50081, _50082, _50083, _50084,
         _50085, _50086, _50087, _50088, _50089, _50090, _50091, _50092,
         _50093, _50094, _50095, _50096, _50097, _50098, _50099, _50100,
         _50101, _50102, _50103, _50104, _50105, _50106, _50107, _50108,
         _50109, _50110, _50111, _50112, _50113, _50114, _50115, _50116,
         _50117, _50118, _50119, _50120, _50121, _50122, _50123, _50124,
         _50125, _50126, _50127, _50128, _50129, _50130, _50131, _50132,
         _50133, _50134, _50135, _50136, _50137, _50138, _50139, _50140,
         _50141, _50142, _50143, _50144, _50145, _50146, _50147, _50148,
         _50149, _50150, _50151, _50152, _50153, _50154, _50155, _50156,
         _50157, _50158, _50159, _50160, _50161, _50162, _50163, _50164,
         _50165, _50166, _50167, _50168, _50169, _50170, _50171, _50172,
         _50173, _50174, _50175, _50176, _50177, _50178, _50179, _50180,
         _50181, _50182, _50183, _50184, _50185, _50186, _50187, _50188,
         _50189, _50190, _50191, _50192, _50193, _50194, _50195, _50196,
         _50197, _50198, _50199, _50200, _50201, _50202, _50203, _50204,
         _50205, _50206, _50207, _50208, _50209, _50210, _50211, _50212,
         _50213, _50214, _50215, _50216, _50217, _50218, _50219, _50220,
         _50221, _50222, _50223, _50224, _50225, _50226, _50227, _50228,
         _50229, _50230, _50231, _50232, _50233, _50234, _50235, _50236,
         _50237, _50238, _50239, _50240, _50241, _50242, _50243, _50244,
         _50245, _50246, _50247, _50248, _50249, _50250, _50251, _50252,
         _50253, _50254, _50255, _50256, _50257, _50258, _50259, _50260,
         _50261, _50262, _50263, _50264, _50265, _50266, _50267, _50268,
         _50269, _50270, _50271, _50272, _50273, _50274, _50275, _50276,
         _50277, _50278, _50279, _50280, _50281, _50282, _50283, _50284,
         _50285, _50286, _50287, _50288, _50289, _50290, _50291, _50292,
         _50293, _50294, _50295, _50296, _50297, _50298, _50299, _50300,
         _50301, _50302, _50303, _50304, _50305, _50306, _50307, _50308,
         _50309, _50310, _50311, _50312, _50313, _50314, _50315, _50316,
         _50317, _50318, _50319, _50320, _50321, _50322, _50323, _50324,
         _50325, _50326, _50327, _50328, _50329, _50330, _50331, _50332,
         _50333, _50334, _50335, _50336, _50337, _50338, _50339, _50340,
         _50341, _50342, _50343, _50344, _50345, _50346, _50347, _50348,
         _50349, _50350, _50351, _50352, _50353, _50354, _50355, _50356,
         _50357, _50358, _50359, _50360, _50361, _50362, _50363, _50364,
         _50365, _50366, _50367, _50368, _50369, _50370, _50371, _50372,
         _50373, _50374, _50375, _50376, _50377, _50378, _50379, _50380,
         _50381, _50382, _50383, _50384, _50385, _50386, _50387, _50388,
         _50389, _50390, _50391, _50392, _50393, _50394, _50395, _50396,
         _50397, _50398, _50399, _50400, _50401, _50402, _50403, _50404,
         _50405, _50406, _50407, _50408, _50409, _50410, _50411, _50412,
         _50413, _50414, _50415, _50416, _50417, _50418, _50419, _50420,
         _50421, _50422, _50423, _50424, _50425, _50426, _50427, _50428,
         _50429, _50430, _50431, _50432, _50433, _50434, _50435, _50436,
         _50437, _50438, _50439, _50440, _50441, _50442, _50443, _50444,
         _50445, _50446, _50447, _50448, _50449, _50450, _50451, _50452,
         _50453, _50454, _50455, _50456, _50457, _50458, _50459, _50460,
         _50461, _50462, _50463, _50464, _50465, _50466, _50467, _50468,
         _50469, _50470, _50471, _50472, _50473, _50474, _50475, _50476,
         _50477, _50478, _50479, _50480, _50481, _50482, _50483, _50484,
         _50485, _50486, _50487, _50488, _50489, _50490, _50491, _50492,
         _50493, _50494, _50495, _50496, _50497, _50498, _50499, _50500,
         _50501, _50502, _50503, _50504, _50505, _50506, _50507, _50508,
         _50509, _50510, _50511, _50512, _50513, _50514, _50515, _50516,
         _50517, _50518, _50519, _50520, _50521, _50522, _50523, _50524,
         _50525, _50526, _50527, _50528, _50529, _50530, _50531, _50532,
         _50533, _50534, _50535, _50536, _50537, _50538, _50539, _50540,
         _50541, _50542, _50543, _50544, _50545, _50546, _50547, _50548,
         _50549, _50550, _50551, _50552, _50553, _50554, _50555, _50556,
         _50557, _50558, _50559, _50560, _50561, _50562, _50563, _50564,
         _50565, _50566, _50567, _50568, _50569, _50570, _50571, _50572,
         _50573, _50574, _50575, _50576, _50577, _50578, _50579, _50580,
         _50581, _50582, _50583, _50584, _50585, _50586, _50587, _50588,
         _50589, _50590, _50591, _50592, _50593, _50594, _50595, _50596,
         _50597, _50598, _50599, _50600, _50601, _50602, _50603, _50604,
         _50605, _50606, _50607, _50608, _50609, _50610, _50611, _50612,
         _50613, _50614, _50615, _50616, _50617, _50618, _50619, _50620,
         _50621, _50622, _50623, _50624, _50625, _50626, _50627, _50628,
         _50629, _50630, _50631, _50632, _50633, _50634, _50635, _50636,
         _50637, _50638, _50639, _50640, _50641, _50642, _50643, _50644,
         _50645, _50646, _50647, _50648, _50649, _50650, _50651, _50652,
         _50653, _50654, _50655, _50656, _50657, _50658, _50659, _50660,
         _50661, _50662, _50663, _50664, _50665, _50666, _50667, _50668,
         _50669, _50670, _50671, _50672, _50673, _50674, _50675, _50676,
         _50677, _50678, _50679, _50680, _50681, _50682, _50683, _50684,
         _50685, _50686, _50687, _50688, _50689, _50690, _50691, _50692,
         _50693, _50694, _50695, _50696, _50697, _50698, _50699, _50700,
         _50701, _50702, _50703, _50704, _50705, _50706, _50707, _50708,
         _50709, _50710, _50711, _50712, _50713, _50714, _50715, _50716,
         _50717, _50718, _50719, _50720, _50721, _50722, _50723, _50724,
         _50725, _50726, _50727, _50728, _50729, _50730, _50731, _50732,
         _50733, _50734, _50735, _50736, _50737, _50738, _50739, _50740,
         _50741, _50742, _50743, _50744, _50745, _50746, _50747, _50748,
         _50749, _50750, _50751, _50752, _50753, _50754, _50755, _50756,
         _50757, _50758, _50759, _50760, _50761, _50762, _50763, _50764,
         _50765, _50766, _50767, _50768, _50769, _50770, _50771, _50772,
         _50773, _50774, _50775, _50776, _50777, _50778, _50779, _50780,
         _50781, _50782, _50783, _50784, _50785, _50786, _50787, _50788,
         _50789, _50790, _50791, _50792, _50793, _50794, _50795, _50796,
         _50797, _50798, _50799, _50800, _50801, _50802, _50803, _50804,
         _50805, _50806, _50807, _50808, _50809, _50810, _50811, _50812,
         _50813, _50814, _50815, _50816, _50817, _50818, _50819, _50820,
         _50821, _50822, _50823, _50824, _50825, _50826, _50827, _50828,
         _50829, _50830, _50831, _50832, _50833, _50834, _50835, _50836,
         _50837, _50838, _50839, _50840, _50841, _50842, _50843, _50844,
         _50845, _50846, _50847, _50848, _50849, _50850, _50851, _50852,
         _50853, _50854, _50855, _50856, _50857, _50858, _50859, _50860,
         _50861, _50862, _50863, _50864, _50865, _50866, _50867, _50868,
         _50869, _50870, _50871, _50872, _50873, _50874, _50875, _50876,
         _50877, _50878, _50879, _50880, _50881, _50882, _50883, _50884,
         _50885, _50886, _50887, _50888, _50889, _50890, _50891, _50892,
         _50893, _50894, _50895, _50896, _50897, _50898, _50899, _50900,
         _50901, _50902, _50903, _50904, _50905, _50906, _50907, _50908,
         _50909, _50910, _50911, _50912, _50913, _50914, _50915, _50916,
         _50917, _50918, _50919, _50920, _50921, _50922, _50923, _50924,
         _50925, _50926, _50927, _50928, _50929, _50930, _50931, _50932,
         _50933, _50934, _50935, _50936, _50937, _50938, _50939, _50940,
         _50941, _50942, _50943, _50944, _50945, _50946, _50947, _50948,
         _50949, _50950, _50951, _50952, _50953, _50954, _50955, _50956,
         _50957, _50958, _50959, _50960, _50961, _50962, _50963, _50964,
         _50965, _50966, _50967, _50968, _50969, _50970, _50971, _50972,
         _50973, _50974, _50975, _50976, _50977, _50978, _50979, _50980,
         _50981, _50982, _50983, _50984, _50985, _50986, _50987, _50988,
         _50989, _50990, _50991, _50992, _50993, _50994, _50995, _50996,
         _50997, _50998, _50999, _51000, _51001, _51002, _51003, _51004,
         _51005, _51006, _51007, _51008, _51009, _51010, _51011, _51012,
         _51013, _51014, _51015, _51016, _51017, _51018, _51019, _51020,
         _51021, _51022, _51023, _51024, _51025, _51026, _51027, _51028,
         _51029, _51030, _51031, _51032, _51033, _51034, _51035, _51036,
         _51037, _51038, _51039, _51040, _51041, _51042, _51043, _51044,
         _51045, _51046, _51047, _51048, _51049, _51050, _51051, _51052,
         _51053, _51054, _51055, _51056, _51057, _51058, _51059, _51060,
         _51061, _51062, _51063, _51064, _51065, _51066, _51067, _51068,
         _51069, _51070, _51071, _51072, _51073, _51074, _51075, _51076,
         _51077, _51078, _51079, _51080, _51081, _51082, _51083, _51084,
         _51085, _51086, _51087, _51088, _51089, _51090, _51091, _51092,
         _51093, _51094, _51095, _51096, _51097, _51098, _51099, _51100,
         _51101, _51102, _51103, _51104, _51105, _51106, _51107, _51108,
         _51109, _51110, _51111, _51112, _51113, _51114, _51115, _51116,
         _51117, _51118, _51119, _51120, _51121, _51122, _51123, _51124,
         _51125, _51126, _51127, _51128, _51129, _51130, _51131, _51132,
         _51133, _51134, _51135, _51136, _51137, _51138, _51139, _51140,
         _51141, _51142, _51143, _51144, _51145, _51146, _51147, _51148,
         _51149, _51150, _51151, _51152, _51153, _51154, _51155, _51156,
         _51157, _51158, _51159, _51160, _51161, _51162, _51163, _51164,
         _51165, _51166, _51167, _51168, _51169, _51170, _51171, _51172,
         _51173, _51174, _51175, _51176, _51177, _51178, _51179, _51180,
         _51181, _51182, _51183, _51184, _51185, _51186, _51187, _51188,
         _51189, _51190, _51191, _51192, _51193, _51194, _51195, _51196,
         _51197, _51198, _51199, _51200, _51201, _51202, _51203, _51204,
         _51205, _51206, _51207, _51208, _51209, _51210, _51211, _51212,
         _51213, _51214, _51215, _51216, _51217, _51218, _51219, _51220,
         _51221, _51222, _51223, _51224, _51225, _51226, _51227, _51228,
         _51229, _51230, _51231, _51232, _51233, _51234, _51235, _51236,
         _51237, _51238, _51239, _51240, _51241, _51242, _51243, _51244,
         _51245, _51246, _51247, _51248, _51249, _51250, _51251, _51252,
         _51253, _51254, _51255, _51256, _51257, _51258, _51259, _51260,
         _51261, _51262, _51263, _51264, _51265, _51266, _51267, _51268,
         _51269, _51270, _51271, _51272, _51273, _51274, _51275, _51276,
         _51277, _51278, _51279, _51280, _51281, _51282, _51283, _51284,
         _51285, _51286, _51287, _51288, _51289, _51290, _51291, _51292,
         _51293, _51294, _51295, _51296, _51297, _51298, _51299, _51300,
         _51301, _51302, _51303, _51304, _51305, _51306, _51307, _51308,
         _51309, _51310, _51311, _51312, _51313, _51314, _51315, _51316,
         _51317, _51318, _51319, _51320, _51321, _51322, _51323, _51324,
         _51325, _51326, _51327, _51328, _51329, _51330, _51331, _51332,
         _51333, _51334, _51335, _51336, _51337, _51338, _51339, _51340,
         _51341, _51342, _51343, _51344, _51345, _51346, _51347, _51348,
         _51349, _51350, _51351, _51352, _51353, _51354, _51355, _51356,
         _51357, _51358, _51359, _51360, _51361, _51362, _51363, _51364,
         _51365, _51366, _51367, _51368, _51369, _51370, _51371, _51372,
         _51373, _51374, _51375, _51376, _51377, _51378, _51379, _51380,
         _51381, _51382, _51383, _51384, _51385, _51386, _51387, _51388,
         _51389, _51390, _51391, _51392, _51393, _51394, _51395, _51396,
         _51397, _51398, _51399, _51400, _51401, _51402, _51403, _51404,
         _51405, _51406, _51407, _51408, _51409, _51410, _51411, _51412,
         _51413, _51414, _51415, _51416, _51417, _51418, _51419, _51420,
         _51421, _51422, _51423, _51424, _51425, _51426, _51427, _51428,
         _51429, _51430, _51431, _51432, _51433, _51434, _51435, _51436,
         _51437, _51438, _51439, _51440, _51441, _51442, _51443, _51444,
         _51445, _51446, _51447, _51448, _51449, _51450, _51451, _51452,
         _51453, _51454, _51455, _51456, _51457, _51458, _51459, _51460,
         _51461, _51462, _51463, _51464, _51465, _51466, _51467, _51468,
         _51469, _51470, _51471, _51472, _51473, _51474, _51475, _51476,
         _51477, _51478, _51479, _51480, _51481, _51482, _51483, _51484,
         _51485, _51486, _51487, _51488, _51489, _51490, _51491, _51492,
         _51493, _51494, _51495, _51496, _51497, _51498, _51499, _51500,
         _51501, _51502, _51503, _51504, _51505, _51506, _51507, _51508,
         _51509, _51510, _51511, _51512, _51513, _51514, _51515, _51516,
         _51517, _51518, _51519, _51520, _51521, _51522, _51523, _51524,
         _51525, _51526, _51527, _51528, _51529, _51530, _51531, _51532,
         _51533, _51534, _51535, _51536, _51537, _51538, _51539, _51540,
         _51541, _51542, _51543, _51544, _51545, _51546, _51547, _51548,
         _51549, _51550, _51551, _51552, _51553, _51554, _51555, _51556,
         _51557, _51558, _51559, _51560, _51561, _51562, _51563, _51564,
         _51565, _51566, _51567, _51568, _51569, _51570, _51571, _51572,
         _51573, _51574, _51575, _51576, _51577, _51578, _51579, _51580,
         _51581, _51582, _51583, _51584, _51585, _51586, _51587, _51588,
         _51589, _51590, _51591, _51592, _51593, _51594, _51595, _51596,
         _51597, _51598, _51599, _51600, _51601, _51602, _51603, _51604,
         _51605, _51606, _51607, _51608, _51609, _51610, _51611, _51612,
         _51613, _51614, _51615, _51616, _51617, _51618, _51619, _51620,
         _51621, _51622, _51623, _51624, _51625, _51626, _51627, _51628,
         _51629, _51630, _51631, _51632, _51633, _51634, _51635, _51636,
         _51637, _51638, _51639, _51640, _51641, _51642, _51643, _51644,
         _51645, _51646, _51647, _51648, _51649, _51650, _51651, _51652,
         _51653, _51654, _51655, _51656, _51657, _51658, _51659, _51660,
         _51661, _51662, _51663, _51664, _51665, _51666, _51667, _51668,
         _51669, _51670, _51671, _51672, _51673, _51674, _51675, _51676,
         _51677, _51678, _51679, _51680, _51681, _51682, _51683, _51684,
         _51685, _51686, _51687, _51688, _51689, _51690, _51691, _51692,
         _51693, _51694, _51695, _51696, _51697, _51698, _51699, _51700,
         _51701, _51702, _51703, _51704, _51705, _51706, _51707, _51708,
         _51709, _51710, _51711, _51712, _51713, _51714, _51715, _51716,
         _51717, _51718, _51719, _51720, _51721, _51722, _51723, _51724,
         _51725, _51726, _51727, _51728, _51729, _51730, _51731, _51732,
         _51733, _51734, _51735, _51736, _51737, _51738, _51739, _51740,
         _51741, _51742, _51743, _51744, _51745, _51746, _51747, _51748,
         _51749, _51750, _51751, _51752, _51753, _51754, _51755, _51756,
         _51757, _51758, _51759, _51760, _51761, _51762, _51763, _51764,
         _51765, _51766, _51767, _51768, _51769, _51770, _51771, _51772,
         _51773, _51774, _51775, _51776, _51777, _51778, _51779, _51780,
         _51781, _51782, _51783, _51784, _51785, _51786, _51787, _51788,
         _51789, _51790, _51791, _51792, _51793, _51794, _51795, _51796,
         _51797, _51798, _51799, _51800, _51801, _51802, _51803, _51804,
         _51805, _51806, _51807, _51808, _51809, _51810, _51811, _51812,
         _51813, _51814, _51815, _51816, _51817, _51818, _51819, _51820,
         _51821, _51822, _51823, _51824, _51825, _51826, _51827, _51828,
         _51829, _51830, _51831, _51832, _51833, _51834, _51835, _51836,
         _51837, _51838, _51839, _51840, _51841, _51842, _51843, _51844,
         _51845, _51846, _51847, _51848, _51849, _51850, _51851, _51852,
         _51853, _51854, _51855, _51856, _51857, _51858, _51859, _51860,
         _51861, _51862, _51863, _51864, _51865, _51866, _51867, _51868,
         _51869, _51870, _51871, _51872, _51873, _51874, _51875, _51876,
         _51877, _51878, _51879, _51880, _51881, _51882, _51883, _51884,
         _51885, _51886, _51887, _51888, _51889, _51890, _51891, _51892,
         _51893, _51894, _51895, _51896, _51897, _51898, _51899, _51900,
         _51901, _51902, _51903, _51904, _51905, _51906, _51907, _51908,
         _51909, _51910, _51911, _51912, _51913, _51914, _51915, _51916,
         _51917, _51918, _51919, _51920, _51921, _51922, _51923, _51924,
         _51925, _51926, _51927, _51928, _51929, _51930, _51931, _51932,
         _51933, _51934, _51935, _51936, _51937, _51938, _51939, _51940,
         _51941, _51942, _51943, _51944, _51945, _51946, _51947, _51948,
         _51949, _51950, _51951, _51952, _51953, _51954, _51955, _51956,
         _51957, _51958, _51959, _51960, _51961, _51962, _51963, _51964,
         _51965, _51966, _51967, _51968, _51969, _51970, _51971, _51972,
         _51973, _51974, _51975, _51976, _51977, _51978, _51979, _51980,
         _51981, _51982, _51983, _51984, _51985, _51986, _51987, _51988,
         _51989, _51990, _51991, _51992, _51993, _51994, _51995, _51996,
         _51997, _51998, _51999, _52000, _52001, _52002, _52003, _52004,
         _52005, _52006, _52007, _52008, _52009, _52010, _52011, _52012,
         _52013, _52014, _52015, _52016, _52017, _52018, _52019, _52020,
         _52021, _52022, _52023, _52024, _52025, _52026, _52027, _52028,
         _52029, _52030, _52031, _52032, _52033, _52034, _52035, _52036,
         _52037, _52038, _52039, _52040, _52041, _52042, _52043, _52044,
         _52045, _52046, _52047, _52048, _52049, _52050, _52051, _52052,
         _52053, _52054, _52055, _52056, _52057, _52058, _52059, _52060,
         _52061, _52062, _52063, _52064, _52065, _52066, _52067, _52068,
         _52069, _52070, _52071, _52072, _52073, _52074, _52075, _52076,
         _52077, _52078, _52079, _52080, _52081, _52082, _52083, _52084,
         _52085, _52086, _52087, _52088, _52089, _52090, _52091, _52092,
         _52093, _52094, _52095, _52096, _52097, _52098, _52099, _52100,
         _52101, _52102, _52103, _52104, _52105, _52106, _52107, _52108,
         _52109, _52110, _52111, _52112, _52113, _52114, _52115, _52116,
         _52117, _52118, _52119, _52120, _52121, _52122, _52123, _52124,
         _52125, _52126, _52127, _52128, _52129, _52130, _52131, _52132,
         _52133, _52134, _52135, _52136, _52137, _52138, _52139, _52140,
         _52141, _52142, _52143, _52144, _52145, _52146, _52147, _52148,
         _52149, _52150, _52151, _52152, _52153, _52154, _52155, _52156,
         _52157, _52158, _52159, _52160, _52161, _52162, _52163, _52164,
         _52165, _52166, _52167, _52168, _52169, _52170, _52171, _52172,
         _52173, _52174, _52175, _52176, _52177, _52178, _52179, _52180,
         _52181, _52182, _52183, _52184, _52185, _52186, _52187, _52188,
         _52189, _52190, _52191, _52192, _52193, _52194, _52195, _52196,
         _52197, _52198, _52199, _52200, _52201, _52202, _52203, _52204,
         _52205, _52206, _52207, _52208, _52209, _52210, _52211, _52212,
         _52213, _52214, _52215, _52216, _52217, _52218, _52219, _52220,
         _52221, _52222, _52223, _52224, _52225, _52226, _52227, _52228,
         _52229, _52230, _52231, _52232, _52233, _52234, _52235, _52236,
         _52237, _52238, _52239, _52240, _52241, _52242, _52243, _52244,
         _52245, _52246, _52247, _52248, _52249, _52250, _52251, _52252,
         _52253, _52254, _52255, _52256, _52257, _52258, _52259, _52260,
         _52261, _52262, _52263, _52264, _52265, _52266, _52267, _52268,
         _52269, _52270, _52271, _52272, _52273, _52274, _52275, _52276,
         _52277, _52278, _52279, _52280, _52281, _52282, _52283, _52284,
         _52285, _52286, _52287, _52288, _52289, _52290, _52291, _52292,
         _52293, _52294, _52295, _52296, _52297, _52298, _52299, _52300,
         _52301, _52302, _52303, _52304, _52305, _52306, _52307, _52308,
         _52309, _52310, _52311, _52312, _52313, _52314, _52315, _52316,
         _52317, _52318, _52319, _52320, _52321, _52322, _52323, _52324,
         _52325, _52326, _52327, _52328, _52329, _52330, _52331, _52332,
         _52333, _52334, _52335, _52336, _52337, _52338, _52339, _52340,
         _52341, _52342, _52343, _52344, _52345, _52346, _52347, _52348,
         _52349, _52350, _52351, _52352, _52353, _52354, _52355, _52356,
         _52357, _52358, _52359, _52360, _52361, _52362, _52363, _52364,
         _52365, _52366, _52367, _52368, _52369, _52370, _52371, _52372,
         _52373, _52374, _52375, _52376, _52377, _52378, _52379, _52380,
         _52381, _52382, _52383, _52384, _52385, _52386, _52387, _52388,
         _52389, _52390, _52391, _52392, _52393, _52394, _52395, _52396,
         _52397, _52398, _52399, _52400, _52401, _52402, _52403, _52404,
         _52405, _52406, _52407, _52408, _52409, _52410, _52411, _52412,
         _52413, _52414, _52415, _52416, _52417, _52418, _52419, _52420,
         _52421, _52422, _52423, _52424, _52425, _52426, _52427, _52428,
         _52429, _52430, _52431, _52432, _52433, _52434, _52435, _52436,
         _52437, _52438, _52439, _52440, _52441, _52442, _52443, _52444,
         _52445, _52446, _52447, _52448, _52449, _52450, _52451, _52452,
         _52453, _52454, _52455, _52456, _52457, _52458, _52459, _52460,
         _52461, _52462, _52463, _52464, _52465, _52466, _52467, _52468,
         _52469, _52470, _52471, _52472, _52473, _52474, _52475, _52476,
         _52477, _52478, _52479, _52480, _52481, _52482, _52483, _52484,
         _52485, _52486, _52487, _52488, _52489, _52490, _52491, _52492,
         _52493, _52494, _52495, _52496, _52497, _52498, _52499, _52500,
         _52501, _52502, _52503, _52504, _52505, _52506, _52507, _52508,
         _52509, _52510, _52511, _52512, _52513, _52514, _52515, _52516,
         _52517, _52518, _52519, _52520, _52521, _52522, _52523, _52524,
         _52525, _52526, _52527, _52528, _52529, _52530, _52531, _52532,
         _52533, _52534, _52535, _52536, _52537, _52538, _52539, _52540,
         _52541, _52542, _52543, _52544, _52545, _52546, _52547, _52548,
         _52549, _52550, _52551, _52552, _52553, _52554, _52555, _52556,
         _52557, _52558, _52559, _52560, _52561, _52562, _52563, _52564,
         _52565, _52566, _52567, _52568, _52569, _52570, _52571, _52572,
         _52573, _52574, _52575, _52576, _52577, _52578, _52579, _52580,
         _52581, _52582, _52583, _52584, _52585, _52586, _52587, _52588,
         _52589, _52590, _52591, _52592, _52593, _52594, _52595, _52596,
         _52597, _52598, _52599, _52600, _52601, _52602, _52603, _52604,
         _52605, _52606, _52607, _52608, _52609, _52610, _52611, _52612,
         _52613, _52614, _52615, _52616, _52617, _52618, _52619, _52620,
         _52621, _52622, _52623, _52624, _52625, _52626, _52627, _52628,
         _52629, _52630, _52631, _52632, _52633, _52634, _52635, _52636,
         _52637, _52638, _52639, _52640, _52641, _52642, _52643, _52644,
         _52645, _52646, _52647, _52648, _52649, _52650, _52651, _52652,
         _52653, _52654, _52655, _52656, _52657, _52658, _52659, _52660,
         _52661, _52662, _52663, _52664, _52665, _52666, _52667, _52668,
         _52669, _52670, _52671, _52672, _52673, _52674, _52675, _52676,
         _52677, _52678, _52679, _52680, _52681, _52682, _52683, _52684,
         _52685, _52686, _52687, _52688, _52689, _52690, _52691, _52692,
         _52693, _52694, _52695, _52696, _52697, _52698, _52699, _52700,
         _52701, _52702, _52703, _52704, _52705, _52706, _52707, _52708,
         _52709, _52710, _52711, _52712, _52713, _52714, _52715, _52716,
         _52717, _52718, _52719, _52720, _52721, _52722, _52723, _52724,
         _52725, _52726, _52727, _52728, _52729, _52730, _52731, _52732,
         _52733, _52734, _52735, _52736, _52737, _52738, _52739, _52740,
         _52741, _52742, _52743, _52744, _52745, _52746, _52747, _52748,
         _52749, _52750, _52751, _52752, _52753, _52754, _52755, _52756,
         _52757, _52758, _52759, _52760, _52761, _52762, _52763, _52764,
         _52765, _52766, _52767, _52768, _52769, _52770, _52771, _52772,
         _52773, _52774, _52775, _52776, _52777, _52778, _52779, _52780,
         _52781, _52782, _52783, _52784, _52785, _52786, _52787, _52788,
         _52789, _52790, _52791, _52792, _52793, _52794, _52795, _52796,
         _52797, _52798, _52799, _52800, _52801, _52802, _52803, _52804,
         _52805, _52806, _52807, _52808, _52809, _52810, _52811, _52812,
         _52813, _52814, _52815, _52816, _52817, _52818, _52819, _52820,
         _52821, _52822, _52823, _52824, _52825, _52826, _52827, _52828,
         _52829, _52830, _52831, _52832, _52833, _52834, _52835, _52836,
         _52837, _52838, _52839, _52840, _52841, _52842, _52843, _52844,
         _52845, _52846, _52847, _52848, _52849, _52850, _52851, _52852,
         _52853, _52854, _52855, _52856, _52857, _52858, _52859, _52860,
         _52861, _52862, _52863, _52864, _52865, _52866, _52867, _52868,
         _52869, _52870, _52871, _52872, _52873, _52874, _52875, _52876,
         _52877, _52878, _52879, _52880, _52881, _52882, _52883, _52884,
         _52885, _52886, _52887, _52888, _52889, _52890, _52891, _52892,
         _52893, _52894, _52895, _52896, _52897, _52898, _52899, _52900,
         _52901, _52902, _52903, _52904, _52905, _52906, _52907, _52908,
         _52909, _52910, _52911, _52912, _52913, _52914, _52915, _52916,
         _52917, _52918, _52919, _52920, _52921, _52922, _52923, _52924,
         _52925, _52926, _52927, _52928, _52929, _52930, _52931, _52932,
         _52933, _52934, _52935, _52936, _52937, _52938, _52939, _52940,
         _52941, _52942, _52943, _52944, _52945, _52946, _52947, _52948,
         _52949, _52950, _52951, _52952, _52953, _52954, _52955, _52956,
         _52957, _52958, _52959, _52960, _52961, _52962, _52963, _52964,
         _52965, _52966, _52967, _52968, _52969, _52970, _52971, _52972,
         _52973, _52974, _52975, _52976, _52977, _52978, _52979, _52980,
         _52981, _52982, _52983, _52984, _52985, _52986, _52987, _52988,
         _52989, _52990, _52991, _52992, _52993, _52994, _52995, _52996,
         _52997, _52998, _52999, _53000, _53001, _53002, _53003, _53004,
         _53005, _53006, _53007, _53008, _53009, _53010, _53011, _53012,
         _53013, _53014, _53015, _53016, _53017, _53018, _53019, _53020,
         _53021, _53022, _53023, _53024, _53025, _53026, _53027, _53028,
         _53029, _53030, _53031, _53032, _53033, _53034, _53035, _53036,
         _53037, _53038, _53039, _53040, _53041, _53042, _53043, _53044,
         _53045, _53046, _53047, _53048, _53049, _53050, _53051, _53052,
         _53053, _53054, _53055, _53056, _53057, _53058, _53059, _53060,
         _53061, _53062, _53063, _53064, _53065, _53066, _53067, _53068,
         _53069, _53070, _53071, _53072, _53073, _53074, _53075, _53076,
         _53077, _53078, _53079, _53080, _53081, _53082, _53083, _53084,
         _53085, _53086, _53087, _53088, _53089, _53090, _53091, _53092,
         _53093, _53094, _53095, _53096, _53097, _53098, _53099, _53100,
         _53101, _53102, _53103, _53104, _53105, _53106, _53107, _53108,
         _53109, _53110, _53111, _53112, _53113, _53114, _53115, _53116,
         _53117, _53118, _53119, _53120, _53121, _53122, _53123, _53124,
         _53125, _53126, _53127, _53128, _53129, _53130, _53131, _53132,
         _53133, _53134, _53135, _53136, _53137, _53138, _53139, _53140,
         _53141, _53142, _53143, _53144, _53145, _53146, _53147, _53148,
         _53149, _53150, _53151, _53152, _53153, _53154, _53155, _53156,
         _53157, _53158, _53159, _53160, _53161, _53162, _53163, _53164,
         _53165, _53166, _53167, _53168, _53169, _53170, _53171, _53172,
         _53173, _53174, _53175, _53176, _53177, _53178, _53179, _53180,
         _53181, _53182, _53183, _53184, _53185, _53186, _53187, _53188,
         _53189, _53190, _53191, _53192, _53193, _53194, _53195, _53196,
         _53197, _53198, _53199, _53200, _53201, _53202, _53203, _53204,
         _53205, _53206, _53207, _53208, _53209, _53210, _53211, _53212,
         _53213, _53214, _53215, _53216, _53217, _53218, _53219, _53220,
         _53221, _53222, _53223, _53224, _53225, _53226, _53227, _53228,
         _53229, _53230, _53231, _53232, _53233, _53234, _53235, _53236,
         _53237, _53238, _53239, _53240, _53241, _53242, _53243, _53244,
         _53245, _53246, _53247, _53248, _53249, _53250, _53251, _53252,
         _53253, _53254, _53255, _53256, _53257, _53258, _53259, _53260,
         _53261, _53262, _53263, _53264, _53265, _53266, _53267, _53268,
         _53269, _53270, _53271, _53272, _53273, _53274, _53275, _53276,
         _53277, _53278, _53279, _53280, _53281, _53282, _53283, _53284,
         _53285, _53286, _53287, _53288, _53289, _53290, _53291, _53292,
         _53293, _53294, _53295, _53296, _53297, _53298, _53299, _53300,
         _53301, _53302, _53303, _53304, _53305, _53306, _53307, _53308,
         _53309, _53310, _53311, _53312, _53313, _53314, _53315, _53316,
         _53317, _53318, _53319, _53320, _53321, _53322, _53323, _53324,
         _53325, _53326, _53327, _53328, _53329, _53330, _53331, _53332,
         _53333, _53334, _53335, _53336, _53337, _53338, _53339, _53340,
         _53341, _53342, _53343, _53344, _53345, _53346, _53347, _53348,
         _53349, _53350, _53351, _53352, _53353, _53354, _53355, _53356,
         _53357, _53358, _53359, _53360, _53361, _53362, _53363, _53364,
         _53365, _53366, _53367, _53368, _53369, _53370, _53371, _53372,
         _53373, _53374, _53375, _53376, _53377, _53378, _53379, _53380,
         _53381, _53382, _53383, _53384, _53385, _53386, _53387, _53388,
         _53389, _53390, _53391, _53392, _53393, _53394, _53395, _53396,
         _53397, _53398, _53399, _53400, _53401, _53402, _53403, _53404,
         _53405, _53406, _53407, _53408, _53409, _53410, _53411, _53412,
         _53413, _53414, _53415, _53416, _53417, _53418, _53419, _53420,
         _53421, _53422, _53423, _53424, _53425, _53426, _53427, _53428,
         _53429, _53430, _53431, _53432, _53433, _53434, _53435, _53436,
         _53437, _53438, _53439, _53440, _53441, _53442, _53443, _53444,
         _53445, _53446, _53447, _53448, _53449, _53450, _53451, _53452,
         _53453, _53454, _53455, _53456, _53457, _53458, _53459, _53460,
         _53461, _53462, _53463, _53464, _53465, _53466, _53467, _53468,
         _53469, _53470, _53471, _53472, _53473, _53474, _53475, _53476,
         _53477, _53478, _53479, _53480, _53481, _53482, _53483, _53484,
         _53485, _53486, _53487, _53488, _53489, _53490, _53491, _53492,
         _53493, _53494, _53495, _53496, _53497, _53498, _53499, _53500,
         _53501, _53502, _53503, _53504, _53505, _53506, _53507, _53508,
         _53509, _53510, _53511, _53512, _53513, _53514, _53515, _53516,
         _53517, _53518, _53519, _53520, _53521, _53522, _53523, _53524,
         _53525, _53526;
  wire   [31:0] ______;
  wire   [31:0] _______;
  wire   [13:0] ____0___________0;
  wire   [15:0] ____1___________0;
  wire   [15:0] ____0___________;
  wire   [11:0] ____1___________;
  wire   [13:0] ____2___________;
  wire   [10:0] ____3___________;
  assign ______[31] = inData[31];
  assign ______[30] = inData[30];
  assign ______[29] = inData[29];
  assign ______[28] = inData[28];
  assign ______[27] = inData[27];
  assign ______[26] = inData[26];
  assign ______[25] = inData[25];
  assign ______[24] = inData[24];
  assign ______[23] = inData[23];
  assign ______[22] = inData[22];
  assign ______[21] = inData[21];
  assign ______[20] = inData[20];
  assign ______[19] = inData[19];
  assign ______[18] = inData[18];
  assign ______[17] = inData[17];
  assign ______[16] = inData[16];
  assign ______[15] = inData[15];
  assign ______[14] = inData[14];
  assign ______[13] = inData[13];
  assign ______[12] = inData[12];
  assign ______[11] = inData[11];
  assign ______[10] = inData[10];
  assign ______[9] = inData[9];
  assign ______[8] = inData[8];
  assign ______[7] = inData[7];
  assign ______[6] = inData[6];
  assign ______[5] = inData[5];
  assign ______[4] = inData[4];
  assign ______[3] = inData[3];
  assign ______[2] = inData[2];
  assign ______[1] = inData[1];
  assign ______[0] = inData[0];
  assign ___ = clk;
  assign _____ = reset;
  assign outData[31] = _______[31];
  assign outData[30] = _______[30];
  assign outData[29] = _______[29];
  assign outData[28] = _______[28];
  assign outData[27] = _______[27];
  assign outData[26] = _______[26];
  assign outData[25] = _______[25];
  assign outData[24] = _______[24];
  assign outData[23] = _______[23];
  assign outData[22] = _______[22];
  assign outData[21] = _______[21];
  assign outData[20] = _______[20];
  assign outData[19] = _______[19];
  assign outData[18] = _______[18];
  assign outData[17] = _______[17];
  assign outData[16] = _______[16];
  assign outData[15] = _______[15];
  assign outData[14] = _______[14];
  assign outData[13] = _______[13];
  assign outData[12] = _______[12];
  assign outData[11] = _______[11];
  assign outData[10] = _______[10];
  assign outData[9] = _______[9];
  assign outData[8] = _______[8];
  assign outData[7] = _______[7];
  assign outData[6] = _______[6];
  assign outData[5] = _______[5];
  assign outData[4] = _______[4];
  assign outData[3] = _______[3];
  assign outData[2] = _______[2];
  assign outData[1] = _______[1];
  assign outData[0] = _______[0];

  dffacs2 _______________1_ ( .DIN(
        _______1____2________________1____________________), .CLK(_26904), 
        .CLRB(_____), .Q(_53366), .QN(_26698) );
  dffacs2 _______________26_ ( .DIN(
        _______26____2________________26____________________), .CLK(_26880), 
        .CLRB(_____), .Q(_53365), .QN(_26331) );
  dffacs2 _______________23_ ( .DIN(
        _______23____2________________23____________________), .CLK(_26913), 
        .CLRB(_____), .Q(_26526), .QN(_53309) );
  dffacs2 _______________22_ ( .DIN(
        _______22____2________________22____________________), .CLK(_26909), 
        .CLRB(_____), .Q(_53314), .QN(_26343) );
  dffacs2 _______________20_ ( .DIN(
        _______20____2________________20____________________), .CLK(_26933), 
        .CLRB(_____), .Q(_53370), .QN(_26778) );
  dffacs2 _______________17_ ( .DIN(
        _______17____2________________17____________________), .CLK(___), 
        .CLRB(_____), .Q(_53373), .QN(_26333) );
  dffacs2 _______________16_ ( .DIN(
        _______16____2________________16____________________), .CLK(_26982), 
        .CLRB(_____), .Q(_53374), .QN(_26322) );
  dffacs2 _______________8_ ( .DIN(
        _______8____2________________8____________________), .CLK(_26981), 
        .CLRB(_____), .Q(_26330), .QN(_53380) );
  dffacs2 _______________5_ ( .DIN(
        _______5____2________________5____________________), .CLK(_26953), 
        .CLRB(_____), .Q(_53357), .QN(_26396) );
  dffacs2 _______________4_ ( .DIN(
        _______4____2________________4____________________), .CLK(_26974), 
        .CLRB(_____), .Q(_53358), .QN(_26448) );
  dffacs2 _______________15_ ( .DIN(
        _______15____2________________15____________________), .CLK(_26982), 
        .CLRB(_____), .Q(_53372), .QN(_26336) );
  dffacs2 _______________7_ ( .DIN(
        _______7____2________________7____________________), .CLK(_26980), 
        .CLRB(_____), .Q(_53350), .QN(_26320) );
  dffacs2 _________________________________________0__1_ ( .DIN(
        _________________________________________2_________), .CLK(_26890), 
        .CLRB(_____), .Q(_53053) );
  dffacs2 _______________14_ ( .DIN(
        _______14____2________________14____________________), .CLK(_26981), 
        .CLRB(_____), .Q(_53338), .QN(_26319) );
  dffacs2 _______________24_ ( .DIN(
        _______24____2________________24____________________), .CLK(_26895), 
        .CLRB(_____), .Q(_26209), .QN(_53367) );
  dffacs2 __________________________________________5__25_ ( .DIN(
        ______________________________154________), .CLK(_26893), .CLRB(_____), 
        .Q(_52934) );
  dffacs2 ____0________________12_ ( .DIN(____0___________0_12_____), .CLK(
        _26895), .CLRB(_____), .Q(_53472), .QN(_26369) );
  dffacs2 ____0________________8_ ( .DIN(____0___________0_8_____), .CLK(
        _26973), .CLRB(_____), .Q(_53478), .QN(_26219) );
  dffacs2 ____0________________1_0 ( .DIN(____0____________1_____), .CLK(
        _26911), .CLRB(_____), .Q(_53448), .QN(_26227) );
  dffacs2 __________________________________________0__13_ ( .DIN(
        __________________________________________13_________), .CLK(_26953), 
        .CLRB(_____), .Q(_53183) );
  dffacs2 _________________________________________5__1_ ( .DIN(
        _____________________________130________), .CLK(_26880), .CLRB(_____), 
        .Q(_53093) );
  dffacs2 _________________________________________6__26_ ( .DIN(
        _____________________________187________), .CLK(_26909), .CLRB(_____), 
        .Q(_53180) );
  dffacs2 _________________________________________9__21_ ( .DIN(
        _____________________________278________), .CLK(_26862), .CLRB(_____), 
        .Q(_53179) );
  dffacs2 __________________________________________6__8_ ( .DIN(
        ______________________________169________), .CLK(_26881), .CLRB(_____), 
        .Q(_52964) );
  dffacs2 ____0________________3_ ( .DIN(____0___________0_3_____), .CLK(
        _26895), .CLRB(_____), .Q(_53479), .QN(_26416) );
  dffacs2 __________________________________________4__31_ ( .DIN(
        ______________________________128________), .CLK(_26899), .CLRB(_____), 
        .Q(_52955) );
  dffacs2 ____0________________0_ ( .DIN(____0___________0_0_____), .CLK(
        _26880), .CLRB(_____), .Q(_53503), .QN(_26364) );
  dffacs2 _______________6_ ( .DIN(
        _______6____2________________6____________________), .CLK(_26925), 
        .CLRB(_____), .Q(_53352), .QN(_26221) );
  dffacs2 _________________________________________2__18_ ( .DIN(
        _____________________________51________), .CLK(_26864), .CLRB(_____), 
        .Q(_53427) );
  dffacs2 __________________________________________3__21_ ( .DIN(
        ______________________________86________), .CLK(_26933), .CLRB(_____), 
        .Q(_53468), .QN(_26745) );
  dffacs2 _______________12_ ( .DIN(
        _______12____2________________12____________________), .CLK(_26913), 
        .CLRB(_____), .Q(_53377), .QN(_26318) );
  dffacs2 _______________31_ ( .DIN(
        _______31____2________________31____________________), .CLK(_26913), 
        .CLRB(_____), .Q(_26803), .QN(_53384) );
  dffacs2 _______________19_ ( .DIN(
        _______19____2________________19____________________), .CLK(_26911), 
        .CLRB(_____), .Q(_53517), .QN(_26323) );
  dffacs2 ____0________________13_ ( .DIN(____0___________0_13_____), .CLK(
        _26895), .CLRB(_____), .Q(_53471), .QN(_26222) );
  dffacs2 ____1________________0_0 ( .DIN(____1___________0[0]), .CLK(_26907), 
        .CLRB(_____), .Q(_26321), .QN(_2064) );
  dffacs2 ____0________________8_1 ( .DIN(____0___________[8]), .CLK(_26968), 
        .CLRB(_____), .Q(_26210), .QN(_2216) );
  dffacs1 _______________21_ ( .DIN(
        _______21____2________________21____________________), .CLK(_26893), 
        .CLRB(_____), .QN(_53371) );
  dffacs1 _______________9_ ( .DIN(
        _______9____2________________9____________________), .CLK(_26981), 
        .CLRB(_____), .QN(_53381) );
  dffacs1 _______________0_ ( .DIN(
        _______0____2________________0____________________), .CLK(_26938), 
        .CLRB(_____), .Q(_26242), .QN(_53369) );
  dffacs1 _______________28_ ( .DIN(
        _______28____2________________28____________________), .CLK(_26937), 
        .CLRB(_____), .Q(_26338), .QN(_53362) );
  dffacs1 _______________27_ ( .DIN(
        _______27____2________________27____________________), .CLK(_26937), 
        .CLRB(_____), .QN(_53361) );
  dffacs1 _______________18_ ( .DIN(
        _______18____2________________18____________________), .CLK(_26982), 
        .CLRB(_____), .QN(_53375) );
  dffacs1 _______________13_ ( .DIN(
        _______13____2________________13____________________), .CLK(_26981), 
        .CLRB(_____), .QN(_53376) );
  dffacs1 _______________10_ ( .DIN(
        _______10____2________________10____________________), .CLK(_26980), 
        .CLRB(_____), .QN(_53346) );
  dffacs1 ____0________________5_ ( .DIN(____0___________0_5_____), .CLK(
        _26973), .CLRB(_____), .Q(_26241), .QN(_53500) );
  dffacs1 ____1________________11_ ( .DIN(____1____________11_____), .CLK(
        _26927), .CLRB(_____), .Q(_26279), .QN(_53419) );
  dffacs1 __________________________________________1__2_ ( .DIN(
        ______________________________3________), .CLK(_26945), .CLRB(_____), 
        .QN(_52896) );
  dffacs1 __________________________________________1__30_ ( .DIN(
        ______________________________31________), .CLK(_26868), .CLRB(_____), 
        .Q(_26653), .QN(_52885) );
  dffacs1 _______________11_ ( .DIN(
        _______11____2________________11____________________), .CLK(_26922), 
        .CLRB(_____), .Q(_26332), .QN(_53379) );
  dffacs1 ___________________________________27_ ( .DIN(
        _________________________________27_________), .CLK(_26861), .CLRB(
        _____), .QN(_52852) );
  dffacs1 ___________________________________24_ ( .DIN(
        _________________________________24_________), .CLK(_26916), .CLRB(
        _____), .QN(_52980) );
  dffacs1 ___________________________________17_ ( .DIN(
        _________________________________17_________), .CLK(_26912), .CLRB(
        _____), .Q(_26314), .QN(_53486) );
  dffacs1 ___________________________________11_ ( .DIN(
        _________________________________11_________), .CLK(_26939), .CLRB(
        _____), .Q(_26598), .QN(_53494) );
  dffacs1 ___________________________________1_ ( .DIN(
        _________________________________1_________), .CLK(_26924), .CLRB(
        _____), .QN(_53511) );
  dffacs1 _________________________________________8__2_ ( .DIN(
        _____________________________227________), .CLK(_26924), .CLRB(_____), 
        .QN(_53116) );
  dffacs1 _________________________________________8__12_ ( .DIN(
        _____________________________237________), .CLK(_26924), .CLRB(_____), 
        .Q(_26574), .QN(_53129) );
  dffacs1 _________________________________________8__24_ ( .DIN(
        _____________________________249________), .CLK(_26862), .CLRB(_____), 
        .Q(_26410), .QN(_53415) );
  dffacs1 _________________________________________8__25_ ( .DIN(
        _____________________________250________), .CLK(_26917), .CLRB(_____), 
        .QN(_53101) );
  dffacs1 _________________________________________8__26_ ( .DIN(
        _____________________________251________), .CLK(_26918), .CLRB(_____), 
        .Q(_26482), .QN(_53172) );
  dffacs1 _________________________________________7__17_ ( .DIN(
        _____________________________210________), .CLK(_26908), .CLRB(_____), 
        .Q(_26609), .QN(_53148) );
  dffacs1 _________________________________________7__18_ ( .DIN(
        _____________________________211________), .CLK(_26957), .CLRB(_____), 
        .Q(_26648), .QN(_53217) );
  dffacs1 _________________________________________7__24_ ( .DIN(
        _____________________________217________), .CLK(_26936), .CLRB(_____), 
        .Q(_26263), .QN(_53219) );
  dffacs1 _________________________________________6__6_ ( .DIN(
        _____________________________167________), .CLK(_26935), .CLRB(_____), 
        .Q(_26716), .QN(_53214) );
  dffacs1 _________________________________________6__7_ ( .DIN(
        _____________________________168________), .CLK(_26908), .CLRB(_____), 
        .Q(_26351), .QN(_53212) );
  dffacs1 _________________________________________6__16_ ( .DIN(
        _____________________________177________), .CLK(_26919), .CLRB(_____), 
        .QN(_53202) );
  dffacs1 _________________________________________6__18_ ( .DIN(
        _____________________________179________), .CLK(_26958), .CLRB(_____), 
        .Q(_26741), .QN(_53201) );
  dffacs1 _________________________________________6__20_ ( .DIN(
        _____________________________181________), .CLK(_26958), .CLRB(_____), 
        .Q(_26489), .QN(_53198) );
  dffacs1 _________________________________________6__22_ ( .DIN(
        _____________________________183________), .CLK(_26884), .CLRB(_____), 
        .Q(_26458), .QN(_53191) );
  dffacs1 _________________________________________6__23_ ( .DIN(
        _____________________________184________), .CLK(_26948), .CLRB(_____), 
        .Q(_26643), .QN(_53270) );
  dffacs1 _________________________________________5__4_ ( .DIN(
        _____________________________133________), .CLK(_26888), .CLRB(_____), 
        .Q(_26664), .QN(_53266) );
  dffacs1 _________________________________________5__6_ ( .DIN(
        _____________________________135________), .CLK(_26889), .CLRB(_____), 
        .QN(_53257) );
  dffacs1 _________________________________________5__11_ ( .DIN(
        _____________________________140________), .CLK(_26925), .CLRB(_____), 
        .Q(_26523), .QN(_53263) );
  dffacs1 _________________________________________5__12_ ( .DIN(
        _____________________________141________), .CLK(_26919), .CLRB(_____), 
        .Q(_26671), .QN(_53262) );
  dffacs1 _________________________________________5__21_ ( .DIN(
        _____________________________150________), .CLK(_26943), .CLRB(_____), 
        .Q(_26557), .QN(_53242) );
  dffacs1 _________________________________________4__2_ ( .DIN(
        _____________________________99________), .CLK(_26881), .CLRB(_____), 
        .Q(_26678), .QN(_53343) );
  dffacs1 _________________________________________4__4_ ( .DIN(
        _____________________________101________), .CLK(_26940), .CLRB(_____), 
        .QN(_53340) );
  dffacs1 _________________________________________4__14_ ( .DIN(
        _____________________________111________), .CLK(_26942), .CLRB(_____), 
        .Q(_26555), .QN(_53304) );
  dffacs1 _________________________________________4__18_ ( .DIN(
        _____________________________115________), .CLK(_26920), .CLRB(_____), 
        .Q(_26309), .QN(_53321) );
  dffacs1 _________________________________________3__6_ ( .DIN(
        _____________________________71________), .CLK(_26890), .CLRB(_____), 
        .QN(_53337) );
  dffacs1 _________________________________________3__9_ ( .DIN(
        _____________________________74________), .CLK(_26946), .CLRB(_____), 
        .Q(_26550), .QN(_53333) );
  dffacs1 _________________________________________3__13_ ( .DIN(
        _____________________________78________), .CLK(_26947), .CLRB(_____), 
        .Q(_26545), .QN(_53313) );
  dffacs1 _________________________________________3__21_ ( .DIN(
        _____________________________86________), .CLK(_26870), .CLRB(_____), 
        .Q(_26269), .QN(_53299) );
  dffacs1 _________________________________________3__25_ ( .DIN(
        _____________________________90________), .CLK(_26870), .CLRB(_____), 
        .Q(_26423), .QN(_53291) );
  dffacs1 _________________________________________2__2_ ( .DIN(
        _____________________________35________), .CLK(_26883), .CLRB(_____), 
        .QN(_53047) );
  dffacs1 _________________________________________2__4_ ( .DIN(
        _____________________________37________), .CLK(_26856), .CLRB(_____), 
        .Q(_26232), .QN(_53048) );
  dffacs1 _________________________________________2__11_ ( .DIN(
        _____________________________44________), .CLK(_26883), .CLRB(_____), 
        .Q(_26590), .QN(_53037) );
  dffacs1 _________________________________________1__12_ ( .DIN(
        _____________________________13________), .CLK(_26949), .CLRB(_____), 
        .Q(_26521), .QN(_53252) );
  dffacs1 _________________________________________1__15_ ( .DIN(
        _____________________________16________), .CLK(_26949), .CLRB(_____), 
        .QN(_53228) );
  dffacs1 _________________________________________1__19_ ( .DIN(
        _____________________________20________), .CLK(_26983), .CLRB(_____), 
        .Q(_26244), .QN(_53196) );
  dffacs1 _________________________________________1__23_ ( .DIN(
        _____________________________24________), .CLK(_26886), .CLRB(_____), 
        .QN(_53026) );
  dffacs1 _________________________________________1__28_ ( .DIN(
        _____________________________29________), .CLK(_26874), .CLRB(_____), 
        .Q(_26253), .QN(_53102) );
  dffacs1 _________________________________________0__2_ ( .DIN(
        _________________________________________3_________), .CLK(_26935), 
        .CLRB(_____), .Q(_26399), .QN(_53318) );
  dffacs1 _________________________________________0__25_ ( .DIN(
        _________________________________________0_________), .CLK(_26954), 
        .CLRB(_____), .Q(_26451), .QN(_53354) );
  dffacs1 _________________________________________0__27_ ( .DIN(
        _________________________________________0________1____________), 
        .CLK(_26954), .CLRB(_____), .Q(_26484), .QN(_53056) );
  dffacs1 __________________________________________5__0_ ( .DIN(
        ______________________________129________), .CLK(_26956), .CLRB(_____), 
        .QN(_52951) );
  dffacs1 __________________________________________5__2_ ( .DIN(
        ______________________________131________), .CLK(_26956), .CLRB(_____), 
        .Q(_26392), .QN(_52950) );
  dffacs1 __________________________________________5__8_ ( .DIN(
        ______________________________137________), .CLK(_26965), .CLRB(_____), 
        .QN(_52939) );
  dffacs1 __________________________________________5__11_ ( .DIN(
        ______________________________140________), .CLK(_26966), .CLRB(_____), 
        .QN(_52948) );
  dffacs1 __________________________________________5__14_ ( .DIN(
        ______________________________143________), .CLK(_26878), .CLRB(_____), 
        .Q(_26354), .QN(_52940) );
  dffacs1 __________________________________________5__17_ ( .DIN(
        ______________________________146________), .CLK(_26920), .CLRB(_____), 
        .Q(_26662), .QN(_52937) );
  dffacs1 __________________________________________5__21_ ( .DIN(
        ______________________________150________), .CLK(_26979), .CLRB(_____), 
        .Q(_26522), .QN(_52935) );
  dffacs1 __________________________________________5__29_ ( .DIN(
        ______________________________158________), .CLK(_26893), .CLRB(_____), 
        .Q(_26584), .QN(_52932) );
  dffacs1 __________________________________________3__13_ ( .DIN(
        ______________________________78________), .CLK(_26977), .CLRB(_____), 
        .Q(_26700), .QN(_52985) );
  dffacs1 __________________________________________3__17_ ( .DIN(
        ______________________________82________), .CLK(_26978), .CLRB(_____), 
        .Q(_26226) );
  dffacs1 __________________________________________3__18_ ( .DIN(
        ______________________________83________), .CLK(_26869), .CLRB(_____), 
        .Q(_26388), .QN(_52977) );
  dffacs1 __________________________________________3__22_ ( .DIN(
        ______________________________87________), .CLK(_26922), .CLRB(_____), 
        .Q(_26257), .QN(_52969) );
  dffacs1 __________________________________________1__1_ ( .DIN(
        ______________________________2________), .CLK(_26869), .CLRB(_____), 
        .Q(_26360), .QN(_52880) );
  dffacs1 __________________________________________1__5_ ( .DIN(
        ______________________________6________), .CLK(_26944), .CLRB(_____), 
        .Q(_26301), .QN(_52965) );
  dffacs1 __________________________________________1__23_ ( .DIN(
        ______________________________24________), .CLK(_26860), .CLRB(_____), 
        .Q(_26389), .QN(_52893) );
  dffacs1 __________________________________________1__25_ ( .DIN(
        ______________________________26________), .CLK(_26892), .CLRB(_____), 
        .QN(_52889) );
  dffacs1 __________________________________________1__26_ ( .DIN(
        ______________________________27________), .CLK(_26976), .CLRB(_____), 
        .Q(_26655), .QN(_52891) );
  dffacs1 __________________________________________1__27_ ( .DIN(
        ______________________________28________), .CLK(_26892), .CLRB(_____), 
        .Q(_26752), .QN(_52890) );
  dffacs1 __________________________________________1__31_ ( .DIN(
        ______________________________32________), .CLK(_26886), .CLRB(_____), 
        .Q(_26618), .QN(_53359) );
  dffacs1 ____________________________________19_ ( .DIN(
        __________________________________19_________), .CLK(_26976), .CLRB(
        _____), .Q(_26726), .QN(_53485) );
  dffacs1 _______________29_ ( .DIN(
        _______29____2________________29____________________), .CLK(_26886), 
        .CLRB(_____), .QN(_53364) );
  dffacs1 _________________________________________9__1_ ( .DIN(
        _____________________________258________), .CLK(_26930), .CLRB(_____), 
        .Q(_26701), .QN(_53090) );
  dffacs1 _________________________________________9__4_ ( .DIN(
        _____________________________261________), .CLK(_26930), .CLRB(_____), 
        .Q(_26355) );
  dffacs1 _________________________________________9__5_ ( .DIN(
        _____________________________262________), .CLK(_26931), .CLRB(_____), 
        .Q(_26256), .QN(_53091) );
  dffacs1 _________________________________________9__10_ ( .DIN(
        _____________________________267________), .CLK(_26896), .CLRB(_____), 
        .QN(_53081) );
  dffacs1 _________________________________________9__15_ ( .DIN(
        _____________________________272________), .CLK(_26940), .CLRB(_____), 
        .QN(_53078) );
  dffacs1 _________________________________________9__27_ ( .DIN(
        _____________________________284________), .CLK(_26861), .CLRB(_____), 
        .Q(_26623) );
  dffacs1 _________________________________________9__30_ ( .DIN(
        _____________________________287________), .CLK(_26951), .CLRB(_____), 
        .QN(_53062) );
  dffacs1 __________________________________________6__1_ ( .DIN(
        ______________________________162________), .CLK(_26929), .CLRB(_____), 
        .Q(_26612), .QN(_53061) );
  dffacs1 __________________________________________4__1_ ( .DIN(
        ______________________________98________), .CLK(_26929), .CLRB(_____), 
        .Q(_26622), .QN(_52953) );
  dffacs1 __________________________________________6__7_ ( .DIN(
        ______________________________168________), .CLK(_26906), .CLRB(_____), 
        .Q(_26614), .QN(_52831) );
  dffacs1 __________________________________________6__11_ ( .DIN(
        ______________________________172________), .CLK(_26877), .CLRB(_____), 
        .QN(_52921) );
  dffacs1 __________________________________________6__12_ ( .DIN(
        ______________________________173________), .CLK(_26877), .CLRB(_____), 
        .Q(_26395), .QN(_52916) );
  dffacs1 __________________________________________6__18_ ( .DIN(
        ______________________________179________), .CLK(_26915), .CLRB(_____), 
        .Q(_26670), .QN(_52911) );
  dffacs1 __________________________________________6__24_ ( .DIN(
        ______________________________185________), .CLK(_26866), .CLRB(_____), 
        .Q(_26282), .QN(_52910) );
  dffacs1 __________________________________________6__27_ ( .DIN(
        ______________________________188________), .CLK(_26867), .CLRB(_____), 
        .QN(_52903) );
  dffacs1 __________________________________________4__2_ ( .DIN(
        ______________________________99________), .CLK(_26956), .CLRB(_____), 
        .QN(_53005) );
  dffacs1 __________________________________________4__20_ ( .DIN(
        ______________________________117________), .CLK(_26916), .CLRB(_____), 
        .Q(_26271), .QN(_52975) );
  dffacs1 __________________________________________4__21_ ( .DIN(
        ______________________________118________), .CLK(_26921), .CLRB(_____), 
        .Q(_26705), .QN(_52973) );
  dffacs1 __________________________________________4__25_ ( .DIN(
        ______________________________122________), .CLK(_26941), .CLRB(_____), 
        .QN(_52963) );
  dffacs1 __________________________________________4__29_ ( .DIN(
        ______________________________126________), .CLK(_26894), .CLRB(_____), 
        .Q(_26461), .QN(_52960) );
  dffacs1 __________________________________________2__0_ ( .DIN(
        ______________________________33________), .CLK(_26872), .CLRB(_____), 
        .QN(_52876) );
  dffacs1 __________________________________________2__5_ ( .DIN(
        ______________________________38________), .CLK(_26872), .CLRB(_____), 
        .Q(_26608), .QN(_52873) );
  dffacs1 __________________________________________2__6_ ( .DIN(
        ______________________________39________), .CLK(_26872), .CLRB(_____), 
        .Q(_26426) );
  dffacs1 __________________________________________2__8_ ( .DIN(
        ______________________________41________), .CLK(_26873), .CLRB(_____), 
        .QN(_52833) );
  dffacs1 __________________________________________2__10_ ( .DIN(
        ______________________________43________), .CLK(_26887), .CLRB(_____), 
        .Q(_26588), .QN(_52870) );
  dffacs1 __________________________________________2__14_ ( .DIN(
        ______________________________47________), .CLK(_26857), .CLRB(_____), 
        .QN(_52868) );
  dffacs1 __________________________________________2__21_ ( .DIN(
        ______________________________54________), .CLK(_26933), .CLRB(_____), 
        .Q(_26293), .QN(_52865) );
  dffacs1 __________________________________________2__24_ ( .DIN(
        ______________________________57________), .CLK(_26945), .CLRB(_____), 
        .QN(_52861) );
  dffacs1 __________________________________________0__2_ ( .DIN(
        __________________________________________2_________), .CLK(_26986), 
        .CLRB(_____), .QN(_52872) );
  dffacs1 __________________________________________0__7_ ( .DIN(
        __________________________________________7_________), .CLK(_26986), 
        .CLRB(_____), .Q(_26620), .QN(_52854) );
  dffacs1 __________________________________________0__14_ ( .DIN(
        __________________________________________14_________), .CLK(_26986), 
        .CLRB(_____), .QN(_52929) );
  dffacs1 __________________________________________0__17_ ( .DIN(
        __________________________________________17_________), .CLK(_26866), 
        .CLRB(_____), .Q(_26264), .QN(_52840) );
  dffacs1 __________________________________________0__23_ ( .DIN(
        __________________________________________23_________), .CLK(_26951), 
        .CLRB(_____), .Q(_26494), .QN(_52892) );
  dffacs1 __________________________________________0__8_ ( .DIN(
        __________________________________________8_________), .CLK(_26901), 
        .CLRB(_____), .Q(_26308), .QN(_53389) );
  dffacs1 ____3________________1_ ( .DIN(____3____________1_____), .CLK(_26901), .CLRB(_____), .Q(_26286), .QN(_53438) );
  dffacs1 ____1________________4_ ( .DIN(____1____________4_____), .CLK(_26961), .CLRB(_____), .Q(_26585), .QN(_53460) );
  dffacs1 ____0________________0_0 ( .DIN(____0____________0_____), .CLK(
        _26870), .CLRB(_____), .Q(_26428), .QN(_53451) );
  dffacs1 ____0________________11_0 ( .DIN(____0____________11_____), .CLK(
        _26902), .CLRB(_____), .Q(_26214), .QN(_53459) );
  dffacs1 ____0________________6_0 ( .DIN(____0____________6_____), .CLK(
        _26902), .CLRB(_____), .Q(_26243), .QN(_53458) );
  dffacs1 ____0________________7_0 ( .DIN(____0____________7_____), .CLK(
        _26977), .CLRB(_____), .Q(_26387), .QN(_53447) );
  dffacs1 ____0________________3_0 ( .DIN(____0____________3_____), .CLK(
        _26977), .CLRB(_____), .Q(_26215), .QN(_53446) );
  dffacs1 ____0________________9_0 ( .DIN(____0____________9_____), .CLK(
        _26911), .CLRB(_____), .Q(_26262), .QN(_53456) );
  dffacs1 ____1________________8_ ( .DIN(____1____________8_____), .CLK(_26859), .CLRB(_____), .Q(_26212), .QN(_53425) );
  dffacs1 ____1________________2_ ( .DIN(____1____________2_____), .CLK(_26980), .CLRB(_____), .Q(_26275), .QN(_53422) );
  dffacs1 ____1________________5_ ( .DIN(____1____________5_____), .CLK(_26980), .CLRB(_____), .Q(_26285), .QN(_53424) );
  dffacs1 ____1________________7_ ( .DIN(____1____________7_____), .CLK(_26980), .CLRB(_____), .Q(_26699), .QN(_53416) );
  dffacs1 ____1________________10_ ( .DIN(____1____________10_____), .CLK(
        _26980), .CLRB(_____), .Q(_26539), .QN(_53418) );
  dffacs1 ____1________________1_ ( .DIN(____1____________1_____), .CLK(_26885), .CLRB(_____), .Q(_26298), .QN(_53420) );
  dffacs1 ____2________________10_ ( .DIN(____2____________10_____), .CLK(
        _26982), .CLRB(_____), .Q(_26274), .QN(_53414) );
  dffacs1 ____2________________7_ ( .DIN(____2____________7_____), .CLK(_26875), .CLRB(_____), .Q(_26283), .QN(_53400) );
  dffacs1 ____2________________11_ ( .DIN(____2____________11_____), .CLK(
        _26982), .CLRB(_____), .Q(_26443), .QN(_53401) );
  dffacs1 ____2________________12_ ( .DIN(____2____________12_____), .CLK(
        _26883), .CLRB(_____), .QN(_53408) );
  dffacs1 _________________________________________6__29_ ( .DIN(
        _____________________________190________), .CLK(_26889), .CLRB(_____), 
        .Q(_26681), .QN(_53140) );
  dffacs1 _________________________________________4__23_ ( .DIN(
        _____________________________120________), .CLK(_26948), .CLRB(_____), 
        .Q(_26445), .QN(_53281) );
  dffacs1 _________________________________________4__30_ ( .DIN(
        _____________________________127________), .CLK(_26885), .CLRB(_____), 
        .Q(_26213) );
  dffacs1 _________________________________________1__6_ ( .DIN(
        _____________________________7________), .CLK(_26925), .CLRB(_____), 
        .Q(_26259), .QN(_53039) );
  dffacs1 __________________________________________3__12_ ( .DIN(
        ______________________________77________), .CLK(_26960), .CLRB(_____), 
        .Q(_26525), .QN(_53030) );
  dffacs1 __________________________________________1__7_ ( .DIN(
        ______________________________8________), .CLK(_26960), .CLRB(_____), 
        .QN(_52871) );
  dffacs1 ____________________________________18_ ( .DIN(
        __________________________________18_________), .CLK(_26976), .CLRB(
        _____), .Q(_26680), .QN(_52990) );
  dffacs1 ___________________________________26_ ( .DIN(
        _________________________________26_________), .CLK(_26899), .CLRB(
        _____), .Q(_26604), .QN(_53176) );
  dffacs1 ___________________________________23_ ( .DIN(
        _________________________________23_________), .CLK(_26916), .CLRB(
        _____), .Q(_26477), .QN(_53504) );
  dffacs1 _________________________________________8__30_ ( .DIN(
        _____________________________255________), .CLK(_26916), .CLRB(_____), 
        .Q(_26514), .QN(_53097) );
  dffacs1 _________________________________________7__29_ ( .DIN(
        _____________________________222________), .CLK(_26916), .CLRB(_____), 
        .QN(_53225) );
  dffacs1 __________________________________________3__25_ ( .DIN(
        ______________________________90________), .CLK(_26985), .CLRB(_____), 
        .Q(_26235), .QN(_53163) );
  dffacs1 __________________________________________1__17_ ( .DIN(
        ______________________________18________), .CLK(_26985), .CLRB(_____), 
        .QN(_53162) );
  dffacs1 _________________________________________7__8_ ( .DIN(
        _____________________________201________), .CLK(_26985), .CLRB(_____), 
        .Q(_26463), .QN(_53154) );
  dffacs1 _________________________________________7__20_ ( .DIN(
        _____________________________213________), .CLK(_26903), .CLRB(_____), 
        .Q(_26460), .QN(_53143) );
  dffacs1 __________________________________________1__16_ ( .DIN(
        ______________________________17________), .CLK(_26932), .CLRB(_____), 
        .Q(_26486), .QN(_53144) );
  dffacs1 ___________________________________30_ ( .DIN(
        _________________________________30_________), .CLK(_26938), .CLRB(
        _____), .QN(_52851) );
  dffacs1 ___________________________________20_ ( .DIN(
        _________________________________20_________), .CLK(_26894), .CLRB(
        _____), .QN(_53483) );
  dffacs1 ___________________________________19_ ( .DIN(
        _________________________________19_________), .CLK(_26931), .CLRB(
        _____), .Q(_26393), .QN(_53484) );
  dffacs1 _________________________________________5__10_ ( .DIN(
        _____________________________139________), .CLK(_26890), .CLRB(_____), 
        .Q(_26651), .QN(_53271) );
  dffacs1 _________________________________________3__11_ ( .DIN(
        _____________________________76________), .CLK(_26889), .CLRB(_____), 
        .Q(_26520), .QN(_53327) );
  dffacs1 _________________________________________3__12_ ( .DIN(
        _____________________________77________), .CLK(_26959), .CLRB(_____), 
        .Q(_26267), .QN(_53320) );
  dffacs1 _________________________________________2__17_ ( .DIN(
        _____________________________50________), .CLK(_26959), .CLRB(_____), 
        .Q(_26380) );
  dffacs1 _________________________________________1__5_ ( .DIN(
        _____________________________6________), .CLK(_26913), .CLRB(_____), 
        .Q(_26673), .QN(_53041) );
  dffacs1 _________________________________________1__10_ ( .DIN(
        _____________________________11________), .CLK(_26935), .CLRB(_____), 
        .Q(_26650), .QN(_53035) );
  dffacs1 _________________________________________0__23_ ( .DIN(
        _________________________________________24_________), .CLK(_26886), 
        .CLRB(_____), .Q(_26657), .QN(_53103) );
  dffacs1 _________________________________________7__16_ ( .DIN(
        _____________________________209________), .CLK(_26957), .CLRB(_____), 
        .Q(_26661), .QN(_53111) );
  dffacs1 _________________________________________6__13_ ( .DIN(
        _____________________________174________), .CLK(_26919), .CLRB(_____), 
        .Q(_26504), .QN(_53200) );
  dffacs1 __________________________________________1__20_ ( .DIN(
        ______________________________21________), .CLK(_26950), .CLRB(_____), 
        .QN(_52930) );
  dffacs1 ____________________________________1_ ( .DIN(
        __________________________________1_________), .CLK(_26929), .CLRB(
        _____), .QN(_52844) );
  dffacs1 _________________________________________6__19_ ( .DIN(
        _____________________________180________), .CLK(_26958), .CLRB(_____), 
        .Q(_26261), .QN(_53150) );
  dffacs1 _________________________________________6__31_ ( .DIN(
        _____________________________192________), .CLK(_26903), .CLRB(_____), 
        .Q(_26524), .QN(_53136) );
  dffacs1 __________________________________________6__10_ ( .DIN(
        ______________________________171________), .CLK(_26912), .CLRB(_____), 
        .QN(_52920) );
  dffacs1 ___________________________________29_ ( .DIN(
        _________________________________29_________), .CLK(_26938), .CLRB(
        _____), .QN(_52971) );
  dffacs1 __________________________________________5__30_ ( .DIN(
        ______________________________159________), .CLK(_26938), .CLRB(_____), 
        .Q(_26472), .QN(_53279) );
  dffacs1 _________________________________________4__31_ ( .DIN(
        _____________________________128________), .CLK(_26903), .CLRB(_____), 
        .Q(_26300), .QN(_53226) );
  dffacs1 __________________________________________3__24_ ( .DIN(
        ______________________________89________), .CLK(_26899), .CLRB(_____), 
        .Q(_26512), .QN(_53009) );
  dffacs1 _________________________________________2__31_ ( .DIN(
        _____________________________64________), .CLK(_26900), .CLRB(_____), 
        .Q(_26487), .QN(_53050) );
  dffacs1 _________________________________________7__30_ ( .DIN(
        _____________________________223________), .CLK(_26889), .CLRB(_____), 
        .Q(_26629), .QN(_53224) );
  dffacs1 _________________________________________4__0_ ( .DIN(
        _____________________________97________), .CLK(_26899), .CLRB(_____), 
        .QN(_53275) );
  dffacs1 ___________________________________13_ ( .DIN(
        _________________________________13_________), .CLK(_26858), .CLRB(
        _____), .Q(_26546), .QN(_52999) );
  dffacs1 _________________________________________1__30_ ( .DIN(
        _____________________________31________), .CLK(_26902), .CLRB(_____), 
        .Q(_26663), .QN(_53018) );
  dffacs1 __________________________________________3__6_ ( .DIN(
        ______________________________71________), .CLK(_26872), .CLRB(_____), 
        .Q(_26405), .QN(_53095) );
  dffacs1 _________________________________________8__16_ ( .DIN(
        _____________________________241________), .CLK(_26957), .CLRB(_____), 
        .QN(_53131) );
  dffacs1 _________________________________________0__30_ ( .DIN(
        _________________________________________0________4____________), 
        .CLK(_26961), .CLRB(_____), .Q(_26690), .QN(_53132) );
  dffacs1 _________________________________________0__0_ ( .DIN(
        _________________________________________1_________), .CLK(_26961), 
        .CLRB(_____), .QN(_53319) );
  dffacs1 _________________________________________0__9_ ( .DIN(
        _________________________________________10_________), .CLK(_26914), 
        .CLRB(_____), .Q(_26462), .QN(_53316) );
  dffacs1 _________________________________________8__7_ ( .DIN(
        _____________________________232________), .CLK(_26915), .CLRB(_____), 
        .Q(_26230) );
  dffacs1 _________________________________________3__30_ ( .DIN(
        _____________________________95________), .CLK(_26900), .CLRB(_____), 
        .Q(_26367), .QN(_53280) );
  dffacs1 _________________________________________6__27_ ( .DIN(
        _____________________________188________), .CLK(_26898), .CLRB(_____), 
        .QN(_53186) );
  dffacs1 ___________________________________22_ ( .DIN(
        _________________________________22_________), .CLK(_26974), .CLRB(
        _____), .QN(_53184) );
  dffacs1 _________________________________________7__2_ ( .DIN(
        _____________________________195________), .CLK(_26937), .CLRB(_____), 
        .QN(_53356) );
  dffacs1 _________________________________________8__17_ ( .DIN(
        _____________________________242________), .CLK(_26908), .CLRB(_____), 
        .Q(_26449), .QN(_53355) );
  dffacs1 ____________________________________20_ ( .DIN(
        __________________________________20_________), .CLK(_26955), .CLRB(
        _____), .Q(_26702), .QN(_52846) );
  dffacs1 ____________________________________17_ ( .DIN(
        __________________________________17_________), .CLK(_26954), .CLRB(
        _____), .Q(_26291), .QN(_53487) );
  dffacs1 ____________________________________16_ ( .DIN(
        __________________________________16_________), .CLK(_26954), .CLRB(
        _____), .QN(_52845) );
  dffacs1 _________________________________________9__29_ ( .DIN(
        _____________________________286________), .CLK(_26963), .CLRB(_____), 
        .QN(_53060) );
  dffacs1 _________________________________________9__28_ ( .DIN(
        _____________________________285________), .CLK(_26922), .CLRB(_____), 
        .QN(_53059) );
  dffacs1 __________________________________________4__9_ ( .DIN(
        ______________________________106________), .CLK(_26877), .CLRB(_____), 
        .Q(_26492), .QN(_52993) );
  dffacs1 __________________________________________0__5_ ( .DIN(
        __________________________________________5_________), .CLK(_26874), 
        .CLRB(_____), .QN(_52838) );
  dffacs1 __________________________________________2__25_ ( .DIN(
        ______________________________58________), .CLK(_26985), .CLRB(_____), 
        .Q(_26299), .QN(_52991) );
  dffacs1 __________________________________________6__19_ ( .DIN(
        ______________________________180________), .CLK(_26874), .CLRB(_____), 
        .QN(_52905) );
  dffacs1 _________________________________________9__14_ ( .DIN(
        _____________________________271________), .CLK(_26858), .CLRB(_____), 
        .QN(_53074) );
  dffacs1 _________________________________________2__29_ ( .DIN(
        _____________________________62________), .CLK(_26856), .CLRB(_____), 
        .QN(_53054) );
  dffacs1 __________________________________________5__27_ ( .DIN(
        ______________________________156________), .CLK(_26857), .CLRB(_____), 
        .QN(_53019) );
  dffacs1 ____________________________________11_ ( .DIN(
        __________________________________11_________), .CLK(_26927), .CLRB(
        _____), .Q(_26755), .QN(_52843) );
  dffacs1 ____________________________________8_ ( .DIN(
        __________________________________8_________), .CLK(_26928), .CLRB(
        _____), .Q(_26411), .QN(_53497) );
  dffacs1 __________________________________________5__4_ ( .DIN(
        ______________________________133________), .CLK(_26953), .CLRB(_____), 
        .QN(_52922) );
  dffacs1 __________________________________________5__20_ ( .DIN(
        ______________________________149________), .CLK(_26978), .CLRB(_____), 
        .Q(_26302), .QN(_52906) );
  dffacs1 _________________________________________9__18_ ( .DIN(
        _____________________________275________), .CLK(_26940), .CLRB(_____), 
        .QN(_53082) );
  dffacs1 _________________________________________9__22_ ( .DIN(
        _____________________________279________), .CLK(_26862), .CLRB(_____), 
        .Q(_26586), .QN(_53083) );
  dffacs1 __________________________________________6__2_ ( .DIN(
        ______________________________163________), .CLK(_26928), .CLRB(_____), 
        .QN(_53238) );
  dffacs1 _________________________________________5__22_ ( .DIN(
        _____________________________151________), .CLK(_26884), .CLRB(_____), 
        .QN(_53190) );
  dffacs1 _________________________________________4__20_ ( .DIN(
        _____________________________117________), .CLK(_26959), .CLRB(_____), 
        .QN(_53300) );
  dffacs1 _________________________________________4__24_ ( .DIN(
        _____________________________121________), .CLK(_26973), .CLRB(_____), 
        .QN(_53236) );
  dffacs1 _________________________________________1__9_ ( .DIN(
        _____________________________10________), .CLK(_26935), .CLRB(_____), 
        .QN(_53036) );
  dffacs1 __________________________________________5__9_ ( .DIN(
        ______________________________138________), .CLK(_26963), .CLRB(_____), 
        .QN(_53292) );
  dffacs1 __________________________________________2__16_ ( .DIN(
        ______________________________49________), .CLK(_26926), .CLRB(_____), 
        .QN(_52867) );
  dffacs1 __________________________________________3__15_ ( .DIN(
        ______________________________80________), .CLK(_26926), .CLRB(_____), 
        .QN(_52982) );
  dffacs1 ____________________________________5_ ( .DIN(
        __________________________________5_________), .CLK(_26867), .CLRB(
        _____), .Q(_26454), .QN(_53513) );
  dffacs1 __________________________________________4__13_ ( .DIN(
        ______________________________110________), .CLK(_26912), .CLRB(_____), 
        .QN(_53000) );
  dffacs1 __________________________________________4__17_ ( .DIN(
        ______________________________114________), .CLK(_26912), .CLRB(_____), 
        .Q(_26711), .QN(_52984) );
  dffacs1 __________________________________________0__31_ ( .DIN(
        __________________________________________25________5____________), 
        .CLK(_26962), .CLRB(_____), .QN(_52979) );
  dffacs1 __________________________________________2__4_ ( .DIN(
        ______________________________37________), .CLK(_26879), .CLRB(_____), 
        .QN(_52878) );
  dffacs1 __________________________________________6__26_ ( .DIN(
        ______________________________187________), .CLK(_26910), .CLRB(_____), 
        .Q(_26679), .QN(_52834) );
  dffacs1 _________________________________________4__16_ ( .DIN(
        _____________________________113________), .CLK(_26879), .CLRB(_____), 
        .Q(_26757), .QN(_53248) );
  dffacs1 __________________________________________0__24_ ( .DIN(
        __________________________________________24_________), .CLK(_26946), 
        .CLRB(_____), .QN(_53311) );
  dffacs1 __________________________________________3__8_ ( .DIN(
        ______________________________73________), .CLK(_26945), .CLRB(_____), 
        .QN(_52994) );
  dffacs1 __________________________________________4__30_ ( .DIN(
        ______________________________127________), .CLK(_26898), .CLRB(_____), 
        .QN(_53181) );
  dffacs1 __________________________________________6__14_ ( .DIN(
        ______________________________175________), .CLK(_26878), .CLRB(_____), 
        .QN(_53182) );
  dffacs1 _________________________________________6__28_ ( .DIN(
        _____________________________189________), .CLK(_26898), .CLRB(_____), 
        .QN(_53185) );
  dffacs1 ____3________________8_ ( .DIN(____3____________8_____), .CLK(_26876), .CLRB(_____), .Q(_26228), .QN(_53441) );
  dffacs1 __________________________________________4__6_ ( .DIN(
        ______________________________103________), .CLK(_26876), .CLRB(_____), 
        .Q(_26493), .QN(_53382) );
  dffacs1 __________________________________________6__29_ ( .DIN(
        ______________________________190________), .CLK(_26893), .CLRB(_____), 
        .QN(_52902) );
  dffacs1 __________________________________________4__15_ ( .DIN(
        ______________________________112________), .CLK(_26878), .CLRB(_____), 
        .QN(_52836) );
  dffacs1 ___________________________________21_ ( .DIN(
        _________________________________21_________), .CLK(_26974), .CLRB(
        _____), .Q(_26457), .QN(_53482) );
  dffacs1 _________________________________________9__16_ ( .DIN(
        _____________________________273________), .CLK(_26957), .CLRB(_____), 
        .Q(_26708), .QN(_53073) );
  dffacs1 ____________________________________22_ ( .DIN(
        __________________________________22_________), .CLK(_26873), .CLRB(
        _____), .Q(_26435), .QN(_53480) );
  dffacs1 _________________________________________3__17_ ( .DIN(
        _____________________________82________), .CLK(_26959), .CLRB(_____), 
        .Q(_26403), .QN(_53306) );
  dffacs1 _________________________________________1__24_ ( .DIN(
        _____________________________25________), .CLK(_26950), .CLRB(_____), 
        .Q(_26480), .QN(_53114) );
  dffacs1 __________________________________________3__4_ ( .DIN(
        ______________________________69________), .CLK(_26878), .CLRB(_____), 
        .QN(_53001) );
  dffacs1 _________________________________________2__28_ ( .DIN(
        _____________________________61________), .CLK(_26878), .CLRB(_____), 
        .Q(_26617), .QN(_53021) );
  dffacs1 __________________________________________5__6_ ( .DIN(
        ______________________________135________), .CLK(_26952), .CLRB(_____), 
        .QN(_53020) );
  dffacs1 _________________________________________5__28_ ( .DIN(
        _____________________________157________), .CLK(_26888), .CLRB(_____), 
        .Q(_26292), .QN(_53234) );
  dffacs1 _________________________________________3__3_ ( .DIN(
        _____________________________68________), .CLK(_26865), .CLRB(_____), 
        .Q(_26519), .QN(_53347) );
  dffacs1 _________________________________________4__26_ ( .DIN(
        _____________________________123________), .CLK(_26910), .CLRB(_____), 
        .Q(_26682), .QN(_53235) );
  dffacs1 __________________________________________2__9_ ( .DIN(
        ______________________________42________), .CLK(_26944), .CLRB(_____), 
        .Q(_26704), .QN(_52987) );
  dffacs1 ____3________________0_ ( .DIN(____3____________0_____), .CLK(_26876), .CLRB(_____), .Q(_26587), .QN(_53439) );
  dffacs1 _________________________________________7__3_ ( .DIN(
        _____________________________196________), .CLK(_26917), .CLRB(_____), 
        .Q(_26386), .QN(_53391) );
  dffacs1 _________________________________________6__17_ ( .DIN(
        _____________________________178________), .CLK(_26917), .CLRB(_____), 
        .Q(_26381) );
  dffacs1 _________________________________________5__18_ ( .DIN(
        _____________________________147________), .CLK(_26958), .CLRB(_____), 
        .Q(_26734), .QN(_53197) );
  dffacs1 _________________________________________4__7_ ( .DIN(
        _____________________________104________), .CLK(_26891), .CLRB(_____), 
        .Q(_26503), .QN(_53261) );
  dffacs1 _________________________________________3__24_ ( .DIN(
        _____________________________89________), .CLK(_26891), .CLRB(_____), 
        .Q(_26570), .QN(_53293) );
  dffacs1 _________________________________________2__9_ ( .DIN(
        _____________________________42________), .CLK(_26947), .CLRB(_____), 
        .Q(_26287), .QN(_53244) );
  dffacs1 _________________________________________2__13_ ( .DIN(
        _____________________________46________), .CLK(_26960), .CLRB(_____), 
        .QN(_53113) );
  dffacs1 __________________________________________1__28_ ( .DIN(
        ______________________________29________), .CLK(_26868), .CLRB(_____), 
        .QN(_53106) );
  dffacs1 _________________________________________2__20_ ( .DIN(
        _____________________________53________), .CLK(_26947), .CLRB(_____), 
        .QN(_53029) );
  dffacs1 _________________________________________8__19_ ( .DIN(
        _____________________________244________), .CLK(_26868), .CLRB(_____), 
        .QN(_53071) );
  dffacs1 _________________________________________5__20_ ( .DIN(
        _____________________________149________), .CLK(_26958), .CLRB(_____), 
        .QN(_53240) );
  dffacs1 _________________________________________4__27_ ( .DIN(
        _____________________________124________), .CLK(_26885), .CLRB(_____), 
        .Q(_26394), .QN(_53285) );
  dffacs1 _________________________________________2__3_ ( .DIN(
        _____________________________36________), .CLK(_26885), .CLRB(_____), 
        .Q(_26658), .QN(_53287) );
  dffacs1 __________________________________________5__13_ ( .DIN(
        ______________________________142________), .CLK(_26962), .CLRB(_____), 
        .Q(_26548), .QN(_52943) );
  dffacs1 __________________________________________3__2_ ( .DIN(
        ______________________________67________), .CLK(_26962), .CLRB(_____), 
        .Q(_26537), .QN(_53007) );
  dffacs1 __________________________________________2__1_ ( .DIN(
        ______________________________34________), .CLK(_26909), .CLRB(_____), 
        .Q(_26621), .QN(_52912) );
  dffacs1 __________________________________________4__11_ ( .DIN(
        ______________________________108________), .CLK(_26909), .CLRB(_____), 
        .Q(_26634), .QN(_53433) );
  dffacs1 _________________________________________9__12_ ( .DIN(
        _____________________________269________), .CLK(_26858), .CLRB(_____), 
        .Q(_26516), .QN(_53121) );
  dffacs1 _________________________________________8__10_ ( .DIN(
        _____________________________235________), .CLK(_26858), .CLRB(_____), 
        .Q(_26720), .QN(_53120) );
  dffacs1 __________________________________________2__15_ ( .DIN(
        ______________________________48________), .CLK(_26926), .CLRB(_____), 
        .Q(_26442), .QN(_53094) );
  dffacs1 __________________________________________2__7_ ( .DIN(
        ______________________________40________), .CLK(_26872), .CLRB(_____), 
        .QN(_52875) );
  dffacs1 _________________________________________9__0_ ( .DIN(
        _____________________________257________), .CLK(_26925), .CLRB(_____), 
        .Q(_26406), .QN(_53351) );
  dffacs1 _________________________________________9__3_ ( .DIN(
        _____________________________260________), .CLK(_26929), .CLRB(_____), 
        .Q(_26239), .QN(_53394) );
  dffacs1 ____2________________4_ ( .DIN(____2____________4_____), .CLK(_26864), .CLRB(_____), .Q(_26578), .QN(_53409) );
  dffacs1 ___________________________________8_ ( .DIN(
        _________________________________8_________), .CLK(_26864), .CLRB(
        _____), .Q(_26747), .QN(_52850) );
  dffacs1 _________________________________________4__3_ ( .DIN(
        _____________________________100________), .CLK(_26864), .CLRB(_____), 
        .Q(_26668), .QN(_53349) );
  dffacs1 _________________________________________3__4_ ( .DIN(
        _____________________________69________), .CLK(_26984), .CLRB(_____), 
        .Q(_26490), .QN(_53341) );
  dffacs1 _________________________________________5__5_ ( .DIN(
        _____________________________134________), .CLK(_26888), .CLRB(_____), 
        .QN(_53268) );
  dffacs1 _________________________________________5__29_ ( .DIN(
        _____________________________158________), .CLK(_26888), .CLRB(_____), 
        .QN(_53267) );
  dffacs1 ___________________________________28_ ( .DIN(
        _________________________________28_________), .CLK(_26934), .CLRB(
        _____), .Q(_26756), .QN(_52972) );
  dffacs1 _________________________________________7__11_ ( .DIN(
        _____________________________204________), .CLK(_26984), .CLRB(_____), 
        .QN(_53157) );
  dffacs1 _________________________________________7__28_ ( .DIN(
        _____________________________221________), .CLK(_26897), .CLRB(_____), 
        .Q(_26455), .QN(_53155) );
  dffacs1 _________________________________________6__21_ ( .DIN(
        _____________________________182________), .CLK(_26943), .CLRB(_____), 
        .QN(_53232) );
  dffacs1 _________________________________________1__14_ ( .DIN(
        _____________________________15________), .CLK(_26861), .CLRB(_____), 
        .QN(_53231) );
  dffacs1 ____2________________3_ ( .DIN(____2____________3_____), .CLK(_26883), .CLRB(_____), .Q(_26707), .QN(_53410) );
  dffacs1 _________________________________________4__6_ ( .DIN(
        _____________________________103________), .CLK(_26890), .CLRB(_____), 
        .Q(_26357) );
  dffacs1 _________________________________________7__19_ ( .DIN(
        _____________________________212________), .CLK(_26958), .CLRB(_____), 
        .QN(_53147) );
  dffacs1 _________________________________________2__24_ ( .DIN(
        _____________________________57________), .CLK(_26891), .CLRB(_____), 
        .Q(_26485), .QN(_53149) );
  dffacs1 __________________________________________0__25_ ( .DIN(
        __________________________________________25_________), .CLK(_26892), 
        .CLRB(_____), .QN(_52888) );
  dffacs1 __________________________________________4__14_ ( .DIN(
        ______________________________111________), .CLK(_26878), .CLRB(_____), 
        .Q(_26270), .QN(_53055) );
  dffacs1 __________________________________________0__1_ ( .DIN(
        __________________________________________1_________), .CLK(_26874), 
        .CLRB(_____), .Q(_26753), .QN(_52837) );
  dffacs1 _________________________________________9__31_ ( .DIN(
        _____________________________288________), .CLK(_26923), .CLRB(_____), 
        .Q(_26712), .QN(_53137) );
  dffacs1 _________________________________________6__8_ ( .DIN(
        _____________________________169________), .CLK(_26930), .CLRB(_____), 
        .QN(_53210) );
  dffacs1 _________________________________________1__13_ ( .DIN(
        _____________________________14________), .CLK(_26949), .CLRB(_____), 
        .QN(_53034) );
  dffacs1 _________________________________________6__25_ ( .DIN(
        _____________________________186________), .CLK(_26898), .CLRB(_____), 
        .Q(_26347), .QN(_53189) );
  dffacs1 _________________________________________8__15_ ( .DIN(
        _____________________________240________), .CLK(_26907), .CLRB(_____), 
        .Q(_26258), .QN(_53523) );
  dffacs1 _________________________________________2__0_ ( .DIN(
        _____________________________33________), .CLK(_26898), .CLRB(_____), 
        .Q(_26554), .QN(_53013) );
  dffacs1 __________________________________________1__8_ ( .DIN(
        ______________________________9________), .CLK(_26873), .CLRB(_____), 
        .Q(_26251), .QN(_53017) );
  dffacs1 __________________________________________1__3_ ( .DIN(
        ______________________________4________), .CLK(_26869), .CLRB(_____), 
        .QN(_52879) );
  dffacs1 _________________________________________0__24_ ( .DIN(
        _________________________________________25_________), .CLK(_26937), 
        .CLRB(_____), .Q(_26644), .QN(_53250) );
  dffacs1 _________________________________________5__15_ ( .DIN(
        _____________________________144________), .CLK(_26869), .CLRB(_____), 
        .Q(_26549), .QN(_53246) );
  dffacs1 _________________________________________7__26_ ( .DIN(
        _____________________________219________), .CLK(_26918), .CLRB(_____), 
        .Q(_26422), .QN(_53466) );
  dffacs1 _________________________________________7__14_ ( .DIN(
        _____________________________207________), .CLK(_26918), .CLRB(_____), 
        .QN(_53152) );
  dffacs1 _________________________________________3__15_ ( .DIN(
        _____________________________80________), .CLK(_26946), .CLRB(_____), 
        .QN(_53331) );
  dffacs1 _________________________________________1__25_ ( .DIN(
        _____________________________26________), .CLK(_26950), .CLRB(_____), 
        .QN(_53330) );
  dffacs1 _________________________________________5__19_ ( .DIN(
        _____________________________148________), .CLK(_26948), .CLRB(_____), 
        .Q(_26676), .QN(_53245) );
  dffacs1 _________________________________________2__22_ ( .DIN(
        _____________________________55________), .CLK(_26936), .CLRB(_____), 
        .QN(_53028) );
  dffacs1 __________________________________________1__18_ ( .DIN(
        ______________________________19________), .CLK(_26932), .CLRB(_____), 
        .Q(_26667), .QN(_52908) );
  dffacs1 __________________________________________5__18_ ( .DIN(
        ______________________________147________), .CLK(_26915), .CLRB(_____), 
        .QN(_52938) );
  dffacs1 _________________________________________7__21_ ( .DIN(
        _____________________________214________), .CLK(_26883), .CLRB(_____), 
        .Q(_26517), .QN(_53146) );
  dffacs1 __________________________________________3__7_ ( .DIN(
        ______________________________72________), .CLK(_26978), .CLRB(_____), 
        .QN(_52995) );
  dffacs1 __________________________________________1__11_ ( .DIN(
        ______________________________12________), .CLK(_26865), .CLRB(_____), 
        .Q(_26365), .QN(_53123) );
  dffacs1 _________________________________________8__8_ ( .DIN(
        _____________________________233________), .CLK(_26915), .CLRB(_____), 
        .Q(_26754), .QN(_53124) );
  dffacs1 __________________________________________6__15_ ( .DIN(
        ______________________________176________), .CLK(_26915), .CLRB(_____), 
        .QN(_53122) );
  dffacs1 __________________________________________0__28_ ( .DIN(
        __________________________________________25________2____________), 
        .CLK(_26962), .CLRB(_____), .Q(_26491), .QN(_52884) );
  dffacs1 _________________________________________0__4_ ( .DIN(
        _________________________________________5_________), .CLK(_26975), 
        .CLRB(_____), .QN(_53023) );
  dffacs1 ____2________________0_ ( .DIN(____2____________0_____), .CLK(_26983), .CLRB(_____), .Q(_26240), .QN(_53405) );
  dffacs1 _________________________________________1__31_ ( .DIN(
        _____________________________32________), .CLK(_26914), .CLRB(_____), 
        .Q(_26600), .QN(_53208) );
  dffacs1 _________________________________________8__9_ ( .DIN(
        _____________________________234________), .CLK(_26859), .CLRB(_____), 
        .Q(_26453), .QN(_53430) );
  dffacs1 ____0________________15_ ( .DIN(____0____________15_____), .CLK(
        _26902), .CLRB(_____), .Q(_26576), .QN(_53453) );
  dffacs1 _________________________________________6__14_ ( .DIN(
        _____________________________175________), .CLK(_26919), .CLRB(_____), 
        .Q(_26606), .QN(_53151) );
  dffacs1 _________________________________________2__26_ ( .DIN(
        _____________________________59________), .CLK(_26937), .CLRB(_____), 
        .QN(_53223) );
  dffacs1 _________________________________________6__0_ ( .DIN(
        _____________________________161________), .CLK(_26938), .CLRB(_____), 
        .QN(_53222) );
  dffacs1 _________________________________________8__28_ ( .DIN(
        _____________________________253________), .CLK(_26923), .CLRB(_____), 
        .Q(_26552), .QN(_53100) );
  dffacs1 __________________________________________1__0_ ( .DIN(
        ______________________________1________), .CLK(_26909), .CLRB(_____), 
        .Q(_26603), .QN(_52881) );
  dffacs1 __________________________________________2__27_ ( .DIN(
        ______________________________60________), .CLK(_26985), .CLRB(_____), 
        .QN(_52859) );
  dffacs1 ____1________________6_ ( .DIN(____1____________6_____), .CLK(_26859), .CLRB(_____), .Q(_26722), .QN(_53423) );
  dffacs1 __________________________________________2__20_ ( .DIN(
        ______________________________53________), .CLK(_26860), .CLRB(_____), 
        .QN(_53413) );
  dffacs1 ____0________________10_0 ( .DIN(____0____________10_____), .CLK(
        _26911), .CLRB(_____), .Q(_26345), .QN(_53450) );
  dffacs1 __________________________________________4__10_ ( .DIN(
        ______________________________107________), .CLK(_26911), .CLRB(_____), 
        .QN(_53434) );
  dffacs1 ____________________________________25_ ( .DIN(
        __________________________________25_________), .CLK(_26975), .CLRB(
        _____), .Q(_26429), .QN(_53045) );
  dffacs1 _________________________________________0__5_ ( .DIN(
        _________________________________________6_________), .CLK(_26975), 
        .CLRB(_____), .QN(_53012) );
  dffacs1 __________________________________________0__12_ ( .DIN(
        __________________________________________12_________), .CLK(_26873), 
        .CLRB(_____), .QN(_53046) );
  dffacs1 __________________________________________0__9_ ( .DIN(
        __________________________________________9_________), .CLK(_26908), 
        .CLRB(_____), .Q(_26640), .QN(_53258) );
  dffacs1 _________________________________________3__5_ ( .DIN(
        _____________________________70________), .CLK(_26984), .CLRB(_____), 
        .Q(_26737), .QN(_53259) );
  dffacs1 _________________________________________5__8_ ( .DIN(
        _____________________________137________), .CLK(_26908), .CLRB(_____), 
        .Q(_26610), .QN(_53260) );
  dffacs1 __________________________________________4__16_ ( .DIN(
        ______________________________113________), .CLK(_26882), .CLRB(_____), 
        .Q(_26645), .QN(_53332) );
  dffacs1 _________________________________________1__17_ ( .DIN(
        _____________________________18________), .CLK(_26862), .CLRB(_____), 
        .Q(_26371), .QN(_53227) );
  dffacs1 _________________________________________9__17_ ( .DIN(
        _____________________________274________), .CLK(_26912), .CLRB(_____), 
        .Q(_26556), .QN(_52901) );
  dffacs1 _________________________________________3__10_ ( .DIN(
        _____________________________75________), .CLK(_26946), .CLRB(_____), 
        .Q(_26605), .QN(_53328) );
  dffacs1 _________________________________________2__5_ ( .DIN(
        _____________________________38________), .CLK(_26912), .CLRB(_____), 
        .QN(_53072) );
  dffacs1 _________________________________________6__9_ ( .DIN(
        _____________________________170________), .CLK(_26880), .CLRB(_____), 
        .Q(_26407), .QN(_53207) );
  dffacs1 _________________________________________8__5_ ( .DIN(
        _____________________________230________), .CLK(_26865), .CLRB(_____), 
        .Q(_26579), .QN(_53431) );
  dffacs1 _________________________________________5__30_ ( .DIN(
        _____________________________159________), .CLK(_26899), .CLRB(_____), 
        .Q(_26518), .QN(_53215) );
  dffacs1 __________________________________________5__7_ ( .DIN(
        ______________________________136________), .CLK(_26953), .CLRB(_____), 
        .Q(_26591), .QN(_53386) );
  dffacs1 __________________________________________3__16_ ( .DIN(
        ______________________________81________), .CLK(_26926), .CLRB(_____), 
        .QN(_53388) );
  dffacs1 ____3________________4_ ( .DIN(____3____________4_____), .CLK(_26875), .CLRB(_____), .Q(_26288), .QN(_53443) );
  dffacs1 _________________________________________1__0_ ( .DIN(
        _____________________________1________), .CLK(_26856), .CLRB(_____), 
        .Q(_26719), .QN(_53049) );
  dffacs1 _________________________________________4__13_ ( .DIN(
        _____________________________110________), .CLK(_26961), .CLRB(_____), 
        .QN(_53325) );
  dffacs1 _________________________________________1__2_ ( .DIN(
        _____________________________3________), .CLK(_26961), .CLRB(_____), 
        .Q(_26602), .QN(_53315) );
  dffacs1 __________________________________________1__24_ ( .DIN(
        ______________________________25________), .CLK(_26945), .CLRB(_____), 
        .QN(_52887) );
  dffacs1 ____2________________2_ ( .DIN(____2____________2_____), .CLK(_26983), .CLRB(_____), .Q(_26696), .QN(_53402) );
  dffacs1 ____0________________4_ ( .DIN(____0___________0_4_____), .CLK(
        _26894), .CLRB(_____), .QN(_53499) );
  dffacs1 ___________________________________18_ ( .DIN(
        _________________________________18_________), .CLK(_26894), .CLRB(
        _____), .Q(_26507), .QN(_53461) );
  dffacs1 ____0________________13_0 ( .DIN(____0____________13_____), .CLK(
        _26887), .CLRB(_____), .QN(_53454) );
  dffacs1 __________________________________________6__13_ ( .DIN(
        ______________________________174________), .CLK(_26877), .CLRB(_____), 
        .Q(_26672), .QN(_52915) );
  dffacs1 __________________________________________4__7_ ( .DIN(
        ______________________________104________), .CLK(_26953), .CLRB(_____), 
        .QN(_52996) );
  dffacs1 ____________________________________14_ ( .DIN(
        __________________________________14_________), .CLK(_26977), .CLRB(
        _____), .Q(_26758), .QN(_53490) );
  dffacs1 _________________________________________4__8_ ( .DIN(
        _____________________________105________), .CLK(_26881), .CLRB(_____), 
        .Q(_26553), .QN(_53336) );
  dffacs1 __________________________________________4__23_ ( .DIN(
        ______________________________120________), .CLK(_26921), .CLRB(_____), 
        .QN(_52968) );
  dffacs1 _________________________________________8__22_ ( .DIN(
        _____________________________247________), .CLK(_26868), .CLRB(_____), 
        .Q(_26547), .QN(_53104) );
  dffacs1 __________________________________________3__30_ ( .DIN(
        ______________________________95________), .CLK(_26922), .CLRB(_____), 
        .Q(_26349), .QN(_52957) );
  dffacs1 _________________________________________3__31_ ( .DIN(
        _____________________________96________), .CLK(_26903), .CLRB(_____), 
        .Q(_26743), .QN(_53276) );
  dffacs1 ____0________________6_ ( .DIN(____0___________0_6_____), .CLK(
        _26963), .CLRB(_____), .Q(_26565), .QN(_53474) );
  dffacs1 ____0________________7_ ( .DIN(____0___________0_7_____), .CLK(
        _26973), .CLRB(_____), .Q(_26233), .QN(_53476) );
  dffacs1 _________________________________________9__8_ ( .DIN(
        _____________________________265________), .CLK(_26981), .CLRB(_____), 
        .Q(_26751), .QN(_53085) );
  dffacs1 ____3________________5_ ( .DIN(____3____________5_____), .CLK(_26901), .CLRB(_____), .QN(_53436) );
  dffacs1 __________________________________________6__30_ ( .DIN(
        ______________________________191________), .CLK(_26895), .CLRB(_____), 
        .QN(_53464) );
  dffacs1 ____________________________________26_ ( .DIN(
        __________________________________26_________), .CLK(_26895), .CLRB(
        _____), .QN(_53463) );
  dffacs1 __________________________________________2__26_ ( .DIN(
        ______________________________59________), .CLK(_26934), .CLRB(_____), 
        .QN(_52860) );
  dffacs1 __________________________________________3__0_ ( .DIN(
        ______________________________65________), .CLK(_26936), .CLRB(_____), 
        .Q(_26359), .QN(_53426) );
  dffacs1 _________________________________________7__25_ ( .DIN(
        _____________________________218________), .CLK(_26936), .CLRB(_____), 
        .Q(_26500), .QN(_53428) );
  dffacs1 ____1________________0_ ( .DIN(____1____________0_____), .CLK(_26864), .CLRB(_____), .Q(_26538), .QN(_53417) );
  dffacs1 _________________________________________2__7_ ( .DIN(
        _____________________________40________), .CLK(_26900), .CLRB(_____), 
        .Q(_26237), .QN(_53383) );
  dffacs1 _________________________________________0__6_ ( .DIN(
        _________________________________________7_________), .CLK(_26913), 
        .CLRB(_____), .QN(_53011) );
  dffacs1 _________________________________________0__11_ ( .DIN(
        _________________________________________12_________), .CLK(_26877), 
        .CLRB(_____), .Q(_26488), .QN(_53272) );
  dffacs1 _________________________________________0__18_ ( .DIN(
        _________________________________________19_________), .CLK(_26935), 
        .CLRB(_____), .Q(_26439), .QN(_53165) );
  dffacs1 _________________________________________0__13_ ( .DIN(
        _________________________________________14_________), .CLK(_26974), 
        .CLRB(_____), .QN(_53241) );
  dffacs1 ____0________________0_1 ( .DIN(____0___________0[0]), .CLK(_26906), 
        .CLRB(_____), .Q(_26409), .QN(_1877) );
  dffacs1 ____0________________1_1 ( .DIN(____0___________0[1]), .CLK(_26905), 
        .CLRB(_____), .QN(_1876) );
  dffacs1 ____0________________6_1 ( .DIN(____0___________0[6]), .CLK(_26905), 
        .CLRB(_____), .Q(_26652), .QN(_1853) );
  dffacs1 ____0________________7_1 ( .DIN(____0___________0[7]), .CLK(_26905), 
        .CLRB(_____), .QN(_1852) );
  dffacs1 ____0________________5_1 ( .DIN(____0___________0[5]), .CLK(_26904), 
        .CLRB(_____), .Q(_26697), .QN(_1860) );
  dffacs1 ____0________________2_1 ( .DIN(____0___________0[2]), .CLK(_26906), 
        .CLRB(_____), .Q(_26245), .QN(_53526) );
  dffacs1 ____0________________12_1 ( .DIN(____0___________0[12]), .CLK(_26904), .CLRB(_____), .QN(_1825) );
  dffacs1 ____0________________9_1 ( .DIN(____0___________0[9]), .CLK(_26906), 
        .CLRB(_____), .Q(_26421), .QN(_53524) );
  dffacs1 ____0________________3_1 ( .DIN(____0___________0[3]), .CLK(_26905), 
        .CLRB(_____), .QN(_1863) );
  dffacs1 ____0________________13_1 ( .DIN(____0___________0[13]), .CLK(_26904), .CLRB(_____), .QN(_1824) );
  dffacs1 ____0________________11_1 ( .DIN(____0___________0[11]), .CLK(_26904), .CLRB(_____), .Q(_26414), .QN(_1826) );
  dffacs1 ____0________________10_1 ( .DIN(____0___________0[10]), .CLK(_26904), .CLRB(_____), .Q(_26438), .QN(_1827) );
  dffacs1 ____0________________4_1 ( .DIN(____0___________0[4]), .CLK(_26905), 
        .CLRB(_____), .Q(_26541), .QN(_53525) );
  dffacs1 ____0________________8_2 ( .DIN(____0___________0[8]), .CLK(_26905), 
        .CLRB(_____), .Q(_26312), .QN(_1851) );
  dffacs1 ____3________________0_0 ( .DIN(____3___________[0]), .CLK(_26882), 
        .CLRB(_____), .Q(_26724), .QN(_2731) );
  dffacs1 ____3________________5_0 ( .DIN(____3___________[5]), .CLK(_26968), 
        .CLRB(_____), .QN(_53521) );
  dffacs1 ____3________________6_0 ( .DIN(____3___________[6]), .CLK(_26969), 
        .CLRB(_____), .QN(_2711) );
  dffacs1 ____3________________7_0 ( .DIN(____3___________[7]), .CLK(_26969), 
        .CLRB(_____), .Q(_26225), .QN(_2699) );
  dffacs1 ____3________________10_0 ( .DIN(____3___________[10]), .CLK(_26969), 
        .CLRB(_____), .Q(_26468), .QN(_2684) );
  dffacs1 ____3________________2_0 ( .DIN(____3___________[2]), .CLK(_26969), 
        .CLRB(_____), .Q(_26249), .QN(_2724) );
  dffacs1 ____3________________1_0 ( .DIN(____3___________[1]), .CLK(_26968), 
        .CLRB(_____), .Q(_26315), .QN(_2730) );
  dffacs1 ____1________________0_1 ( .DIN(____1___________[0]), .CLK(_26966), 
        .CLRB(_____), .Q(_26303), .QN(_2474) );
  dffacs1 ____1________________7_0 ( .DIN(____1___________[7]), .CLK(_26964), 
        .CLRB(_____), .Q(_26725), .QN(_2432) );
  dffacs1 ____1________________12_ ( .DIN(____1___________0[12]), .CLK(_26871), 
        .CLRB(_____), .QN(_2022) );
  dffacs1 ____1________________3_0 ( .DIN(____1___________0[3]), .CLK(_26907), 
        .CLRB(_____), .Q(_26254), .QN(_2061) );
  dffacs1 ____1________________7_1 ( .DIN(____1___________0[7]), .CLK(_26907), 
        .CLRB(_____), .Q(_26327), .QN(_2030) );
  dffacs1 ____1________________6_0 ( .DIN(____1___________0[6]), .CLK(_26914), 
        .CLRB(_____), .QN(_2031) );
  dffacs1 ____1________________5_0 ( .DIN(____1___________0[5]), .CLK(_26906), 
        .CLRB(_____), .Q(_26280), .QN(_2056) );
  dffacs1 ____1________________1_0 ( .DIN(____1___________0[1]), .CLK(_26871), 
        .CLRB(_____), .Q(_26444), .QN(_2063) );
  dffacs1 ____1________________8_0 ( .DIN(____1___________0[8]), .CLK(_26923), 
        .CLRB(_____), .Q(_26413), .QN(_2027) );
  dffacs1 ____1________________14_ ( .DIN(____1___________0[14]), .CLK(_26872), 
        .CLRB(_____), .Q(_26415), .QN(_2006) );
  dffacs1 ____1________________11_0 ( .DIN(____1___________0[11]), .CLK(_26871), .CLRB(_____), .Q(_26641), .QN(_2023) );
  dffacs1 ____1________________10_0 ( .DIN(____1___________0[10]), .CLK(_26871), .CLRB(_____), .QN(_2025) );
  dffacs1 ____1________________2_0 ( .DIN(____1___________0[2]), .CLK(_26907), 
        .CLRB(_____), .Q(_26647), .QN(_2062) );
  dffacs1 ____1________________13_ ( .DIN(____1___________0[13]), .CLK(_26871), 
        .CLRB(_____), .Q(_26277), .QN(_2015) );
  dffacs1 ____1________________4_0 ( .DIN(____1___________0[4]), .CLK(_26907), 
        .CLRB(_____), .QN(_2057) );
  dffacs1 ____1________________15_ ( .DIN(____1___________0[15]), .CLK(_26906), 
        .CLRB(_____), .Q(_26326), .QN(_1986) );
  dffacs1 ____1________________9_0 ( .DIN(____1___________0[9]), .CLK(_26906), 
        .CLRB(_____), .QN(_2026) );
  dffacs1 ____2________________0_0 ( .DIN(____2___________[0]), .CLK(_26972), 
        .CLRB(_____), .Q(_26310), .QN(_2643) );
  dffacs1 ____2________________7_0 ( .DIN(____2___________[7]), .CLK(_26971), 
        .CLRB(_____), .Q(_26665), .QN(_2599) );
  dffacs1 ____2________________13_0 ( .DIN(____2___________[13]), .CLK(_26972), 
        .CLRB(_____), .Q(_26358), .QN(_53516) );
  dffacs1 ____2________________3_0 ( .DIN(____2___________[3]), .CLK(_26970), 
        .CLRB(_____), .Q(_26273), .QN(_2628) );
  dffacs1 ____2________________8_0 ( .DIN(____2___________[8]), .CLK(_26971), 
        .CLRB(_____), .Q(_26398), .QN(_2598) );
  dffacs1 ____2________________5_0 ( .DIN(____2___________[5]), .CLK(_26972), 
        .CLRB(_____), .Q(_26417), .QN(_2625) );
  dffacs1 ____2________________2_0 ( .DIN(____2___________[2]), .CLK(_26971), 
        .CLRB(_____), .Q(_26573), .QN(_2637) );
  dffacs1 ____2________________9_0 ( .DIN(____2___________[9]), .CLK(_26972), 
        .CLRB(_____), .Q(_26246), .QN(_2590) );
  dffacs1 ____2________________6_0 ( .DIN(____2___________[6]), .CLK(_26971), 
        .CLRB(_____), .QN(_2624) );
  dffacs1 ____2________________12_0 ( .DIN(____2___________[12]), .CLK(_26970), 
        .CLRB(_____), .Q(_26247), .QN(_2571) );
  dffacs1 ____2________________4_0 ( .DIN(____2___________[4]), .CLK(_26971), 
        .CLRB(_____), .Q(_26340), .QN(_2627) );
  dffacs1 ____2________________11_0 ( .DIN(____2___________[11]), .CLK(_26970), 
        .CLRB(_____), .Q(_26567), .QN(_2575) );
  dffacs1 ____2________________10_0 ( .DIN(____2___________[10]), .CLK(_26970), 
        .CLRB(_____), .Q(_26229), .QN(_2576) );
  dffacs1 ____2________________1_0 ( .DIN(____2___________[1]), .CLK(_26971), 
        .CLRB(_____), .Q(_26216), .QN(_2642) );
  dffacs1 ____3________________9_0 ( .DIN(____3___________[9]), .CLK(_26970), 
        .CLRB(_____), .Q(_26363), .QN(_2697) );
  dffacs1 ____3________________3_0 ( .DIN(____3___________[3]), .CLK(_26969), 
        .CLRB(_____), .Q(_26575), .QN(_2722) );
  dffacs1 ____3________________8_0 ( .DIN(____3___________[8]), .CLK(_26970), 
        .CLRB(_____), .Q(_26328), .QN(_2698) );
  dffacs1 ____3________________4_0 ( .DIN(____3___________[4]), .CLK(_26969), 
        .CLRB(_____), .Q(_26692), .QN(_2718) );
  dffacs1 ____0________________7_2 ( .DIN(____0___________[7]), .CLK(_26967), 
        .CLRB(_____), .Q(_26370), .QN(_2217) );
  dffacs1 ____0________________6_2 ( .DIN(____0___________[6]), .CLK(_26968), 
        .CLRB(_____), .Q(_26294), .QN(_2238) );
  dffacs1 ____0________________5_2 ( .DIN(____0___________[5]), .CLK(_26967), 
        .CLRB(_____), .Q(_26311), .QN(_2251) );
  dffacs1 ____0________________0_2 ( .DIN(____0___________[0]), .CLK(_26887), 
        .CLRB(_____), .Q(_26646), .QN(_2274) );
  dffacs1 ____0________________2_2 ( .DIN(____0___________[2]), .CLK(_26966), 
        .CLRB(_____), .Q(_26217), .QN(_53522) );
  dffacs1 ____0________________9_2 ( .DIN(____0___________[9]), .CLK(_26966), 
        .CLRB(_____), .Q(_26433), .QN(_2214) );
  dffacs1 ____0________________12_2 ( .DIN(____0___________[12]), .CLK(_26967), 
        .CLRB(_____), .QN(_2181) );
  dffacs1 ____0________________1_2 ( .DIN(____0___________[1]), .CLK(_26968), 
        .CLRB(_____), .QN(_2273) );
  dffacs1 ____0________________11_2 ( .DIN(____0___________[11]), .CLK(_26966), 
        .CLRB(_____), .Q(_26509), .QN(_2182) );
  dffacs1 ____0________________10_2 ( .DIN(____0___________[10]), .CLK(_26966), 
        .CLRB(_____), .Q(_26248), .QN(_2203) );
  dffacs1 ____0________________13_2 ( .DIN(____0___________[13]), .CLK(_26967), 
        .CLRB(_____), .QN(_2180) );
  dffacs1 ____0________________14_0 ( .DIN(____0___________[14]), .CLK(_26967), 
        .CLRB(_____), .Q(_26223), .QN(_2179) );
  dffacs1 ____0________________15_0 ( .DIN(____0___________[15]), .CLK(_26966), 
        .CLRB(_____), .Q(_26419), .QN(_2175) );
  dffacs1 ____0________________4_2 ( .DIN(____0___________[4]), .CLK(_26968), 
        .CLRB(_____), .Q(_26706), .QN(_2252) );
  dffacs1 ____0________________3_2 ( .DIN(____0___________[3]), .CLK(_26967), 
        .CLRB(_____), .Q(_26709), .QN(_2253) );
  dffacs1 ____1________________4_1 ( .DIN(____1___________[4]), .CLK(_26964), 
        .CLRB(_____), .Q(_26316), .QN(_2440) );
  dffacs1 ____1________________10_1 ( .DIN(____1___________[10]), .CLK(_26964), 
        .CLRB(_____), .Q(_26633), .QN(_2395) );
  dffacs1 ____1________________1_1 ( .DIN(____1___________[1]), .CLK(_26965), 
        .CLRB(_____), .Q(_26580), .QN(_2473) );
  dffacs1 ____1________________5_1 ( .DIN(____1___________[5]), .CLK(_26963), 
        .CLRB(_____), .QN(_2439) );
  dffacs1 ____1________________3_1 ( .DIN(____1___________[3]), .CLK(_26964), 
        .CLRB(_____), .QN(_53518) );
  dffacs1 ____1________________11_1 ( .DIN(____1___________[11]), .CLK(_26964), 
        .CLRB(_____), .Q(_26430), .QN(_2320) );
  dffacs1 ____1________________9_1 ( .DIN(____1___________[9]), .CLK(_26965), 
        .CLRB(_____), .Q(_26278), .QN(_53520) );
  dffacs1 ____1________________6_1 ( .DIN(____1___________[6]), .CLK(_26965), 
        .CLRB(_____), .Q(_26714), .QN(_53519) );
  dffacs1 ____1________________2_1 ( .DIN(____1___________[2]), .CLK(_26964), 
        .CLRB(_____), .Q(_26642), .QN(_2472) );
  dffacs1 ____1________________8_1 ( .DIN(____1___________[8]), .CLK(_26965), 
        .CLRB(_____), .Q(_26324), .QN(_2429) );
  dffacs1 _________________________________________7__4_ ( .DIN(
        _____________________________197________), .CLK(_26880), .CLRB(_____), 
        .QN(_26483) );
  dffacs1 _________________________________________5__24_ ( .DIN(
        _____________________________153________), .CLK(_26973), .CLRB(_____), 
        .QN(_26656) );
  dffacs1 __________________________________________5__23_ ( .DIN(
        ______________________________152________), .CLK(_26979), .CLRB(_____), 
        .QN(_26511) );
  dffacs1 _________________________________________5__2_ ( .DIN(
        _____________________________131________), .CLK(_26890), .CLRB(_____), 
        .QN(_26375) );
  dffacs1 __________________________________________6__22_ ( .DIN(
        ______________________________183________), .CLK(_26874), .CLRB(_____), 
        .QN(_26481) );
  dffacs1 _________________________________________5__0_ ( .DIN(
        _____________________________129________), .CLK(_26893), .CLRB(_____), 
        .QN(_26569) );
  dffacs1 _________________________________________2__12_ ( .DIN(
        _____________________________45________), .CLK(_26960), .CLRB(_____), 
        .QN(_26374) );
  dffacs1 _________________________________________4__10_ ( .DIN(
        _____________________________107________), .CLK(_26890), .CLRB(_____), 
        .QN(_26284) );
  dffacs1 _________________________________________5__14_ ( .DIN(
        _____________________________143________), .CLK(_26879), .CLRB(_____), 
        .QN(_26342) );
  dffacs1 _________________________________________6__2_ ( .DIN(
        _____________________________163________), .CLK(_26974), .CLRB(_____), 
        .QN(_26268) );
  dffacs1 ____3________________6_ ( .DIN(____3____________6_____), .CLK(_26900), .CLRB(_____), .QN(_26211) );
  dffacs1 _________________________________________3__27_ ( .DIN(
        _____________________________92________), .CLK(_26870), .CLRB(_____), 
        .Q(_53284), .QN(_26224) );
  dffacs1 __________________________________________3__23_ ( .DIN(
        ______________________________88________), .CLK(_26921), .CLRB(_____), 
        .Q(_53339), .QN(_26401) );
  dffacs1 _________________________________________9__19_ ( .DIN(
        _____________________________276________), .CLK(_26981), .CLRB(_____), 
        .Q(_53070), .QN(_26432) );
  dffacs1 _________________________________________8__11_ ( .DIN(
        _____________________________236________), .CLK(_26923), .CLRB(_____), 
        .Q(_53130), .QN(_26373) );
  dffacs1 _________________________________________1__16_ ( .DIN(
        _____________________________17________), .CLK(_26949), .CLRB(_____), 
        .Q(_53195), .QN(_26379) );
  dffacs1 _________________________________________1__18_ ( .DIN(
        _____________________________19________), .CLK(_26899), .CLRB(_____), 
        .Q(_53194), .QN(_26404) );
  dffacs1 _________________________________________1__21_ ( .DIN(
        _____________________________22________), .CLK(_26983), .CLRB(_____), 
        .Q(_53166), .QN(_26348) );
  dffacs1 _________________________________________2__6_ ( .DIN(
        _____________________________39________), .CLK(_26985), .CLRB(_____), 
        .Q(_53161), .QN(_26384) );
  dffacs1 _________________________________________3__2_ ( .DIN(
        _____________________________67________), .CLK(_26914), .CLRB(_____), 
        .Q(_53345), .QN(_26220) );
  dffacs1 _________________________________________2__14_ ( .DIN(
        _____________________________47________), .CLK(_26907), .CLRB(_____), 
        .Q(_53033), .QN(_26307) );
  dffacs1 _________________________________________7__22_ ( .DIN(
        _____________________________215________), .CLK(_26884), .CLRB(_____), 
        .Q(_53145), .QN(_26236) );
  dffacs1 _________________________________________5__7_ ( .DIN(
        _____________________________136________), .CLK(_26908), .CLRB(_____), 
        .Q(_53265), .QN(_26255) );
  dffacs1 _________________________________________0__12_ ( .DIN(
        _________________________________________13_________), .CLK(_26982), 
        .CLRB(_____), .Q(_53254) );
  dffacs1 _________________________________________5__17_ ( .DIN(
        _____________________________146________), .CLK(_26941), .CLRB(_____), 
        .Q(_53249), .QN(_26649) );
  dffacs1 __________________________________________0__27_ ( .DIN(
        __________________________________________25________1____________), 
        .CLK(_26892), .CLRB(_____), .Q(_53274), .QN(_26377) );
  dffacs1 _________________________________________1__11_ ( .DIN(
        _____________________________12________), .CLK(_26949), .CLRB(_____), 
        .Q(_53253), .QN(_26290) );
  dffacs1 _________________________________________7__9_ ( .DIN(
        _____________________________202________), .CLK(_26859), .CLRB(_____), 
        .Q(_53164), .QN(_26390) );
  dffacs1 _________________________________________8__3_ ( .DIN(
        _____________________________228________), .CLK(_26865), .CLRB(_____), 
        .Q(_53088), .QN(_26424) );
  dffacs1 _________________________________________6__12_ ( .DIN(
        _____________________________173________), .CLK(_26859), .CLRB(_____), 
        .Q(_53213), .QN(_26372) );
  dffacs1 _________________________________________0__3_ ( .DIN(
        _________________________________________4_________), .CLK(_26885), 
        .CLRB(_____), .Q(_53317), .QN(_26479) );
  dffacs1 __________________________________________3__9_ ( .DIN(
        ______________________________74________), .CLK(_26869), .CLRB(_____), 
        .Q(_52992), .QN(_26478) );
  dffacs1 _________________________________________2__21_ ( .DIN(
        _____________________________54________), .CLK(_26947), .CLRB(_____), 
        .Q(_53203), .QN(_26505) );
  dffacs1 __________________________________________1__15_ ( .DIN(
        ______________________________16________), .CLK(_26860), .CLRB(_____), 
        .Q(_52928), .QN(_26475) );
  dffacs1 _________________________________________7__7_ ( .DIN(
        _____________________________200________), .CLK(_26863), .CLRB(_____), 
        .Q(_53169), .QN(_26252) );
  dffacs1 __________________________________________3__14_ ( .DIN(
        ______________________________79________), .CLK(_26978), .CLRB(_____), 
        .Q(_52983) );
  dffacs1 _________________________________________0__14_ ( .DIN(
        _________________________________________15_________), .CLK(_26980), 
        .CLRB(_____), .Q(_53229) );
  dffacs1 ____2________________13_ ( .DIN(____2____________13_____), .CLK(
        _26875), .CLRB(_____), .Q(_53403), .QN(_26515) );
  dffacs1 _________________________________________7__0_ ( .DIN(
        _____________________________193________), .CLK(_26917), .CLRB(_____), 
        .Q(_52835) );
  dffacs1 __________________________________________6__21_ ( .DIN(
        ______________________________182________), .CLK(_26957), .CLRB(_____), 
        .Q(_52907), .QN(_26459) );
  dffacs1 _________________________________________5__26_ ( .DIN(
        _____________________________155________), .CLK(_26910), .CLRB(_____), 
        .Q(_53255), .QN(_26476) );
  dffacs1 _________________________________________3__0_ ( .DIN(
        _____________________________65________), .CLK(_26898), .CLRB(_____), 
        .Q(_53014), .QN(_26441) );
  dffacs1 __________________________________________0__20_ ( .DIN(
        __________________________________________20_________), .CLK(_26950), 
        .CLRB(_____), .Q(_52899), .QN(_26502) );
  dffacs1 _________________________________________5__27_ ( .DIN(
        _____________________________156________), .CLK(_26888), .CLRB(_____), 
        .Q(_53323), .QN(_26260) );
  dffacs1 _________________________________________8__13_ ( .DIN(
        _____________________________238________), .CLK(_26923), .CLRB(_____), 
        .Q(_53118), .QN(_26452) );
  dffacs1 __________________________________________4__22_ ( .DIN(
        ______________________________119________), .CLK(_26921), .CLRB(_____), 
        .Q(_52962) );
  dffacs1 __________________________________________4__5_ ( .DIN(
        ______________________________102________), .CLK(_26897), .CLRB(_____), 
        .Q(_52946) );
  dffacs1 _________________________________________0__16_ ( .DIN(
        _________________________________________17_________), .CLK(_26973), 
        .CLRB(_____), .Q(_53193) );
  dffacs1 __________________________________________1__22_ ( .DIN(
        ______________________________23________), .CLK(_26933), .CLRB(_____), 
        .Q(_52894), .QN(_26234) );
  dffacs1 __________________________________________0__19_ ( .DIN(
        __________________________________________19_________), .CLK(_26932), 
        .CLRB(_____), .Q(_52895), .QN(_26544) );
  dffacs1 _________________________________________5__13_ ( .DIN(
        _____________________________142________), .CLK(_26919), .CLRB(_____), 
        .Q(_53204), .QN(_26597) );
  dffacs1 _________________________________________4__19_ ( .DIN(
        _____________________________116________), .CLK(_26920), .CLRB(_____), 
        .Q(_53303), .QN(_26601) );
  dffacs1 __________________________________________0__4_ ( .DIN(
        __________________________________________4_________), .CLK(_26951), 
        .CLRB(_____), .Q(_52858), .QN(_26572) );
  dffacs1 _________________________________________7__6_ ( .DIN(
        _____________________________199________), .CLK(_26892), .CLRB(_____), 
        .Q(_53167), .QN(_26501) );
  dffacs1 __________________________________________4__28_ ( .DIN(
        ______________________________125________), .CLK(_26867), .CLRB(_____), 
        .Q(_53395), .QN(_26440) );
  dffacs1 _________________________________________1__20_ ( .DIN(
        _____________________________21________), .CLK(_26983), .CLRB(_____), 
        .Q(_53399), .QN(_26362) );
  dffacs1 _________________________________________3__18_ ( .DIN(
        _____________________________83________), .CLK(_26950), .CLRB(_____), 
        .Q(_53305), .QN(_26378) );
  dffacs1 _________________________________________5__25_ ( .DIN(
        _____________________________154________), .CLK(_26942), .CLRB(_____), 
        .Q(_53187) );
  dffacs1 _________________________________________9__6_ ( .DIN(
        _____________________________263________), .CLK(_26931), .CLRB(_____), 
        .Q(_53086) );
  dffacs1 _________________________________________2__8_ ( .DIN(
        _____________________________41________), .CLK(_26882), .CLRB(_____), 
        .Q(_53044), .QN(_26350) );
  dffacs1 __________________________________________6__17_ ( .DIN(
        ______________________________178________), .CLK(_26915), .CLRB(_____), 
        .Q(_52914), .QN(_26571) );
  dffacs1 _________________________________________2__25_ ( .DIN(
        _____________________________58________), .CLK(_26879), .CLRB(_____), 
        .Q(_53322), .QN(_26376) );
  dffacs1 __________________________________________4__8_ ( .DIN(
        ______________________________105________), .CLK(_26877), .CLRB(_____), 
        .Q(_52997), .QN(_26391) );
  dffacs1 _________________________________________3__23_ ( .DIN(
        _____________________________88________), .CLK(_26936), .CLRB(_____), 
        .Q(_53294), .QN(_26412) );
  dffacs1 _________________________________________3__28_ ( .DIN(
        _____________________________93________), .CLK(_26939), .CLRB(_____), 
        .Q(_53283), .QN(_26420) );
  dffacs1 _________________________________________1__7_ ( .DIN(
        _____________________________8________), .CLK(_26913), .CLRB(_____), 
        .Q(_53038), .QN(_26695) );
  dffacs1 _________________________________________7__23_ ( .DIN(
        _____________________________216________), .CLK(_26883), .CLRB(_____), 
        .Q(_53398), .QN(_26543) );
  dffacs1 _________________________________________1__29_ ( .DIN(
        _____________________________30________), .CLK(_26875), .CLRB(_____), 
        .Q(_53139), .QN(_26639) );
  dffacs1 _________________________________________3__1_ ( .DIN(
        _____________________________66________), .CLK(_26881), .CLRB(_____), 
        .Q(_53015), .QN(_26513) );
  dffacs1 __________________________________________3__1_ ( .DIN(
        ______________________________66________), .CLK(_26975), .CLRB(_____), 
        .Q(_52853), .QN(_26732) );
  dffacs1 __________________________________________4__18_ ( .DIN(
        ______________________________115________), .CLK(_26916), .CLRB(_____), 
        .Q(_53211), .QN(_26718) );
  dffacs1 _________________________________________2__19_ ( .DIN(
        _____________________________52________), .CLK(_26947), .CLRB(_____), 
        .Q(_53031), .QN(_26352) );
  dffacs1 __________________________________________5__28_ ( .DIN(
        ______________________________157________), .CLK(_26867), .CLRB(_____), 
        .Q(_52927), .QN(_26583) );
  dffacs1 _________________________________________2__30_ ( .DIN(
        _____________________________63________), .CLK(_26902), .CLRB(_____), 
        .Q(_53069), .QN(_26339) );
  dffacs1 __________________________________________0__16_ ( .DIN(
        __________________________________________16_________), .CLK(_26873), 
        .CLRB(_____), .Q(_52909), .QN(_26599) );
  dffacs1 ____________________________________29_ ( .DIN(
        __________________________________29_________), .CLK(_26882), .CLRB(
        _____), .Q(_52970), .QN(_26425) );
  dffacs1 _________________________________________2__27_ ( .DIN(
        _____________________________60________), .CLK(_26871), .CLRB(_____), 
        .Q(_53024), .QN(_26346) );
  dffacs1 __________________________________________1__29_ ( .DIN(
        ______________________________30________), .CLK(_26892), .CLRB(_____), 
        .Q(_52886), .QN(_26402) );
  dffacs1 ____________________________________0_ ( .DIN(
        __________________________________0_________), .CLK(_26928), .CLRB(
        _____), .Q(_53512), .QN(_26562) );
  dffacs1 __________________________________________6__31_ ( .DIN(
        ______________________________192________), .CLK(_26896), .CLRB(_____), 
        .Q(_52900) );
  dffacs1 __________________________________________6__9_ ( .DIN(
        ______________________________170________), .CLK(_26881), .CLRB(_____), 
        .Q(_52917) );
  dffacs1 _________________________________________4__22_ ( .DIN(
        _____________________________119________), .CLK(_26884), .CLRB(_____), 
        .Q(_53282) );
  dffacs1 __________________________________________3__11_ ( .DIN(
        ______________________________76________), .CLK(_26948), .CLRB(_____), 
        .Q(_52989) );
  dffacs1 __________________________________________5__15_ ( .DIN(
        ______________________________144________), .CLK(_26942), .CLRB(_____), 
        .Q(_52913) );
  dffacs1 _________________________________________0__17_ ( .DIN(
        _________________________________________18_________), .CLK(_26935), 
        .CLRB(_____), .Q(_53178), .QN(_26499) );
  dffacs1 __________________________________________6__4_ ( .DIN(
        ______________________________165________), .CLK(_26953), .CLRB(_____), 
        .Q(_52923), .QN(_26581) );
  dffacs1 __________________________________________2__30_ ( .DIN(
        ______________________________63________), .CLK(_26922), .CLRB(_____), 
        .Q(_53058), .QN(_26630) );
  dffacs1 ____________________________________3_ ( .DIN(
        __________________________________3_________), .CLK(_26928), .CLRB(
        _____), .Q(_53509), .QN(_26542) );
  dffacs1 _________________________________________4__25_ ( .DIN(
        _____________________________122________), .CLK(_26942), .CLRB(_____), 
        .Q(_53298), .QN(_26510) );
  dffacs1 __________________________________________0__15_ ( .DIN(
        __________________________________________15_________), .CLK(_26943), 
        .CLRB(_____), .Q(_52919), .QN(_26693) );
  dffacs1 _________________________________________3__26_ ( .DIN(
        _____________________________91________), .CLK(_26870), .CLRB(_____), 
        .Q(_53290), .QN(_26281) );
  dffacs1 __________________________________________5__31_ ( .DIN(
        ______________________________160________), .CLK(_26962), .CLRB(_____), 
        .Q(_52941), .QN(_26498) );
  dffacs1 _________________________________________3__8_ ( .DIN(
        _____________________________73________), .CLK(_26864), .CLRB(_____), 
        .Q(_53334), .QN(_26582) );
  dffacs1 __________________________________________2__28_ ( .DIN(
        ______________________________61________), .CLK(_26986), .CLRB(_____), 
        .Q(_52857) );
  dffacs1 _________________________________________6__4_ ( .DIN(
        _____________________________165________), .CLK(_26863), .CLRB(_____), 
        .Q(_53216), .QN(_26533) );
  dffacs1 __________________________________________1__19_ ( .DIN(
        ______________________________20________), .CLK(_26932), .CLRB(_____), 
        .Q(_52897), .QN(_26637) );
  dffacs1 _________________________________________3__7_ ( .DIN(
        _____________________________72________), .CLK(_26890), .CLRB(_____), 
        .Q(_53335), .QN(_26474) );
  dffacs1 _________________________________________4__17_ ( .DIN(
        _____________________________114________), .CLK(_26945), .CLRB(_____), 
        .Q(_53247), .QN(_26750) );
  dffacs1 _________________________________________0__19_ ( .DIN(
        _________________________________________20_________), .CLK(_26984), 
        .CLRB(_____), .Q(_53233), .QN(_26638) );
  dffacs1 ____________________________________23_ ( .DIN(
        __________________________________23_________), .CLK(_26866), .CLRB(
        _____), .Q(_53505), .QN(_26560) );
  dffacs1 __________________________________________0__10_ ( .DIN(
        __________________________________________10_________), .CLK(_26917), 
        .CLRB(_____), .Q(_53199) );
  dffacs1 __________________________________________2__13_ ( .DIN(
        ______________________________46________), .CLK(_26857), .CLRB(_____), 
        .Q(_52931) );
  dffacs1 _________________________________________0__28_ ( .DIN(
        _________________________________________0________2____________), 
        .CLK(_26955), .CLRB(_____), .Q(_53141), .QN(_26636) );
  dffacs1 __________________________________________1__4_ ( .DIN(
        ______________________________5________), .CLK(_26961), .CLRB(_____), 
        .Q(_52877), .QN(_26635) );
  dffacs1 ___________________________________12_ ( .DIN(
        _________________________________12_________), .CLK(_26939), .CLRB(
        _____), .Q(_53492), .QN(_26749) );
  dffacs1 _________________________________________3__19_ ( .DIN(
        _____________________________84________), .CLK(_26920), .CLRB(_____), 
        .Q(_53302) );
  dffacs1 _________________________________________1__26_ ( .DIN(
        _____________________________27________), .CLK(_26900), .CLRB(_____), 
        .Q(_53066), .QN(_26563) );
  dffacs1 _________________________________________0__8_ ( .DIN(
        _________________________________________9_________), .CLK(_26914), 
        .CLRB(_____), .Q(_53008) );
  dffacs1 _________________________________________4__12_ ( .DIN(
        _____________________________109________), .CLK(_26920), .CLRB(_____), 
        .Q(_53324), .QN(_26456) );
  dffacs1 ___________________________________5_ ( .DIN(
        _________________________________5_________), .CLK(_26931), .CLRB(
        _____), .Q(_53514), .QN(_26559) );
  dffacs1 ____3________________3_ ( .DIN(____3____________3_____), .CLK(_26876), .CLRB(_____), .Q(_53435), .QN(_26686) );
  dffacs1 _________________________________________9__7_ ( .DIN(
        _____________________________264________), .CLK(_26896), .CLRB(_____), 
        .Q(_53079) );
  dffacs1 __________________________________________2__29_ ( .DIN(
        ______________________________62________), .CLK(_26952), .CLRB(_____), 
        .Q(_52956) );
  dffacs1 __________________________________________0__6_ ( .DIN(
        __________________________________________6_________), .CLK(_26986), 
        .CLRB(_____), .Q(_52856) );
  dffacs1 _________________________________________1__3_ ( .DIN(
        _____________________________4________), .CLK(_26885), .CLRB(_____), 
        .Q(_53043) );
  dffacs1 _________________________________________9__11_ ( .DIN(
        _____________________________268________), .CLK(_26858), .CLRB(_____), 
        .Q(_53075) );
  dffacs1 __________________________________________0__29_ ( .DIN(
        __________________________________________25________3____________), 
        .CLK(_26891), .CLRB(_____), .Q(_53393), .QN(_26564) );
  dffacs1 _________________________________________9__9_ ( .DIN(
        _____________________________266________), .CLK(_26896), .CLRB(_____), 
        .Q(_53084), .QN(_26313) );
  dffacs1 __________________________________________1__10_ ( .DIN(
        ______________________________11________), .CLK(_26944), .CLRB(_____), 
        .Q(_52986), .QN(_26506) );
  dffacs1 _________________________________________5__9_ ( .DIN(
        _____________________________138________), .CLK(_26889), .CLRB(_____), 
        .Q(_53264), .QN(_26566) );
  dffacs1 __________________________________________2__31_ ( .DIN(
        ______________________________64________), .CLK(_26865), .CLRB(_____), 
        .Q(_53126) );
  dffacs1 _________________________________________7__10_ ( .DIN(
        _____________________________203________), .CLK(_26984), .CLRB(_____), 
        .Q(_53397), .QN(_26469) );
  dffacs1 _________________________________________6__30_ ( .DIN(
        _____________________________191________), .CLK(_26899), .CLRB(_____), 
        .Q(_53177), .QN(_26632) );
  dffacs1 __________________________________________3__26_ ( .DIN(
        ______________________________91________), .CLK(_26934), .CLRB(_____), 
        .Q(_52855), .QN(_26496) );
  dffacs1 _________________________________________4__11_ ( .DIN(
        _____________________________108________), .CLK(_26888), .CLRB(_____), 
        .Q(_53326), .QN(_26400) );
  dffacs1 _________________________________________9__26_ ( .DIN(
        _____________________________283________), .CLK(_26974), .CLRB(_____), 
        .Q(_53515), .QN(_26540) );
  dffacs1 _________________________________________3__16_ ( .DIN(
        _____________________________81________), .CLK(_26959), .CLRB(_____), 
        .Q(_53308), .QN(_26689) );
  dffacs1 _________________________________________4__29_ ( .DIN(
        _____________________________126________), .CLK(_26884), .CLRB(_____), 
        .Q(_53286), .QN(_26436) );
  dffacs1 __________________________________________6__3_ ( .DIN(
        ______________________________164________), .CLK(_26929), .CLRB(_____), 
        .Q(_52924), .QN(_26688) );
  dffacs1 _________________________________________9__25_ ( .DIN(
        _____________________________282________), .CLK(_26934), .CLRB(_____), 
        .Q(_53063) );
  dffacs1 _________________________________________4__15_ ( .DIN(
        _____________________________112________), .CLK(_26946), .CLRB(_____), 
        .Q(_53310) );
  dffacs1 __________________________________________2__17_ ( .DIN(
        ______________________________50________), .CLK(_26860), .CLRB(_____), 
        .Q(_52864) );
  dffacs1 __________________________________________4__26_ ( .DIN(
        ______________________________123________), .CLK(_26941), .CLRB(_____), 
        .Q(_52961) );
  dffacs1 __________________________________________5__19_ ( .DIN(
        ______________________________148________), .CLK(_26921), .CLRB(_____), 
        .Q(_52936) );
  dffacs1 _________________________________________0__21_ ( .DIN(
        _________________________________________22_________), .CLK(_26954), 
        .CLRB(_____), .Q(_53127), .QN(_26535) );
  dffacs1 _________________________________________0__15_ ( .DIN(
        _________________________________________16_________), .CLK(_26935), 
        .CLRB(_____), .Q(_53470), .QN(_26534) );
  dffacs1 _________________________________________5__3_ ( .DIN(
        _____________________________132________), .CLK(_26947), .CLRB(_____), 
        .Q(_53269), .QN(_26385) );
  dffacs1 __________________________________________1__13_ ( .DIN(
        ______________________________14________), .CLK(_26943), .CLRB(_____), 
        .Q(_53192), .QN(_26628) );
  dffacs1 __________________________________________1__12_ ( .DIN(
        ______________________________13________), .CLK(_26873), .CLRB(_____), 
        .Q(_53016), .QN(_26473) );
  dffacs1 __________________________________________5__3_ ( .DIN(
        ______________________________132________), .CLK(_26910), .CLRB(_____), 
        .Q(_52949), .QN(_26532) );
  dffacs1 __________________________________________0__3_ ( .DIN(
        __________________________________________3_________), .CLK(_26986), 
        .CLRB(_____), .Q(_52866), .QN(_26715) );
  dffacs1 __________________________________________2__19_ ( .DIN(
        ______________________________52________), .CLK(_26926), .CLRB(_____), 
        .Q(_53396), .QN(_26305) );
  dffacs1 _________________________________________9__13_ ( .DIN(
        _____________________________270________), .CLK(_26858), .CLRB(_____), 
        .Q(_53076), .QN(_26631) );
  dffacs1 ____2________________5_ ( .DIN(____2____________5_____), .CLK(_26891), .CLRB(_____), .Q(_53412) );
  dffacs1 __________________________________________4__19_ ( .DIN(
        ______________________________116________), .CLK(_26921), .CLRB(_____), 
        .Q(_52976), .QN(_26687) );
  dffacs1 _________________________________________8__1_ ( .DIN(
        _____________________________226________), .CLK(_26961), .CLRB(_____), 
        .Q(_53133), .QN(_26450) );
  dffacs1 __________________________________________0__11_ ( .DIN(
        __________________________________________11_________), .CLK(_26866), 
        .CLRB(_____), .Q(_52839) );
  dffacs1 __________________________________________5__24_ ( .DIN(
        ______________________________153________), .CLK(_26975), .CLRB(_____), 
        .Q(_52904), .QN(_26368) );
  dffacs1 _________________________________________4__5_ ( .DIN(
        _____________________________102________), .CLK(_26972), .CLRB(_____), 
        .Q(_53348), .QN(_26344) );
  dffacs1 __________________________________________6__5_ ( .DIN(
        ______________________________166________), .CLK(_26923), .CLRB(_____), 
        .Q(_52926), .QN(_26527) );
  dffacs1 __________________________________________4__27_ ( .DIN(
        ______________________________124________), .CLK(_26941), .CLRB(_____), 
        .Q(_52959), .QN(_26536) );
  dffacs1 ____________________________________12_ ( .DIN(
        __________________________________12_________), .CLK(_26877), .CLRB(
        _____), .Q(_53493), .QN(_26611) );
  dffacs1 __________________________________________3__31_ ( .DIN(
        ______________________________96________), .CLK(_26922), .CLRB(_____), 
        .Q(_52954), .QN(_26471) );
  dffacs1 __________________________________________0__26_ ( .DIN(
        __________________________________________25________0____________), 
        .CLK(_26892), .CLRB(_____), .Q(_53390), .QN(_26508) );
  dffacs1 __________________________________________0__18_ ( .DIN(
        __________________________________________18_________), .CLK(_26932), 
        .CLRB(_____), .Q(_52849), .QN(_26306) );
  dffacs1 __________________________________________5__26_ ( .DIN(
        ______________________________155________), .CLK(_26893), .CLRB(_____), 
        .Q(_52933), .QN(_26250) );
  dffacs1 _________________________________________4__28_ ( .DIN(
        _____________________________125________), .CLK(_26884), .CLRB(_____), 
        .Q(_53297), .QN(_26266) );
  dffacs1 _________________________________________8__14_ ( .DIN(
        _____________________________239________), .CLK(_26924), .CLRB(_____), 
        .Q(_53117), .QN(_26694) );
  dffacs1 _________________________________________3__14_ ( .DIN(
        _____________________________79________), .CLK(_26946), .CLRB(_____), 
        .Q(_53312), .QN(_26531) );
  dffacs1 ____________________________________31_ ( .DIN(
        __________________________________31_________), .CLK(_26891), .CLRB(
        _____), .Q(_52883), .QN(_26730) );
  dffacs1 __________________________________________3__28_ ( .DIN(
        ______________________________93________), .CLK(_26952), .CLRB(_____), 
        .Q(_53107), .QN(_26731) );
  dffacs1 _________________________________________2__23_ ( .DIN(
        _____________________________56________), .CLK(_26939), .CLRB(_____), 
        .Q(_53243), .QN(_26366) );
  dffacs1 _________________________________________7__12_ ( .DIN(
        _____________________________205________), .CLK(_26859), .CLRB(_____), 
        .Q(_53160), .QN(_26627) );
  dffacs1 _________________________________________0__20_ ( .DIN(
        _________________________________________21_________), .CLK(_26955), 
        .CLRB(_____), .Q(_53142), .QN(_26397) );
  dffacs1 __________________________________________4__3_ ( .DIN(
        ______________________________100________), .CLK(_26910), .CLRB(_____), 
        .Q(_53003), .QN(_26691) );
  dffacs1 _________________________________________9__23_ ( .DIN(
        _____________________________280________), .CLK(_26904), .CLRB(_____), 
        .Q(_53065) );
  dffacs1 __________________________________________2__22_ ( .DIN(
        ______________________________55________), .CLK(_26933), .CLRB(_____), 
        .Q(_52863) );
  dffacs1 __________________________________________3__3_ ( .DIN(
        ______________________________68________), .CLK(_26911), .CLRB(_____), 
        .Q(_53006), .QN(_26744) );
  dffacs1 _________________________________________8__31_ ( .DIN(
        _____________________________256________), .CLK(_26902), .CLRB(_____), 
        .Q(_53138), .QN(_26276) );
  dffacs1 __________________________________________5__16_ ( .DIN(
        ______________________________145________), .CLK(_26920), .CLRB(_____), 
        .Q(_53089) );
  dffacs1 __________________________________________6__16_ ( .DIN(
        ______________________________177________), .CLK(_26909), .CLRB(_____), 
        .Q(_52988), .QN(_26418) );
  dffacs1 _________________________________________8__18_ ( .DIN(
        _____________________________243________), .CLK(_26863), .CLRB(_____), 
        .Q(_53110), .QN(_26713) );
  dffacs1 _________________________________________6__5_ ( .DIN(
        _____________________________166________), .CLK(_26880), .CLRB(_____), 
        .Q(_53256), .QN(_26272) );
  dffacs1 __________________________________________5__12_ ( .DIN(
        ______________________________141________), .CLK(_26942), .CLRB(_____), 
        .Q(_52942) );
  dffacs1 _________________________________________9__24_ ( .DIN(
        _____________________________281________), .CLK(_26862), .CLRB(_____), 
        .Q(_53068) );
  dffacs1 __________________________________________6__20_ ( .DIN(
        ______________________________181________), .CLK(_26955), .CLRB(_____), 
        .Q(_52832) );
  dffacs1 _________________________________________8__27_ ( .DIN(
        _____________________________252________), .CLK(_26861), .CLRB(_____), 
        .Q(_53230), .QN(_26683) );
  dffacs1 __________________________________________4__0_ ( .DIN(
        ______________________________97________), .CLK(_26897), .CLRB(_____), 
        .Q(_53002), .QN(_26736) );
  dffacs1 ___________________________________4_ ( .DIN(
        _________________________________4_________), .CLK(_26897), .CLRB(
        _____), .Q(_53508), .QN(_26723) );
  dffacs1 ____________________________________15_ ( .DIN(
        __________________________________15_________), .CLK(_26977), .CLRB(
        _____), .Q(_53488), .QN(_26742) );
  dffacs1 _________________________________________0__29_ ( .DIN(
        _________________________________________0________3____________), 
        .CLK(_26955), .CLRB(_____), .Q(_53052), .QN(_26530) );
  dffacs1 __________________________________________3__29_ ( .DIN(
        ______________________________94________), .CLK(_26952), .CLRB(_____), 
        .Q(_52958), .QN(_26383) );
  dffacs1 __________________________________________2__12_ ( .DIN(
        ______________________________45________), .CLK(_26857), .CLRB(_____), 
        .Q(_53128), .QN(_26561) );
  dffacs1 ____0________________12_0 ( .DIN(____0____________12_____), .CLK(
        _26909), .CLRB(_____), .Q(_53452), .QN(_26297) );
  dffacs1 ___________________________________16_ ( .DIN(
        _________________________________16_________), .CLK(_26957), .CLRB(
        _____), .Q(_53387), .QN(_26470) );
  dffacs1 ____3________________7_ ( .DIN(____3____________7_____), .CLK(_26876), .CLRB(_____), .Q(_53437), .QN(_26356) );
  dffacs1 __________________________________________5__5_ ( .DIN(
        ______________________________134________), .CLK(_26897), .CLRB(_____), 
        .Q(_52947) );
  dffacs1 _________________________________________6__10_ ( .DIN(
        _____________________________171________), .CLK(_26925), .CLRB(_____), 
        .Q(_53158) );
  dffacs1 __________________________________________2__2_ ( .DIN(
        ______________________________35________), .CLK(_26945), .CLRB(_____), 
        .Q(_53025) );
  dffacs1 __________________________________________6__25_ ( .DIN(
        ______________________________186________), .CLK(_26910), .CLRB(_____), 
        .Q(_53289), .QN(_26382) );
  dffacs1 ____1________________3_ ( .DIN(____1____________3_____), .CLK(_26930), .CLRB(_____), .Q(_53421), .QN(_26626) );
  dffacs1 ____0________________1_ ( .DIN(____0___________0_1_____), .CLK(
        _26918), .CLRB(_____), .Q(_53502), .QN(_26467) );
  dffacs1 ____2________________1_ ( .DIN(____2____________1_____), .CLK(_26984), .CLRB(_____), .Q(_53404), .QN(_26218) );
  dffacs1 ____0________________10_ ( .DIN(____0___________0_10_____), .CLK(
        _26894), .CLRB(_____), .Q(_53475), .QN(_26231) );
  dffacs1 __________________________________________1__6_ ( .DIN(
        ______________________________7________), .CLK(_26944), .CLRB(_____), 
        .Q(_52874), .QN(_26568) );
  dffacs1 ___________________________________14_ ( .DIN(
        _________________________________14_________), .CLK(_26974), .CLRB(
        _____), .Q(_53491), .QN(_26721) );
  dffacs1 _________________________________________5__23_ ( .DIN(
        _____________________________152________), .CLK(_26948), .CLRB(_____), 
        .Q(_53301) );
  dffacs1 __________________________________________3__5_ ( .DIN(
        ______________________________70________), .CLK(_26979), .CLRB(_____), 
        .Q(_52998) );
  dffacs1 _________________________________________7__15_ ( .DIN(
        _____________________________208________), .CLK(_26925), .CLRB(_____), 
        .Q(_53159), .QN(_26495) );
  dffacs1 _________________________________________7__1_ ( .DIN(
        _____________________________194________), .CLK(_26917), .CLRB(_____), 
        .Q(_53170) );
  dffacs1 __________________________________________3__19_ ( .DIN(
        ______________________________84________), .CLK(_26869), .CLRB(_____), 
        .Q(_52974) );
  dffacs1 __________________________________________4__12_ ( .DIN(
        ______________________________109________), .CLK(_26912), .CLRB(_____), 
        .Q(_53288), .QN(_26497) );
  dffacs1 _________________________________________6__1_ ( .DIN(
        _____________________________162________), .CLK(_26863), .CLRB(_____), 
        .Q(_53218), .QN(_26595) );
  dffacs1 __________________________________________3__20_ ( .DIN(
        ______________________________85________), .CLK(_26933), .CLRB(_____), 
        .Q(_53027), .QN(_26729) );
  dffacs1 _________________________________________2__10_ ( .DIN(
        _____________________________43________), .CLK(_26938), .CLRB(_____), 
        .Q(_53278), .QN(_26529) );
  dffacs1 _________________________________________5__16_ ( .DIN(
        _____________________________145________), .CLK(_26879), .CLRB(_____), 
        .Q(_53251) );
  dffacs1 _________________________________________2__15_ ( .DIN(
        _____________________________48________), .CLK(_26960), .CLRB(_____), 
        .Q(_53032), .QN(_26675) );
  dffacs1 _________________________________________8__4_ ( .DIN(
        _____________________________229________), .CLK(_26879), .CLRB(_____), 
        .Q(_53307), .QN(_26427) );
  dffacs1 __________________________________________5__10_ ( .DIN(
        ______________________________139________), .CLK(_26978), .CLRB(_____), 
        .Q(_52945) );
  dffacs1 ____________________________________28_ ( .DIN(
        __________________________________28_________), .CLK(_26975), .CLRB(
        _____), .Q(_53188), .QN(_26434) );
  dffacs1 __________________________________________6__23_ ( .DIN(
        ______________________________184________), .CLK(_26866), .CLRB(_____), 
        .Q(_53173) );
  dffacs1 _________________________________________1__4_ ( .DIN(
        _____________________________5________), .CLK(_26913), .CLRB(_____), 
        .Q(_53042), .QN(_26446) );
  dffacs1 _________________________________________7__5_ ( .DIN(
        _____________________________198________), .CLK(_26880), .CLRB(_____), 
        .Q(_53168), .QN(_26625) );
  dffacs1 __________________________________________6__0_ ( .DIN(
        ______________________________161________), .CLK(_26928), .CLRB(_____), 
        .Q(_52925), .QN(_26296) );
  dffacs1 _________________________________________7__31_ ( .DIN(
        _____________________________224________), .CLK(_26903), .CLRB(_____), 
        .Q(_53096), .QN(_26596) );
  dffacs1 __________________________________________6__28_ ( .DIN(
        ______________________________189________), .CLK(_26867), .CLRB(_____), 
        .Q(_53040), .QN(_26728) );
  dffacs1 ___________________________________0_ ( .DIN(
        _________________________________0_________), .CLK(_26924), .CLRB(
        _____), .Q(_53135) );
  dffacs1 _________________________________________9__2_ ( .DIN(
        _____________________________259________), .CLK(_26930), .CLRB(_____), 
        .Q(_53087), .QN(_26677) );
  dffacs1 __________________________________________4__24_ ( .DIN(
        ______________________________121________), .CLK(_26882), .CLRB(_____), 
        .Q(_52967), .QN(_26685) );
  dffacs1 __________________________________________3__27_ ( .DIN(
        ______________________________92________), .CLK(_26959), .CLRB(_____), 
        .Q(_53174) );
  dffacs1 __________________________________________5__22_ ( .DIN(
        ______________________________151________), .CLK(_26978), .CLRB(_____), 
        .Q(_52944), .QN(_26710) );
  dffacs1 _________________________________________8__21_ ( .DIN(
        _____________________________246________), .CLK(_26868), .CLRB(_____), 
        .Q(_53105), .QN(_26735) );
  dffacs1 __________________________________________4__4_ ( .DIN(
        ______________________________101________), .CLK(_26897), .CLRB(_____), 
        .Q(_53004) );
  dffacs1 _________________________________________1__8_ ( .DIN(
        _____________________________9________), .CLK(_26949), .CLRB(_____), 
        .Q(_53209) );
  dffacs1 ___________________________________9_ ( .DIN(
        _________________________________9_________), .CLK(_26896), .CLRB(
        _____), .Q(_53496), .QN(_26431) );
  dffacs1 ____0________________11_ ( .DIN(____0___________0_11_____), .CLK(
        _26963), .CLRB(_____), .Q(_53473), .QN(_26558) );
  dffacs1 ____3________________10_ ( .DIN(____3____________10_____), .CLK(
        _26876), .CLRB(_____), .Q(_53392), .QN(_26437) );
  dffacs1 ____3________________9_ ( .DIN(____3____________9_____), .CLK(_26901), .CLRB(_____), .Q(_53440), .QN(_26238) );
  dffacs1 __________________________________________0__21_ ( .DIN(
        __________________________________________21_________), .CLK(_26861), 
        .CLRB(_____), .Q(_53385) );
  dffacs1 ____________________________________4_ ( .DIN(
        __________________________________4_________), .CLK(_26952), .CLRB(
        _____), .Q(_53507) );
  dffacs1 _________________________________________3__22_ ( .DIN(
        _____________________________87________), .CLK(_26973), .CLRB(_____), 
        .Q(_53296) );
  dffacs1 _________________________________________0__31_ ( .DIN(
        _________________________________________0________5____________), 
        .CLK(_26962), .CLRB(_____), .Q(_53051), .QN(_26669) );
  dffacs1 _________________________________________0__7_ ( .DIN(
        _________________________________________8_________), .CLK(_26918), 
        .CLRB(_____), .Q(_53465), .QN(_26528) );
  dffacs1 ____3________________2_ ( .DIN(____3____________2_____), .CLK(_26901), .CLRB(_____), .Q(_53442), .QN(_26466) );
  dffacs1 _________________________________________6__3_ ( .DIN(
        _____________________________164________), .CLK(_26863), .CLRB(_____), 
        .Q(_53220), .QN(_26594) );
  dffacs1 ____________________________________27_ ( .DIN(
        __________________________________27_________), .CLK(_26942), .CLRB(
        _____), .Q(_53099) );
  dffacs1 _________________________________________4__1_ ( .DIN(
        _____________________________98________), .CLK(_26881), .CLRB(_____), 
        .Q(_53344), .QN(_26613) );
  dffacs1 __________________________________________6__6_ ( .DIN(
        ______________________________167________), .CLK(_26893), .CLRB(_____), 
        .Q(_53273) );
  dffacs1 _________________________________________8__0_ ( .DIN(
        _____________________________225________), .CLK(_26924), .CLRB(_____), 
        .Q(_53092) );
  dffacs1 ____________________________________30_ ( .DIN(
        __________________________________30_________), .CLK(_26886), .CLRB(
        _____), .Q(_53175), .QN(_26295) );
  dffacs1 _________________________________________1__22_ ( .DIN(
        _____________________________23________), .CLK(_26885), .CLRB(_____), 
        .Q(_53112) );
  dffacs1 _________________________________________4__9_ ( .DIN(
        _____________________________106________), .CLK(_26882), .CLRB(_____), 
        .Q(_53329), .QN(_26447) );
  dffacs1 _________________________________________8__6_ ( .DIN(
        _____________________________231________), .CLK(_26865), .CLRB(_____), 
        .Q(_53119) );
  dffacs1 _________________________________________6__11_ ( .DIN(
        _____________________________172________), .CLK(_26925), .CLRB(_____), 
        .Q(_53206), .QN(_26265) );
  dffacs1 _________________________________________3__29_ ( .DIN(
        _____________________________94________), .CLK(_26895), .CLRB(_____), 
        .Q(_53462), .QN(_26740) );
  dffacs1 _________________________________________2__1_ ( .DIN(
        _____________________________34________), .CLK(_26856), .CLRB(_____), 
        .Q(_52841) );
  dffacs1 _________________________________________9__20_ ( .DIN(
        _____________________________277________), .CLK(_26862), .CLRB(_____), 
        .Q(_53077) );
  dffacs1 ___________________________________6_ ( .DIN(
        _________________________________6_________), .CLK(_26931), .CLRB(
        _____), .Q(_53498) );
  dffacs1 ____0________________5_0 ( .DIN(____0____________5_____), .CLK(
        _26886), .CLRB(_____), .Q(_53445), .QN(_26207) );
  dffacs1 _________________________________________5__31_ ( .DIN(
        _____________________________160________), .CLK(_26903), .CLRB(_____), 
        .Q(_53277), .QN(_26619) );
  dffacs1 ___________________________________31_ ( .DIN(
        _________________________________31_________), .CLK(_26923), .CLRB(
        _____), .Q(_53378) );
  dffacs1 ____________________________________10_ ( .DIN(
        __________________________________10_________), .CLK(_26931), .CLRB(
        _____), .Q(_52848), .QN(_26660) );
  dffacs1 __________________________________________2__18_ ( .DIN(
        ______________________________51________), .CLK(_26926), .CLRB(_____), 
        .Q(_52898) );
  dffacs1 ____2________________6_ ( .DIN(____2____________6_____), .CLK(_26983), .CLRB(_____), .Q(_53411) );
  dffacs1 _________________________________________2__16_ ( .DIN(
        _____________________________49________), .CLK(_26960), .CLRB(_____), 
        .Q(_53010) );
  dffacs1 _________________________________________4__21_ ( .DIN(
        _____________________________118________), .CLK(_26959), .CLRB(_____), 
        .Q(_53239) );
  dffacs1 ___________________________________7_ ( .DIN(
        _________________________________7_________), .CLK(_26930), .CLRB(
        _____), .Q(_53057), .QN(_26739) );
  dffacs1 ____________________________________13_ ( .DIN(
        __________________________________13_________), .CLK(_26976), .CLRB(
        _____), .Q(_52847) );
  dffacs1 __________________________________________1__14_ ( .DIN(
        ______________________________15________), .CLK(_26943), .CLRB(_____), 
        .Q(_53469), .QN(_26592) );
  dffacs1 ____1________________9_ ( .DIN(____1____________9_____), .CLK(_26979), .CLRB(_____), .Q(_53429), .QN(_26334) );
  dffacs1 ___________________________________2_ ( .DIN(
        _________________________________2_________), .CLK(_26887), .CLRB(
        _____), .Q(_53134), .QN(_26727) );
  dffacs1 ____0________________9_ ( .DIN(____0___________0_9_____), .CLK(
        _26889), .CLRB(_____), .Q(_53477), .QN(_26325) );
  dffacs1 _________________________________________6__15_ ( .DIN(
        _____________________________176________), .CLK(_26919), .CLRB(_____), 
        .Q(_53205) );
  dffacs1 ____0________________2_0 ( .DIN(____0____________2_____), .CLK(
        _26979), .CLRB(_____), .Q(_53444), .QN(_26624) );
  dffacs1 __________________________________________2__23_ ( .DIN(
        ______________________________56________), .CLK(_26860), .CLRB(_____), 
        .Q(_52862), .QN(_26666) );
  dffacs1 _________________________________________7__27_ ( .DIN(
        _____________________________220________), .CLK(_26936), .CLRB(_____), 
        .Q(_53098), .QN(_26616) );
  dffacs1 __________________________________________1__9_ ( .DIN(
        ______________________________10________), .CLK(_26944), .CLRB(_____), 
        .Q(_52966), .QN(_26304) );
  dffacs1 ___________________________________10_ ( .DIN(
        _________________________________10_________), .CLK(_26979), .CLRB(
        _____), .Q(_53495), .QN(_26577) );
  dffacs1 ____________________________________21_ ( .DIN(
        __________________________________21_________), .CLK(_26956), .CLRB(
        _____), .Q(_53481), .QN(_26703) );
  dffacs1 _________________________________________3__20_ ( .DIN(
        _____________________________85________), .CLK(_26870), .CLRB(_____), 
        .Q(_53221) );
  dffacs1 ____0________________2_ ( .DIN(____0___________0_2_____), .CLK(
        _26963), .CLRB(_____), .Q(_53501) );
  dffacs1 ____0________________8_0 ( .DIN(____0____________8_____), .CLK(
        _26911), .CLRB(_____), .Q(_53457), .QN(_26353) );
  dffacs1 ____2________________8_ ( .DIN(____2____________8_____), .CLK(_26875), .CLRB(_____), .Q(_53407), .QN(_26208) );
  dffacs1 ___________________________________3_ ( .DIN(
        _________________________________3_________), .CLK(_26929), .CLRB(
        _____), .Q(_53510), .QN(_26551) );
  dffacs1 ____0________________4_0 ( .DIN(____0____________4_____), .CLK(
        _26977), .CLRB(_____), .Q(_53449), .QN(_26408) );
  dffacs1 _________________________________________6__24_ ( .DIN(
        _____________________________185________), .CLK(_26972), .CLRB(_____), 
        .Q(_53342) );
  dffacs1 __________________________________________3__10_ ( .DIN(
        ______________________________75________), .CLK(_26887), .CLRB(_____), 
        .Q(_53432) );
  dffacs1 ____________________________________7_ ( .DIN(
        __________________________________7_________), .CLK(_26976), .CLRB(
        _____), .Q(_53360) );
  dffacs1 ____________________________________24_ ( .DIN(
        __________________________________24_________), .CLK(_26866), .CLRB(
        _____), .Q(_52981), .QN(_26659) );
  dffacs1 __________________________________________2__11_ ( .DIN(
        ______________________________44________), .CLK(_26857), .CLRB(_____), 
        .Q(_52869) );
  dffacs1 ___________________________________25_ ( .DIN(
        _________________________________25_________), .CLK(_26934), .CLRB(
        _____), .Q(_52978) );
  dffacs1 __________________________________________1__21_ ( .DIN(
        ______________________________22________), .CLK(_26860), .CLRB(_____), 
        .Q(_52918), .QN(_26674) );
  dffacs1 _________________________________________1__27_ ( .DIN(
        _____________________________28________), .CLK(_26874), .CLRB(_____), 
        .Q(_53022) );
  dffacs1 __________________________________________5__1_ ( .DIN(
        ______________________________130________), .CLK(_26956), .CLRB(_____), 
        .Q(_52952), .QN(_26733) );
  dffacs1 _________________________________________8__23_ ( .DIN(
        _____________________________248________), .CLK(_26881), .CLRB(_____), 
        .Q(_53109), .QN(_26738) );
  dffacs1 ____________________________________2_ ( .DIN(
        __________________________________2_________), .CLK(_26928), .CLRB(
        _____), .Q(_53506) );
  dffacs1 _________________________________________0__26_ ( .DIN(
        _________________________________________0________0____________), 
        .CLK(_26900), .CLRB(_____), .Q(_53067), .QN(_26593) );
  dffacs1 ____0________________14_ ( .DIN(____0____________14_____), .CLK(
        _26901), .CLRB(_____), .Q(_53455), .QN(_26465) );
  dffacs1 _________________________________________1__1_ ( .DIN(
        _____________________________2________), .CLK(_26856), .CLRB(_____), 
        .Q(_53080) );
  dffacs1 __________________________________________2__3_ ( .DIN(
        ______________________________36________), .CLK(_26944), .CLRB(_____), 
        .Q(_52882) );
  dffacs1 __________________________________________0__22_ ( .DIN(
        __________________________________________22_________), .CLK(_26934), 
        .CLRB(_____), .Q(_53237) );
  dffacs1 __________________________________________0__30_ ( .DIN(
        __________________________________________25________4____________), 
        .CLK(_26868), .CLRB(_____), .Q(_52842) );
  dffacs1 ___________________________________15_ ( .DIN(
        _________________________________15_________), .CLK(_26863), .CLRB(
        _____), .Q(_53489), .QN(_26464) );
  dffacs1 ____2________________9_ ( .DIN(____2____________9_____), .CLK(_26875), .CLRB(_____), .Q(_53406), .QN(_26615) );
  dffacs1 ____________________________________9_ ( .DIN(
        __________________________________9_________), .CLK(_26914), .CLRB(
        _____), .Q(_53125), .QN(_26607) );
  dffacs1 __________________________________________0__0_ ( .DIN(
        __________________________________________0_________), .CLK(_26951), 
        .CLRB(_____), .Q(_53064), .QN(_26654) );
  dffacs1 ____________________________________6_ ( .DIN(
        __________________________________6_________), .CLK(_26976), .CLRB(
        _____), .Q(_53156) );
  dffacs1 _____________23_ ( .DIN(_26787), .CLK(_26940), .CLRB(_____), .Q(
        _______[23]) );
  dffacs1 _____________4_ ( .DIN(_640), .CLK(_26951), .CLRB(_____), .Q(
        _______[4]) );
  dffacs1 _____________2_ ( .DIN(_26795), .CLK(_26951), .CLRB(_____), .Q(
        _______[2]) );
  dffacs1 _____________29_ ( .DIN(_359), .CLK(_26940), .CLRB(_____), .Q(
        _______[29]) );
  dffacs1 _____________25_ ( .DIN(_26823), .CLK(_26950), .CLRB(_____), .Q(
        _______[25]) );
  dffacs1 _____________14_ ( .DIN(_26791), .CLK(_26927), .CLRB(_____), .Q(
        _______[14]) );
  dffacs1 _____________11_ ( .DIN(_26824), .CLK(_26952), .CLRB(_____), .Q(
        _______[11]) );
  dffacs1 _____________7_ ( .DIN(_438), .CLK(_26930), .CLRB(_____), .Q(
        _______[7]) );
  dffacs1 _____________6_ ( .DIN(_26794), .CLK(_26956), .CLRB(_____), .Q(
        _______[6]) );
  dffacs1 _____________16_ ( .DIN(_408), .CLK(_26943), .CLRB(_____), .Q(
        _______[16]) );
  dffacs1 _____________12_ ( .DIN(_420), .CLK(_26941), .CLRB(_____), .Q(
        _______[12]) );
  dffacs1 _____________1_ ( .DIN(_26820), .CLK(_26955), .CLRB(_____), .Q(
        _______[1]) );
  dffacs1 _____________26_ ( .DIN(_356), .CLK(_26856), .CLRB(_____), .Q(
        _______[26]) );
  dffacs1 _____________5_ ( .DIN(_14172), .CLK(_26867), .CLRB(_____), .Q(
        _______[5]) );
  dffacs1 _____________30_ ( .DIN(_15544), .CLK(_26940), .CLRB(_____), .Q(
        _______[30]) );
  dffacs1 _____________28_ ( .DIN(_15546), .CLK(_26933), .CLRB(_____), .Q(
        _______[28]) );
  dffacs1 _____________22_ ( .DIN(_15550), .CLK(_26941), .CLRB(_____), .Q(
        _______[22]) );
  dffacs1 _____________21_ ( .DIN(_15551), .CLK(_26965), .CLRB(_____), .Q(
        _______[21]) );
  dffacs1 _____________18_ ( .DIN(_15553), .CLK(_26927), .CLRB(_____), .Q(
        _______[18]) );
  dffacs1 _____________15_ ( .DIN(_15555), .CLK(_26927), .CLRB(_____), .Q(
        _______[15]) );
  dffacs1 _____________10_ ( .DIN(_15560), .CLK(_26927), .CLRB(_____), .Q(
        _______[10]) );
  dffacs1 _____________9_ ( .DIN(_15561), .CLK(_26896), .CLRB(_____), .Q(
        _______[9]) );
  dffacs1 _____________8_ ( .DIN(_433), .CLK(_26927), .CLRB(_____), .Q(
        _______[8]) );
  dffacs1 _____________3_ ( .DIN(_15563), .CLK(_26887), .CLRB(_____), .Q(
        _______[3]) );
  dffacs1 _____________31_ ( .DIN(_922), .CLK(_26948), .CLRB(_____), .Q(
        _______[31]) );
  dffacs1 _____________17_ ( .DIN(_26204), .CLK(_26939), .CLRB(_____), .Q(
        _______[17]) );
  dffacs1 _____________0_ ( .DIN(_654), .CLK(_26932), .CLRB(_____), .Q(
        _______[0]) );
  dffacs1 _____________24_ ( .DIN(_353), .CLK(_26939), .CLRB(_____), .Q(
        _______[24]) );
  dffacs1 _____________20_ ( .DIN(_26205), .CLK(_26894), .CLRB(_____), .Q(
        _______[20]) );
  dffacs1 _____________19_ ( .DIN(_398), .CLK(_26953), .CLRB(_____), .Q(
        _______[19]) );
  dffacs1 _____________27_ ( .DIN(_15547), .CLK(_26861), .CLRB(_____), .Q(
        _______[27]) );
  dffacs1 _____________13_ ( .DIN(_26206), .CLK(_26857), .CLRB(_____), .Q(
        _______[13]) );
  dffacs1 _______________25_ ( .DIN(
        _______25____2________________25____________________), .CLK(___), 
        .CLRB(_____), .Q(_53368), .QN(_26780) );
  dffacs1 _________________________________________8__20_ ( .DIN(
        _____________________________245________), .CLK(_26910), .CLRB(_____), 
        .Q(_53108), .QN(_26748) );
  dffacs1 _________________________________________8__29_ ( .DIN(
        _____________________________254________), .CLK(_26918), .CLRB(_____), 
        .Q(_53171), .QN(_26746) );
  dffacs1 _________________________________________0__22_ ( .DIN(
        _________________________________________23_________), .CLK(_26954), 
        .CLRB(_____), .Q(_53115), .QN(_26717) );
  dffacs1 _________________________________________7__13_ ( .DIN(
        _____________________________206________), .CLK(_26968), .CLRB(_____), 
        .Q(_26684), .QN(_53153) );
  dffacs1 _______________3_ ( .DIN(
        _______3____2________________3____________________), .CLK(_26981), 
        .CLRB(_____), .Q(_26341), .QN(_53467) );
  dffacs1 _______________30_ ( .DIN(
        _______30____2________________30____________________), .CLK(_26937), 
        .CLRB(_____), .Q(_53363), .QN(_26335) );
  dffacs1 _______________2_ ( .DIN(
        _______2____2________________2____________________), .CLK(_26982), 
        .CLRB(_____), .Q(_53353), .QN(_26329) );
  dffacs1 _________________________________________0__10_ ( .DIN(
        _________________________________________11_________), .CLK(___), 
        .CLRB(_____), .Q(_53295) );
  nnd2s1 _26868_inst ( .DIN1(_26772), .DIN2(_39002), .Q(_26289) );
  hi1s1 _26869_inst ( .DIN(_48218), .Q(_26844) );
  xnr2s1 _26870_inst ( .DIN1(_29579), .DIN2(_46010), .Q(_26317) );
  and2s1 _26871_inst ( .DIN1(_46052), .DIN2(_46053), .Q(_26337) );
  nnd2s1 _26872_inst ( .DIN1(_48117), .DIN2(_26792), .Q(_26361) );
  ib1s1 _26873_inst ( .DIN(_51796), .Q(_26847) );
  xnr2s1 _26874_inst ( .DIN1(_15550), .DIN2(_31884), .Q(_26589) );
  xor2s1 _26875_inst ( .DIN1(_34515), .DIN2(_38354), .Q(_26759) );
  xor2s1 _26876_inst ( .DIN1(_27620), .DIN2(_38304), .Q(_26760) );
  xor2s1 _26877_inst ( .DIN1(_26526), .DIN2(_35860), .Q(_26761) );
  xor2s1 _26878_inst ( .DIN1(_34515), .DIN2(_34517), .Q(_26762) );
  xor2s1 _26879_inst ( .DIN1(_34515), .DIN2(_35168), .Q(_26763) );
  hi1s1 _26880_inst ( .DIN(_26589), .Q(_26764) );
  hi1s1 _26881_inst ( .DIN(_26317), .Q(_26765) );
  hi1s1 _26882_inst ( .DIN(_26852), .Q(_26766) );
  hi1s1 _26883_inst ( .DIN(_26851), .Q(_26767) );
  hi1s1 _26884_inst ( .DIN(_26783), .Q(_26768) );
  hi1s1 _26885_inst ( .DIN(_26783), .Q(_26769) );
  ib1s1 _26886_inst ( .DIN(_26337), .Q(_26770) );
  ib1s1 _26887_inst ( .DIN(______[16]), .Q(_26771) );
  ib1s1 _26888_inst ( .DIN(______[16]), .Q(_26772) );
  ib1s1 _26889_inst ( .DIN(______[28]), .Q(_26773) );
  ib1s1 _26890_inst ( .DIN(______[28]), .Q(_26774) );
  ib1s1 _26891_inst ( .DIN(_33225), .Q(_26775) );
  xnr2s1 _26892_inst ( .DIN1(_29231), .DIN2(_38185), .Q(_38207) );
  ib1s1 _26893_inst ( .DIN(_38207), .Q(_26776) );
  ib1s1 _26894_inst ( .DIN(_53361), .Q(_34515) );
  xnr2s1 _26895_inst ( .DIN1(_31802), .DIN2(_31803), .Q(_31723) );
  ib1s1 _26896_inst ( .DIN(_31723), .Q(_26777) );
  ib1s1 _26897_inst ( .DIN(_32979), .Q(_26779) );
  ib1s1 _26898_inst ( .DIN(_26780), .Q(_26781) );
  and2s1 _26899_inst ( .DIN1(______[21]), .DIN2(_46127), .Q(_46227) );
  ib1s1 _26900_inst ( .DIN(_46227), .Q(_26782) );
  ib1s1 _26901_inst ( .DIN(______[7]), .Q(_39015) );
  ib1s1 _26902_inst ( .DIN(_51281), .Q(_50605) );
  and2s1 _26903_inst ( .DIN1(______[24]), .DIN2(_48130), .Q(_48179) );
  ib1s1 _26904_inst ( .DIN(_48179), .Q(_26783) );
  xnr2s1 _26905_inst ( .DIN1(_26318), .DIN2(_38875), .Q(_38906) );
  ib1s1 _26906_inst ( .DIN(_38906), .Q(_26784) );
  xnr2s1 _26907_inst ( .DIN1(_34787), .DIN2(_38276), .Q(_38598) );
  ib1s1 _26908_inst ( .DIN(_38598), .Q(_26785) );
  xnr2s1 _26909_inst ( .DIN1(_26780), .DIN2(_38407), .Q(_38420) );
  ib1s1 _26910_inst ( .DIN(_38420), .Q(_26786) );
  ib1s1 _26911_inst ( .DIN(_53364), .Q(_27620) );
  ib1s1 _26912_inst ( .DIN(_29332), .Q(_26787) );
  ib1s1 _26913_inst ( .DIN(_382), .Q(_29332) );
  hi1s1 _26914_inst ( .DIN(_31718), .Q(_26788) );
  ib1s1 _26915_inst ( .DIN(_26788), .Q(_26789) );
  ib1s1 _26916_inst ( .DIN(_359), .Q(_31483) );
  ib1s1 _26917_inst ( .DIN(_33333), .Q(_26790) );
  ib1s1 _26918_inst ( .DIN(_29580), .Q(_26791) );
  ib1s1 _26919_inst ( .DIN(_414), .Q(_29580) );
  ib1s1 _26920_inst ( .DIN(_46961), .Q(_26792) );
  ib1s1 _26921_inst ( .DIN(_41360), .Q(_26793) );
  ib1s1 _26922_inst ( .DIN(_32715), .Q(_26794) );
  ib1s1 _26923_inst ( .DIN(_441), .Q(_32715) );
  ib1s1 _26924_inst ( .DIN(_32713), .Q(_26795) );
  ib1s1 _26925_inst ( .DIN(_27175), .Q(_26796) );
  ib1s1 _26926_inst ( .DIN(_33123), .Q(_26797) );
  ib1s1 _26927_inst ( .DIN(_29752), .Q(_26798) );
  ib1s1 _26928_inst ( .DIN(_44715), .Q(_26799) );
  ib1s1 _26929_inst ( .DIN(_44771), .Q(_44715) );
  ib1s1 _26930_inst ( .DIN(_33082), .Q(_26800) );
  ib1s1 _26931_inst ( .DIN(_34034), .Q(_26801) );
  ib1s1 _26932_inst ( .DIN(_33396), .Q(_26802) );
  ib1s1 _26933_inst ( .DIN(______[14]), .Q(_27651) );
  ib1s1 _26934_inst ( .DIN(______[24]), .Q(_27082) );
  ib1s1 _26935_inst ( .DIN(_44725), .Q(_26804) );
  ib1s1 _26936_inst ( .DIN(_26804), .Q(_26805) );
  hi1s1 _26937_inst ( .DIN(_48130), .Q(_26806) );
  ib1s1 _26938_inst ( .DIN(_48130), .Q(_48332) );
  and2s1 _26939_inst ( .DIN1(______[9]), .DIN2(_26772), .Q(_51816) );
  ib1s1 _26940_inst ( .DIN(_51816), .Q(_26807) );
  ib1s1 _26941_inst ( .DIN(_26807), .Q(_51818) );
  ib1s1 _26942_inst ( .DIN(______[30]), .Q(_26808) );
  ib1s1 _26943_inst ( .DIN(______[30]), .Q(_28100) );
  ib1s1 _26944_inst ( .DIN(______[26]), .Q(_26809) );
  ib1s1 _26945_inst ( .DIN(______[26]), .Q(_27365) );
  xnr2s1 _26946_inst ( .DIN1(_26319), .DIN2(_37979), .Q(_38272) );
  ib1s1 _26947_inst ( .DIN(_38272), .Q(_26810) );
  xnr2s1 _26948_inst ( .DIN1(_26332), .DIN2(_38595), .Q(_38594) );
  ib1s1 _26949_inst ( .DIN(_38594), .Q(_26811) );
  ib1s1 _26950_inst ( .DIN(_31976), .Q(_26205) );
  xnr2s1 _26951_inst ( .DIN1(_34787), .DIN2(_38846), .Q(_38871) );
  ib1s1 _26952_inst ( .DIN(_38871), .Q(_26812) );
  ib1s1 _26953_inst ( .DIN(_31515), .Q(_15544) );
  xnr2s1 _26954_inst ( .DIN1(_26322), .DIN2(_37591), .Q(_37786) );
  ib1s1 _26955_inst ( .DIN(_37786), .Q(_26813) );
  xnr2s1 _26956_inst ( .DIN1(_36332), .DIN2(_36334), .Q(_36538) );
  ib1s1 _26957_inst ( .DIN(_36538), .Q(_26814) );
  xnr2s1 _26958_inst ( .DIN1(_26318), .DIN2(_38597), .Q(_38596) );
  ib1s1 _26959_inst ( .DIN(_38596), .Q(_26815) );
  xor2s1 _26960_inst ( .DIN1(_27338), .DIN2(_42653), .Q(_26816) );
  ib1s1 _26961_inst ( .DIN(_27329), .Q(_27338) );
  ib1s1 _26962_inst ( .DIN(_53346), .Q(_27558) );
  xnr2s1 _26963_inst ( .DIN1(_398), .DIN2(_15551), .Q(_31993) );
  ib1s1 _26964_inst ( .DIN(_31993), .Q(_26817) );
  xnr2s1 _26965_inst ( .DIN1(_15563), .DIN2(_14172), .Q(_32654) );
  ib1s1 _26966_inst ( .DIN(_32654), .Q(_26818) );
  ib1s1 _26967_inst ( .DIN(_32169), .Q(_15553) );
  xnr2s1 _26968_inst ( .DIN1(_15555), .DIN2(_26204), .Q(_32204) );
  ib1s1 _26969_inst ( .DIN(_32204), .Q(_26819) );
  ib1s1 _26970_inst ( .DIN(_32219), .Q(_26204) );
  ib1s1 _26971_inst ( .DIN(_32707), .Q(_26820) );
  ib1s1 _26972_inst ( .DIN(_652), .Q(_32707) );
  xnr2s1 _26973_inst ( .DIN1(_433), .DIN2(_15560), .Q(_32670) );
  ib1s1 _26974_inst ( .DIN(_32670), .Q(_26821) );
  ib1s1 _26975_inst ( .DIN(_33315), .Q(_26822) );
  ib1s1 _26976_inst ( .DIN(_29304), .Q(_26823) );
  ib1s1 _26977_inst ( .DIN(_355), .Q(_29304) );
  ib1s1 _26978_inst ( .DIN(_32473), .Q(_26824) );
  ib1s1 _26979_inst ( .DIN(_43336), .Q(_26825) );
  ib1s1 _26980_inst ( .DIN(_32211), .Q(_26826) );
  ib1s1 _26981_inst ( .DIN(_408), .Q(_32211) );
  ib1s1 _26982_inst ( .DIN(_29871), .Q(_26827) );
  ib1s1 _26983_inst ( .DIN(_640), .Q(_29871) );
  ib1s1 _26984_inst ( .DIN(_33029), .Q(_26828) );
  ib1s1 _26985_inst ( .DIN(_32479), .Q(_26829) );
  ib1s1 _26986_inst ( .DIN(_31670), .Q(_26830) );
  xnr2s1 _26987_inst ( .DIN1(_37171), .DIN2(_37182), .Q(_33435) );
  ib1s1 _26988_inst ( .DIN(_33435), .Q(_26831) );
  ib1s1 _26989_inst ( .DIN(_33172), .Q(_26832) );
  xnr2s1 _26990_inst ( .DIN1(_37238), .DIN2(_37254), .Q(_33480) );
  ib1s1 _26991_inst ( .DIN(_33480), .Q(_26833) );
  xnr2s1 _26992_inst ( .DIN1(_36921), .DIN2(_36942), .Q(_33246) );
  ib1s1 _26993_inst ( .DIN(_33246), .Q(_26834) );
  ib1s1 _26994_inst ( .DIN(______[22]), .Q(_27039) );
  ib1s1 _26995_inst ( .DIN(______[10]), .Q(_27614) );
  ib1s1 _26996_inst ( .DIN(______[4]), .Q(_28684) );
  ib1s1 _26997_inst ( .DIN(_51888), .Q(_26835) );
  ib1s1 _26998_inst ( .DIN(_51802), .Q(_51888) );
  ib1s1 _26999_inst ( .DIN(_47228), .Q(_46961) );
  xor2s1 _27000_inst ( .DIN1(_31233), .DIN2(_29231), .Q(_29169) );
  ib1s1 _27001_inst ( .DIN(_29169), .Q(_26836) );
  ib1s1 _27002_inst ( .DIN(_26836), .Q(_29166) );
  ib1s1 _27003_inst ( .DIN(______[12]), .Q(_27774) );
  ib1s1 _27004_inst ( .DIN(______[2]), .Q(_27393) );
  ib1s1 _27005_inst ( .DIN(_41903), .Q(_26837) );
  ib1s1 _27006_inst ( .DIN(_42312), .Q(_41903) );
  ib1s1 _27007_inst ( .DIN(_39383), .Q(_26838) );
  ib1s1 _27008_inst ( .DIN(_39537), .Q(_39383) );
  ib1s1 _27009_inst ( .DIN(_46112), .Q(_26839) );
  ib1s1 _27010_inst ( .DIN(_26839), .Q(_26840) );
  ib1s1 _27011_inst ( .DIN(_40581), .Q(_26841) );
  ib1s1 _27012_inst ( .DIN(_26841), .Q(_26842) );
  ib1s1 _27013_inst ( .DIN(______[18]), .Q(_27291) );
  and2s1 _27014_inst ( .DIN1(_48130), .DIN2(_27082), .Q(_48218) );
  ib1s1 _27015_inst ( .DIN(_48218), .Q(_26843) );
  ib1s1 _27016_inst ( .DIN(_26843), .Q(_48137) );
  and2s1 _27017_inst ( .DIN1(______[7]), .DIN2(_26774), .Q(_44760) );
  ib1s1 _27018_inst ( .DIN(_44760), .Q(_26845) );
  ib1s1 _27019_inst ( .DIN(_26845), .Q(_44951) );
  ib1s1 _27020_inst ( .DIN(______[6]), .Q(_26846) );
  ib1s1 _27021_inst ( .DIN(______[6]), .Q(_28646) );
  ib1s1 _27022_inst ( .DIN(_26847), .Q(_26848) );
  ib1s1 _27023_inst ( .DIN(_26803), .Q(_26849) );
  ib1s1 _27024_inst ( .DIN(_26849), .Q(_26850) );
  and2s1 _27025_inst ( .DIN1(_26774), .DIN2(_39015), .Q(_45044) );
  ib1s1 _27026_inst ( .DIN(_45044), .Q(_26851) );
  ib1s1 _27027_inst ( .DIN(_45044), .Q(_26852) );
  ib1s1 _27028_inst ( .DIN(______[20]), .Q(_26853) );
  ib1s1 _27029_inst ( .DIN(______[20]), .Q(_27448) );
  ib1s1 _27030_inst ( .DIN(______[8]), .Q(_26854) );
  ib1s1 _27031_inst ( .DIN(______[8]), .Q(_27066) );
  ib1s1 _27032_inst ( .DIN(______[0]), .Q(_26855) );
  ib1s1 _27033_inst ( .DIN(______[0]), .Q(_27241) );
  hi1s1 _27034_inst ( .DIN(_26988), .Q(_26856) );
  hi1s1 _27035_inst ( .DIN(_26988), .Q(_26857) );
  hi1s1 _27036_inst ( .DIN(_26988), .Q(_26858) );
  hi1s1 _27037_inst ( .DIN(_26988), .Q(_26859) );
  hi1s1 _27038_inst ( .DIN(_26988), .Q(_26860) );
  hi1s1 _27039_inst ( .DIN(_26987), .Q(_26861) );
  hi1s1 _27040_inst ( .DIN(_26990), .Q(_26862) );
  hi1s1 _27041_inst ( .DIN(_26990), .Q(_26863) );
  hi1s1 _27042_inst ( .DIN(_26988), .Q(_26864) );
  hi1s1 _27043_inst ( .DIN(_26988), .Q(_26865) );
  hi1s1 _27044_inst ( .DIN(_26989), .Q(_26866) );
  hi1s1 _27045_inst ( .DIN(_26990), .Q(_26867) );
  hi1s1 _27046_inst ( .DIN(_26989), .Q(_26868) );
  hi1s1 _27047_inst ( .DIN(_26991), .Q(_26869) );
  hi1s1 _27048_inst ( .DIN(_26987), .Q(_26870) );
  hi1s1 _27049_inst ( .DIN(_26991), .Q(_26871) );
  hi1s1 _27050_inst ( .DIN(_26987), .Q(_26872) );
  hi1s1 _27051_inst ( .DIN(_26989), .Q(_26873) );
  hi1s1 _27052_inst ( .DIN(_26991), .Q(_26874) );
  hi1s1 _27053_inst ( .DIN(_26988), .Q(_26875) );
  hi1s1 _27054_inst ( .DIN(_26988), .Q(_26876) );
  hi1s1 _27055_inst ( .DIN(_26991), .Q(_26877) );
  hi1s1 _27056_inst ( .DIN(_26988), .Q(_26878) );
  hi1s1 _27057_inst ( .DIN(_26989), .Q(_26879) );
  hi1s1 _27058_inst ( .DIN(_26990), .Q(_26880) );
  hi1s1 _27059_inst ( .DIN(_26987), .Q(_26881) );
  hi1s1 _27060_inst ( .DIN(_26990), .Q(_26882) );
  hi1s1 _27061_inst ( .DIN(_26988), .Q(_26883) );
  hi1s1 _27062_inst ( .DIN(_26989), .Q(_26884) );
  hi1s1 _27063_inst ( .DIN(_26990), .Q(_26885) );
  hi1s1 _27064_inst ( .DIN(_26988), .Q(_26886) );
  hi1s1 _27065_inst ( .DIN(_26991), .Q(_26887) );
  hi1s1 _27066_inst ( .DIN(_26987), .Q(_26888) );
  hi1s1 _27067_inst ( .DIN(_26991), .Q(_26889) );
  hi1s1 _27068_inst ( .DIN(_26991), .Q(_26890) );
  hi1s1 _27069_inst ( .DIN(_26989), .Q(_26891) );
  hi1s1 _27070_inst ( .DIN(_26990), .Q(_26892) );
  hi1s1 _27071_inst ( .DIN(_26988), .Q(_26893) );
  hi1s1 _27072_inst ( .DIN(_26991), .Q(_26894) );
  hi1s1 _27073_inst ( .DIN(_26988), .Q(_26895) );
  hi1s1 _27074_inst ( .DIN(_26987), .Q(_26896) );
  hi1s1 _27075_inst ( .DIN(_26991), .Q(_26897) );
  hi1s1 _27076_inst ( .DIN(_26988), .Q(_26898) );
  hi1s1 _27077_inst ( .DIN(_26987), .Q(_26899) );
  hi1s1 _27078_inst ( .DIN(_26991), .Q(_26900) );
  hi1s1 _27079_inst ( .DIN(_26987), .Q(_26901) );
  hi1s1 _27080_inst ( .DIN(_26989), .Q(_26902) );
  hi1s1 _27081_inst ( .DIN(_26989), .Q(_26903) );
  hi1s1 _27082_inst ( .DIN(_26987), .Q(_26904) );
  hi1s1 _27083_inst ( .DIN(_26989), .Q(_26905) );
  hi1s1 _27084_inst ( .DIN(_26990), .Q(_26906) );
  hi1s1 _27085_inst ( .DIN(_26988), .Q(_26907) );
  hi1s1 _27086_inst ( .DIN(_26991), .Q(_26908) );
  hi1s1 _27087_inst ( .DIN(_26987), .Q(_26909) );
  hi1s1 _27088_inst ( .DIN(_26990), .Q(_26910) );
  hi1s1 _27089_inst ( .DIN(_26989), .Q(_26911) );
  hi1s1 _27090_inst ( .DIN(_26990), .Q(_26912) );
  hi1s1 _27091_inst ( .DIN(_26988), .Q(_26913) );
  hi1s1 _27092_inst ( .DIN(_26987), .Q(_26914) );
  hi1s1 _27093_inst ( .DIN(_26988), .Q(_26915) );
  hi1s1 _27094_inst ( .DIN(_26987), .Q(_26916) );
  hi1s1 _27095_inst ( .DIN(_26989), .Q(_26917) );
  hi1s1 _27096_inst ( .DIN(_26990), .Q(_26918) );
  hi1s1 _27097_inst ( .DIN(_26988), .Q(_26919) );
  hi1s1 _27098_inst ( .DIN(_26991), .Q(_26920) );
  hi1s1 _27099_inst ( .DIN(_26987), .Q(_26921) );
  hi1s1 _27100_inst ( .DIN(_26989), .Q(_26922) );
  hi1s1 _27101_inst ( .DIN(_26990), .Q(_26923) );
  hi1s1 _27102_inst ( .DIN(_26988), .Q(_26924) );
  hi1s1 _27103_inst ( .DIN(_26991), .Q(_26925) );
  hi1s1 _27104_inst ( .DIN(_26989), .Q(_26926) );
  hi1s1 _27105_inst ( .DIN(_26990), .Q(_26927) );
  hi1s1 _27106_inst ( .DIN(_26991), .Q(_26928) );
  hi1s1 _27107_inst ( .DIN(_26987), .Q(_26929) );
  hi1s1 _27108_inst ( .DIN(_26990), .Q(_26930) );
  hi1s1 _27109_inst ( .DIN(_26987), .Q(_26931) );
  hi1s1 _27110_inst ( .DIN(_26987), .Q(_26932) );
  hi1s1 _27111_inst ( .DIN(_26988), .Q(_26933) );
  hi1s1 _27112_inst ( .DIN(_26988), .Q(_26934) );
  hi1s1 _27113_inst ( .DIN(_26990), .Q(_26935) );
  hi1s1 _27114_inst ( .DIN(_26989), .Q(_26936) );
  hi1s1 _27115_inst ( .DIN(_26989), .Q(_26937) );
  hi1s1 _27116_inst ( .DIN(_26989), .Q(_26938) );
  hi1s1 _27117_inst ( .DIN(_26989), .Q(_26939) );
  hi1s1 _27118_inst ( .DIN(_26989), .Q(_26940) );
  hi1s1 _27119_inst ( .DIN(_26989), .Q(_26941) );
  hi1s1 _27120_inst ( .DIN(_26989), .Q(_26942) );
  hi1s1 _27121_inst ( .DIN(_26989), .Q(_26943) );
  hi1s1 _27122_inst ( .DIN(_26989), .Q(_26944) );
  hi1s1 _27123_inst ( .DIN(_26989), .Q(_26945) );
  hi1s1 _27124_inst ( .DIN(_26989), .Q(_26946) );
  hi1s1 _27125_inst ( .DIN(_26990), .Q(_26947) );
  hi1s1 _27126_inst ( .DIN(_26990), .Q(_26948) );
  hi1s1 _27127_inst ( .DIN(_26990), .Q(_26949) );
  hi1s1 _27128_inst ( .DIN(_26990), .Q(_26950) );
  hi1s1 _27129_inst ( .DIN(_26990), .Q(_26951) );
  hi1s1 _27130_inst ( .DIN(_26990), .Q(_26952) );
  hi1s1 _27131_inst ( .DIN(_26990), .Q(_26953) );
  hi1s1 _27132_inst ( .DIN(_26990), .Q(_26954) );
  hi1s1 _27133_inst ( .DIN(_26990), .Q(_26955) );
  hi1s1 _27134_inst ( .DIN(_26990), .Q(_26956) );
  hi1s1 _27135_inst ( .DIN(_26990), .Q(_26957) );
  hi1s1 _27136_inst ( .DIN(_26989), .Q(_26958) );
  hi1s1 _27137_inst ( .DIN(_26990), .Q(_26959) );
  hi1s1 _27138_inst ( .DIN(_26989), .Q(_26960) );
  hi1s1 _27139_inst ( .DIN(_26990), .Q(_26961) );
  hi1s1 _27140_inst ( .DIN(_26988), .Q(_26962) );
  hi1s1 _27141_inst ( .DIN(_26991), .Q(_26963) );
  hi1s1 _27142_inst ( .DIN(_26987), .Q(_26964) );
  hi1s1 _27143_inst ( .DIN(_26991), .Q(_26965) );
  hi1s1 _27144_inst ( .DIN(_26990), .Q(_26966) );
  hi1s1 _27145_inst ( .DIN(_26989), .Q(_26967) );
  hi1s1 _27146_inst ( .DIN(_26990), .Q(_26968) );
  hi1s1 _27147_inst ( .DIN(_26988), .Q(_26969) );
  hi1s1 _27148_inst ( .DIN(_26987), .Q(_26970) );
  hi1s1 _27149_inst ( .DIN(_26989), .Q(_26971) );
  hi1s1 _27150_inst ( .DIN(_26990), .Q(_26972) );
  hi1s1 _27151_inst ( .DIN(_26991), .Q(_26973) );
  hi1s1 _27152_inst ( .DIN(_26987), .Q(_26974) );
  hi1s1 _27153_inst ( .DIN(_26989), .Q(_26975) );
  hi1s1 _27154_inst ( .DIN(_26988), .Q(_26976) );
  hi1s1 _27155_inst ( .DIN(_26991), .Q(_26977) );
  hi1s1 _27156_inst ( .DIN(_26991), .Q(_26978) );
  hi1s1 _27157_inst ( .DIN(_26991), .Q(_26979) );
  hi1s1 _27158_inst ( .DIN(_26991), .Q(_26980) );
  hi1s1 _27159_inst ( .DIN(_26991), .Q(_26981) );
  hi1s1 _27160_inst ( .DIN(_26991), .Q(_26982) );
  hi1s1 _27161_inst ( .DIN(_26991), .Q(_26983) );
  hi1s1 _27162_inst ( .DIN(_26991), .Q(_26984) );
  hi1s1 _27163_inst ( .DIN(_26991), .Q(_26985) );
  hi1s1 _27164_inst ( .DIN(_26987), .Q(_26986) );
  ib1s1 _27165_inst ( .DIN(___), .Q(_26987) );
  ib1s1 _27166_inst ( .DIN(___), .Q(_26988) );
  ib1s1 _27167_inst ( .DIN(___), .Q(_26989) );
  ib1s1 _27168_inst ( .DIN(___), .Q(_26990) );
  ib1s1 _27169_inst ( .DIN(___), .Q(_26991) );
  nnd2s1 _27170_inst ( .DIN1(_26992), .DIN2(_26993), .Q(
        __________________________________________9_________) );
  nor2s1 _27171_inst ( .DIN1(_26994), .DIN2(_26995), .Q(_26992) );
  nor2s1 _27172_inst ( .DIN1(_26996), .DIN2(_26997), .Q(_26995) );
  xor2s1 _27173_inst ( .DIN1(_26998), .DIN2(_26999), .Q(_26997) );
  nnd2s1 _27174_inst ( .DIN1(_27000), .DIN2(_27001), .Q(_26999) );
  nnd2s1 _27175_inst ( .DIN1(_27002), .DIN2(_27003), .Q(_27001) );
  and2s1 _27176_inst ( .DIN1(_27004), .DIN2(_53199), .Q(_27002) );
  nnd2s1 _27177_inst ( .DIN1(_27005), .DIN2(_27006), .Q(_27000) );
  nor2s1 _27178_inst ( .DIN1(_53259), .DIN2(_27007), .Q(_26994) );
  nnd2s1 _27179_inst ( .DIN1(_27008), .DIN2(_27009), .Q(
        __________________________________________8_________) );
  nnd2s1 _27180_inst ( .DIN1(_27010), .DIN2(_27011), .Q(_27009) );
  nnd2s1 _27181_inst ( .DIN1(_27012), .DIN2(_27013), .Q(_27011) );
  xor2s1 _27182_inst ( .DIN1(_53064), .DIN2(_53311), .Q(_27012) );
  nor2s1 _27183_inst ( .DIN1(_27014), .DIN2(_27015), .Q(_27008) );
  nor2s1 _27184_inst ( .DIN1(_27016), .DIN2(_27017), .Q(_27015) );
  nnd2s1 _27185_inst ( .DIN1(_27018), .DIN2(_27019), .Q(_27017) );
  nor2s1 _27186_inst ( .DIN1(_26772), .DIN2(_27020), .Q(_27014) );
  nnd2s1 _27187_inst ( .DIN1(_27021), .DIN2(_27022), .Q(_27020) );
  xor2s1 _27188_inst ( .DIN1(_53390), .DIN2(_53438), .Q(_27022) );
  nnd2s1 _27189_inst ( .DIN1(_27023), .DIN2(_27024), .Q(
        __________________________________________7_________) );
  nor2s1 _27190_inst ( .DIN1(_27025), .DIN2(_27026), .Q(_27024) );
  nor2s1 _27191_inst ( .DIN1(_27027), .DIN2(_27028), .Q(_27026) );
  nor2s1 _27192_inst ( .DIN1(_27029), .DIN2(_27030), .Q(_27023) );
  nor2s1 _27193_inst ( .DIN1(_53258), .DIN2(_27031), .Q(_27030) );
  nor2s1 _27194_inst ( .DIN1(_27032), .DIN2(_27033), .Q(_27029) );
  nnd2s1 _27195_inst ( .DIN1(_27034), .DIN2(_27035), .Q(
        __________________________________________6_________) );
  nor2s1 _27196_inst ( .DIN1(_27025), .DIN2(_27036), .Q(_27035) );
  nor2s1 _27197_inst ( .DIN1(_27037), .DIN2(_27031), .Q(_27036) );
  nor2s1 _27198_inst ( .DIN1(_27038), .DIN2(_27039), .Q(_27037) );
  xor2s1 _27199_inst ( .DIN1(_26620), .DIN2(_53258), .Q(_27038) );
  nor2s1 _27200_inst ( .DIN1(_27040), .DIN2(_27041), .Q(_27034) );
  nor2s1 _27201_inst ( .DIN1(_27042), .DIN2(_27028), .Q(_27041) );
  nor2s1 _27202_inst ( .DIN1(_27043), .DIN2(_27044), .Q(_27040) );
  nor2s1 _27203_inst ( .DIN1(_27045), .DIN2(_27046), .Q(_27044) );
  nnd2s1 _27204_inst ( .DIN1(______[2]), .DIN2(_27047), .Q(_27046) );
  xor2s1 _27205_inst ( .DIN1(_52857), .DIN2(_27048), .Q(_27045) );
  nnd2s1 _27206_inst ( .DIN1(_27049), .DIN2(_27050), .Q(
        __________________________________________5_________) );
  nor2s1 _27207_inst ( .DIN1(_27051), .DIN2(_27052), .Q(_27049) );
  nor2s1 _27208_inst ( .DIN1(_27053), .DIN2(_27054), .Q(_27052) );
  nnd2s1 _27209_inst ( .DIN1(_27055), .DIN2(_27056), .Q(_27054) );
  nnd2s1 _27210_inst ( .DIN1(_27057), .DIN2(_27058), .Q(_27056) );
  nnd2s1 _27211_inst ( .DIN1(_27059), .DIN2(_27060), .Q(_27055) );
  xnr2s1 _27212_inst ( .DIN1(_27061), .DIN2(_27062), .Q(_27060) );
  xor2s1 _27213_inst ( .DIN1(_52837), .DIN2(_52866), .Q(_27062) );
  nor2s1 _27214_inst ( .DIN1(_26772), .DIN2(_27063), .Q(_27059) );
  nor2s1 _27215_inst ( .DIN1(_27064), .DIN2(_27065), .Q(_27051) );
  nor2s1 _27216_inst ( .DIN1(_26854), .DIN2(_26299), .Q(_27065) );
  nnd2s1 _27217_inst ( .DIN1(_27067), .DIN2(_27068), .Q(
        __________________________________________4_________) );
  nnd2s1 _27218_inst ( .DIN1(_27010), .DIN2(_27069), .Q(_27068) );
  nnd2s1 _27219_inst ( .DIN1(_27070), .DIN2(______[12]), .Q(_27069) );
  nor2s1 _27220_inst ( .DIN1(_27071), .DIN2(_27072), .Q(_27070) );
  nor2s1 _27221_inst ( .DIN1(_26308), .DIN2(_27073), .Q(_27072) );
  nnd2s1 _27222_inst ( .DIN1(_53064), .DIN2(_26572), .Q(_27073) );
  nor2s1 _27223_inst ( .DIN1(_53389), .DIN2(_26572), .Q(_27071) );
  nor2s1 _27224_inst ( .DIN1(_27074), .DIN2(_27075), .Q(_27010) );
  nor2s1 _27225_inst ( .DIN1(_27076), .DIN2(_27077), .Q(_27067) );
  nor2s1 _27226_inst ( .DIN1(_27078), .DIN2(_27074), .Q(_27077) );
  nor2s1 _27227_inst ( .DIN1(_27079), .DIN2(_27080), .Q(_27078) );
  and2s1 _27228_inst ( .DIN1(_27081), .DIN2(_27075), .Q(_27079) );
  nor2s1 _27229_inst ( .DIN1(_27082), .DIN2(_27083), .Q(_27076) );
  nnd2s1 _27230_inst ( .DIN1(_27021), .DIN2(_27084), .Q(_27083) );
  xnr2s1 _27231_inst ( .DIN1(_27085), .DIN2(_27086), .Q(_27084) );
  xor2s1 _27232_inst ( .DIN1(_52840), .DIN2(_52892), .Q(_27086) );
  nnd2s1 _27233_inst ( .DIN1(_27087), .DIN2(_27088), .Q(
        __________________________________________3_________) );
  nnd2s1 _27234_inst ( .DIN1(_27089), .DIN2(_27090), .Q(_27088) );
  xor2s1 _27235_inst ( .DIN1(_27091), .DIN2(_52856), .Q(_27089) );
  nnd2s1 _27236_inst ( .DIN1(_27043), .DIN2(_27092), .Q(_27087) );
  xor2s1 _27237_inst ( .DIN1(_27093), .DIN2(_27094), .Q(_27092) );
  nor2s1 _27238_inst ( .DIN1(_27095), .DIN2(_27096), .Q(_27094) );
  nnd2s1 _27239_inst ( .DIN1(_27097), .DIN2(_27098), .Q(_27096) );
  nnd2s1 _27240_inst ( .DIN1(_27058), .DIN2(_27099), .Q(_27098) );
  nnd2s1 _27241_inst ( .DIN1(_27100), .DIN2(_27101), .Q(_27097) );
  nnd2s1 _27242_inst ( .DIN1(_52838), .DIN2(_26861), .Q(_27100) );
  nnd2s1 _27243_inst ( .DIN1(_27102), .DIN2(_27103), .Q(
        __________________________________________2_________) );
  nnd2s1 _27244_inst ( .DIN1(_27104), .DIN2(_26715), .Q(_27103) );
  nnd2s1 _27245_inst ( .DIN1(_27105), .DIN2(_27106), .Q(_27104) );
  nnd2s1 _27246_inst ( .DIN1(_27107), .DIN2(______[4]), .Q(_27106) );
  nor2s1 _27247_inst ( .DIN1(_27095), .DIN2(_27058), .Q(_27107) );
  hi1s1 _27248_inst ( .DIN(_27108), .Q(_27095) );
  nor2s1 _27249_inst ( .DIN1(_27109), .DIN2(_27110), .Q(_27102) );
  nor2s1 _27250_inst ( .DIN1(_27111), .DIN2(_27112), .Q(_27110) );
  nnd2s1 _27251_inst ( .DIN1(_27105), .DIN2(_27058), .Q(_27112) );
  hi1s1 _27252_inst ( .DIN(_27113), .Q(_27109) );
  nnd2s1 _27253_inst ( .DIN1(_27114), .DIN2(_27115), .Q(
        __________________________________________25_________) );
  nnd2s1 _27254_inst ( .DIN1(_27116), .DIN2(_27117), .Q(_27115) );
  nnd2s1 _27255_inst ( .DIN1(_27118), .DIN2(_27119), .Q(_27117) );
  nnd2s1 _27256_inst ( .DIN1(_27120), .DIN2(_26508), .Q(_27119) );
  nnd2s1 _27257_inst ( .DIN1(_27121), .DIN2(_27122), .Q(_27114) );
  nor2s1 _27258_inst ( .DIN1(_27123), .DIN2(_27124), .Q(_27121) );
  xor2s1 _27259_inst ( .DIN1(_26270), .DIN2(_53022), .Q(_27124) );
  nnd2s1 _27260_inst ( .DIN1(_27125), .DIN2(_27126), .Q(
        __________________________________________25________5____________) );
  nor2s1 _27261_inst ( .DIN1(_27127), .DIN2(_27128), .Q(_27125) );
  nor2s1 _27262_inst ( .DIN1(_27129), .DIN2(_27130), .Q(_27128) );
  xor2s1 _27263_inst ( .DIN1(_52946), .DIN2(_53000), .Q(_27130) );
  nor2s1 _27264_inst ( .DIN1(_27131), .DIN2(_27132), .Q(_27127) );
  nor2s1 _27265_inst ( .DIN1(_27133), .DIN2(_27134), .Q(_27131) );
  nor2s1 _27266_inst ( .DIN1(_27135), .DIN2(_27136), .Q(_27133) );
  xnr2s1 _27267_inst ( .DIN1(_27137), .DIN2(_27138), .Q(_27136) );
  xor2s1 _27268_inst ( .DIN1(_26491), .DIN2(_52842), .Q(_27137) );
  nnd2s1 _27269_inst ( .DIN1(_27139), .DIN2(_27140), .Q(
        __________________________________________25________4____________) );
  nor2s1 _27270_inst ( .DIN1(_27141), .DIN2(_27142), .Q(_27140) );
  nor2s1 _27271_inst ( .DIN1(_27143), .DIN2(_27144), .Q(_27142) );
  nor2s1 _27272_inst ( .DIN1(_27145), .DIN2(_27134), .Q(_27143) );
  nor2s1 _27273_inst ( .DIN1(_52979), .DIN2(_27135), .Q(_27145) );
  nor2s1 _27274_inst ( .DIN1(_27146), .DIN2(_27147), .Q(_27141) );
  nnd2s1 _27275_inst ( .DIN1(_52842), .DIN2(_26549), .Q(_27147) );
  nor2s1 _27276_inst ( .DIN1(_27148), .DIN2(_27149), .Q(_27139) );
  nor2s1 _27277_inst ( .DIN1(_52842), .DIN2(_27150), .Q(_27148) );
  nnd2s1 _27278_inst ( .DIN1(_27151), .DIN2(_27152), .Q(
        __________________________________________25________3____________) );
  nnd2s1 _27279_inst ( .DIN1(_27153), .DIN2(_27154), .Q(_27152) );
  nor2s1 _27280_inst ( .DIN1(_27155), .DIN2(_27156), .Q(_27153) );
  nor2s1 _27281_inst ( .DIN1(_27157), .DIN2(_27158), .Q(_27156) );
  nor2s1 _27282_inst ( .DIN1(_27135), .DIN2(_27159), .Q(_27155) );
  nor2s1 _27283_inst ( .DIN1(_52842), .DIN2(_27160), .Q(_27159) );
  nnd2s1 _27284_inst ( .DIN1(_53394), .DIN2(_27161), .Q(_27151) );
  nnd2s1 _27285_inst ( .DIN1(_27162), .DIN2(_27163), .Q(
        __________________________________________25________2____________) );
  nnd2s1 _27286_inst ( .DIN1(_27164), .DIN2(_27165), .Q(_27163) );
  nnd2s1 _27287_inst ( .DIN1(_27166), .DIN2(_27167), .Q(_27165) );
  nnd2s1 _27288_inst ( .DIN1(_27168), .DIN2(_27158), .Q(_27167) );
  nnd2s1 _27289_inst ( .DIN1(_27169), .DIN2(______[6]), .Q(_27168) );
  nor2s1 _27290_inst ( .DIN1(_27170), .DIN2(_27171), .Q(_27169) );
  nor2s1 _27291_inst ( .DIN1(_26491), .DIN2(_27138), .Q(_27171) );
  or2s1 _27292_inst ( .DIN1(_26564), .DIN2(_52842), .Q(_27138) );
  nor2s1 _27293_inst ( .DIN1(_53393), .DIN2(_27172), .Q(_27170) );
  nor2s1 _27294_inst ( .DIN1(_52842), .DIN2(_26491), .Q(_27172) );
  hi1s1 _27295_inst ( .DIN(_27134), .Q(_27166) );
  nnd2s1 _27296_inst ( .DIN1(_27173), .DIN2(_27174), .Q(_27134) );
  nnd2s1 _27297_inst ( .DIN1(_27160), .DIN2(_27158), .Q(_27174) );
  nnd2s1 _27298_inst ( .DIN1(_27135), .DIN2(_27175), .Q(_27173) );
  nnd2s1 _27299_inst ( .DIN1(_27176), .DIN2(_27177), .Q(_27162) );
  xor2s1 _27300_inst ( .DIN1(_53080), .DIN2(_53084), .Q(_27176) );
  nnd2s1 _27301_inst ( .DIN1(_27178), .DIN2(_27179), .Q(
        __________________________________________25________1____________) );
  nnd2s1 _27302_inst ( .DIN1(_27180), .DIN2(______[0]), .Q(_27179) );
  nor2s1 _27303_inst ( .DIN1(_27181), .DIN2(_27182), .Q(_27180) );
  xor2s1 _27304_inst ( .DIN1(_26569), .DIN2(_53273), .Q(_27181) );
  nnd2s1 _27305_inst ( .DIN1(_27183), .DIN2(_27184), .Q(_27178) );
  nnd2s1 _27306_inst ( .DIN1(_27118), .DIN2(_27185), .Q(_27184) );
  nnd2s1 _27307_inst ( .DIN1(_27186), .DIN2(_27120), .Q(_27185) );
  xor2s1 _27308_inst ( .DIN1(_27187), .DIN2(_27188), .Q(_27186) );
  xor2s1 _27309_inst ( .DIN1(_53237), .DIN2(_53390), .Q(_27188) );
  nor2s1 _27310_inst ( .DIN1(_52888), .DIN2(_26377), .Q(_27187) );
  nnd2s1 _27311_inst ( .DIN1(_27189), .DIN2(_26796), .Q(_27118) );
  nnd2s1 _27312_inst ( .DIN1(_27190), .DIN2(_27191), .Q(
        __________________________________________25________0____________) );
  nnd2s1 _27313_inst ( .DIN1(_27192), .DIN2(_27018), .Q(_27191) );
  nor2s1 _27314_inst ( .DIN1(_27193), .DIN2(_27194), .Q(_27192) );
  nor2s1 _27315_inst ( .DIN1(_27175), .DIN2(_27195), .Q(_27194) );
  nor2s1 _27316_inst ( .DIN1(_26377), .DIN2(_27196), .Q(_27193) );
  nnd2s1 _27317_inst ( .DIN1(______[6]), .DIN2(_27120), .Q(_27196) );
  nnd2s1 _27318_inst ( .DIN1(_27021), .DIN2(_53438), .Q(_27190) );
  nnd2s1 _27319_inst ( .DIN1(_27197), .DIN2(_27198), .Q(
        __________________________________________24_________) );
  nor2s1 _27320_inst ( .DIN1(_27199), .DIN2(_27200), .Q(_27197) );
  nor2s1 _27321_inst ( .DIN1(_27201), .DIN2(_27202), .Q(_27200) );
  and2s1 _27322_inst ( .DIN1(______[26]), .DIN2(_53310), .Q(_27202) );
  nor2s1 _27323_inst ( .DIN1(_27203), .DIN2(_27204), .Q(_27199) );
  nor2s1 _27324_inst ( .DIN1(_27080), .DIN2(_27205), .Q(_27203) );
  nnd2s1 _27325_inst ( .DIN1(_27206), .DIN2(_27207), .Q(_27205) );
  nnd2s1 _27326_inst ( .DIN1(_27208), .DIN2(_27016), .Q(_27207) );
  nor2s1 _27327_inst ( .DIN1(_26654), .DIN2(_26308), .Q(_27208) );
  or2s1 _27328_inst ( .DIN1(_27209), .DIN2(_27016), .Q(_27206) );
  and2s1 _27329_inst ( .DIN1(_27210), .DIN2(_27016), .Q(_27080) );
  nnd2s1 _27330_inst ( .DIN1(_27013), .DIN2(_27211), .Q(_27210) );
  nnd2s1 _27331_inst ( .DIN1(_26308), .DIN2(_26654), .Q(_27211) );
  nnd2s1 _27332_inst ( .DIN1(_27212), .DIN2(_27213), .Q(
        __________________________________________23_________) );
  nnd2s1 _27333_inst ( .DIN1(_27214), .DIN2(_27074), .Q(_27213) );
  nnd2s1 _27334_inst ( .DIN1(_52858), .DIN2(_27215), .Q(_27214) );
  nnd2s1 _27335_inst ( .DIN1(_27216), .DIN2(_27018), .Q(_27212) );
  nor2s1 _27336_inst ( .DIN1(_27217), .DIN2(_27218), .Q(_27216) );
  nor2s1 _27337_inst ( .DIN1(_27219), .DIN2(_27220), .Q(_27218) );
  xor2s1 _27338_inst ( .DIN1(_26306), .DIN2(_27221), .Q(_27220) );
  nor2s1 _27339_inst ( .DIN1(_27222), .DIN2(_27223), .Q(_27217) );
  nnd2s1 _27340_inst ( .DIN1(_27224), .DIN2(_27225), .Q(
        __________________________________________22_________) );
  nnd2s1 _27341_inst ( .DIN1(_27226), .DIN2(_27227), .Q(_27225) );
  nor2s1 _27342_inst ( .DIN1(_27228), .DIN2(_27229), .Q(_27226) );
  nor2s1 _27343_inst ( .DIN1(_27230), .DIN2(_27231), .Q(_27229) );
  xor2s1 _27344_inst ( .DIN1(_52888), .DIN2(_26508), .Q(_27231) );
  nor2s1 _27345_inst ( .DIN1(_27195), .DIN2(_27232), .Q(_27228) );
  nnd2s1 _27346_inst ( .DIN1(_53075), .DIN2(_27233), .Q(_27224) );
  nor2s1 _27347_inst ( .DIN1(_27234), .DIN2(_27235), .Q(
        __________________________________________21_________) );
  nor2s1 _27348_inst ( .DIN1(_27236), .DIN2(_27237), .Q(_27234) );
  nor2s1 _27349_inst ( .DIN1(_27222), .DIN2(_27238), .Q(_27237) );
  nor2s1 _27350_inst ( .DIN1(_27239), .DIN2(_27219), .Q(_27236) );
  or2s1 _27351_inst ( .DIN1(_27240), .DIN2(_26855), .Q(_27219) );
  xor2s1 _27352_inst ( .DIN1(_26494), .DIN2(_27242), .Q(_27239) );
  nnd2s1 _27353_inst ( .DIN1(_27243), .DIN2(_27244), .Q(
        __________________________________________20_________) );
  nnd2s1 _27354_inst ( .DIN1(_27245), .DIN2(_52898), .Q(_27244) );
  and2s1 _27355_inst ( .DIN1(______[2]), .DIN2(_27246), .Q(_27245) );
  nnd2s1 _27356_inst ( .DIN1(_27247), .DIN2(_27248), .Q(_27243) );
  nnd2s1 _27357_inst ( .DIN1(_27249), .DIN2(_27250), .Q(_27248) );
  nnd2s1 _27358_inst ( .DIN1(_27251), .DIN2(_27120), .Q(_27250) );
  xor2s1 _27359_inst ( .DIN1(_27252), .DIN2(_27253), .Q(_27251) );
  xor2s1 _27360_inst ( .DIN1(_52909), .DIN2(_53046), .Q(_27253) );
  nnd2s1 _27361_inst ( .DIN1(_52899), .DIN2(_53183), .Q(_27252) );
  nnd2s1 _27362_inst ( .DIN1(_27254), .DIN2(_27189), .Q(_27249) );
  nnd2s1 _27363_inst ( .DIN1(_27255), .DIN2(_27256), .Q(
        __________________________________________1_________) );
  nor2s1 _27364_inst ( .DIN1(_27257), .DIN2(_27258), .Q(_27255) );
  nor2s1 _27365_inst ( .DIN1(_27122), .DIN2(_27259), .Q(_27258) );
  nnd2s1 _27366_inst ( .DIN1(_27260), .DIN2(_27261), .Q(_27259) );
  or2s1 _27367_inst ( .DIN1(_27262), .DIN2(_27101), .Q(_27261) );
  nnd2s1 _27368_inst ( .DIN1(_27263), .DIN2(_27264), .Q(_27260) );
  nor2s1 _27369_inst ( .DIN1(_27048), .DIN2(_27063), .Q(_27264) );
  nor2s1 _27370_inst ( .DIN1(_27082), .DIN2(_27265), .Q(_27263) );
  nnd2s1 _27371_inst ( .DIN1(_27266), .DIN2(_27267), .Q(_27265) );
  nnd2s1 _27372_inst ( .DIN1(_52872), .DIN2(_26753), .Q(_27267) );
  nnd2s1 _27373_inst ( .DIN1(_27061), .DIN2(_52837), .Q(_27266) );
  nor2s1 _27374_inst ( .DIN1(_27116), .DIN2(_27268), .Q(_27257) );
  xor2s1 _27375_inst ( .DIN1(_27269), .DIN2(_52888), .Q(_27268) );
  nnd2s1 _27376_inst ( .DIN1(_53055), .DIN2(_53022), .Q(_27269) );
  nnd2s1 _27377_inst ( .DIN1(_27270), .DIN2(_27271), .Q(
        __________________________________________19_________) );
  nnd2s1 _27378_inst ( .DIN1(_27018), .DIN2(_27272), .Q(_27271) );
  nnd2s1 _27379_inst ( .DIN1(_27273), .DIN2(_27274), .Q(_27272) );
  nor2s1 _27380_inst ( .DIN1(_27275), .DIN2(_27276), .Q(_27273) );
  nor2s1 _27381_inst ( .DIN1(_27222), .DIN2(_27277), .Q(_27276) );
  nor2s1 _27382_inst ( .DIN1(_53385), .DIN2(_27278), .Q(_27275) );
  nnd2s1 _27383_inst ( .DIN1(_52892), .DIN2(_27021), .Q(_27270) );
  nor2s1 _27384_inst ( .DIN1(_27279), .DIN2(_27018), .Q(_27021) );
  nnd2s1 _27385_inst ( .DIN1(_27280), .DIN2(_27281), .Q(
        __________________________________________18_________) );
  nor2s1 _27386_inst ( .DIN1(_27282), .DIN2(_27283), .Q(_27280) );
  nor2s1 _27387_inst ( .DIN1(_27284), .DIN2(_27285), .Q(_27283) );
  nnd2s1 _27388_inst ( .DIN1(_27286), .DIN2(_27287), .Q(_27285) );
  nnd2s1 _27389_inst ( .DIN1(_27288), .DIN2(_27289), .Q(_27287) );
  nor2s1 _27390_inst ( .DIN1(_27242), .DIN2(_27290), .Q(_27289) );
  nor2s1 _27391_inst ( .DIN1(_53385), .DIN2(_26544), .Q(_27290) );
  hi1s1 _27392_inst ( .DIN(_27221), .Q(_27242) );
  nnd2s1 _27393_inst ( .DIN1(_53385), .DIN2(_26544), .Q(_27221) );
  nor2s1 _27394_inst ( .DIN1(_27240), .DIN2(_27291), .Q(_27288) );
  nnd2s1 _27395_inst ( .DIN1(_27222), .DIN2(_27292), .Q(_27240) );
  nnd2s1 _27396_inst ( .DIN1(_27293), .DIN2(_27294), .Q(_27292) );
  nor2s1 _27397_inst ( .DIN1(_27295), .DIN2(_27296), .Q(_27294) );
  nnd2s1 _27398_inst ( .DIN1(_27278), .DIN2(_27297), .Q(_27286) );
  nor2s1 _27399_inst ( .DIN1(_27298), .DIN2(_26660), .Q(_27282) );
  nnd2s1 _27400_inst ( .DIN1(_27299), .DIN2(_27300), .Q(
        __________________________________________17_________) );
  nnd2s1 _27401_inst ( .DIN1(_27301), .DIN2(_27074), .Q(_27300) );
  nnd2s1 _27402_inst ( .DIN1(_27302), .DIN2(_27303), .Q(_27301) );
  nor2s1 _27403_inst ( .DIN1(_27279), .DIN2(_27304), .Q(_27303) );
  nor2s1 _27404_inst ( .DIN1(_52895), .DIN2(_27305), .Q(_27304) );
  nor2s1 _27405_inst ( .DIN1(_26494), .DIN2(_26264), .Q(_27305) );
  hi1s1 _27406_inst ( .DIN(_27215), .Q(_27279) );
  nnd2s1 _27407_inst ( .DIN1(_27306), .DIN2(_27307), .Q(_27215) );
  nor2s1 _27408_inst ( .DIN1(_27308), .DIN2(_27309), .Q(_27307) );
  nor2s1 _27409_inst ( .DIN1(_27310), .DIN2(_27311), .Q(_27306) );
  nor2s1 _27410_inst ( .DIN1(_27312), .DIN2(_26987), .Q(_27302) );
  nor2s1 _27411_inst ( .DIN1(_26264), .DIN2(_27085), .Q(_27312) );
  nnd2s1 _27412_inst ( .DIN1(_52892), .DIN2(_52895), .Q(_27085) );
  nnd2s1 _27413_inst ( .DIN1(_27313), .DIN2(_27018), .Q(_27299) );
  hi1s1 _27414_inst ( .DIN(_27074), .Q(_27018) );
  nnd2s1 _27415_inst ( .DIN1(_27314), .DIN2(_27315), .Q(_27074) );
  nor2s1 _27416_inst ( .DIN1(_27308), .DIN2(_27316), .Q(_27315) );
  nor2s1 _27417_inst ( .DIN1(_27317), .DIN2(_27318), .Q(_27314) );
  nor2s1 _27418_inst ( .DIN1(_27319), .DIN2(_27320), .Q(_27313) );
  nnd2s1 _27419_inst ( .DIN1(_27321), .DIN2(_27322), .Q(_27320) );
  nnd2s1 _27420_inst ( .DIN1(_27278), .DIN2(_27323), .Q(_27322) );
  nnd2s1 _27421_inst ( .DIN1(_27032), .DIN2(_27222), .Q(_27321) );
  xnr2s1 _27422_inst ( .DIN1(_52839), .DIN2(_52929), .Q(_27032) );
  hi1s1 _27423_inst ( .DIN(_27274), .Q(_27319) );
  nnd2s1 _27424_inst ( .DIN1(_27324), .DIN2(_27325), .Q(
        __________________________________________16_________) );
  nor2s1 _27425_inst ( .DIN1(_27326), .DIN2(_27327), .Q(_27324) );
  nor2s1 _27426_inst ( .DIN1(_27328), .DIN2(_27329), .Q(_27327) );
  nor2s1 _27427_inst ( .DIN1(_27330), .DIN2(_27331), .Q(_27328) );
  nor2s1 _27428_inst ( .DIN1(_27230), .DIN2(_26502), .Q(_27331) );
  hi1s1 _27429_inst ( .DIN(_27120), .Q(_27230) );
  nnd2s1 _27430_inst ( .DIN1(_27332), .DIN2(_27333), .Q(_27120) );
  nor2s1 _27431_inst ( .DIN1(_27295), .DIN2(_27334), .Q(_27333) );
  nnd2s1 _27432_inst ( .DIN1(_27335), .DIN2(_27336), .Q(_27334) );
  nor2s1 _27433_inst ( .DIN1(_27337), .DIN2(_27195), .Q(_27330) );
  nor2s1 _27434_inst ( .DIN1(_27338), .DIN2(_27339), .Q(_27326) );
  nnd2s1 _27435_inst ( .DIN1(_27189), .DIN2(_27337), .Q(_27339) );
  hi1s1 _27436_inst ( .DIN(_27195), .Q(_27189) );
  nnd2s1 _27437_inst ( .DIN1(_27340), .DIN2(_27341), .Q(_27195) );
  nor2s1 _27438_inst ( .DIN1(_27342), .DIN2(_27343), .Q(_27341) );
  nor2s1 _27439_inst ( .DIN1(_27344), .DIN2(_27345), .Q(_27340) );
  xor2s1 _27440_inst ( .DIN1(_27346), .DIN2(_27347), .Q(_27345) );
  nnd2s1 _27441_inst ( .DIN1(_27348), .DIN2(_27349), .Q(_27347) );
  nnd2s1 _27442_inst ( .DIN1(_27350), .DIN2(_27351), .Q(
        __________________________________________15_________) );
  nnd2s1 _27443_inst ( .DIN1(_27352), .DIN2(_27090), .Q(_27351) );
  xor2s1 _27444_inst ( .DIN1(_27353), .DIN2(_52854), .Q(_27352) );
  nnd2s1 _27445_inst ( .DIN1(_52929), .DIN2(_52839), .Q(_27353) );
  nnd2s1 _27446_inst ( .DIN1(_27043), .DIN2(_27354), .Q(_27350) );
  nnd2s1 _27447_inst ( .DIN1(_27355), .DIN2(_27274), .Q(_27354) );
  nnd2s1 _27448_inst ( .DIN1(_27293), .DIN2(_27356), .Q(_27274) );
  nor2s1 _27449_inst ( .DIN1(_27278), .DIN2(_27357), .Q(_27356) );
  nnd2s1 _27450_inst ( .DIN1(_27358), .DIN2(_27359), .Q(_27357) );
  nor2s1 _27451_inst ( .DIN1(_27360), .DIN2(_27361), .Q(_27293) );
  nor2s1 _27452_inst ( .DIN1(_27362), .DIN2(_27363), .Q(_27355) );
  nor2s1 _27453_inst ( .DIN1(_27278), .DIN2(_27364), .Q(_27363) );
  nor2s1 _27454_inst ( .DIN1(_26809), .DIN2(_27366), .Q(_27364) );
  xor2s1 _27455_inst ( .DIN1(_52840), .DIN2(_27367), .Q(_27366) );
  nor2s1 _27456_inst ( .DIN1(_52929), .DIN2(_52919), .Q(_27367) );
  and2s1 _27457_inst ( .DIN1(_27368), .DIN2(_27278), .Q(_27362) );
  hi1s1 _27458_inst ( .DIN(_27222), .Q(_27278) );
  nnd2s1 _27459_inst ( .DIN1(_27369), .DIN2(_27370), .Q(_27222) );
  nor2s1 _27460_inst ( .DIN1(_27371), .DIN2(_27372), .Q(_27370) );
  nnd2s1 _27461_inst ( .DIN1(_27358), .DIN2(_27373), .Q(_27372) );
  nor2s1 _27462_inst ( .DIN1(_27374), .DIN2(_27375), .Q(_27371) );
  nor2s1 _27463_inst ( .DIN1(_27376), .DIN2(_27377), .Q(_27369) );
  nnd2s1 _27464_inst ( .DIN1(_27378), .DIN2(_27379), .Q(
        __________________________________________14_________) );
  nnd2s1 _27465_inst ( .DIN1(_27380), .DIN2(_27381), .Q(_27379) );
  hi1s1 _27466_inst ( .DIN(_27028), .Q(_27381) );
  nor2s1 _27467_inst ( .DIN1(_27382), .DIN2(_27383), .Q(_27378) );
  nor2s1 _27468_inst ( .DIN1(_27043), .DIN2(_27384), .Q(_27383) );
  nor2s1 _27469_inst ( .DIN1(_27291), .DIN2(_27385), .Q(_27384) );
  nnd2s1 _27470_inst ( .DIN1(_27386), .DIN2(_27047), .Q(_27385) );
  xor2s1 _27471_inst ( .DIN1(_52839), .DIN2(_52919), .Q(_27386) );
  nor2s1 _27472_inst ( .DIN1(_27387), .DIN2(_27388), .Q(_27382) );
  or2s1 _27473_inst ( .DIN1(_27031), .DIN2(_26772), .Q(_27388) );
  nnd2s1 _27474_inst ( .DIN1(_27004), .DIN2(_26693), .Q(_27387) );
  nnd2s1 _27475_inst ( .DIN1(_27389), .DIN2(_27390), .Q(
        __________________________________________13_________) );
  nnd2s1 _27476_inst ( .DIN1(_27391), .DIN2(_27392), .Q(_27390) );
  nor2s1 _27477_inst ( .DIN1(_27393), .DIN2(_27394), .Q(_27391) );
  nnd2s1 _27478_inst ( .DIN1(_27395), .DIN2(_27396), .Q(_27394) );
  xor2s1 _27479_inst ( .DIN1(_53182), .DIN2(_53185), .Q(_27395) );
  nnd2s1 _27480_inst ( .DIN1(_27397), .DIN2(_27398), .Q(_27389) );
  nnd2s1 _27481_inst ( .DIN1(_27399), .DIN2(_27400), .Q(_27398) );
  nnd2s1 _27482_inst ( .DIN1(_27401), .DIN2(_27016), .Q(_27400) );
  nor2s1 _27483_inst ( .DIN1(_26774), .DIN2(_27402), .Q(_27401) );
  nnd2s1 _27484_inst ( .DIN1(_52909), .DIN2(_27013), .Q(_27402) );
  nnd2s1 _27485_inst ( .DIN1(_27403), .DIN2(_27075), .Q(_27399) );
  nnd2s1 _27486_inst ( .DIN1(_27404), .DIN2(_27405), .Q(
        __________________________________________12_________) );
  nor2s1 _27487_inst ( .DIN1(_27406), .DIN2(_27407), .Q(_27404) );
  nor2s1 _27488_inst ( .DIN1(_27408), .DIN2(_27409), .Q(_27407) );
  nnd2s1 _27489_inst ( .DIN1(_27410), .DIN2(_27411), .Q(_27409) );
  nnd2s1 _27490_inst ( .DIN1(_27412), .DIN2(_27016), .Q(_27411) );
  xor2s1 _27491_inst ( .DIN1(_27413), .DIN2(_27414), .Q(_27410) );
  nor2s1 _27492_inst ( .DIN1(_27415), .DIN2(_27416), .Q(_27414) );
  xor2s1 _27493_inst ( .DIN1(_27417), .DIN2(_27418), .Q(_27416) );
  nnd2s1 _27494_inst ( .DIN1(_27419), .DIN2(_27016), .Q(_27417) );
  xor2s1 _27495_inst ( .DIN1(_26599), .DIN2(_53183), .Q(_27419) );
  nor2s1 _27496_inst ( .DIN1(_27016), .DIN2(_27420), .Q(_27415) );
  nor2s1 _27497_inst ( .DIN1(_27421), .DIN2(_27422), .Q(_27406) );
  xor2s1 _27498_inst ( .DIN1(_52841), .DIN2(_53045), .Q(_27422) );
  nnd2s1 _27499_inst ( .DIN1(_27423), .DIN2(_27424), .Q(
        __________________________________________11_________) );
  nor2s1 _27500_inst ( .DIN1(_27025), .DIN2(_27425), .Q(_27424) );
  nor2s1 _27501_inst ( .DIN1(_27291), .DIN2(_27426), .Q(_27425) );
  nnd2s1 _27502_inst ( .DIN1(_27090), .DIN2(_52929), .Q(_27426) );
  hi1s1 _27503_inst ( .DIN(_27033), .Q(_27090) );
  nnd2s1 _27504_inst ( .DIN1(_27047), .DIN2(_27427), .Q(_27033) );
  nnd2s1 _27505_inst ( .DIN1(_27428), .DIN2(_27429), .Q(_27047) );
  nor2s1 _27506_inst ( .DIN1(_27430), .DIN2(_27431), .Q(_27429) );
  nor2s1 _27507_inst ( .DIN1(_27432), .DIN2(_27433), .Q(_27428) );
  nor2s1 _27508_inst ( .DIN1(_27031), .DIN2(_27004), .Q(_27025) );
  nor2s1 _27509_inst ( .DIN1(_27434), .DIN2(_27435), .Q(_27423) );
  nor2s1 _27510_inst ( .DIN1(_27436), .DIN2(_27028), .Q(_27435) );
  nnd2s1 _27511_inst ( .DIN1(_27043), .DIN2(_27005), .Q(_27028) );
  nor2s1 _27512_inst ( .DIN1(_27437), .DIN2(_27031), .Q(_27434) );
  nnd2s1 _27513_inst ( .DIN1(_27043), .DIN2(_27003), .Q(_27031) );
  hi1s1 _27514_inst ( .DIN(_27427), .Q(_27043) );
  nnd2s1 _27515_inst ( .DIN1(_27438), .DIN2(_27439), .Q(_27427) );
  nor2s1 _27516_inst ( .DIN1(_27309), .DIN2(_27440), .Q(_27439) );
  nnd2s1 _27517_inst ( .DIN1(_27441), .DIN2(_27442), .Q(_27440) );
  nor2s1 _27518_inst ( .DIN1(_27443), .DIN2(_27444), .Q(_27438) );
  nnd2s1 _27519_inst ( .DIN1(_27445), .DIN2(_27446), .Q(_27444) );
  nor2s1 _27520_inst ( .DIN1(_27447), .DIN2(_27448), .Q(_27437) );
  xor2s1 _27521_inst ( .DIN1(_52929), .DIN2(_26264), .Q(_27447) );
  nnd2s1 _27522_inst ( .DIN1(_27449), .DIN2(_27450), .Q(
        __________________________________________10_________) );
  nor2s1 _27523_inst ( .DIN1(_27451), .DIN2(_27452), .Q(_27449) );
  nor2s1 _27524_inst ( .DIN1(_27453), .DIN2(_27454), .Q(_27452) );
  nor2s1 _27525_inst ( .DIN1(_27455), .DIN2(_27456), .Q(_27454) );
  nor2s1 _27526_inst ( .DIN1(_27003), .DIN2(_27457), .Q(_27456) );
  nor2s1 _27527_inst ( .DIN1(_27005), .DIN2(_27458), .Q(_27455) );
  nnd2s1 _27528_inst ( .DIN1(_27459), .DIN2(_27004), .Q(_27458) );
  xor2s1 _27529_inst ( .DIN1(_27460), .DIN2(_27461), .Q(_27459) );
  xor2s1 _27530_inst ( .DIN1(_52856), .DIN2(_53258), .Q(_27461) );
  nnd2s1 _27531_inst ( .DIN1(_52854), .DIN2(_53199), .Q(_27460) );
  hi1s1 _27532_inst ( .DIN(_27003), .Q(_27005) );
  nnd2s1 _27533_inst ( .DIN1(_27462), .DIN2(_27463), .Q(_27003) );
  nor2s1 _27534_inst ( .DIN1(_27464), .DIN2(_27465), .Q(_27463) );
  nnd2s1 _27535_inst ( .DIN1(_27359), .DIN2(_27373), .Q(_27465) );
  nnd2s1 _27536_inst ( .DIN1(_27466), .DIN2(_27467), .Q(_27464) );
  nor2s1 _27537_inst ( .DIN1(_27468), .DIN2(_27469), .Q(_27462) );
  nnd2s1 _27538_inst ( .DIN1(_27470), .DIN2(_27471), .Q(_27469) );
  nnd2s1 _27539_inst ( .DIN1(_27472), .DIN2(_27473), .Q(_27468) );
  or2s1 _27540_inst ( .DIN1(_27474), .DIN2(_27475), .Q(_27472) );
  nor2s1 _27541_inst ( .DIN1(_27476), .DIN2(_27477), .Q(_27451) );
  nor2s1 _27542_inst ( .DIN1(_26853), .DIN2(_27478), .Q(_27477) );
  nnd2s1 _27543_inst ( .DIN1(_27479), .DIN2(_27480), .Q(_27478) );
  nnd2s1 _27544_inst ( .DIN1(_53439), .DIN2(_26386), .Q(_27479) );
  nnd2s1 _27545_inst ( .DIN1(_27481), .DIN2(_27482), .Q(
        __________________________________________0_________) );
  nnd2s1 _27546_inst ( .DIN1(_27483), .DIN2(_27421), .Q(_27482) );
  nor2s1 _27547_inst ( .DIN1(_27484), .DIN2(_27485), .Q(_27483) );
  nor2s1 _27548_inst ( .DIN1(_27016), .DIN2(_27486), .Q(_27485) );
  nor2s1 _27549_inst ( .DIN1(_27075), .DIN2(_27487), .Q(_27484) );
  nor2s1 _27550_inst ( .DIN1(_52858), .DIN2(_27412), .Q(_27487) );
  hi1s1 _27551_inst ( .DIN(_27016), .Q(_27075) );
  nnd2s1 _27552_inst ( .DIN1(_27488), .DIN2(_27489), .Q(_27016) );
  nor2s1 _27553_inst ( .DIN1(_27490), .DIN2(_27491), .Q(_27489) );
  nnd2s1 _27554_inst ( .DIN1(_27492), .DIN2(_27493), .Q(_27491) );
  nnd2s1 _27555_inst ( .DIN1(_27335), .DIN2(_27494), .Q(_27490) );
  nor2s1 _27556_inst ( .DIN1(_27376), .DIN2(_27495), .Q(_27488) );
  nnd2s1 _27557_inst ( .DIN1(_27496), .DIN2(_27497), .Q(_27495) );
  nnd2s1 _27558_inst ( .DIN1(_27498), .DIN2(_26378), .Q(_27481) );
  nor2s1 _27559_inst ( .DIN1(_27499), .DIN2(_27500), .Q(
        _________________________________________9_________) );
  nor2s1 _27560_inst ( .DIN1(_27501), .DIN2(_27502), .Q(_27499) );
  nor2s1 _27561_inst ( .DIN1(_27503), .DIN2(_26319), .Q(_27502) );
  nor2s1 _27562_inst ( .DIN1(_26462), .DIN2(_27504), .Q(_27501) );
  nnd2s1 _27563_inst ( .DIN1(_27505), .DIN2(______[6]), .Q(_27504) );
  nnd2s1 _27564_inst ( .DIN1(_27506), .DIN2(_27507), .Q(
        _________________________________________8_________) );
  nnd2s1 _27565_inst ( .DIN1(_27508), .DIN2(_27509), .Q(_27507) );
  nnd2s1 _27566_inst ( .DIN1(_27510), .DIN2(_26467), .Q(_27508) );
  nnd2s1 _27567_inst ( .DIN1(_27511), .DIN2(_27512), .Q(_27506) );
  nor2s1 _27568_inst ( .DIN1(_27513), .DIN2(_27514), .Q(_27511) );
  nor2s1 _27569_inst ( .DIN1(_27515), .DIN2(_27516), .Q(_27514) );
  xor2s1 _27570_inst ( .DIN1(_53008), .DIN2(_26462), .Q(_27515) );
  nor2s1 _27571_inst ( .DIN1(_53376), .DIN2(_27503), .Q(_27513) );
  nnd2s1 _27572_inst ( .DIN1(_27517), .DIN2(_27518), .Q(
        _________________________________________7_________) );
  nnd2s1 _27573_inst ( .DIN1(_27519), .DIN2(_27520), .Q(_27518) );
  nnd2s1 _27574_inst ( .DIN1(_27521), .DIN2(_53272), .Q(_27519) );
  nor2s1 _27575_inst ( .DIN1(_27522), .DIN2(_26771), .Q(_27521) );
  nnd2s1 _27576_inst ( .DIN1(_27523), .DIN2(_27524), .Q(_27517) );
  nor2s1 _27577_inst ( .DIN1(_27525), .DIN2(_27526), .Q(_27523) );
  nor2s1 _27578_inst ( .DIN1(_27527), .DIN2(_27528), .Q(_27526) );
  xor2s1 _27579_inst ( .DIN1(_26479), .DIN2(_27529), .Q(_27528) );
  nor2s1 _27580_inst ( .DIN1(_27503), .DIN2(_26318), .Q(_27525) );
  nnd2s1 _27581_inst ( .DIN1(_27530), .DIN2(_27405), .Q(
        _________________________________________6_________) );
  nor2s1 _27582_inst ( .DIN1(_27531), .DIN2(_27532), .Q(_27530) );
  nor2s1 _27583_inst ( .DIN1(_27408), .DIN2(_27533), .Q(_27532) );
  nnd2s1 _27584_inst ( .DIN1(_27534), .DIN2(_27535), .Q(_27533) );
  nnd2s1 _27585_inst ( .DIN1(_53379), .DIN2(_27536), .Q(_27535) );
  nnd2s1 _27586_inst ( .DIN1(_27537), .DIN2(_27538), .Q(_27534) );
  xor2s1 _27587_inst ( .DIN1(_53011), .DIN2(_27539), .Q(_27538) );
  hi1s1 _27588_inst ( .DIN(_27516), .Q(_27537) );
  nnd2s1 _27589_inst ( .DIN1(______[10]), .DIN2(_27505), .Q(_27516) );
  nor2s1 _27590_inst ( .DIN1(_27421), .DIN2(_27540), .Q(_27531) );
  nor2s1 _27591_inst ( .DIN1(_27541), .DIN2(_27241), .Q(_27540) );
  xor2s1 _27592_inst ( .DIN1(_27542), .DIN2(_53046), .Q(_27541) );
  nnd2s1 _27593_inst ( .DIN1(_53012), .DIN2(_53045), .Q(_27542) );
  nnd2s1 _27594_inst ( .DIN1(_27543), .DIN2(_27544), .Q(
        _________________________________________5_________) );
  nnd2s1 _27595_inst ( .DIN1(_27545), .DIN2(_27546), .Q(_27544) );
  nnd2s1 _27596_inst ( .DIN1(_27547), .DIN2(_27548), .Q(_27545) );
  xor2s1 _27597_inst ( .DIN1(_27549), .DIN2(_27550), .Q(_27548) );
  xor2s1 _27598_inst ( .DIN1(_52884), .DIN2(_53080), .Q(_27550) );
  nnd2s1 _27599_inst ( .DIN1(_53023), .DIN2(_53084), .Q(_27549) );
  nor2s1 _27600_inst ( .DIN1(_27551), .DIN2(_26990), .Q(_27547) );
  nnd2s1 _27601_inst ( .DIN1(_27552), .DIN2(_27164), .Q(_27543) );
  nor2s1 _27602_inst ( .DIN1(_27553), .DIN2(_27554), .Q(_27552) );
  nor2s1 _27603_inst ( .DIN1(_27555), .DIN2(_27556), .Q(_27554) );
  nnd2s1 _27604_inst ( .DIN1(_53012), .DIN2(______[6]), .Q(_27556) );
  nor2s1 _27605_inst ( .DIN1(_27557), .DIN2(_27558), .Q(_27553) );
  nnd2s1 _27606_inst ( .DIN1(_27559), .DIN2(_27560), .Q(
        _________________________________________4_________) );
  nor2s1 _27607_inst ( .DIN1(_27561), .DIN2(_27562), .Q(_27559) );
  nor2s1 _27608_inst ( .DIN1(_27563), .DIN2(_27564), .Q(_27562) );
  nnd2s1 _27609_inst ( .DIN1(_27565), .DIN2(_27566), .Q(_27564) );
  nnd2s1 _27610_inst ( .DIN1(_53381), .DIN2(_27567), .Q(_27566) );
  nnd2s1 _27611_inst ( .DIN1(_27568), .DIN2(_27569), .Q(_27565) );
  nor2s1 _27612_inst ( .DIN1(_27539), .DIN2(_27570), .Q(_27568) );
  nor2s1 _27613_inst ( .DIN1(_53012), .DIN2(_53023), .Q(_27570) );
  hi1s1 _27614_inst ( .DIN(_27529), .Q(_27539) );
  nnd2s1 _27615_inst ( .DIN1(_53012), .DIN2(_53023), .Q(_27529) );
  nor2s1 _27616_inst ( .DIN1(_27571), .DIN2(_27572), .Q(_27561) );
  nor2s1 _27617_inst ( .DIN1(_26854), .DIN2(_27573), .Q(_27572) );
  xor2s1 _27618_inst ( .DIN1(_26374), .DIN2(_27574), .Q(_27573) );
  nnd2s1 _27619_inst ( .DIN1(_27575), .DIN2(_27576), .Q(
        _________________________________________3_________) );
  nor2s1 _27620_inst ( .DIN1(_27577), .DIN2(_27578), .Q(_27575) );
  nor2s1 _27621_inst ( .DIN1(_27579), .DIN2(_27580), .Q(_27578) );
  nor2s1 _27622_inst ( .DIN1(_27581), .DIN2(_27582), .Q(_27580) );
  nor2s1 _27623_inst ( .DIN1(_27557), .DIN2(_26330), .Q(_27582) );
  nor2s1 _27624_inst ( .DIN1(_27567), .DIN2(_27583), .Q(_27581) );
  nnd2s1 _27625_inst ( .DIN1(_27584), .DIN2(_27585), .Q(_27583) );
  nor2s1 _27626_inst ( .DIN1(_27586), .DIN2(_26771), .Q(_27584) );
  xor2s1 _27627_inst ( .DIN1(_27587), .DIN2(_27588), .Q(_27586) );
  and2s1 _27628_inst ( .DIN1(_26399), .DIN2(_53319), .Q(_27588) );
  xor2s1 _27629_inst ( .DIN1(_26663), .DIN2(_53053), .Q(_27587) );
  nor2s1 _27630_inst ( .DIN1(_27589), .DIN2(_27590), .Q(_27577) );
  nor2s1 _27631_inst ( .DIN1(_27591), .DIN2(_26771), .Q(_27590) );
  xor2s1 _27632_inst ( .DIN1(_26499), .DIN2(_53102), .Q(_27591) );
  nor2s1 _27633_inst ( .DIN1(_27592), .DIN2(_27593), .Q(
        _________________________________________2_________) );
  nor2s1 _27634_inst ( .DIN1(_27594), .DIN2(_27595), .Q(_27592) );
  nor2s1 _27635_inst ( .DIN1(_27557), .DIN2(_26320), .Q(_27595) );
  and2s1 _27636_inst ( .DIN1(_26399), .DIN2(_27569), .Q(_27594) );
  nor2s1 _27637_inst ( .DIN1(_27596), .DIN2(_27393), .Q(_27569) );
  nnd2s1 _27638_inst ( .DIN1(_27597), .DIN2(_27598), .Q(
        _________________________________________25_________) );
  nnd2s1 _27639_inst ( .DIN1(_27146), .DIN2(_27599), .Q(_27598) );
  nnd2s1 _27640_inst ( .DIN1(_27600), .DIN2(_27601), .Q(_27599) );
  nnd2s1 _27641_inst ( .DIN1(_27602), .DIN2(_53067), .Q(_27601) );
  nor2s1 _27642_inst ( .DIN1(_26809), .DIN2(_27603), .Q(_27602) );
  nnd2s1 _27643_inst ( .DIN1(_53363), .DIN2(_27604), .Q(_27600) );
  nnd2s1 _27644_inst ( .DIN1(_27605), .DIN2(_27144), .Q(_27597) );
  nor2s1 _27645_inst ( .DIN1(_52842), .DIN2(_27606), .Q(_27605) );
  nnd2s1 _27646_inst ( .DIN1(_27607), .DIN2(_27608), .Q(
        _________________________________________24_________) );
  nor2s1 _27647_inst ( .DIN1(_27609), .DIN2(_27610), .Q(_27607) );
  nor2s1 _27648_inst ( .DIN1(_27611), .DIN2(_27612), .Q(_27610) );
  nor2s1 _27649_inst ( .DIN1(_27613), .DIN2(_27614), .Q(_27612) );
  xor2s1 _27650_inst ( .DIN1(_26673), .DIN2(_53035), .Q(_27613) );
  nor2s1 _27651_inst ( .DIN1(_27615), .DIN2(_27616), .Q(_27609) );
  nor2s1 _27652_inst ( .DIN1(_27617), .DIN2(_27618), .Q(_27615) );
  nor2s1 _27653_inst ( .DIN1(_27619), .DIN2(_27620), .Q(_27618) );
  nor2s1 _27654_inst ( .DIN1(_27603), .DIN2(_27621), .Q(_27617) );
  xor2s1 _27655_inst ( .DIN1(_53067), .DIN2(_53250), .Q(_27621) );
  nnd2s1 _27656_inst ( .DIN1(_27622), .DIN2(_27623), .Q(
        _________________________________________23_________) );
  or2s1 _27657_inst ( .DIN1(_26451), .DIN2(_27624), .Q(_27623) );
  nor2s1 _27658_inst ( .DIN1(_27625), .DIN2(_27626), .Q(_27622) );
  and2s1 _27659_inst ( .DIN1(_27627), .DIN2(_53362), .Q(_27626) );
  nor2s1 _27660_inst ( .DIN1(_27628), .DIN2(_27629), .Q(_27625) );
  nor2s1 _27661_inst ( .DIN1(_27630), .DIN2(_27631), .Q(_27628) );
  xor2s1 _27662_inst ( .DIN1(_53142), .DIN2(_53233), .Q(_27631) );
  nnd2s1 _27663_inst ( .DIN1(_27632), .DIN2(_27633), .Q(
        _________________________________________22_________) );
  nnd2s1 _27664_inst ( .DIN1(_53361), .DIN2(_27627), .Q(_27633) );
  nor2s1 _27665_inst ( .DIN1(_27634), .DIN2(_27635), .Q(_27632) );
  nor2s1 _27666_inst ( .DIN1(_27636), .DIN2(_27629), .Q(_27635) );
  nor2s1 _27667_inst ( .DIN1(_27637), .DIN2(_27638), .Q(_27636) );
  nnd2s1 _27668_inst ( .DIN1(_27639), .DIN2(_27640), .Q(_27638) );
  nnd2s1 _27669_inst ( .DIN1(_27641), .DIN2(_26717), .Q(_27640) );
  nor2s1 _27670_inst ( .DIN1(_53127), .DIN2(_26397), .Q(_27641) );
  nnd2s1 _27671_inst ( .DIN1(_53127), .DIN2(_53115), .Q(_27639) );
  nor2s1 _27672_inst ( .DIN1(_27624), .DIN2(_27642), .Q(_27634) );
  xor2s1 _27673_inst ( .DIN1(_26484), .DIN2(_53115), .Q(_27642) );
  nnd2s1 _27674_inst ( .DIN1(_27643), .DIN2(_27644), .Q(
        _________________________________________21_________) );
  nor2s1 _27675_inst ( .DIN1(_27645), .DIN2(_27646), .Q(_27643) );
  nor2s1 _27676_inst ( .DIN1(_27647), .DIN2(_27648), .Q(_27646) );
  nor2s1 _27677_inst ( .DIN1(_27649), .DIN2(_27650), .Q(_27647) );
  nor2s1 _27678_inst ( .DIN1(_27651), .DIN2(_27652), .Q(_27650) );
  nnd2s1 _27679_inst ( .DIN1(_27653), .DIN2(_26535), .Q(_27652) );
  nor2s1 _27680_inst ( .DIN1(_27654), .DIN2(_26331), .Q(_27649) );
  nor2s1 _27681_inst ( .DIN1(_27655), .DIN2(_27656), .Q(_27645) );
  nor2s1 _27682_inst ( .DIN1(_27657), .DIN2(_27658), .Q(_27656) );
  nor2s1 _27683_inst ( .DIN1(_52846), .DIN2(_53487), .Q(_27657) );
  nnd2s1 _27684_inst ( .DIN1(_27659), .DIN2(_27660), .Q(
        _________________________________________20_________) );
  nor2s1 _27685_inst ( .DIN1(_27661), .DIN2(_27662), .Q(_27659) );
  nor2s1 _27686_inst ( .DIN1(_27663), .DIN2(_27664), .Q(_27662) );
  nnd2s1 _27687_inst ( .DIN1(_27665), .DIN2(_27666), .Q(_27664) );
  nnd2s1 _27688_inst ( .DIN1(_26781), .DIN2(_27667), .Q(_27666) );
  nnd2s1 _27689_inst ( .DIN1(_27668), .DIN2(_27669), .Q(_27665) );
  hi1s1 _27690_inst ( .DIN(_27637), .Q(_27669) );
  nnd2s1 _27691_inst ( .DIN1(_27653), .DIN2(_27670), .Q(_27637) );
  nnd2s1 _27692_inst ( .DIN1(_53115), .DIN2(_26397), .Q(_27670) );
  nor2s1 _27693_inst ( .DIN1(_27671), .DIN2(_26773), .Q(_27668) );
  nor2s1 _27694_inst ( .DIN1(_53115), .DIN2(_26397), .Q(_27671) );
  nor2s1 _27695_inst ( .DIN1(_27672), .DIN2(_27673), .Q(_27661) );
  xor2s1 _27696_inst ( .DIN1(_27674), .DIN2(_53341), .Q(_27673) );
  nnd2s1 _27697_inst ( .DIN1(_27675), .DIN2(_27676), .Q(
        _________________________________________1_________) );
  nor2s1 _27698_inst ( .DIN1(_27677), .DIN2(_27678), .Q(_27675) );
  nor2s1 _27699_inst ( .DIN1(_27679), .DIN2(_27680), .Q(_27678) );
  nnd2s1 _27700_inst ( .DIN1(_27681), .DIN2(_27682), .Q(_27680) );
  nnd2s1 _27701_inst ( .DIN1(_53352), .DIN2(_27567), .Q(_27682) );
  nnd2s1 _27702_inst ( .DIN1(_53053), .DIN2(_27683), .Q(_27681) );
  nor2s1 _27703_inst ( .DIN1(_27684), .DIN2(_27685), .Q(_27677) );
  xor2s1 _27704_inst ( .DIN1(_26450), .DIN2(_27686), .Q(_27685) );
  nnd2s1 _27705_inst ( .DIN1(_53131), .DIN2(_53132), .Q(_27686) );
  nnd2s1 _27706_inst ( .DIN1(_27687), .DIN2(_27688), .Q(
        _________________________________________19_________) );
  nor2s1 _27707_inst ( .DIN1(_27689), .DIN2(_27690), .Q(_27687) );
  nor2s1 _27708_inst ( .DIN1(_27691), .DIN2(_27692), .Q(_27690) );
  nor2s1 _27709_inst ( .DIN1(_27693), .DIN2(_27694), .Q(_27691) );
  nor2s1 _27710_inst ( .DIN1(_27630), .DIN2(_27695), .Q(_27694) );
  nnd2s1 _27711_inst ( .DIN1(______[18]), .DIN2(_27696), .Q(_27695) );
  xor2s1 _27712_inst ( .DIN1(_27697), .DIN2(_27698), .Q(_27696) );
  xor2s1 _27713_inst ( .DIN1(_53178), .DIN2(_53470), .Q(_27698) );
  and2s1 _27714_inst ( .DIN1(_26439), .DIN2(_53193), .Q(_27697) );
  nor2s1 _27715_inst ( .DIN1(_27654), .DIN2(_26209), .Q(_27693) );
  nor2s1 _27716_inst ( .DIN1(_27699), .DIN2(_27700), .Q(_27689) );
  xor2s1 _27717_inst ( .DIN1(_27701), .DIN2(_52885), .Q(_27700) );
  nnd2s1 _27718_inst ( .DIN1(_53011), .DIN2(_53272), .Q(_27701) );
  nnd2s1 _27719_inst ( .DIN1(_27702), .DIN2(_27703), .Q(
        _________________________________________18_________) );
  nnd2s1 _27720_inst ( .DIN1(_27627), .DIN2(_26526), .Q(_27703) );
  nor2s1 _27721_inst ( .DIN1(_27654), .DIN2(_27579), .Q(_27627) );
  nor2s1 _27722_inst ( .DIN1(_27704), .DIN2(_27705), .Q(_27702) );
  nor2s1 _27723_inst ( .DIN1(_27706), .DIN2(_27629), .Q(_27705) );
  nnd2s1 _27724_inst ( .DIN1(_27589), .DIN2(_27654), .Q(_27629) );
  hi1s1 _27725_inst ( .DIN(_27667), .Q(_27654) );
  nor2s1 _27726_inst ( .DIN1(_27707), .DIN2(_27708), .Q(_27667) );
  nor2s1 _27727_inst ( .DIN1(_53165), .DIN2(_27630), .Q(_27706) );
  nor2s1 _27728_inst ( .DIN1(_27624), .DIN2(_27709), .Q(_27704) );
  xnr2s1 _27729_inst ( .DIN1(_53026), .DIN2(_27710), .Q(_27709) );
  nnd2s1 _27730_inst ( .DIN1(_53318), .DIN2(_53102), .Q(_27710) );
  nnd2s1 _27731_inst ( .DIN1(_27711), .DIN2(_27712), .Q(
        _________________________________________17_________) );
  nnd2s1 _27732_inst ( .DIN1(_53314), .DIN2(_27713), .Q(_27712) );
  nnd2s1 _27733_inst ( .DIN1(_27714), .DIN2(_27715), .Q(
        _________________________________________16_________) );
  nnd2s1 _27734_inst ( .DIN1(_27716), .DIN2(_27717), .Q(_27715) );
  nor2s1 _27735_inst ( .DIN1(_27718), .DIN2(_26771), .Q(_27716) );
  xor2s1 _27736_inst ( .DIN1(_27719), .DIN2(_53103), .Q(_27718) );
  nnd2s1 _27737_inst ( .DIN1(_53470), .DIN2(_53035), .Q(_27719) );
  nnd2s1 _27738_inst ( .DIN1(_27611), .DIN2(_27720), .Q(_27714) );
  nnd2s1 _27739_inst ( .DIN1(_53371), .DIN2(_27721), .Q(_27720) );
  nor2s1 _27740_inst ( .DIN1(_26778), .DIN2(_27722), .Q(
        _________________________________________15_________) );
  nnd2s1 _27741_inst ( .DIN1(_27721), .DIN2(_27723), .Q(_27722) );
  nnd2s1 _27742_inst ( .DIN1(_27724), .DIN2(_27688), .Q(
        _________________________________________14_________) );
  hi1s1 _27743_inst ( .DIN(_27725), .Q(_27688) );
  nor2s1 _27744_inst ( .DIN1(_27726), .DIN2(_27727), .Q(_27724) );
  nor2s1 _27745_inst ( .DIN1(_27728), .DIN2(_27692), .Q(_27727) );
  nor2s1 _27746_inst ( .DIN1(_27729), .DIN2(_26323), .Q(_27728) );
  nor2s1 _27747_inst ( .DIN1(______[13]), .DIN2(_27699), .Q(_27726) );
  nnd2s1 _27748_inst ( .DIN1(_27711), .DIN2(_27730), .Q(
        _________________________________________13_________) );
  nnd2s1 _27749_inst ( .DIN1(_27713), .DIN2(_27731), .Q(_27730) );
  nnd2s1 _27750_inst ( .DIN1(_27732), .DIN2(_27692), .Q(_27711) );
  nnd2s1 _27751_inst ( .DIN1(_27733), .DIN2(_27734), .Q(
        _________________________________________12_________) );
  nnd2s1 _27752_inst ( .DIN1(_53373), .DIN2(_27713), .Q(_27734) );
  nor2s1 _27753_inst ( .DIN1(_27729), .DIN2(_27692), .Q(_27713) );
  hi1s1 _27754_inst ( .DIN(_27721), .Q(_27729) );
  nor2s1 _27755_inst ( .DIN1(_27725), .DIN2(_27735), .Q(_27733) );
  nor2s1 _27756_inst ( .DIN1(_27699), .DIN2(_27736), .Q(_27735) );
  nor2s1 _27757_inst ( .DIN1(_27737), .DIN2(_27241), .Q(_27736) );
  xor2s1 _27758_inst ( .DIN1(_26439), .DIN2(_53011), .Q(_27737) );
  nor2s1 _27759_inst ( .DIN1(_27732), .DIN2(_27699), .Q(_27725) );
  hi1s1 _27760_inst ( .DIN(_27692), .Q(_27699) );
  nnd2s1 _27761_inst ( .DIN1(_27738), .DIN2(_27739), .Q(_27692) );
  nor2s1 _27762_inst ( .DIN1(_27740), .DIN2(_27741), .Q(_27739) );
  or2s1 _27763_inst ( .DIN1(_27742), .DIN2(_27743), .Q(_27741) );
  nor2s1 _27764_inst ( .DIN1(_27744), .DIN2(_27745), .Q(_27738) );
  or2s1 _27765_inst ( .DIN1(_27746), .DIN2(_27747), .Q(_27732) );
  nor2s1 _27766_inst ( .DIN1(_27748), .DIN2(_27749), .Q(
        _________________________________________11_________) );
  nor2s1 _27767_inst ( .DIN1(_27750), .DIN2(_27751), .Q(_27748) );
  nor2s1 _27768_inst ( .DIN1(_27503), .DIN2(_26322), .Q(_27751) );
  nor2s1 _27769_inst ( .DIN1(_27527), .DIN2(_27752), .Q(_27750) );
  xor2s1 _27770_inst ( .DIN1(_27753), .DIN2(_27754), .Q(_27752) );
  xor2s1 _27771_inst ( .DIN1(_53316), .DIN2(_53465), .Q(_27754) );
  and2s1 _27772_inst ( .DIN1(_53008), .DIN2(_53295), .Q(_27753) );
  hi1s1 _27773_inst ( .DIN(_27505), .Q(_27527) );
  nnd2s1 _27774_inst ( .DIN1(_27755), .DIN2(_27676), .Q(
        _________________________________________10_________) );
  nor2s1 _27775_inst ( .DIN1(_27756), .DIN2(_27757), .Q(_27755) );
  nor2s1 _27776_inst ( .DIN1(_27679), .DIN2(_27758), .Q(_27757) );
  nnd2s1 _27777_inst ( .DIN1(_27759), .DIN2(_27760), .Q(_27758) );
  nnd2s1 _27778_inst ( .DIN1(_53295), .DIN2(_27505), .Q(_27760) );
  nor2s1 _27779_inst ( .DIN1(_27536), .DIN2(_27761), .Q(_27505) );
  nnd2s1 _27780_inst ( .DIN1(_53372), .DIN2(_27536), .Q(_27759) );
  nor2s1 _27781_inst ( .DIN1(_27684), .DIN2(_27762), .Q(_27756) );
  xor2s1 _27782_inst ( .DIN1(_26220), .DIN2(_27763), .Q(_27762) );
  nnd2s1 _27783_inst ( .DIN1(_53316), .DIN2(_53125), .Q(_27763) );
  nnd2s1 _27784_inst ( .DIN1(_27764), .DIN2(_27576), .Q(
        _________________________________________0_________) );
  nor2s1 _27785_inst ( .DIN1(_27765), .DIN2(_27766), .Q(_27764) );
  nor2s1 _27786_inst ( .DIN1(_27579), .DIN2(_27767), .Q(_27766) );
  nor2s1 _27787_inst ( .DIN1(_27768), .DIN2(_27769), .Q(_27767) );
  nor2s1 _27788_inst ( .DIN1(_26850), .DIN2(_27158), .Q(_27769) );
  nor2s1 _27789_inst ( .DIN1(_27135), .DIN2(_27770), .Q(_27768) );
  nnd2s1 _27790_inst ( .DIN1(_27771), .DIN2(_53208), .Q(_27770) );
  nor2s1 _27791_inst ( .DIN1(_27160), .DIN2(_26771), .Q(_27771) );
  nor2s1 _27792_inst ( .DIN1(_27589), .DIN2(_27772), .Q(_27765) );
  nor2s1 _27793_inst ( .DIN1(_27773), .DIN2(_27774), .Q(_27772) );
  xor2s1 _27794_inst ( .DIN1(_27775), .DIN2(_53056), .Q(_27773) );
  nnd2s1 _27795_inst ( .DIN1(_53115), .DIN2(_53354), .Q(_27775) );
  nnd2s1 _27796_inst ( .DIN1(_27776), .DIN2(_27777), .Q(
        _________________________________________0________5____________) );
  nnd2s1 _27797_inst ( .DIN1(_27778), .DIN2(_27779), .Q(_27777) );
  nnd2s1 _27798_inst ( .DIN1(_26537), .DIN2(_27780), .Q(_27778) );
  nnd2s1 _27799_inst ( .DIN1(_27781), .DIN2(_27782), .Q(_27776) );
  nnd2s1 _27800_inst ( .DIN1(_27783), .DIN2(_27784), .Q(_27781) );
  nnd2s1 _27801_inst ( .DIN1(_27785), .DIN2(_27786), .Q(_27784) );
  nor2s1 _27802_inst ( .DIN1(_27787), .DIN2(_27788), .Q(_27785) );
  xor2s1 _27803_inst ( .DIN1(_27789), .DIN2(_53141), .Q(_27788) );
  nnd2s1 _27804_inst ( .DIN1(_53132), .DIN2(_26530), .Q(_27789) );
  nnd2s1 _27805_inst ( .DIN1(_27790), .DIN2(_27676), .Q(
        _________________________________________0________4____________) );
  nor2s1 _27806_inst ( .DIN1(_27791), .DIN2(_27792), .Q(_27790) );
  nor2s1 _27807_inst ( .DIN1(_27679), .DIN2(_27793), .Q(_27792) );
  nnd2s1 _27808_inst ( .DIN1(_27794), .DIN2(_27783), .Q(_27793) );
  nnd2s1 _27809_inst ( .DIN1(_27795), .DIN2(_26849), .Q(_27783) );
  nnd2s1 _27810_inst ( .DIN1(_27796), .DIN2(_27797), .Q(_27794) );
  xor2s1 _27811_inst ( .DIN1(_26530), .DIN2(_53051), .Q(_27796) );
  nor2s1 _27812_inst ( .DIN1(_27684), .DIN2(_27798), .Q(_27791) );
  nor2s1 _27813_inst ( .DIN1(_27799), .DIN2(_27241), .Q(_27798) );
  xnr2s1 _27814_inst ( .DIN1(_53319), .DIN2(_53131), .Q(_27799) );
  nnd2s1 _27815_inst ( .DIN1(_27800), .DIN2(_27801), .Q(
        _________________________________________0________3____________) );
  nnd2s1 _27816_inst ( .DIN1(_27802), .DIN2(_27803), .Q(_27801) );
  xor2s1 _27817_inst ( .DIN1(_52951), .DIN2(_52952), .Q(_27803) );
  hi1s1 _27818_inst ( .DIN(_27804), .Q(_27802) );
  nnd2s1 _27819_inst ( .DIN1(_27805), .DIN2(_27806), .Q(_27800) );
  nor2s1 _27820_inst ( .DIN1(_27807), .DIN2(_27808), .Q(_27805) );
  nor2s1 _27821_inst ( .DIN1(_27604), .DIN2(_27809), .Q(_27808) );
  nnd2s1 _27822_inst ( .DIN1(_53132), .DIN2(_27810), .Q(_27809) );
  nor2s1 _27823_inst ( .DIN1(_26850), .DIN2(_27619), .Q(_27807) );
  nnd2s1 _27824_inst ( .DIN1(_27811), .DIN2(_27660), .Q(
        _________________________________________0________2____________) );
  nor2s1 _27825_inst ( .DIN1(_27812), .DIN2(_27813), .Q(_27811) );
  nor2s1 _27826_inst ( .DIN1(_27672), .DIN2(_27814), .Q(_27813) );
  xor2s1 _27827_inst ( .DIN1(_27815), .DIN2(_52972), .Q(_27814) );
  nor2s1 _27828_inst ( .DIN1(_27816), .DIN2(_27663), .Q(_27812) );
  nor2s1 _27829_inst ( .DIN1(_27817), .DIN2(_27818), .Q(_27816) );
  nor2s1 _27830_inst ( .DIN1(_27603), .DIN2(_27819), .Q(_27817) );
  xor2s1 _27831_inst ( .DIN1(_53052), .DIN2(_53132), .Q(_27819) );
  nnd2s1 _27832_inst ( .DIN1(_27820), .DIN2(_27576), .Q(
        _________________________________________0________1____________) );
  nnd2s1 _27833_inst ( .DIN1(_27624), .DIN2(_27579), .Q(_27576) );
  nor2s1 _27834_inst ( .DIN1(_27821), .DIN2(_27822), .Q(_27624) );
  nor2s1 _27835_inst ( .DIN1(_27823), .DIN2(_27824), .Q(_27820) );
  nor2s1 _27836_inst ( .DIN1(_27589), .DIN2(_27825), .Q(_27824) );
  xor2s1 _27837_inst ( .DIN1(_53115), .DIN2(_53127), .Q(_27825) );
  hi1s1 _27838_inst ( .DIN(_27579), .Q(_27589) );
  nor2s1 _27839_inst ( .DIN1(_27826), .DIN2(_27579), .Q(_27823) );
  nnd2s1 _27840_inst ( .DIN1(_27827), .DIN2(_27828), .Q(_27579) );
  nor2s1 _27841_inst ( .DIN1(_27829), .DIN2(_27818), .Q(_27826) );
  hi1s1 _27842_inst ( .DIN(_27830), .Q(_27818) );
  nor2s1 _27843_inst ( .DIN1(_27603), .DIN2(_27831), .Q(_27829) );
  xor2s1 _27844_inst ( .DIN1(_27832), .DIN2(_27833), .Q(_27831) );
  xor2s1 _27845_inst ( .DIN1(_53067), .DIN2(_53103), .Q(_27833) );
  nor2s1 _27846_inst ( .DIN1(_53250), .DIN2(_53056), .Q(_27832) );
  nnd2s1 _27847_inst ( .DIN1(_27834), .DIN2(_27835), .Q(
        _________________________________________0________0____________) );
  nnd2s1 _27848_inst ( .DIN1(_27836), .DIN2(_27837), .Q(_27835) );
  nnd2s1 _27849_inst ( .DIN1(_27830), .DIN2(_27838), .Q(_27837) );
  or2s1 _27850_inst ( .DIN1(_27603), .DIN2(_53056), .Q(_27838) );
  nnd2s1 _27851_inst ( .DIN1(_27619), .DIN2(_27810), .Q(_27603) );
  hi1s1 _27852_inst ( .DIN(_27604), .Q(_27619) );
  nnd2s1 _27853_inst ( .DIN1(_53384), .DIN2(_27604), .Q(_27830) );
  xor2s1 _27854_inst ( .DIN1(_27839), .DIN2(_27840), .Q(_27604) );
  nnd2s1 _27855_inst ( .DIN1(_27841), .DIN2(_27842), .Q(_27839) );
  nor2s1 _27856_inst ( .DIN1(_27653), .DIN2(_27843), .Q(_27841) );
  nnd2s1 _27857_inst ( .DIN1(_27844), .DIN2(_27845), .Q(_27834) );
  nor2s1 _27858_inst ( .DIN1(_27846), .DIN2(_27847), .Q(_27844) );
  nnd2s1 _27859_inst ( .DIN1(_27848), .DIN2(_27849), .Q(_27847) );
  nnd2s1 _27860_inst ( .DIN1(_27850), .DIN2(_26367), .Q(_27848) );
  nnd2s1 _27861_inst ( .DIN1(_53186), .DIN2(_53067), .Q(_27850) );
  nor2s1 _27862_inst ( .DIN1(_26593), .DIN2(_27851), .Q(_27846) );
  nnd2s1 _27863_inst ( .DIN1(_27852), .DIN2(_27853), .Q(
        __________________________________9_________) );
  nnd2s1 _27864_inst ( .DIN1(_27854), .DIN2(_27845), .Q(_27853) );
  nor2s1 _27865_inst ( .DIN1(_27855), .DIN2(_26230), .Q(_27854) );
  nnd2s1 _27866_inst ( .DIN1(_27856), .DIN2(_27836), .Q(_27852) );
  nnd2s1 _27867_inst ( .DIN1(_27857), .DIN2(_27858), .Q(_27856) );
  nnd2s1 _27868_inst ( .DIN1(_27859), .DIN2(_27860), .Q(_27858) );
  nor2s1 _27869_inst ( .DIN1(_27861), .DIN2(_27862), .Q(_27859) );
  xor2s1 _27870_inst ( .DIN1(_27863), .DIN2(_53497), .Q(_27861) );
  nnd2s1 _27871_inst ( .DIN1(_27864), .DIN2(_52917), .Q(_27857) );
  nnd2s1 _27872_inst ( .DIN1(_27865), .DIN2(_27866), .Q(
        __________________________________8_________) );
  nnd2s1 _27873_inst ( .DIN1(_27867), .DIN2(_27868), .Q(_27866) );
  nor2s1 _27874_inst ( .DIN1(_27869), .DIN2(_27870), .Q(_27867) );
  and2s1 _27875_inst ( .DIN1(_52964), .DIN2(_27864), .Q(_27870) );
  nor2s1 _27876_inst ( .DIN1(_27864), .DIN2(_27871), .Q(_27869) );
  nnd2s1 _27877_inst ( .DIN1(_27872), .DIN2(______[26]), .Q(_27871) );
  nor2s1 _27878_inst ( .DIN1(_27873), .DIN2(_27874), .Q(_27872) );
  xor2s1 _27879_inst ( .DIN1(_27863), .DIN2(_52843), .Q(_27874) );
  nnd2s1 _27880_inst ( .DIN1(_27875), .DIN2(_26542), .Q(_27865) );
  nnd2s1 _27881_inst ( .DIN1(_27876), .DIN2(_27877), .Q(
        __________________________________7_________) );
  nnd2s1 _27882_inst ( .DIN1(_27878), .DIN2(_27879), .Q(_27877) );
  xor2s1 _27883_inst ( .DIN1(_27880), .DIN2(_53364), .Q(_27879) );
  nor2s1 _27884_inst ( .DIN1(_26854), .DIN2(_27881), .Q(_27878) );
  nnd2s1 _27885_inst ( .DIN1(_27882), .DIN2(_27883), .Q(_27876) );
  nnd2s1 _27886_inst ( .DIN1(_27884), .DIN2(_27885), .Q(_27883) );
  nor2s1 _27887_inst ( .DIN1(_27886), .DIN2(_27887), .Q(_27884) );
  nor2s1 _27888_inst ( .DIN1(_27888), .DIN2(_26614), .Q(_27887) );
  nor2s1 _27889_inst ( .DIN1(_27889), .DIN2(_27890), .Q(_27886) );
  xor2s1 _27890_inst ( .DIN1(_26454), .DIN2(_53156), .Q(_27890) );
  nnd2s1 _27891_inst ( .DIN1(_27891), .DIN2(_27892), .Q(
        __________________________________6_________) );
  nnd2s1 _27892_inst ( .DIN1(_27893), .DIN2(_27894), .Q(_27892) );
  nor2s1 _27893_inst ( .DIN1(_53404), .DIN2(_26989), .Q(_27893) );
  nnd2s1 _27894_inst ( .DIN1(_27895), .DIN2(_27896), .Q(_27891) );
  nnd2s1 _27895_inst ( .DIN1(_27897), .DIN2(_27885), .Q(_27896) );
  nor2s1 _27896_inst ( .DIN1(_27898), .DIN2(_27899), .Q(_27897) );
  nor2s1 _27897_inst ( .DIN1(_27889), .DIN2(_27900), .Q(_27899) );
  nor2s1 _27898_inst ( .DIN1(_53273), .DIN2(_27888), .Q(_27898) );
  nnd2s1 _27899_inst ( .DIN1(_27901), .DIN2(_27902), .Q(
        __________________________________5_________) );
  nnd2s1 _27900_inst ( .DIN1(_27903), .DIN2(_27904), .Q(_27902) );
  xor2s1 _27901_inst ( .DIN1(_52848), .DIN2(_52849), .Q(_27904) );
  nnd2s1 _27902_inst ( .DIN1(_27298), .DIN2(_27905), .Q(_27901) );
  nnd2s1 _27903_inst ( .DIN1(_27906), .DIN2(_27885), .Q(_27905) );
  nor2s1 _27904_inst ( .DIN1(_27907), .DIN2(_27908), .Q(_27906) );
  nor2s1 _27905_inst ( .DIN1(_27889), .DIN2(_27909), .Q(_27908) );
  nor2s1 _27906_inst ( .DIN1(_53507), .DIN2(_27614), .Q(_27909) );
  nor2s1 _27907_inst ( .DIN1(_27888), .DIN2(_26527), .Q(_27907) );
  nnd2s1 _27908_inst ( .DIN1(_27910), .DIN2(_27911), .Q(
        __________________________________4_________) );
  nnd2s1 _27909_inst ( .DIN1(_27912), .DIN2(______[26]), .Q(_27911) );
  nor2s1 _27910_inst ( .DIN1(_27913), .DIN2(_27914), .Q(_27912) );
  xor2s1 _27911_inst ( .DIN1(_53506), .DIN2(_26465), .Q(_27914) );
  nnd2s1 _27912_inst ( .DIN1(_27915), .DIN2(_27916), .Q(_27910) );
  nnd2s1 _27913_inst ( .DIN1(_27917), .DIN2(_27885), .Q(_27916) );
  nor2s1 _27914_inst ( .DIN1(_27918), .DIN2(_27919), .Q(_27917) );
  nor2s1 _27915_inst ( .DIN1(_27889), .DIN2(_27920), .Q(_27919) );
  nor2s1 _27916_inst ( .DIN1(_27921), .DIN2(_27291), .Q(_27920) );
  xor2s1 _27917_inst ( .DIN1(_27922), .DIN2(_27923), .Q(_27921) );
  xor2s1 _27918_inst ( .DIN1(_27924), .DIN2(_27925), .Q(_27923) );
  nor2s1 _27919_inst ( .DIN1(_53507), .DIN2(_53156), .Q(_27925) );
  xor2s1 _27920_inst ( .DIN1(_26454), .DIN2(_53360), .Q(_27922) );
  nor2s1 _27921_inst ( .DIN1(_27888), .DIN2(_26581), .Q(_27918) );
  nnd2s1 _27922_inst ( .DIN1(_27926), .DIN2(_27927), .Q(
        __________________________________3_________) );
  nnd2s1 _27923_inst ( .DIN1(_27928), .DIN2(_27929), .Q(_27927) );
  nnd2s1 _27924_inst ( .DIN1(_27930), .DIN2(_27931), .Q(_27928) );
  xnr2s1 _27925_inst ( .DIN1(_52922), .DIN2(_27932), .Q(_27931) );
  nor2s1 _27926_inst ( .DIN1(_53509), .DIN2(_53497), .Q(_27932) );
  nor2s1 _27927_inst ( .DIN1(_27933), .DIN2(_27241), .Q(_27930) );
  nor2s1 _27928_inst ( .DIN1(_27934), .DIN2(_27935), .Q(_27933) );
  or2s1 _27929_inst ( .DIN1(_27936), .DIN2(_27937), .Q(_27935) );
  nnd2s1 _27930_inst ( .DIN1(_27938), .DIN2(_27868), .Q(_27926) );
  nor2s1 _27931_inst ( .DIN1(_27939), .DIN2(_27940), .Q(_27938) );
  nnd2s1 _27932_inst ( .DIN1(_27941), .DIN2(_27942), .Q(_27940) );
  nnd2s1 _27933_inst ( .DIN1(_27889), .DIN2(_26688), .Q(_27942) );
  nnd2s1 _27934_inst ( .DIN1(_27943), .DIN2(_27888), .Q(_27941) );
  xor2s1 _27935_inst ( .DIN1(_26562), .DIN2(_53506), .Q(_27943) );
  hi1s1 _27936_inst ( .DIN(_27885), .Q(_27939) );
  nnd2s1 _27937_inst ( .DIN1(_27944), .DIN2(_27945), .Q(
        __________________________________31_________) );
  nnd2s1 _27938_inst ( .DIN1(_27246), .DIN2(_27946), .Q(_27945) );
  xor2s1 _27939_inst ( .DIN1(_26502), .DIN2(_27947), .Q(_27946) );
  nnd2s1 _27940_inst ( .DIN1(_52898), .DIN2(_52883), .Q(_27947) );
  nnd2s1 _27941_inst ( .DIN1(_27247), .DIN2(_27948), .Q(_27944) );
  nnd2s1 _27942_inst ( .DIN1(_27949), .DIN2(_27950), .Q(_27948) );
  nnd2s1 _27943_inst ( .DIN1(_52900), .DIN2(_27951), .Q(_27950) );
  nnd2s1 _27944_inst ( .DIN1(_27952), .DIN2(_27953), .Q(_27949) );
  xnr2s1 _27945_inst ( .DIN1(_53106), .DIN2(_27954), .Q(_27953) );
  nnd2s1 _27946_inst ( .DIN1(_52885), .DIN2(_26402), .Q(_27954) );
  xor2s1 _27947_inst ( .DIN1(_27955), .DIN2(_27956), .Q(_27952) );
  nnd2s1 _27948_inst ( .DIN1(_27957), .DIN2(_27958), .Q(
        __________________________________30_________) );
  nnd2s1 _27949_inst ( .DIN1(_27959), .DIN2(_27960), .Q(_27958) );
  nor2s1 _27950_inst ( .DIN1(_27961), .DIN2(_27962), .Q(_27960) );
  nor2s1 _27951_inst ( .DIN1(_27963), .DIN2(_27964), .Q(_27962) );
  nor2s1 _27952_inst ( .DIN1(_26425), .DIN2(_27241), .Q(_27964) );
  nor2s1 _27953_inst ( .DIN1(_53464), .DIN2(_27965), .Q(_27961) );
  nor2s1 _27954_inst ( .DIN1(_27966), .DIN2(_27967), .Q(_27959) );
  nnd2s1 _27955_inst ( .DIN1(_52920), .DIN2(_27968), .Q(_27957) );
  nnd2s1 _27956_inst ( .DIN1(_27969), .DIN2(_27970), .Q(
        __________________________________2_________) );
  nor2s1 _27957_inst ( .DIN1(_27971), .DIN2(_27972), .Q(_27969) );
  nor2s1 _27958_inst ( .DIN1(_27973), .DIN2(_27974), .Q(_27972) );
  nnd2s1 _27959_inst ( .DIN1(_27975), .DIN2(_27885), .Q(_27974) );
  nnd2s1 _27960_inst ( .DIN1(_27976), .DIN2(_27873), .Q(_27885) );
  nor2s1 _27961_inst ( .DIN1(_27977), .DIN2(_27889), .Q(_27976) );
  nor2s1 _27962_inst ( .DIN1(_27978), .DIN2(_27979), .Q(_27975) );
  nor2s1 _27963_inst ( .DIN1(_53512), .DIN2(_27889), .Q(_27979) );
  and2s1 _27964_inst ( .DIN1(_27889), .DIN2(_53238), .Q(_27978) );
  nor2s1 _27965_inst ( .DIN1(_27915), .DIN2(_27980), .Q(_27971) );
  nor2s1 _27966_inst ( .DIN1(_26855), .DIN2(_27981), .Q(_27980) );
  xor2s1 _27967_inst ( .DIN1(_53455), .DIN2(_53507), .Q(_27981) );
  nnd2s1 _27968_inst ( .DIN1(_27982), .DIN2(_27983), .Q(
        __________________________________29_________) );
  nor2s1 _27969_inst ( .DIN1(_27984), .DIN2(_27985), .Q(_27982) );
  nor2s1 _27970_inst ( .DIN1(_27500), .DIN2(_27986), .Q(_27985) );
  nnd2s1 _27971_inst ( .DIN1(_27987), .DIN2(_27988), .Q(_27986) );
  nor2s1 _27972_inst ( .DIN1(_27989), .DIN2(_27990), .Q(_27988) );
  nor2s1 _27973_inst ( .DIN1(_53188), .DIN2(_27991), .Q(_27990) );
  nor2s1 _27974_inst ( .DIN1(_26434), .DIN2(_27992), .Q(_27989) );
  nor2s1 _27975_inst ( .DIN1(_27966), .DIN2(_27993), .Q(_27987) );
  nor2s1 _27976_inst ( .DIN1(_52902), .DIN2(_27965), .Q(_27993) );
  nor2s1 _27977_inst ( .DIN1(_27994), .DIN2(_27995), .Q(_27984) );
  nor2s1 _27978_inst ( .DIN1(_26853), .DIN2(_27996), .Q(_27995) );
  xor2s1 _27979_inst ( .DIN1(_53104), .DIN2(_53206), .Q(_27996) );
  nnd2s1 _27980_inst ( .DIN1(_27997), .DIN2(_27998), .Q(
        __________________________________28_________) );
  nor2s1 _27981_inst ( .DIN1(_27999), .DIN2(_28000), .Q(_27997) );
  nor2s1 _27982_inst ( .DIN1(_27749), .DIN2(_28001), .Q(_28000) );
  nnd2s1 _27983_inst ( .DIN1(_28002), .DIN2(_28003), .Q(_28001) );
  nor2s1 _27984_inst ( .DIN1(_28004), .DIN2(_28005), .Q(_28003) );
  nor2s1 _27985_inst ( .DIN1(_53359), .DIN2(_27991), .Q(_28005) );
  nnd2s1 _27986_inst ( .DIN1(_27965), .DIN2(_28006), .Q(_27991) );
  nor2s1 _27987_inst ( .DIN1(_26618), .DIN2(_27992), .Q(_28004) );
  nnd2s1 _27988_inst ( .DIN1(_28007), .DIN2(_27965), .Q(_27992) );
  hi1s1 _27989_inst ( .DIN(_28006), .Q(_28007) );
  nor2s1 _27990_inst ( .DIN1(_27966), .DIN2(_28008), .Q(_28002) );
  nor2s1 _27991_inst ( .DIN1(_53040), .DIN2(_27965), .Q(_28008) );
  hi1s1 _27992_inst ( .DIN(_28009), .Q(_27966) );
  nor2s1 _27993_inst ( .DIN1(_28010), .DIN2(_28011), .Q(_27999) );
  xor2s1 _27994_inst ( .DIN1(_26554), .DIN2(_53523), .Q(_28011) );
  nnd2s1 _27995_inst ( .DIN1(_28012), .DIN2(_28013), .Q(
        __________________________________27_________) );
  nor2s1 _27996_inst ( .DIN1(_28014), .DIN2(_28015), .Q(_28013) );
  nor2s1 _27997_inst ( .DIN1(_28016), .DIN2(_28017), .Q(_28015) );
  nnd2s1 _27998_inst ( .DIN1(_28018), .DIN2(_28009), .Q(_28017) );
  nor2s1 _27999_inst ( .DIN1(_28019), .DIN2(_28020), .Q(_28018) );
  nor2s1 _28000_inst ( .DIN1(_27963), .DIN2(_28021), .Q(_28020) );
  nor2s1 _28001_inst ( .DIN1(_28022), .DIN2(_28023), .Q(_28021) );
  and2s1 _28002_inst ( .DIN1(_53045), .DIN2(_53463), .Q(_28023) );
  and2s1 _28003_inst ( .DIN1(_27963), .DIN2(_52903), .Q(_28019) );
  nor2s1 _28004_inst ( .DIN1(_28024), .DIN2(_28025), .Q(_28014) );
  or2s1 _28005_inst ( .DIN1(_53232), .DIN2(_53231), .Q(_28025) );
  and2s1 _28006_inst ( .DIN1(_28026), .DIN2(_28027), .Q(_28012) );
  nnd2s1 _28007_inst ( .DIN1(_28028), .DIN2(_28029), .Q(
        __________________________________26_________) );
  nor2s1 _28008_inst ( .DIN1(_28030), .DIN2(_28031), .Q(_28029) );
  nor2s1 _28009_inst ( .DIN1(_28032), .DIN2(_28033), .Q(_28031) );
  nnd2s1 _28010_inst ( .DIN1(_28034), .DIN2(_28009), .Q(_28033) );
  nor2s1 _28011_inst ( .DIN1(_28035), .DIN2(_28036), .Q(_28034) );
  nor2s1 _28012_inst ( .DIN1(_27963), .DIN2(_26429), .Q(_28036) );
  nor2s1 _28013_inst ( .DIN1(_52834), .DIN2(_27965), .Q(_28035) );
  nor2s1 _28014_inst ( .DIN1(_28037), .DIN2(_28038), .Q(_28030) );
  nor2s1 _28015_inst ( .DIN1(_28039), .DIN2(_27774), .Q(_28038) );
  and2s1 _28016_inst ( .DIN1(_28040), .DIN2(_53479), .Q(_28039) );
  nor2s1 _28017_inst ( .DIN1(_28041), .DIN2(_28042), .Q(_28028) );
  nor2s1 _28018_inst ( .DIN1(_53479), .DIN2(_28043), .Q(_28042) );
  nnd2s1 _28019_inst ( .DIN1(_28044), .DIN2(_28045), .Q(
        __________________________________25_________) );
  nor2s1 _28020_inst ( .DIN1(_28046), .DIN2(_28047), .Q(_28044) );
  nor2s1 _28021_inst ( .DIN1(_28048), .DIN2(_28049), .Q(_28047) );
  nor2s1 _28022_inst ( .DIN1(_28050), .DIN2(_28051), .Q(_28048) );
  nor2s1 _28023_inst ( .DIN1(_28052), .DIN2(_26382), .Q(_28051) );
  nor2s1 _28024_inst ( .DIN1(_27066), .DIN2(_28053), .Q(_28050) );
  nnd2s1 _28025_inst ( .DIN1(_28054), .DIN2(_28055), .Q(_28053) );
  xor2s1 _28026_inst ( .DIN1(_52981), .DIN2(_28022), .Q(_28054) );
  nor2s1 _28027_inst ( .DIN1(_28056), .DIN2(_28057), .Q(_28046) );
  and2s1 _28028_inst ( .DIN1(______[8]), .DIN2(_53012), .Q(_28057) );
  nnd2s1 _28029_inst ( .DIN1(_28058), .DIN2(_28059), .Q(
        __________________________________24_________) );
  nnd2s1 _28030_inst ( .DIN1(_28060), .DIN2(_28061), .Q(_28059) );
  nnd2s1 _28031_inst ( .DIN1(_28062), .DIN2(_28063), .Q(_28061) );
  nnd2s1 _28032_inst ( .DIN1(_28064), .DIN2(______[22]), .Q(_28063) );
  nor2s1 _28033_inst ( .DIN1(_28065), .DIN2(_28066), .Q(_28064) );
  xnr2s1 _28034_inst ( .DIN1(_53099), .DIN2(_28022), .Q(_28066) );
  nor2s1 _28035_inst ( .DIN1(_53045), .DIN2(_53463), .Q(_28022) );
  nnd2s1 _28036_inst ( .DIN1(_28067), .DIN2(_26282), .Q(_28062) );
  nnd2s1 _28037_inst ( .DIN1(_28068), .DIN2(_28069), .Q(_28058) );
  nor2s1 _28038_inst ( .DIN1(_26459), .DIN2(_28070), .Q(_28068) );
  nnd2s1 _28039_inst ( .DIN1(______[30]), .DIN2(_28071), .Q(_28070) );
  nnd2s1 _28040_inst ( .DIN1(_28072), .DIN2(_28073), .Q(
        __________________________________23_________) );
  nor2s1 _28041_inst ( .DIN1(_28074), .DIN2(_28075), .Q(_28072) );
  nor2s1 _28042_inst ( .DIN1(_27235), .DIN2(_28076), .Q(_28075) );
  nnd2s1 _28043_inst ( .DIN1(_28077), .DIN2(_28078), .Q(_28076) );
  nnd2s1 _28044_inst ( .DIN1(_53173), .DIN2(_28067), .Q(_28078) );
  nnd2s1 _28045_inst ( .DIN1(_28079), .DIN2(______[16]), .Q(_28077) );
  nor2s1 _28046_inst ( .DIN1(_28065), .DIN2(_28080), .Q(_28079) );
  xor2s1 _28047_inst ( .DIN1(_26435), .DIN2(_53481), .Q(_28080) );
  nor2s1 _28048_inst ( .DIN1(_27325), .DIN2(_28081), .Q(_28074) );
  xor2s1 _28049_inst ( .DIN1(_28082), .DIN2(_53454), .Q(_28081) );
  nor2s1 _28050_inst ( .DIN1(_28083), .DIN2(_28084), .Q(
        __________________________________22_________) );
  nor2s1 _28051_inst ( .DIN1(_28085), .DIN2(_28086), .Q(_28083) );
  xor2s1 _28052_inst ( .DIN1(_28087), .DIN2(_28088), .Q(_28086) );
  nnd2s1 _28053_inst ( .DIN1(_28052), .DIN2(_28089), .Q(_28087) );
  nnd2s1 _28054_inst ( .DIN1(_53481), .DIN2(_28055), .Q(_28089) );
  nor2s1 _28055_inst ( .DIN1(_28052), .DIN2(_26481), .Q(_28085) );
  nnd2s1 _28056_inst ( .DIN1(_28090), .DIN2(_28091), .Q(
        __________________________________21_________) );
  nor2s1 _28057_inst ( .DIN1(_28092), .DIN2(_28093), .Q(_28090) );
  nor2s1 _28058_inst ( .DIN1(_28094), .DIN2(_28095), .Q(_28093) );
  nor2s1 _28059_inst ( .DIN1(_28096), .DIN2(_28097), .Q(_28094) );
  nor2s1 _28060_inst ( .DIN1(_52846), .DIN2(_28065), .Q(_28097) );
  hi1s1 _28061_inst ( .DIN(_28055), .Q(_28065) );
  nor2s1 _28062_inst ( .DIN1(_28052), .DIN2(_26459), .Q(_28096) );
  nor2s1 _28063_inst ( .DIN1(_28098), .DIN2(_28099), .Q(_28092) );
  nor2s1 _28064_inst ( .DIN1(_26808), .DIN2(_28101), .Q(_28099) );
  xor2s1 _28065_inst ( .DIN1(_28102), .DIN2(_28103), .Q(_28101) );
  xor2s1 _28066_inst ( .DIN1(_53468), .DIN2(_53475), .Q(_28103) );
  nor2s1 _28067_inst ( .DIN1(_53481), .DIN2(_26592), .Q(_28102) );
  nnd2s1 _28068_inst ( .DIN1(_28104), .DIN2(_27644), .Q(
        __________________________________20_________) );
  nor2s1 _28069_inst ( .DIN1(_28105), .DIN2(_28106), .Q(_28104) );
  nor2s1 _28070_inst ( .DIN1(_28107), .DIN2(_27648), .Q(_28106) );
  nor2s1 _28071_inst ( .DIN1(_28108), .DIN2(_28109), .Q(_28107) );
  nor2s1 _28072_inst ( .DIN1(_52832), .DIN2(_28052), .Q(_28109) );
  hi1s1 _28073_inst ( .DIN(_28067), .Q(_28052) );
  nor2s1 _28074_inst ( .DIN1(_28055), .DIN2(_28110), .Q(_28067) );
  nor2s1 _28075_inst ( .DIN1(_28111), .DIN2(_28112), .Q(_28108) );
  nnd2s1 _28076_inst ( .DIN1(______[8]), .DIN2(_28055), .Q(_28112) );
  nnd2s1 _28077_inst ( .DIN1(_28113), .DIN2(_28114), .Q(_28055) );
  nor2s1 _28078_inst ( .DIN1(_28115), .DIN2(_28116), .Q(_28113) );
  xor2s1 _28079_inst ( .DIN1(_28117), .DIN2(_28118), .Q(_28111) );
  xor2s1 _28080_inst ( .DIN1(_53481), .DIN2(_53505), .Q(_28118) );
  nor2s1 _28081_inst ( .DIN1(_52846), .DIN2(_26435), .Q(_28117) );
  nor2s1 _28082_inst ( .DIN1(_27655), .DIN2(_28119), .Q(_28105) );
  nor2s1 _28083_inst ( .DIN1(_26291), .DIN2(_27291), .Q(_28119) );
  nnd2s1 _28084_inst ( .DIN1(_28120), .DIN2(_28121), .Q(
        __________________________________1_________) );
  nnd2s1 _28085_inst ( .DIN1(_28122), .DIN2(_28069), .Q(_28121) );
  nnd2s1 _28086_inst ( .DIN1(_28123), .DIN2(_28124), .Q(_28122) );
  xor2s1 _28087_inst ( .DIN1(_26391), .DIN2(_28125), .Q(_28124) );
  nnd2s1 _28088_inst ( .DIN1(_53150), .DIN2(_52844), .Q(_28125) );
  nnd2s1 _28089_inst ( .DIN1(_28126), .DIN2(_28060), .Q(_28120) );
  nor2s1 _28090_inst ( .DIN1(_28127), .DIN2(_28128), .Q(_28126) );
  nor2s1 _28091_inst ( .DIN1(_28129), .DIN2(_28130), .Q(_28128) );
  xor2s1 _28092_inst ( .DIN1(_28131), .DIN2(_28132), .Q(_28130) );
  xor2s1 _28093_inst ( .DIN1(_53509), .DIN2(_53512), .Q(_28132) );
  nnd2s1 _28094_inst ( .DIN1(_53506), .DIN2(_52844), .Q(_28131) );
  nor2s1 _28095_inst ( .DIN1(_53061), .DIN2(_28133), .Q(_28127) );
  nnd2s1 _28096_inst ( .DIN1(_28134), .DIN2(_28135), .Q(
        __________________________________19_________) );
  nnd2s1 _28097_inst ( .DIN1(_28136), .DIN2(_28137), .Q(_28135) );
  nnd2s1 _28098_inst ( .DIN1(_28138), .DIN2(______[6]), .Q(_28136) );
  and2s1 _28099_inst ( .DIN1(_28139), .DIN2(_53360), .Q(_28138) );
  nnd2s1 _28100_inst ( .DIN1(_28140), .DIN2(_27882), .Q(_28134) );
  nor2s1 _28101_inst ( .DIN1(_52905), .DIN2(_27888), .Q(_28140) );
  nnd2s1 _28102_inst ( .DIN1(_28141), .DIN2(_28142), .Q(
        __________________________________18_________) );
  nnd2s1 _28103_inst ( .DIN1(_28143), .DIN2(_28144), .Q(_28142) );
  nor2s1 _28104_inst ( .DIN1(_52911), .DIN2(_27888), .Q(_28143) );
  nnd2s1 _28105_inst ( .DIN1(_28145), .DIN2(_28146), .Q(_28141) );
  xor2s1 _28106_inst ( .DIN1(_53177), .DIN2(_53493), .Q(_28145) );
  nnd2s1 _28107_inst ( .DIN1(_28147), .DIN2(_28148), .Q(
        __________________________________17_________) );
  nor2s1 _28108_inst ( .DIN1(_28149), .DIN2(_28150), .Q(_28147) );
  nor2s1 _28109_inst ( .DIN1(_28151), .DIN2(_28152), .Q(_28150) );
  nnd2s1 _28110_inst ( .DIN1(_27889), .DIN2(_26571), .Q(_28152) );
  nor2s1 _28111_inst ( .DIN1(_28153), .DIN2(_28154), .Q(_28149) );
  xnr2s1 _28112_inst ( .DIN1(_27658), .DIN2(_52845), .Q(_28154) );
  nnd2s1 _28113_inst ( .DIN1(_28155), .DIN2(_28156), .Q(
        __________________________________16_________) );
  nnd2s1 _28114_inst ( .DIN1(_28153), .DIN2(_28157), .Q(_28156) );
  nnd2s1 _28115_inst ( .DIN1(_52988), .DIN2(_27889), .Q(_28157) );
  nnd2s1 _28116_inst ( .DIN1(_28158), .DIN2(_28151), .Q(_28155) );
  nor2s1 _28117_inst ( .DIN1(_28159), .DIN2(_28160), .Q(_28158) );
  xor2s1 _28118_inst ( .DIN1(_53142), .DIN2(_27658), .Q(_28160) );
  nor2s1 _28119_inst ( .DIN1(_26702), .DIN2(_26291), .Q(_27658) );
  nnd2s1 _28120_inst ( .DIN1(_28161), .DIN2(_26993), .Q(
        __________________________________15_________) );
  nor2s1 _28121_inst ( .DIN1(_28162), .DIN2(_28163), .Q(_28161) );
  nor2s1 _28122_inst ( .DIN1(_26996), .DIN2(_28164), .Q(_28163) );
  or2s1 _28123_inst ( .DIN1(_27888), .DIN2(_53122), .Q(_28164) );
  hi1s1 _28124_inst ( .DIN(_27889), .Q(_27888) );
  nor2s1 _28125_inst ( .DIN1(_27007), .DIN2(_28165), .Q(_28162) );
  xor2s1 _28126_inst ( .DIN1(_52967), .DIN2(_53329), .Q(_28165) );
  nnd2s1 _28127_inst ( .DIN1(_27994), .DIN2(_28166), .Q(
        __________________________________14_________) );
  nnd2s1 _28128_inst ( .DIN1(_27889), .DIN2(_53182), .Q(_28166) );
  nor2s1 _28129_inst ( .DIN1(_28167), .DIN2(_28168), .Q(_27889) );
  nnd2s1 _28130_inst ( .DIN1(_28169), .DIN2(_28170), .Q(_28167) );
  nnd2s1 _28131_inst ( .DIN1(_28171), .DIN2(_28172), .Q(
        __________________________________13_________) );
  nnd2s1 _28132_inst ( .DIN1(_28173), .DIN2(_28010), .Q(_28172) );
  nor2s1 _28133_inst ( .DIN1(_28174), .DIN2(_28175), .Q(_28173) );
  nor2s1 _28134_inst ( .DIN1(_26672), .DIN2(_27860), .Q(_28175) );
  nor2s1 _28135_inst ( .DIN1(_27864), .DIN2(_28176), .Q(_28174) );
  or2s1 _28136_inst ( .DIN1(_27862), .DIN2(_26611), .Q(_28176) );
  nnd2s1 _28137_inst ( .DIN1(______[6]), .DIN2(_28177), .Q(_27862) );
  nnd2s1 _28138_inst ( .DIN1(_28178), .DIN2(_53156), .Q(_28171) );
  nnd2s1 _28139_inst ( .DIN1(_28179), .DIN2(_28180), .Q(
        __________________________________12_________) );
  nnd2s1 _28140_inst ( .DIN1(_28181), .DIN2(_53177), .Q(_28180) );
  nor2s1 _28141_inst ( .DIN1(_28182), .DIN2(_27241), .Q(_28181) );
  nnd2s1 _28142_inst ( .DIN1(_28183), .DIN2(_28144), .Q(_28179) );
  nor2s1 _28143_inst ( .DIN1(_28184), .DIN2(_28185), .Q(_28183) );
  nor2s1 _28144_inst ( .DIN1(_27864), .DIN2(_28186), .Q(_28185) );
  nor2s1 _28145_inst ( .DIN1(_27873), .DIN2(_28187), .Q(_28186) );
  xor2s1 _28146_inst ( .DIN1(_28188), .DIN2(_28189), .Q(_28187) );
  xor2s1 _28147_inst ( .DIN1(_52847), .DIN2(_53488), .Q(_28189) );
  nor2s1 _28148_inst ( .DIN1(_53490), .DIN2(_52847), .Q(_28188) );
  nor2s1 _28149_inst ( .DIN1(_26395), .DIN2(_27860), .Q(_28184) );
  nnd2s1 _28150_inst ( .DIN1(_28190), .DIN2(_28191), .Q(
        __________________________________11_________) );
  nnd2s1 _28151_inst ( .DIN1(_28192), .DIN2(_27875), .Q(_28191) );
  nor2s1 _28152_inst ( .DIN1(_28193), .DIN2(_27393), .Q(_28192) );
  xor2s1 _28153_inst ( .DIN1(_52922), .DIN2(_26411), .Q(_28193) );
  nnd2s1 _28154_inst ( .DIN1(_28194), .DIN2(_27868), .Q(_28190) );
  xor2s1 _28155_inst ( .DIN1(_28195), .DIN2(_28196), .Q(_28194) );
  nor2s1 _28156_inst ( .DIN1(_28197), .DIN2(_28198), .Q(_28196) );
  nor2s1 _28157_inst ( .DIN1(_27864), .DIN2(_28199), .Q(_28198) );
  nor2s1 _28158_inst ( .DIN1(_28200), .DIN2(_28201), .Q(_28199) );
  nnd2s1 _28159_inst ( .DIN1(_28177), .DIN2(_27863), .Q(_28201) );
  nnd2s1 _28160_inst ( .DIN1(_52848), .DIN2(_53125), .Q(_27863) );
  nor2s1 _28161_inst ( .DIN1(_53125), .DIN2(_52848), .Q(_28200) );
  nor2s1 _28162_inst ( .DIN1(_52921), .DIN2(_27860), .Q(_28197) );
  nnd2s1 _28163_inst ( .DIN1(_28202), .DIN2(_27281), .Q(
        __________________________________10_________) );
  nor2s1 _28164_inst ( .DIN1(_28203), .DIN2(_28204), .Q(_28202) );
  nor2s1 _28165_inst ( .DIN1(_27284), .DIN2(_28205), .Q(_28204) );
  nor2s1 _28166_inst ( .DIN1(_28206), .DIN2(_28207), .Q(_28205) );
  and2s1 _28167_inst ( .DIN1(_52920), .DIN2(_27864), .Q(_28207) );
  nor2s1 _28168_inst ( .DIN1(_27864), .DIN2(_28208), .Q(_28206) );
  nnd2s1 _28169_inst ( .DIN1(_28209), .DIN2(_53125), .Q(_28208) );
  hi1s1 _28170_inst ( .DIN(_27860), .Q(_27864) );
  nnd2s1 _28171_inst ( .DIN1(_28210), .DIN2(_28211), .Q(_27860) );
  nor2s1 _28172_inst ( .DIN1(_28212), .DIN2(_28213), .Q(_28211) );
  nnd2s1 _28173_inst ( .DIN1(_28214), .DIN2(_28169), .Q(_28213) );
  nor2s1 _28174_inst ( .DIN1(_28215), .DIN2(_28110), .Q(_28210) );
  nor2s1 _28175_inst ( .DIN1(_27298), .DIN2(_28216), .Q(_28203) );
  nor2s1 _28176_inst ( .DIN1(_27774), .DIN2(_28217), .Q(_28216) );
  xor2s1 _28177_inst ( .DIN1(_52849), .DIN2(_53086), .Q(_28217) );
  nor2s1 _28178_inst ( .DIN1(_28218), .DIN2(_28219), .Q(
        __________________________________0_________) );
  nor2s1 _28179_inst ( .DIN1(_28220), .DIN2(_28221), .Q(_28219) );
  nor2s1 _28180_inst ( .DIN1(_52925), .DIN2(_28133), .Q(_28221) );
  nor2s1 _28181_inst ( .DIN1(_27291), .DIN2(_28222), .Q(_28220) );
  nnd2s1 _28182_inst ( .DIN1(_52844), .DIN2(_28223), .Q(_28222) );
  nnd2s1 _28183_inst ( .DIN1(_28224), .DIN2(_28225), .Q(
        _________________________________9_________) );
  nnd2s1 _28184_inst ( .DIN1(_28226), .DIN2(_26313), .Q(_28225) );
  nor2s1 _28185_inst ( .DIN1(_28227), .DIN2(_28228), .Q(_28224) );
  nor2s1 _28186_inst ( .DIN1(_28229), .DIN2(_28230), .Q(_28228) );
  nor2s1 _28187_inst ( .DIN1(_28231), .DIN2(_28232), .Q(_28229) );
  nnd2s1 _28188_inst ( .DIN1(______[8]), .DIN2(_28233), .Q(_28232) );
  xor2s1 _28189_inst ( .DIN1(_53492), .DIN2(_53494), .Q(_28231) );
  nor2s1 _28190_inst ( .DIN1(_28234), .DIN2(_28235), .Q(_28227) );
  nnd2s1 _28191_inst ( .DIN1(______[2]), .DIN2(_28236), .Q(_28235) );
  xor2s1 _28192_inst ( .DIN1(_53495), .DIN2(_53514), .Q(_28236) );
  nnd2s1 _28193_inst ( .DIN1(_28237), .DIN2(_28238), .Q(
        _________________________________8_________) );
  nor2s1 _28194_inst ( .DIN1(_28239), .DIN2(_28240), .Q(_28237) );
  nor2s1 _28195_inst ( .DIN1(_28241), .DIN2(_28242), .Q(_28240) );
  nor2s1 _28196_inst ( .DIN1(_28243), .DIN2(_28244), .Q(_28242) );
  nor2s1 _28197_inst ( .DIN1(_28245), .DIN2(_28246), .Q(_28244) );
  nor2s1 _28198_inst ( .DIN1(_28247), .DIN2(_28248), .Q(_28246) );
  nor2s1 _28199_inst ( .DIN1(_53057), .DIN2(_53498), .Q(_28247) );
  nor2s1 _28200_inst ( .DIN1(_53085), .DIN2(_28249), .Q(_28243) );
  nor2s1 _28201_inst ( .DIN1(_28250), .DIN2(_28251), .Q(_28239) );
  nor2s1 _28202_inst ( .DIN1(_27614), .DIN2(_26668), .Q(_28251) );
  nnd2s1 _28203_inst ( .DIN1(_28252), .DIN2(_28253), .Q(
        _________________________________7_________) );
  nor2s1 _28204_inst ( .DIN1(_28254), .DIN2(_28255), .Q(_28252) );
  nor2s1 _28205_inst ( .DIN1(_28249), .DIN2(_28256), .Q(_28255) );
  xor2s1 _28206_inst ( .DIN1(_27346), .DIN2(_53079), .Q(_28256) );
  nor2s1 _28207_inst ( .DIN1(_28245), .DIN2(_28257), .Q(_28254) );
  nnd2s1 _28208_inst ( .DIN1(_28258), .DIN2(_28233), .Q(_28257) );
  xor2s1 _28209_inst ( .DIN1(_27346), .DIN2(_53498), .Q(_28258) );
  nor2s1 _28210_inst ( .DIN1(_27593), .DIN2(_28259), .Q(
        _________________________________6_________) );
  nnd2s1 _28211_inst ( .DIN1(_28260), .DIN2(_28261), .Q(_28259) );
  or2s1 _28212_inst ( .DIN1(_28249), .DIN2(_53086), .Q(_28261) );
  nnd2s1 _28213_inst ( .DIN1(_28262), .DIN2(_28249), .Q(_28260) );
  nnd2s1 _28214_inst ( .DIN1(_28263), .DIN2(______[20]), .Q(_28262) );
  nor2s1 _28215_inst ( .DIN1(_28264), .DIN2(_28265), .Q(_28263) );
  nor2s1 _28216_inst ( .DIN1(_53514), .DIN2(_28266), .Q(_28265) );
  and2s1 _28217_inst ( .DIN1(_28233), .DIN2(_28267), .Q(_28266) );
  and2s1 _28218_inst ( .DIN1(_28248), .DIN2(_53514), .Q(_28264) );
  nnd2s1 _28219_inst ( .DIN1(_28268), .DIN2(_28269), .Q(
        _________________________________5_________) );
  nnd2s1 _28220_inst ( .DIN1(_28226), .DIN2(_26256), .Q(_28269) );
  hi1s1 _28221_inst ( .DIN(_28270), .Q(_28226) );
  nor2s1 _28222_inst ( .DIN1(_28271), .DIN2(_28272), .Q(_28268) );
  nor2s1 _28223_inst ( .DIN1(_28273), .DIN2(_28274), .Q(_28272) );
  nnd2s1 _28224_inst ( .DIN1(_28275), .DIN2(______[6]), .Q(_28274) );
  xor2s1 _28225_inst ( .DIN1(_26598), .DIN2(_28276), .Q(_28273) );
  nnd2s1 _28226_inst ( .DIN1(_53495), .DIN2(_53496), .Q(_28276) );
  nor2s1 _28227_inst ( .DIN1(_28277), .DIN2(_28278), .Q(_28271) );
  or2s1 _28228_inst ( .DIN1(_28230), .DIN2(_26772), .Q(_28278) );
  nnd2s1 _28229_inst ( .DIN1(_28279), .DIN2(_28280), .Q(_28277) );
  nnd2s1 _28230_inst ( .DIN1(_52850), .DIN2(_28248), .Q(_28280) );
  nnd2s1 _28231_inst ( .DIN1(_28233), .DIN2(_28281), .Q(_28248) );
  nnd2s1 _28232_inst ( .DIN1(_28282), .DIN2(_26747), .Q(_28279) );
  nnd2s1 _28233_inst ( .DIN1(_28267), .DIN2(_28233), .Q(_28282) );
  hi1s1 _28234_inst ( .DIN(_28281), .Q(_28267) );
  nnd2s1 _28235_inst ( .DIN1(_53057), .DIN2(_53498), .Q(_28281) );
  nnd2s1 _28236_inst ( .DIN1(_28283), .DIN2(_28284), .Q(
        _________________________________4_________) );
  nor2s1 _28237_inst ( .DIN1(_28285), .DIN2(_28286), .Q(_28283) );
  nor2s1 _28238_inst ( .DIN1(_27144), .DIN2(_28287), .Q(_28286) );
  nnd2s1 _28239_inst ( .DIN1(_28288), .DIN2(_28289), .Q(_28287) );
  nor2s1 _28240_inst ( .DIN1(_28290), .DIN2(_28291), .Q(_28288) );
  nor2s1 _28241_inst ( .DIN1(_28292), .DIN2(_26355), .Q(_28291) );
  nor2s1 _28242_inst ( .DIN1(_28293), .DIN2(_28294), .Q(_28290) );
  xor2s1 _28243_inst ( .DIN1(_26727), .DIN2(_53510), .Q(_28294) );
  nor2s1 _28244_inst ( .DIN1(_27146), .DIN2(_28295), .Q(_28285) );
  xor2s1 _28245_inst ( .DIN1(_28296), .DIN2(_26441), .Q(_28295) );
  nnd2s1 _28246_inst ( .DIN1(_28297), .DIN2(_28298), .Q(
        _________________________________3_________) );
  nor2s1 _28247_inst ( .DIN1(_28299), .DIN2(_28300), .Q(_28297) );
  nor2s1 _28248_inst ( .DIN1(_28301), .DIN2(_28302), .Q(_28300) );
  nor2s1 _28249_inst ( .DIN1(_28303), .DIN2(_28304), .Q(_28301) );
  nnd2s1 _28250_inst ( .DIN1(_28305), .DIN2(_28306), .Q(_28304) );
  nnd2s1 _28251_inst ( .DIN1(_28293), .DIN2(_26239), .Q(_28306) );
  nnd2s1 _28252_inst ( .DIN1(_28307), .DIN2(_28292), .Q(_28305) );
  nnd2s1 _28253_inst ( .DIN1(______[20]), .DIN2(_53134), .Q(_28307) );
  nor2s1 _28254_inst ( .DIN1(_28308), .DIN2(_26464), .Q(_28299) );
  nnd2s1 _28255_inst ( .DIN1(_28309), .DIN2(_28310), .Q(
        _________________________________31_________) );
  nor2s1 _28256_inst ( .DIN1(_28311), .DIN2(_28312), .Q(_28309) );
  nor2s1 _28257_inst ( .DIN1(_28313), .DIN2(_28314), .Q(_28312) );
  nnd2s1 _28258_inst ( .DIN1(_28315), .DIN2(_28316), .Q(_28314) );
  nnd2s1 _28259_inst ( .DIN1(_53137), .DIN2(_28317), .Q(_28316) );
  nnd2s1 _28260_inst ( .DIN1(_28318), .DIN2(_28319), .Q(_28315) );
  xor2s1 _28261_inst ( .DIN1(_28320), .DIN2(_26596), .Q(_28319) );
  nor2s1 _28262_inst ( .DIN1(_28321), .DIN2(_28100), .Q(_28318) );
  nor2s1 _28263_inst ( .DIN1(_28322), .DIN2(_28323), .Q(_28311) );
  xor2s1 _28264_inst ( .DIN1(_26319), .DIN2(_28324), .Q(_28323) );
  nnd2s1 _28265_inst ( .DIN1(_28325), .DIN2(_28326), .Q(
        _________________________________30_________) );
  nor2s1 _28266_inst ( .DIN1(_28327), .DIN2(_28328), .Q(_28325) );
  nor2s1 _28267_inst ( .DIN1(_28329), .DIN2(_28330), .Q(_28328) );
  nor2s1 _28268_inst ( .DIN1(_28331), .DIN2(_28332), .Q(_28330) );
  nor2s1 _28269_inst ( .DIN1(_28333), .DIN2(_28334), .Q(_28332) );
  nor2s1 _28270_inst ( .DIN1(_26855), .DIN2(_28335), .Q(_28334) );
  or2s1 _28271_inst ( .DIN1(_28336), .DIN2(_52971), .Q(_28335) );
  nor2s1 _28272_inst ( .DIN1(_53062), .DIN2(_28337), .Q(_28331) );
  nor2s1 _28273_inst ( .DIN1(_53483), .DIN2(_28338), .Q(_28327) );
  nnd2s1 _28274_inst ( .DIN1(_28339), .DIN2(_28340), .Q(
        _________________________________2_________) );
  nnd2s1 _28275_inst ( .DIN1(_28341), .DIN2(_28342), .Q(_28340) );
  nor2s1 _28276_inst ( .DIN1(_28343), .DIN2(_28344), .Q(_28341) );
  nor2s1 _28277_inst ( .DIN1(_28293), .DIN2(_28345), .Q(_28344) );
  nor2s1 _28278_inst ( .DIN1(_53511), .DIN2(_26988), .Q(_28345) );
  nor2s1 _28279_inst ( .DIN1(_28292), .DIN2(_26677), .Q(_28343) );
  nnd2s1 _28280_inst ( .DIN1(_28346), .DIN2(_28347), .Q(_28339) );
  nnd2s1 _28281_inst ( .DIN1(_28348), .DIN2(_28349), .Q(_28346) );
  and2s1 _28282_inst ( .DIN1(_28350), .DIN2(_28351), .Q(_28349) );
  nor2s1 _28283_inst ( .DIN1(_28352), .DIN2(_26773), .Q(_28348) );
  nor2s1 _28284_inst ( .DIN1(_53135), .DIN2(_53511), .Q(_28352) );
  nnd2s1 _28285_inst ( .DIN1(_28353), .DIN2(_28354), .Q(
        _________________________________29_________) );
  nnd2s1 _28286_inst ( .DIN1(_28355), .DIN2(_28356), .Q(_28354) );
  nor2s1 _28287_inst ( .DIN1(_28357), .DIN2(_28358), .Q(_28355) );
  nor2s1 _28288_inst ( .DIN1(_28333), .DIN2(_28359), .Q(_28358) );
  nor2s1 _28289_inst ( .DIN1(_28336), .DIN2(_28360), .Q(_28359) );
  xor2s1 _28290_inst ( .DIN1(_28361), .DIN2(_28362), .Q(_28360) );
  xor2s1 _28291_inst ( .DIN1(_52851), .DIN2(_53366), .Q(_28362) );
  nor2s1 _28292_inst ( .DIN1(_52971), .DIN2(_26242), .Q(_28361) );
  nor2s1 _28293_inst ( .DIN1(_53060), .DIN2(_28337), .Q(_28357) );
  nnd2s1 _28294_inst ( .DIN1(_28363), .DIN2(_28364), .Q(_28353) );
  xor2s1 _28295_inst ( .DIN1(_53278), .DIN2(_53279), .Q(_28363) );
  nnd2s1 _28296_inst ( .DIN1(_28365), .DIN2(_28366), .Q(
        _________________________________28_________) );
  nnd2s1 _28297_inst ( .DIN1(_27672), .DIN2(_28367), .Q(_28366) );
  nnd2s1 _28298_inst ( .DIN1(_28368), .DIN2(_28369), .Q(_28367) );
  nor2s1 _28299_inst ( .DIN1(_28370), .DIN2(_28371), .Q(_28368) );
  nor2s1 _28300_inst ( .DIN1(_28372), .DIN2(_28373), .Q(_28371) );
  nor2s1 _28301_inst ( .DIN1(_28374), .DIN2(_28100), .Q(_28373) );
  nor2s1 _28302_inst ( .DIN1(_53059), .DIN2(_28375), .Q(_28370) );
  nnd2s1 _28303_inst ( .DIN1(_28376), .DIN2(_27663), .Q(_28365) );
  nor2s1 _28304_inst ( .DIN1(_28377), .DIN2(_28378), .Q(_28376) );
  nnd2s1 _28305_inst ( .DIN1(_28379), .DIN2(_27815), .Q(_28378) );
  nnd2s1 _28306_inst ( .DIN1(_28380), .DIN2(_28381), .Q(_28379) );
  nor2s1 _28307_inst ( .DIN1(_53155), .DIN2(_53157), .Q(_28377) );
  nnd2s1 _28308_inst ( .DIN1(_28382), .DIN2(_28383), .Q(
        _________________________________27_________) );
  nor2s1 _28309_inst ( .DIN1(_28384), .DIN2(_28385), .Q(_28383) );
  nor2s1 _28310_inst ( .DIN1(_28386), .DIN2(_28387), .Q(_28385) );
  or2s1 _28311_inst ( .DIN1(_28388), .DIN2(_26809), .Q(_28387) );
  nnd2s1 _28312_inst ( .DIN1(_53176), .DIN2(_28389), .Q(_28386) );
  nor2s1 _28313_inst ( .DIN1(_28390), .DIN2(_28391), .Q(_28382) );
  nor2s1 _28314_inst ( .DIN1(_28392), .DIN2(_26623), .Q(_28391) );
  nor2s1 _28315_inst ( .DIN1(_28322), .DIN2(_28393), .Q(_28390) );
  nor2s1 _28316_inst ( .DIN1(_28394), .DIN2(_27241), .Q(_28393) );
  xor2s1 _28317_inst ( .DIN1(_28395), .DIN2(_52978), .Q(_28394) );
  nnd2s1 _28318_inst ( .DIN1(_52852), .DIN2(_52980), .Q(_28395) );
  nnd2s1 _28319_inst ( .DIN1(_28396), .DIN2(_28397), .Q(
        _________________________________26_________) );
  nnd2s1 _28320_inst ( .DIN1(_28398), .DIN2(_28399), .Q(_28397) );
  nor2s1 _28321_inst ( .DIN1(_28400), .DIN2(_28401), .Q(_28398) );
  nor2s1 _28322_inst ( .DIN1(_28374), .DIN2(_26604), .Q(_28401) );
  nor2s1 _28323_inst ( .DIN1(_52852), .DIN2(_52978), .Q(_28374) );
  nor2s1 _28324_inst ( .DIN1(_52978), .DIN2(_53176), .Q(_28400) );
  nor2s1 _28325_inst ( .DIN1(_28402), .DIN2(_28403), .Q(_28396) );
  nor2s1 _28326_inst ( .DIN1(_28404), .DIN2(_28405), .Q(_28403) );
  nor2s1 _28327_inst ( .DIN1(_28406), .DIN2(_28407), .Q(_28404) );
  hi1s1 _28328_inst ( .DIN(_28369), .Q(_28407) );
  nnd2s1 _28329_inst ( .DIN1(_28408), .DIN2(_28375), .Q(_28369) );
  nnd2s1 _28330_inst ( .DIN1(_28389), .DIN2(_28409), .Q(_28408) );
  nnd2s1 _28331_inst ( .DIN1(_52852), .DIN2(_52978), .Q(_28409) );
  nor2s1 _28332_inst ( .DIN1(_28375), .DIN2(_26540), .Q(_28406) );
  nor2s1 _28333_inst ( .DIN1(_28144), .DIN2(_28410), .Q(_28402) );
  nor2s1 _28334_inst ( .DIN1(_28411), .DIN2(_28412), .Q(_28410) );
  xor2s1 _28335_inst ( .DIN1(_26680), .DIN2(_28413), .Q(_28412) );
  nnd2s1 _28336_inst ( .DIN1(_28414), .DIN2(_28415), .Q(
        _________________________________25_________) );
  nor2s1 _28337_inst ( .DIN1(_28416), .DIN2(_28417), .Q(_28415) );
  nor2s1 _28338_inst ( .DIN1(_28418), .DIN2(_28419), .Q(_28417) );
  nnd2s1 _28339_inst ( .DIN1(______[18]), .DIN2(_52980), .Q(_28419) );
  nnd2s1 _28340_inst ( .DIN1(_28420), .DIN2(_28313), .Q(_28418) );
  nor2s1 _28341_inst ( .DIN1(_28421), .DIN2(_28422), .Q(_28414) );
  nor2s1 _28342_inst ( .DIN1(_53063), .DIN2(_28392), .Q(_28422) );
  nor2s1 _28343_inst ( .DIN1(_28423), .DIN2(_28388), .Q(_28421) );
  nor2s1 _28344_inst ( .DIN1(_27039), .DIN2(_28424), .Q(_28423) );
  xor2s1 _28345_inst ( .DIN1(_52852), .DIN2(_52972), .Q(_28424) );
  nnd2s1 _28346_inst ( .DIN1(_28425), .DIN2(_28426), .Q(
        _________________________________24_________) );
  nor2s1 _28347_inst ( .DIN1(_28427), .DIN2(_28428), .Q(_28426) );
  or2s1 _28348_inst ( .DIN1(_28416), .DIN2(_28384), .Q(_28428) );
  nor2s1 _28349_inst ( .DIN1(_28388), .DIN2(_28389), .Q(_28416) );
  nor2s1 _28350_inst ( .DIN1(_28322), .DIN2(_28429), .Q(_28427) );
  nor2s1 _28351_inst ( .DIN1(_26314), .DIN2(_26987), .Q(_28429) );
  nor2s1 _28352_inst ( .DIN1(_28430), .DIN2(_28431), .Q(_28425) );
  nor2s1 _28353_inst ( .DIN1(_53068), .DIN2(_28392), .Q(_28431) );
  nnd2s1 _28354_inst ( .DIN1(_28372), .DIN2(_28322), .Q(_28392) );
  nor2s1 _28355_inst ( .DIN1(_28432), .DIN2(_28388), .Q(_28430) );
  nnd2s1 _28356_inst ( .DIN1(_28322), .DIN2(_28375), .Q(_28388) );
  nor2s1 _28357_inst ( .DIN1(_28433), .DIN2(_26773), .Q(_28432) );
  xor2s1 _28358_inst ( .DIN1(_26477), .DIN2(_53184), .Q(_28433) );
  nnd2s1 _28359_inst ( .DIN1(_28434), .DIN2(_28435), .Q(
        _________________________________23_________) );
  nnd2s1 _28360_inst ( .DIN1(_28399), .DIN2(_28436), .Q(_28435) );
  nnd2s1 _28361_inst ( .DIN1(_28437), .DIN2(______[0]), .Q(_28436) );
  and2s1 _28362_inst ( .DIN1(_28389), .DIN2(_53184), .Q(_28437) );
  nor2s1 _28363_inst ( .DIN1(_28405), .DIN2(_28372), .Q(_28399) );
  nor2s1 _28364_inst ( .DIN1(_28438), .DIN2(_28439), .Q(_28434) );
  nor2s1 _28365_inst ( .DIN1(_28405), .DIN2(_28440), .Q(_28439) );
  nnd2s1 _28366_inst ( .DIN1(_53065), .DIN2(_28372), .Q(_28440) );
  hi1s1 _28367_inst ( .DIN(_28375), .Q(_28372) );
  nnd2s1 _28368_inst ( .DIN1(_28441), .DIN2(_28442), .Q(_28375) );
  nor2s1 _28369_inst ( .DIN1(_28144), .DIN2(_28443), .Q(_28438) );
  nor2s1 _28370_inst ( .DIN1(_28182), .DIN2(_26514), .Q(_28443) );
  nnd2s1 _28371_inst ( .DIN1(_28444), .DIN2(_28445), .Q(
        _________________________________22_________) );
  nor2s1 _28372_inst ( .DIN1(_28446), .DIN2(_28447), .Q(_28444) );
  nor2s1 _28373_inst ( .DIN1(_27845), .DIN2(_28448), .Q(_28447) );
  nnd2s1 _28374_inst ( .DIN1(_28449), .DIN2(_28450), .Q(_28448) );
  or2s1 _28375_inst ( .DIN1(_28451), .DIN2(_53482), .Q(_28450) );
  nnd2s1 _28376_inst ( .DIN1(_53083), .DIN2(_28452), .Q(_28449) );
  nor2s1 _28377_inst ( .DIN1(_27836), .DIN2(_28453), .Q(_28446) );
  nor2s1 _28378_inst ( .DIN1(_28454), .DIN2(_27365), .Q(_28453) );
  xor2s1 _28379_inst ( .DIN1(_27851), .DIN2(_28455), .Q(_28454) );
  xor2s1 _28380_inst ( .DIN1(_53067), .DIN2(_53186), .Q(_28455) );
  nnd2s1 _28381_inst ( .DIN1(_53280), .DIN2(_53186), .Q(_27851) );
  nnd2s1 _28382_inst ( .DIN1(_28456), .DIN2(_28457), .Q(
        _________________________________21_________) );
  nnd2s1 _28383_inst ( .DIN1(_28458), .DIN2(_28452), .Q(_28457) );
  nor2s1 _28384_inst ( .DIN1(_53179), .DIN2(_28084), .Q(_28458) );
  nnd2s1 _28385_inst ( .DIN1(_28459), .DIN2(_28460), .Q(_28456) );
  nor2s1 _28386_inst ( .DIN1(_28461), .DIN2(_27241), .Q(_28460) );
  xor2s1 _28387_inst ( .DIN1(_28462), .DIN2(_28463), .Q(_28461) );
  xor2s1 _28388_inst ( .DIN1(_52980), .DIN2(_53184), .Q(_28463) );
  nnd2s1 _28389_inst ( .DIN1(_53504), .DIN2(_26457), .Q(_28462) );
  nor2s1 _28390_inst ( .DIN1(_28084), .DIN2(_28451), .Q(_28459) );
  nnd2s1 _28391_inst ( .DIN1(_28464), .DIN2(_28465), .Q(
        _________________________________20_________) );
  nnd2s1 _28392_inst ( .DIN1(_28466), .DIN2(_28467), .Q(_28465) );
  nnd2s1 _28393_inst ( .DIN1(_28468), .DIN2(_28146), .Q(_28466) );
  xor2s1 _28394_inst ( .DIN1(_26393), .DIN2(_28469), .Q(_28468) );
  nnd2s1 _28395_inst ( .DIN1(_52851), .DIN2(_53483), .Q(_28469) );
  nnd2s1 _28396_inst ( .DIN1(_28470), .DIN2(_28471), .Q(_28464) );
  nnd2s1 _28397_inst ( .DIN1(_28472), .DIN2(_28473), .Q(_28471) );
  nnd2s1 _28398_inst ( .DIN1(_28474), .DIN2(_28475), .Q(_28473) );
  nor2s1 _28399_inst ( .DIN1(_28476), .DIN2(_28477), .Q(_28474) );
  nor2s1 _28400_inst ( .DIN1(_53484), .DIN2(_26507), .Q(_28477) );
  or2s1 _28401_inst ( .DIN1(_28478), .DIN2(_53077), .Q(_28472) );
  nnd2s1 _28402_inst ( .DIN1(_28479), .DIN2(_28480), .Q(
        _________________________________1_________) );
  nnd2s1 _28403_inst ( .DIN1(_28481), .DIN2(_28342), .Q(_28480) );
  nor2s1 _28404_inst ( .DIN1(_28347), .DIN2(_28303), .Q(_28342) );
  nor2s1 _28405_inst ( .DIN1(_28482), .DIN2(_28483), .Q(_28481) );
  nor2s1 _28406_inst ( .DIN1(_28293), .DIN2(_28484), .Q(_28483) );
  xor2s1 _28407_inst ( .DIN1(_28485), .DIN2(_28486), .Q(_28484) );
  xor2s1 _28408_inst ( .DIN1(_53134), .DIN2(_53508), .Q(_28486) );
  nor2s1 _28409_inst ( .DIN1(_53511), .DIN2(_53510), .Q(_28485) );
  nor2s1 _28410_inst ( .DIN1(_28292), .DIN2(_26701), .Q(_28482) );
  nnd2s1 _28411_inst ( .DIN1(_28487), .DIN2(_28347), .Q(_28479) );
  nnd2s1 _28412_inst ( .DIN1(_28488), .DIN2(______[20]), .Q(_28487) );
  and2s1 _28413_inst ( .DIN1(_28350), .DIN2(_53135), .Q(_28488) );
  nnd2s1 _28414_inst ( .DIN1(_28489), .DIN2(_28490), .Q(
        _________________________________19_________) );
  nnd2s1 _28415_inst ( .DIN1(_28491), .DIN2(_28467), .Q(_28490) );
  nnd2s1 _28416_inst ( .DIN1(_28492), .DIN2(_28493), .Q(_28491) );
  xor2s1 _28417_inst ( .DIN1(_52851), .DIN2(_52897), .Q(_28493) );
  hi1s1 _28418_inst ( .DIN(_28411), .Q(_28492) );
  nnd2s1 _28419_inst ( .DIN1(______[28]), .DIN2(_28146), .Q(_28411) );
  nnd2s1 _28420_inst ( .DIN1(_28494), .DIN2(_28470), .Q(_28489) );
  nor2s1 _28421_inst ( .DIN1(_28495), .DIN2(_28496), .Q(_28494) );
  nor2s1 _28422_inst ( .DIN1(_28451), .DIN2(_28497), .Q(_28496) );
  nnd2s1 _28423_inst ( .DIN1(______[30]), .DIN2(_26507), .Q(_28497) );
  nor2s1 _28424_inst ( .DIN1(_28478), .DIN2(_26432), .Q(_28495) );
  nnd2s1 _28425_inst ( .DIN1(_28498), .DIN2(_28073), .Q(
        _________________________________18_________) );
  nor2s1 _28426_inst ( .DIN1(_28499), .DIN2(_28500), .Q(_28498) );
  nor2s1 _28427_inst ( .DIN1(_27325), .DIN2(_28501), .Q(_28500) );
  xor2s1 _28428_inst ( .DIN1(_28502), .DIN2(_26346), .Q(_28501) );
  nor2s1 _28429_inst ( .DIN1(_28503), .DIN2(_27235), .Q(_28499) );
  nor2s1 _28430_inst ( .DIN1(_28504), .DIN2(_28505), .Q(_28503) );
  and2s1 _28431_inst ( .DIN1(_28452), .DIN2(_53082), .Q(_28505) );
  nor2s1 _28432_inst ( .DIN1(_28506), .DIN2(_28507), .Q(_28504) );
  nnd2s1 _28433_inst ( .DIN1(______[30]), .DIN2(_28508), .Q(_28507) );
  xor2s1 _28434_inst ( .DIN1(_53486), .DIN2(_28476), .Q(_28508) );
  nnd2s1 _28435_inst ( .DIN1(_28509), .DIN2(_28510), .Q(
        _________________________________17_________) );
  nnd2s1 _28436_inst ( .DIN1(_28511), .DIN2(_28313), .Q(_28510) );
  nnd2s1 _28437_inst ( .DIN1(______[28]), .DIN2(_28512), .Q(_28511) );
  xor2s1 _28438_inst ( .DIN1(_28513), .DIN2(_28514), .Q(_28512) );
  xor2s1 _28439_inst ( .DIN1(_52852), .DIN2(_52980), .Q(_28514) );
  and2s1 _28440_inst ( .DIN1(_52980), .DIN2(_52978), .Q(_28513) );
  nor2s1 _28441_inst ( .DIN1(_28384), .DIN2(_28515), .Q(_28509) );
  nor2s1 _28442_inst ( .DIN1(_28516), .DIN2(_28517), .Q(_28515) );
  nor2s1 _28443_inst ( .DIN1(_28518), .DIN2(_26773), .Q(_28517) );
  nor2s1 _28444_inst ( .DIN1(_28519), .DIN2(_28313), .Q(_28518) );
  nor2s1 _28445_inst ( .DIN1(_28451), .DIN2(_28520), .Q(_28519) );
  xor2s1 _28446_inst ( .DIN1(_53483), .DIN2(_28476), .Q(_28520) );
  nor2s1 _28447_inst ( .DIN1(_26393), .DIN2(_53461), .Q(_28476) );
  xor2s1 _28448_inst ( .DIN1(_28506), .DIN2(_28521), .Q(_28451) );
  hi1s1 _28449_inst ( .DIN(_28475), .Q(_28506) );
  nor2s1 _28450_inst ( .DIN1(_28522), .DIN2(_28452), .Q(_28475) );
  hi1s1 _28451_inst ( .DIN(_28478), .Q(_28452) );
  nor2s1 _28452_inst ( .DIN1(_28478), .DIN2(_26556), .Q(_28516) );
  nnd2s1 _28453_inst ( .DIN1(_28523), .DIN2(_28524), .Q(_28478) );
  nor2s1 _28454_inst ( .DIN1(_28525), .DIN2(_28526), .Q(_28524) );
  nor2s1 _28455_inst ( .DIN1(_28527), .DIN2(_28528), .Q(_28523) );
  nnd2s1 _28456_inst ( .DIN1(_28529), .DIN2(_28530), .Q(
        _________________________________16_________) );
  nor2s1 _28457_inst ( .DIN1(_28531), .DIN2(_28532), .Q(_28529) );
  nor2s1 _28458_inst ( .DIN1(_28533), .DIN2(_28534), .Q(_28532) );
  nor2s1 _28459_inst ( .DIN1(_28535), .DIN2(_28536), .Q(_28534) );
  nor2s1 _28460_inst ( .DIN1(_28537), .DIN2(_28538), .Q(_28536) );
  nor2s1 _28461_inst ( .DIN1(_28539), .DIN2(_28540), .Q(_28538) );
  nor2s1 _28462_inst ( .DIN1(_53489), .DIN2(_26546), .Q(_28539) );
  nor2s1 _28463_inst ( .DIN1(_28541), .DIN2(_26708), .Q(_28535) );
  nor2s1 _28464_inst ( .DIN1(_28542), .DIN2(_28543), .Q(_28531) );
  nor2s1 _28465_inst ( .DIN1(_26808), .DIN2(_28544), .Q(_28543) );
  xor2s1 _28466_inst ( .DIN1(_53443), .DIN2(_28545), .Q(_28544) );
  nnd2s1 _28467_inst ( .DIN1(_28546), .DIN2(_28298), .Q(
        _________________________________15_________) );
  nor2s1 _28468_inst ( .DIN1(_28547), .DIN2(_28548), .Q(_28546) );
  nor2s1 _28469_inst ( .DIN1(_28308), .DIN2(_28549), .Q(_28548) );
  xor2s1 _28470_inst ( .DIN1(_53220), .DIN2(_53510), .Q(_28549) );
  nor2s1 _28471_inst ( .DIN1(_28550), .DIN2(_28302), .Q(_28547) );
  nor2s1 _28472_inst ( .DIN1(_28551), .DIN2(_28552), .Q(_28550) );
  nnd2s1 _28473_inst ( .DIN1(_28553), .DIN2(_28554), .Q(_28552) );
  nnd2s1 _28474_inst ( .DIN1(_28537), .DIN2(_53078), .Q(_28554) );
  nnd2s1 _28475_inst ( .DIN1(_28555), .DIN2(_28541), .Q(_28553) );
  nnd2s1 _28476_inst ( .DIN1(______[24]), .DIN2(_53491), .Q(_28555) );
  nnd2s1 _28477_inst ( .DIN1(_28556), .DIN2(_27723), .Q(
        _________________________________14_________) );
  nor2s1 _28478_inst ( .DIN1(_28557), .DIN2(_28558), .Q(_28556) );
  nor2s1 _28479_inst ( .DIN1(_28537), .DIN2(_28559), .Q(_28558) );
  nnd2s1 _28480_inst ( .DIN1(_28560), .DIN2(_28561), .Q(_28559) );
  nor2s1 _28481_inst ( .DIN1(_28562), .DIN2(_28563), .Q(_28561) );
  nor2s1 _28482_inst ( .DIN1(_26546), .DIN2(_28564), .Q(_28563) );
  nnd2s1 _28483_inst ( .DIN1(_53491), .DIN2(_26464), .Q(_28564) );
  nor2s1 _28484_inst ( .DIN1(_52999), .DIN2(_53491), .Q(_28562) );
  hi1s1 _28485_inst ( .DIN(_28540), .Q(_28560) );
  nnd2s1 _28486_inst ( .DIN1(_28565), .DIN2(_28566), .Q(_28540) );
  nnd2s1 _28487_inst ( .DIN1(_28522), .DIN2(_28567), .Q(_28566) );
  nnd2s1 _28488_inst ( .DIN1(_53489), .DIN2(_26546), .Q(_28565) );
  nor2s1 _28489_inst ( .DIN1(_53074), .DIN2(_28541), .Q(_28557) );
  nnd2s1 _28490_inst ( .DIN1(_28568), .DIN2(_28569), .Q(
        _________________________________13_________) );
  nor2s1 _28491_inst ( .DIN1(_28570), .DIN2(_28571), .Q(_28568) );
  nor2s1 _28492_inst ( .DIN1(_28572), .DIN2(_28573), .Q(_28571) );
  xor2s1 _28493_inst ( .DIN1(_53018), .DIN2(_53138), .Q(_28573) );
  nor2s1 _28494_inst ( .DIN1(_28574), .DIN2(_28575), .Q(_28570) );
  nor2s1 _28495_inst ( .DIN1(_28551), .DIN2(_28576), .Q(_28574) );
  nnd2s1 _28496_inst ( .DIN1(_28577), .DIN2(_28578), .Q(_28576) );
  nnd2s1 _28497_inst ( .DIN1(_28537), .DIN2(_26631), .Q(_28578) );
  nnd2s1 _28498_inst ( .DIN1(_28579), .DIN2(_28541), .Q(_28577) );
  xor2s1 _28499_inst ( .DIN1(_26470), .DIN2(_53489), .Q(_28579) );
  nor2s1 _28500_inst ( .DIN1(_28580), .DIN2(_27235), .Q(
        _________________________________12_________) );
  nor2s1 _28501_inst ( .DIN1(_28551), .DIN2(_28581), .Q(_28580) );
  nnd2s1 _28502_inst ( .DIN1(_28582), .DIN2(_28583), .Q(_28581) );
  nnd2s1 _28503_inst ( .DIN1(_28537), .DIN2(_26516), .Q(_28583) );
  nnd2s1 _28504_inst ( .DIN1(_28584), .DIN2(_28541), .Q(_28582) );
  xor2s1 _28505_inst ( .DIN1(_53494), .DIN2(_53496), .Q(_28584) );
  hi1s1 _28506_inst ( .DIN(_28585), .Q(_28551) );
  nnd2s1 _28507_inst ( .DIN1(_28586), .DIN2(_28587), .Q(
        _________________________________11_________) );
  nnd2s1 _28508_inst ( .DIN1(_28275), .DIN2(_28588), .Q(_28587) );
  xor2s1 _28509_inst ( .DIN1(_53495), .DIN2(_53496), .Q(_28588) );
  hi1s1 _28510_inst ( .DIN(_28234), .Q(_28275) );
  nnd2s1 _28511_inst ( .DIN1(_28589), .DIN2(_28590), .Q(_28586) );
  nnd2s1 _28512_inst ( .DIN1(_28591), .DIN2(_28585), .Q(_28590) );
  nnd2s1 _28513_inst ( .DIN1(_28592), .DIN2(_28522), .Q(_28585) );
  and2s1 _28514_inst ( .DIN1(_28593), .DIN2(_28594), .Q(_28522) );
  nor2s1 _28515_inst ( .DIN1(_28595), .DIN2(_28596), .Q(_28594) );
  nor2s1 _28516_inst ( .DIN1(_28597), .DIN2(_28598), .Q(_28593) );
  nor2s1 _28517_inst ( .DIN1(_28599), .DIN2(_28537), .Q(_28592) );
  nor2s1 _28518_inst ( .DIN1(_28600), .DIN2(_28601), .Q(_28591) );
  and2s1 _28519_inst ( .DIN1(_53075), .DIN2(_28537), .Q(_28601) );
  nor2s1 _28520_inst ( .DIN1(_28537), .DIN2(_26577), .Q(_28600) );
  hi1s1 _28521_inst ( .DIN(_28541), .Q(_28537) );
  nnd2s1 _28522_inst ( .DIN1(_28602), .DIN2(_28441), .Q(_28541) );
  nor2s1 _28523_inst ( .DIN1(_28595), .DIN2(_28603), .Q(_28602) );
  nnd2s1 _28524_inst ( .DIN1(_28604), .DIN2(_28605), .Q(
        _________________________________10_________) );
  nor2s1 _28525_inst ( .DIN1(_28606), .DIN2(_28607), .Q(_28605) );
  nor2s1 _28526_inst ( .DIN1(_27093), .DIN2(_28608), .Q(_28607) );
  nnd2s1 _28527_inst ( .DIN1(_28609), .DIN2(_28610), .Q(_28608) );
  nnd2s1 _28528_inst ( .DIN1(_28230), .DIN2(_28611), .Q(_28609) );
  nnd2s1 _28529_inst ( .DIN1(_53081), .DIN2(_28589), .Q(_28611) );
  nor2s1 _28530_inst ( .DIN1(_28612), .DIN2(_28613), .Q(_28606) );
  nor2s1 _28531_inst ( .DIN1(_28614), .DIN2(_28615), .Q(_28612) );
  nor2s1 _28532_inst ( .DIN1(_28347), .DIN2(_28610), .Q(_28615) );
  nnd2s1 _28533_inst ( .DIN1(_28249), .DIN2(_28616), .Q(_28610) );
  nnd2s1 _28534_inst ( .DIN1(_28617), .DIN2(______[16]), .Q(_28616) );
  xor2s1 _28535_inst ( .DIN1(_26431), .DIN2(_28618), .Q(_28617) );
  nor2s1 _28536_inst ( .DIN1(_53495), .DIN2(_26598), .Q(_28618) );
  nor2s1 _28537_inst ( .DIN1(_53081), .DIN2(_28270), .Q(_28614) );
  nnd2s1 _28538_inst ( .DIN1(_28245), .DIN2(_28589), .Q(_28270) );
  hi1s1 _28539_inst ( .DIN(_28249), .Q(_28245) );
  nor2s1 _28540_inst ( .DIN1(_28619), .DIN2(_28620), .Q(_28604) );
  nor2s1 _28541_inst ( .DIN1(_28230), .DIN2(_28233), .Q(_28620) );
  nnd2s1 _28542_inst ( .DIN1(_28589), .DIN2(_28249), .Q(_28230) );
  nnd2s1 _28543_inst ( .DIN1(_28621), .DIN2(_28622), .Q(_28249) );
  nor2s1 _28544_inst ( .DIN1(_28527), .DIN2(_28389), .Q(_28621) );
  nor2s1 _28545_inst ( .DIN1(_26431), .DIN2(_28234), .Q(_28619) );
  nnd2s1 _28546_inst ( .DIN1(_28347), .DIN2(_28350), .Q(_28234) );
  nnd2s1 _28547_inst ( .DIN1(_28623), .DIN2(_28624), .Q(
        _________________________________0_________) );
  nnd2s1 _28548_inst ( .DIN1(_28625), .DIN2(_53092), .Q(_28624) );
  nor2s1 _28549_inst ( .DIN1(_28626), .DIN2(_28627), .Q(_28623) );
  nor2s1 _28550_inst ( .DIN1(_28628), .DIN2(_28629), .Q(_28627) );
  nor2s1 _28551_inst ( .DIN1(_28303), .DIN2(_28630), .Q(_28628) );
  nnd2s1 _28552_inst ( .DIN1(_28631), .DIN2(_28632), .Q(_28630) );
  nnd2s1 _28553_inst ( .DIN1(_28293), .DIN2(_26406), .Q(_28632) );
  nnd2s1 _28554_inst ( .DIN1(_28633), .DIN2(_28292), .Q(_28631) );
  nor2s1 _28555_inst ( .DIN1(_53092), .DIN2(_53133), .Q(_28633) );
  hi1s1 _28556_inst ( .DIN(_28289), .Q(_28303) );
  nor2s1 _28557_inst ( .DIN1(_28634), .DIN2(_28635), .Q(_28626) );
  nnd2s1 _28558_inst ( .DIN1(______[4]), .DIN2(_28350), .Q(_28635) );
  xnr2s1 _28559_inst ( .DIN1(_53092), .DIN2(_28351), .Q(_28634) );
  nnd2s1 _28560_inst ( .DIN1(_28636), .DIN2(_27998), .Q(
        ______________________________9________) );
  nor2s1 _28561_inst ( .DIN1(_28637), .DIN2(_28638), .Q(_28636) );
  nor2s1 _28562_inst ( .DIN1(_27749), .DIN2(_28639), .Q(_28638) );
  nnd2s1 _28563_inst ( .DIN1(_28640), .DIN2(_28641), .Q(_28639) );
  nnd2s1 _28564_inst ( .DIN1(_28642), .DIN2(_53389), .Q(_28641) );
  nnd2s1 _28565_inst ( .DIN1(_28643), .DIN2(_28644), .Q(_28640) );
  nnd2s1 _28566_inst ( .DIN1(_52966), .DIN2(_52986), .Q(_28644) );
  nor2s1 _28567_inst ( .DIN1(_28010), .DIN2(_28645), .Q(_28637) );
  nor2s1 _28568_inst ( .DIN1(_28646), .DIN2(_26473), .Q(_28645) );
  nnd2s1 _28569_inst ( .DIN1(_28647), .DIN2(_28648), .Q(
        ______________________________99________) );
  nnd2s1 _28570_inst ( .DIN1(_28649), .DIN2(_26691), .Q(_28648) );
  nnd2s1 _28571_inst ( .DIN1(_28650), .DIN2(_28651), .Q(_28649) );
  or2s1 _28572_inst ( .DIN1(_28652), .DIN2(_28653), .Q(_28651) );
  nor2s1 _28573_inst ( .DIN1(_28654), .DIN2(_28655), .Q(_28647) );
  nor2s1 _28574_inst ( .DIN1(_28656), .DIN2(_28657), .Q(_28655) );
  nor2s1 _28575_inst ( .DIN1(_28658), .DIN2(_28659), .Q(_28656) );
  nor2s1 _28576_inst ( .DIN1(_28660), .DIN2(_28661), .Q(_28659) );
  xor2s1 _28577_inst ( .DIN1(_28662), .DIN2(_28663), .Q(_28661) );
  xor2s1 _28578_inst ( .DIN1(_26537), .DIN2(_28664), .Q(_28663) );
  nor2s1 _28579_inst ( .DIN1(_26691), .DIN2(_28665), .Q(_28658) );
  nnd2s1 _28580_inst ( .DIN1(_28666), .DIN2(_28653), .Q(_28665) );
  nor2s1 _28581_inst ( .DIN1(_53004), .DIN2(_53005), .Q(_28653) );
  hi1s1 _28582_inst ( .DIN(_28652), .Q(_28666) );
  nnd2s1 _28583_inst ( .DIN1(_28667), .DIN2(_28668), .Q(
        ______________________________98________) );
  nnd2s1 _28584_inst ( .DIN1(_28669), .DIN2(_28670), .Q(_28668) );
  nnd2s1 _28585_inst ( .DIN1(_28671), .DIN2(_28672), .Q(_28669) );
  xor2s1 _28586_inst ( .DIN1(_26623), .DIN2(_28673), .Q(_28671) );
  nor2s1 _28587_inst ( .DIN1(_53062), .DIN2(_26612), .Q(_28673) );
  nor2s1 _28588_inst ( .DIN1(_28674), .DIN2(_28675), .Q(_28667) );
  nor2s1 _28589_inst ( .DIN1(_28676), .DIN2(_28677), .Q(_28675) );
  xor2s1 _28590_inst ( .DIN1(_28678), .DIN2(_28679), .Q(_28676) );
  xor2s1 _28591_inst ( .DIN1(_28680), .DIN2(_52853), .Q(_28678) );
  nor2s1 _28592_inst ( .DIN1(_28681), .DIN2(_28682), .Q(_28674) );
  or2s1 _28593_inst ( .DIN1(_28683), .DIN2(_28684), .Q(_28682) );
  xor2s1 _28594_inst ( .DIN1(_53061), .DIN2(_53464), .Q(_28681) );
  nnd2s1 _28595_inst ( .DIN1(_28685), .DIN2(_28686), .Q(
        ______________________________97________) );
  nnd2s1 _28596_inst ( .DIN1(_28687), .DIN2(_28657), .Q(_28686) );
  nnd2s1 _28597_inst ( .DIN1(_28688), .DIN2(_28689), .Q(_28687) );
  nor2s1 _28598_inst ( .DIN1(_28690), .DIN2(_28691), .Q(_28688) );
  nor2s1 _28599_inst ( .DIN1(_53003), .DIN2(_53005), .Q(_28691) );
  nor2s1 _28600_inst ( .DIN1(_28692), .DIN2(_28693), .Q(_28685) );
  nor2s1 _28601_inst ( .DIN1(_28694), .DIN2(_28695), .Q(_28693) );
  xor2s1 _28602_inst ( .DIN1(_52903), .DIN2(_53040), .Q(_28695) );
  nor2s1 _28603_inst ( .DIN1(_28696), .DIN2(_28697), .Q(_28692) );
  nnd2s1 _28604_inst ( .DIN1(_28698), .DIN2(_28680), .Q(_28697) );
  hi1s1 _28605_inst ( .DIN(_28699), .Q(_28680) );
  nnd2s1 _28606_inst ( .DIN1(_28700), .DIN2(_26359), .Q(_28698) );
  nnd2s1 _28607_inst ( .DIN1(_28701), .DIN2(_28702), .Q(
        ______________________________96________) );
  nnd2s1 _28608_inst ( .DIN1(_28703), .DIN2(_53126), .Q(_28702) );
  nor2s1 _28609_inst ( .DIN1(_28704), .DIN2(_28705), .Q(_28703) );
  nor2s1 _28610_inst ( .DIN1(_28706), .DIN2(_28707), .Q(_28701) );
  nor2s1 _28611_inst ( .DIN1(_26360), .DIN2(_28708), .Q(_28707) );
  or2s1 _28612_inst ( .DIN1(_28709), .DIN2(_26774), .Q(_28708) );
  nor2s1 _28613_inst ( .DIN1(_28710), .DIN2(_28711), .Q(_28706) );
  nnd2s1 _28614_inst ( .DIN1(______[30]), .DIN2(_28712), .Q(_28711) );
  xor2s1 _28615_inst ( .DIN1(_53107), .DIN2(_28713), .Q(_28712) );
  nnd2s1 _28616_inst ( .DIN1(_28714), .DIN2(_28715), .Q(
        ______________________________95________) );
  nnd2s1 _28617_inst ( .DIN1(_28716), .DIN2(_28717), .Q(_28715) );
  nor2s1 _28618_inst ( .DIN1(_28718), .DIN2(_27614), .Q(_28716) );
  xor2s1 _28619_inst ( .DIN1(_28719), .DIN2(_28720), .Q(_28718) );
  xor2s1 _28620_inst ( .DIN1(_52970), .DIN2(_53206), .Q(_28720) );
  nnd2s1 _28621_inst ( .DIN1(_53104), .DIN2(_26349), .Q(_28719) );
  nnd2s1 _28622_inst ( .DIN1(_28721), .DIN2(_27994), .Q(_28714) );
  nor2s1 _28623_inst ( .DIN1(_28722), .DIN2(_28723), .Q(_28721) );
  nor2s1 _28624_inst ( .DIN1(_28705), .DIN2(_26630), .Q(_28723) );
  nor2s1 _28625_inst ( .DIN1(_28724), .DIN2(_28725), .Q(_28722) );
  nnd2s1 _28626_inst ( .DIN1(_28726), .DIN2(______[28]), .Q(_28725) );
  nor2s1 _28627_inst ( .DIN1(_28727), .DIN2(_28728), .Q(_28726) );
  xor2s1 _28628_inst ( .DIN1(_26471), .DIN2(_28713), .Q(_28728) );
  nor2s1 _28629_inst ( .DIN1(_26349), .DIN2(_52958), .Q(_28713) );
  nnd2s1 _28630_inst ( .DIN1(_28729), .DIN2(_28730), .Q(
        ______________________________94________) );
  nor2s1 _28631_inst ( .DIN1(_28731), .DIN2(_28732), .Q(_28730) );
  nor2s1 _28632_inst ( .DIN1(_28733), .DIN2(_28734), .Q(_28732) );
  nor2s1 _28633_inst ( .DIN1(_28735), .DIN2(_28736), .Q(_28734) );
  nor2s1 _28634_inst ( .DIN1(_28724), .DIN2(_28737), .Q(_28736) );
  and2s1 _28635_inst ( .DIN1(_28724), .DIN2(_52956), .Q(_28735) );
  nor2s1 _28636_inst ( .DIN1(______[2]), .DIN2(_28738), .Q(_28731) );
  nor2s1 _28637_inst ( .DIN1(_28739), .DIN2(_28740), .Q(_28729) );
  nnd2s1 _28638_inst ( .DIN1(_28741), .DIN2(_28742), .Q(
        ______________________________93________) );
  nnd2s1 _28639_inst ( .DIN1(_28743), .DIN2(______[16]), .Q(_28742) );
  nor2s1 _28640_inst ( .DIN1(_28744), .DIN2(_28745), .Q(_28743) );
  xnr2s1 _28641_inst ( .DIN1(_53071), .DIN2(_53106), .Q(_28745) );
  nnd2s1 _28642_inst ( .DIN1(_28746), .DIN2(_27571), .Q(_28741) );
  nor2s1 _28643_inst ( .DIN1(_28747), .DIN2(_28748), .Q(_28746) );
  nor2s1 _28644_inst ( .DIN1(_28724), .DIN2(_28749), .Q(_28748) );
  nor2s1 _28645_inst ( .DIN1(_28750), .DIN2(_28751), .Q(_28749) );
  nor2s1 _28646_inst ( .DIN1(_52958), .DIN2(_28752), .Q(_28751) );
  nor2s1 _28647_inst ( .DIN1(_52957), .DIN2(_28727), .Q(_28752) );
  nor2s1 _28648_inst ( .DIN1(_28737), .DIN2(_26383), .Q(_28750) );
  nor2s1 _28649_inst ( .DIN1(_26349), .DIN2(_28727), .Q(_28737) );
  nor2s1 _28650_inst ( .DIN1(_52857), .DIN2(_28705), .Q(_28747) );
  nnd2s1 _28651_inst ( .DIN1(_28753), .DIN2(_28754), .Q(
        ______________________________92________) );
  nnd2s1 _28652_inst ( .DIN1(_28755), .DIN2(_28756), .Q(_28754) );
  nnd2s1 _28653_inst ( .DIN1(_28757), .DIN2(_28758), .Q(_28756) );
  nor2s1 _28654_inst ( .DIN1(_28759), .DIN2(_28760), .Q(_28758) );
  nor2s1 _28655_inst ( .DIN1(_28761), .DIN2(_28762), .Q(_28760) );
  nor2s1 _28656_inst ( .DIN1(_28763), .DIN2(_28646), .Q(_28762) );
  nor2s1 _28657_inst ( .DIN1(_28764), .DIN2(_26512), .Q(_28763) );
  nor2s1 _28658_inst ( .DIN1(_26235), .DIN2(_26496), .Q(_28764) );
  nor2s1 _28659_inst ( .DIN1(_52859), .DIN2(_28765), .Q(_28759) );
  nor2s1 _28660_inst ( .DIN1(_28766), .DIN2(_28767), .Q(_28757) );
  nor2s1 _28661_inst ( .DIN1(_53009), .DIN2(_28768), .Q(_28767) );
  nnd2s1 _28662_inst ( .DIN1(_27968), .DIN2(_53175), .Q(_28753) );
  nnd2s1 _28663_inst ( .DIN1(_28769), .DIN2(_28770), .Q(
        ______________________________91________) );
  nnd2s1 _28664_inst ( .DIN1(_28771), .DIN2(_28772), .Q(_28770) );
  hi1s1 _28665_inst ( .DIN(_28773), .Q(_28772) );
  nor2s1 _28666_inst ( .DIN1(_28774), .DIN2(_28775), .Q(_28771) );
  nor2s1 _28667_inst ( .DIN1(_28776), .DIN2(_28777), .Q(_28775) );
  nor2s1 _28668_inst ( .DIN1(_28778), .DIN2(_28779), .Q(_28777) );
  and2s1 _28669_inst ( .DIN1(_28765), .DIN2(_53174), .Q(_28779) );
  nor2s1 _28670_inst ( .DIN1(_52860), .DIN2(_28765), .Q(_28778) );
  hi1s1 _28671_inst ( .DIN(_28768), .Q(_28776) );
  nor2s1 _28672_inst ( .DIN1(_53174), .DIN2(_28768), .Q(_28774) );
  nnd2s1 _28673_inst ( .DIN1(_28780), .DIN2(_52855), .Q(_28768) );
  nor2s1 _28674_inst ( .DIN1(_28761), .DIN2(_26235), .Q(_28780) );
  nnd2s1 _28675_inst ( .DIN1(_28781), .DIN2(_28782), .Q(
        ______________________________90________) );
  nor2s1 _28676_inst ( .DIN1(_28783), .DIN2(_28784), .Q(_28781) );
  nor2s1 _28677_inst ( .DIN1(_28785), .DIN2(_28786), .Q(_28784) );
  nor2s1 _28678_inst ( .DIN1(_28773), .DIN2(_28787), .Q(_28785) );
  nnd2s1 _28679_inst ( .DIN1(_28788), .DIN2(_28789), .Q(_28787) );
  nnd2s1 _28680_inst ( .DIN1(_28761), .DIN2(_52991), .Q(_28789) );
  nnd2s1 _28681_inst ( .DIN1(_28765), .DIN2(_26496), .Q(_28788) );
  nnd2s1 _28682_inst ( .DIN1(_28790), .DIN2(_28791), .Q(_28773) );
  nnd2s1 _28683_inst ( .DIN1(_28765), .DIN2(_26774), .Q(_28791) );
  nor2s1 _28684_inst ( .DIN1(_53162), .DIN2(_28792), .Q(_28783) );
  nnd2s1 _28685_inst ( .DIN1(_28793), .DIN2(_28794), .Q(
        ______________________________8________) );
  nor2s1 _28686_inst ( .DIN1(_28795), .DIN2(_28796), .Q(_28793) );
  nor2s1 _28687_inst ( .DIN1(_28797), .DIN2(_28798), .Q(_28796) );
  xnr2s1 _28688_inst ( .DIN1(_28799), .DIN2(_53010), .Q(_28798) );
  nor2s1 _28689_inst ( .DIN1(_28800), .DIN2(_28801), .Q(_28795) );
  nor2s1 _28690_inst ( .DIN1(_28802), .DIN2(_28803), .Q(_28800) );
  nor2s1 _28691_inst ( .DIN1(_26620), .DIN2(_28804), .Q(_28803) );
  nor2s1 _28692_inst ( .DIN1(_28805), .DIN2(_28806), .Q(_28802) );
  nnd2s1 _28693_inst ( .DIN1(______[30]), .DIN2(_28807), .Q(_28806) );
  xor2s1 _28694_inst ( .DIN1(_52877), .DIN2(_28808), .Q(_28807) );
  hi1s1 _28695_inst ( .DIN(_28809), .Q(_28805) );
  nnd2s1 _28696_inst ( .DIN1(_28810), .DIN2(_28811), .Q(
        ______________________________89________) );
  nor2s1 _28697_inst ( .DIN1(_28812), .DIN2(_28813), .Q(_28810) );
  nor2s1 _28698_inst ( .DIN1(_28814), .DIN2(_28815), .Q(_28813) );
  nnd2s1 _28699_inst ( .DIN1(_28816), .DIN2(_28790), .Q(_28815) );
  nor2s1 _28700_inst ( .DIN1(_28817), .DIN2(_28818), .Q(_28816) );
  nor2s1 _28701_inst ( .DIN1(_28761), .DIN2(_28819), .Q(_28818) );
  xor2s1 _28702_inst ( .DIN1(_52855), .DIN2(_53163), .Q(_28819) );
  nor2s1 _28703_inst ( .DIN1(_52861), .DIN2(_28765), .Q(_28817) );
  nor2s1 _28704_inst ( .DIN1(_28356), .DIN2(_28820), .Q(_28812) );
  xor2s1 _28705_inst ( .DIN1(_26487), .DIN2(_28821), .Q(_28820) );
  nnd2s1 _28706_inst ( .DIN1(_53224), .DIN2(_53009), .Q(_28821) );
  nnd2s1 _28707_inst ( .DIN1(_28822), .DIN2(_28026), .Q(
        ______________________________88________) );
  nor2s1 _28708_inst ( .DIN1(_28823), .DIN2(_28824), .Q(_28822) );
  nor2s1 _28709_inst ( .DIN1(_28825), .DIN2(_28016), .Q(_28824) );
  nor2s1 _28710_inst ( .DIN1(_28766), .DIN2(_28826), .Q(_28825) );
  nnd2s1 _28711_inst ( .DIN1(_28827), .DIN2(_28828), .Q(_28826) );
  nnd2s1 _28712_inst ( .DIN1(_28761), .DIN2(_52862), .Q(_28828) );
  nnd2s1 _28713_inst ( .DIN1(_28829), .DIN2(_28765), .Q(_28827) );
  nnd2s1 _28714_inst ( .DIN1(_28830), .DIN2(______[0]), .Q(_28829) );
  xor2s1 _28715_inst ( .DIN1(_28831), .DIN2(_53027), .Q(_28830) );
  nnd2s1 _28716_inst ( .DIN1(_53468), .DIN2(_26257), .Q(_28831) );
  hi1s1 _28717_inst ( .DIN(_28790), .Q(_28766) );
  nor2s1 _28718_inst ( .DIN1(_28024), .DIN2(_28832), .Q(_28823) );
  nor2s1 _28719_inst ( .DIN1(_28833), .DIN2(_28834), .Q(_28832) );
  hi1s1 _28720_inst ( .DIN(_28835), .Q(_28834) );
  nor2s1 _28721_inst ( .DIN1(_53410), .DIN2(_53437), .Q(_28833) );
  nnd2s1 _28722_inst ( .DIN1(_28836), .DIN2(_28837), .Q(
        ______________________________87________) );
  nor2s1 _28723_inst ( .DIN1(_28838), .DIN2(_28839), .Q(_28836) );
  nor2s1 _28724_inst ( .DIN1(_28704), .DIN2(_28840), .Q(_28839) );
  nnd2s1 _28725_inst ( .DIN1(_28841), .DIN2(_28790), .Q(_28840) );
  nnd2s1 _28726_inst ( .DIN1(_28842), .DIN2(_28843), .Q(_28790) );
  nor2s1 _28727_inst ( .DIN1(_28761), .DIN2(_28844), .Q(_28842) );
  nor2s1 _28728_inst ( .DIN1(_28845), .DIN2(_28846), .Q(_28841) );
  nor2s1 _28729_inst ( .DIN1(_28761), .DIN2(_28847), .Q(_28846) );
  xor2s1 _28730_inst ( .DIN1(_26401), .DIN2(_53468), .Q(_28847) );
  hi1s1 _28731_inst ( .DIN(_28765), .Q(_28761) );
  nor2s1 _28732_inst ( .DIN1(_52863), .DIN2(_28765), .Q(_28845) );
  nnd2s1 _28733_inst ( .DIN1(_28848), .DIN2(_28727), .Q(_28765) );
  nor2s1 _28734_inst ( .DIN1(_28849), .DIN2(_28850), .Q(_28848) );
  nor2s1 _28735_inst ( .DIN1(_28851), .DIN2(_28852), .Q(_28838) );
  nor2s1 _28736_inst ( .DIN1(_26855), .DIN2(_26471), .Q(_28852) );
  nnd2s1 _28737_inst ( .DIN1(_28853), .DIN2(_28854), .Q(
        ______________________________86________) );
  nnd2s1 _28738_inst ( .DIN1(_28855), .DIN2(_28095), .Q(_28854) );
  nor2s1 _28739_inst ( .DIN1(_28646), .DIN2(_28856), .Q(_28855) );
  nnd2s1 _28740_inst ( .DIN1(_28857), .DIN2(_26703), .Q(_28856) );
  nnd2s1 _28741_inst ( .DIN1(_28858), .DIN2(_28098), .Q(_28853) );
  xor2s1 _28742_inst ( .DIN1(_28859), .DIN2(_28860), .Q(_28858) );
  nor2s1 _28743_inst ( .DIN1(_28861), .DIN2(_28862), .Q(_28859) );
  nor2s1 _28744_inst ( .DIN1(_28863), .DIN2(_26293), .Q(_28862) );
  nor2s1 _28745_inst ( .DIN1(_52969), .DIN2(_28864), .Q(_28861) );
  nnd2s1 _28746_inst ( .DIN1(_28865), .DIN2(_28866), .Q(
        ______________________________85________) );
  nnd2s1 _28747_inst ( .DIN1(_27717), .DIN2(_28867), .Q(_28866) );
  xor2s1 _28748_inst ( .DIN1(_26661), .DIN2(_28868), .Q(_28867) );
  nnd2s1 _28749_inst ( .DIN1(_53200), .DIN2(_53027), .Q(_28868) );
  nnd2s1 _28750_inst ( .DIN1(_28869), .DIN2(_27611), .Q(_28865) );
  nor2s1 _28751_inst ( .DIN1(_28870), .DIN2(_28871), .Q(_28869) );
  nor2s1 _28752_inst ( .DIN1(_53413), .DIN2(_28863), .Q(_28871) );
  nor2s1 _28753_inst ( .DIN1(_28864), .DIN2(_28872), .Q(_28870) );
  xor2s1 _28754_inst ( .DIN1(_52969), .DIN2(_53468), .Q(_28872) );
  nnd2s1 _28755_inst ( .DIN1(_28873), .DIN2(_28874), .Q(
        ______________________________84________) );
  nnd2s1 _28756_inst ( .DIN1(_28875), .DIN2(_26305), .Q(_28874) );
  nor2s1 _28757_inst ( .DIN1(_28876), .DIN2(_28877), .Q(_28873) );
  nor2s1 _28758_inst ( .DIN1(_28878), .DIN2(_28879), .Q(_28877) );
  nor2s1 _28759_inst ( .DIN1(_28880), .DIN2(_28864), .Q(_28878) );
  xnr2s1 _28760_inst ( .DIN1(_28881), .DIN2(_28882), .Q(_28880) );
  xor2s1 _28761_inst ( .DIN1(_53388), .DIN2(_26388), .Q(_28881) );
  nor2s1 _28762_inst ( .DIN1(_28709), .DIN2(_28883), .Q(_28876) );
  nnd2s1 _28763_inst ( .DIN1(______[30]), .DIN2(_28884), .Q(_28883) );
  xor2s1 _28764_inst ( .DIN1(_26257), .DIN2(_28885), .Q(_28884) );
  nnd2s1 _28765_inst ( .DIN1(_52974), .DIN2(_52954), .Q(_28885) );
  nnd2s1 _28766_inst ( .DIN1(_28704), .DIN2(_28886), .Q(_28709) );
  nnd2s1 _28767_inst ( .DIN1(_28887), .DIN2(_28888), .Q(_28886) );
  nnd2s1 _28768_inst ( .DIN1(_28889), .DIN2(_28890), .Q(
        ______________________________83________) );
  nor2s1 _28769_inst ( .DIN1(_28891), .DIN2(_28892), .Q(_28890) );
  nor2s1 _28770_inst ( .DIN1(_28893), .DIN2(_28894), .Q(_28892) );
  or2s1 _28771_inst ( .DIN1(_28879), .DIN2(_28864), .Q(_28894) );
  or2s1 _28772_inst ( .DIN1(_26991), .DIN2(_52974), .Q(_28893) );
  nor2s1 _28773_inst ( .DIN1(_28895), .DIN2(_28896), .Q(_28889) );
  and2s1 _28774_inst ( .DIN1(_52898), .DIN2(_28875), .Q(_28896) );
  nor2s1 _28775_inst ( .DIN1(_28851), .DIN2(_28897), .Q(_28895) );
  nor2s1 _28776_inst ( .DIN1(_28898), .DIN2(_28684), .Q(_28897) );
  xor2s1 _28777_inst ( .DIN1(_26478), .DIN2(_52985), .Q(_28898) );
  nnd2s1 _28778_inst ( .DIN1(_28899), .DIN2(_28900), .Q(
        ______________________________82________) );
  nor2s1 _28779_inst ( .DIN1(_28901), .DIN2(_28902), .Q(_28900) );
  nor2s1 _28780_inst ( .DIN1(_26388), .DIN2(_28903), .Q(_28902) );
  nnd2s1 _28781_inst ( .DIN1(_28904), .DIN2(_28704), .Q(_28903) );
  nor2s1 _28782_inst ( .DIN1(_52977), .DIN2(_28905), .Q(_28901) );
  nor2s1 _28783_inst ( .DIN1(_28906), .DIN2(_28907), .Q(_28905) );
  nor2s1 _28784_inst ( .DIN1(_28851), .DIN2(_28904), .Q(_28907) );
  nor2s1 _28785_inst ( .DIN1(_26226), .DIN2(_26700), .Q(_28904) );
  nor2s1 _28786_inst ( .DIN1(_28879), .DIN2(_28908), .Q(_28906) );
  nnd2s1 _28787_inst ( .DIN1(_28909), .DIN2(______[26]), .Q(_28908) );
  nnd2s1 _28788_inst ( .DIN1(_28851), .DIN2(_28863), .Q(_28879) );
  nor2s1 _28789_inst ( .DIN1(_28891), .DIN2(_28910), .Q(_28899) );
  nor2s1 _28790_inst ( .DIN1(_52864), .DIN2(_28911), .Q(_28910) );
  hi1s1 _28791_inst ( .DIN(_28875), .Q(_28911) );
  nor2s1 _28792_inst ( .DIN1(_28863), .DIN2(_28704), .Q(_28875) );
  nnd2s1 _28793_inst ( .DIN1(_28912), .DIN2(_28913), .Q(
        ______________________________81________) );
  nnd2s1 _28794_inst ( .DIN1(_28308), .DIN2(_28914), .Q(_28913) );
  nnd2s1 _28795_inst ( .DIN1(_28915), .DIN2(_28916), .Q(_28914) );
  nnd2s1 _28796_inst ( .DIN1(_28917), .DIN2(_28909), .Q(_28916) );
  nor2s1 _28797_inst ( .DIN1(_28918), .DIN2(_28919), .Q(_28917) );
  nor2s1 _28798_inst ( .DIN1(_28920), .DIN2(_26226), .Q(_28919) );
  nor2s1 _28799_inst ( .DIN1(_52977), .DIN2(_53388), .Q(_28920) );
  nor2s1 _28800_inst ( .DIN1(_53388), .DIN2(_28882), .Q(_28918) );
  nnd2s1 _28801_inst ( .DIN1(_26388), .DIN2(_26226), .Q(_28882) );
  nnd2s1 _28802_inst ( .DIN1(_52867), .DIN2(_28921), .Q(_28915) );
  hi1s1 _28803_inst ( .DIN(_28863), .Q(_28921) );
  nnd2s1 _28804_inst ( .DIN1(_28922), .DIN2(_28864), .Q(_28863) );
  nnd2s1 _28805_inst ( .DIN1(_28923), .DIN2(_26470), .Q(_28912) );
  nnd2s1 _28806_inst ( .DIN1(_28924), .DIN2(_53094), .Q(
        ______________________________80________) );
  nor2s1 _28807_inst ( .DIN1(_28925), .DIN2(_28926), .Q(_28924) );
  nnd2s1 _28808_inst ( .DIN1(_28927), .DIN2(_28928), .Q(
        ______________________________7________) );
  nnd2s1 _28809_inst ( .DIN1(_28929), .DIN2(_52966), .Q(_28928) );
  nor2s1 _28810_inst ( .DIN1(_28930), .DIN2(_27241), .Q(_28929) );
  nnd2s1 _28811_inst ( .DIN1(_28931), .DIN2(_28932), .Q(_28927) );
  nor2s1 _28812_inst ( .DIN1(_28933), .DIN2(_28934), .Q(_28931) );
  nor2s1 _28813_inst ( .DIN1(_28935), .DIN2(_28936), .Q(_28934) );
  nnd2s1 _28814_inst ( .DIN1(_28937), .DIN2(______[22]), .Q(_28936) );
  nor2s1 _28815_inst ( .DIN1(_28938), .DIN2(_28939), .Q(_28937) );
  xor2s1 _28816_inst ( .DIN1(_52871), .DIN2(_28808), .Q(_28939) );
  nor2s1 _28817_inst ( .DIN1(_52856), .DIN2(_28804), .Q(_28933) );
  nnd2s1 _28818_inst ( .DIN1(_28940), .DIN2(_28941), .Q(
        ______________________________79________) );
  nor2s1 _28819_inst ( .DIN1(_28942), .DIN2(_28943), .Q(_28940) );
  nor2s1 _28820_inst ( .DIN1(_28944), .DIN2(_28945), .Q(_28943) );
  xnr2s1 _28821_inst ( .DIN1(_28946), .DIN2(_28947), .Q(_28945) );
  xor2s1 _28822_inst ( .DIN1(_52944), .DIN2(_52945), .Q(_28947) );
  nor2s1 _28823_inst ( .DIN1(_28948), .DIN2(_28949), .Q(_28942) );
  nor2s1 _28824_inst ( .DIN1(_52868), .DIN2(_28926), .Q(_28948) );
  nnd2s1 _28825_inst ( .DIN1(_28950), .DIN2(_28951), .Q(
        ______________________________78________) );
  nor2s1 _28826_inst ( .DIN1(_28952), .DIN2(_28953), .Q(_28950) );
  nor2s1 _28827_inst ( .DIN1(_28954), .DIN2(_28955), .Q(_28953) );
  nnd2s1 _28828_inst ( .DIN1(_52931), .DIN2(_28956), .Q(_28955) );
  nor2s1 _28829_inst ( .DIN1(_28957), .DIN2(_28958), .Q(_28952) );
  nor2s1 _28830_inst ( .DIN1(_26774), .DIN2(_26226), .Q(_28958) );
  nnd2s1 _28831_inst ( .DIN1(_28959), .DIN2(_28794), .Q(
        ______________________________77________) );
  nor2s1 _28832_inst ( .DIN1(_28960), .DIN2(_28961), .Q(_28959) );
  nor2s1 _28833_inst ( .DIN1(_28801), .DIN2(_28962), .Q(_28961) );
  nnd2s1 _28834_inst ( .DIN1(_53128), .DIN2(_28956), .Q(_28962) );
  nor2s1 _28835_inst ( .DIN1(_28797), .DIN2(_28963), .Q(_28960) );
  nor2s1 _28836_inst ( .DIN1(_28964), .DIN2(_28100), .Q(_28963) );
  xor2s1 _28837_inst ( .DIN1(_26259), .DIN2(_52871), .Q(_28964) );
  nnd2s1 _28838_inst ( .DIN1(_28965), .DIN2(_28966), .Q(
        ______________________________76________) );
  nnd2s1 _28839_inst ( .DIN1(_28967), .DIN2(_28968), .Q(_28966) );
  nor2s1 _28840_inst ( .DIN1(_28969), .DIN2(_27393), .Q(_28967) );
  xnr2s1 _28841_inst ( .DIN1(_53301), .DIN2(_53239), .Q(_28969) );
  nnd2s1 _28842_inst ( .DIN1(_28970), .DIN2(_28971), .Q(_28965) );
  nor2s1 _28843_inst ( .DIN1(_52869), .DIN2(_28926), .Q(_28970) );
  nnd2s1 _28844_inst ( .DIN1(_28972), .DIN2(_28973), .Q(
        ______________________________75________) );
  nnd2s1 _28845_inst ( .DIN1(_28974), .DIN2(_28975), .Q(_28973) );
  xor2s1 _28846_inst ( .DIN1(_28082), .DIN2(_53505), .Q(_28975) );
  nnd2s1 _28847_inst ( .DIN1(_52915), .DIN2(_53432), .Q(_28082) );
  nor2s1 _28848_inst ( .DIN1(_28100), .DIN2(_28976), .Q(_28974) );
  nnd2s1 _28849_inst ( .DIN1(_27325), .DIN2(_28977), .Q(_28972) );
  nnd2s1 _28850_inst ( .DIN1(_28956), .DIN2(_26588), .Q(_28977) );
  nnd2s1 _28851_inst ( .DIN1(_28978), .DIN2(_28979), .Q(
        ______________________________74________) );
  nnd2s1 _28852_inst ( .DIN1(_28980), .DIN2(_28981), .Q(_28979) );
  xor2s1 _28853_inst ( .DIN1(_52977), .DIN2(_52985), .Q(_28981) );
  nnd2s1 _28854_inst ( .DIN1(_28982), .DIN2(_28957), .Q(_28978) );
  nor2s1 _28855_inst ( .DIN1(_28983), .DIN2(_28984), .Q(_28982) );
  nor2s1 _28856_inst ( .DIN1(_53432), .DIN2(_28985), .Q(_28984) );
  nor2s1 _28857_inst ( .DIN1(_28986), .DIN2(_26704), .Q(_28983) );
  nnd2s1 _28858_inst ( .DIN1(_28987), .DIN2(_28988), .Q(
        ______________________________73________) );
  nnd2s1 _28859_inst ( .DIN1(_28989), .DIN2(_28990), .Q(_28988) );
  xor2s1 _28860_inst ( .DIN1(_28991), .DIN2(_53247), .Q(_28990) );
  and2s1 _28861_inst ( .DIN1(______[8]), .DIN2(_28992), .Q(_28989) );
  nnd2s1 _28862_inst ( .DIN1(_27201), .DIN2(_28993), .Q(_28987) );
  nnd2s1 _28863_inst ( .DIN1(_28994), .DIN2(_28995), .Q(_28993) );
  nnd2s1 _28864_inst ( .DIN1(_28849), .DIN2(_28996), .Q(_28995) );
  xor2s1 _28865_inst ( .DIN1(_52992), .DIN2(_53432), .Q(_28996) );
  nnd2s1 _28866_inst ( .DIN1(_52833), .DIN2(_28922), .Q(_28994) );
  nor2s1 _28867_inst ( .DIN1(_28997), .DIN2(_28998), .Q(
        ______________________________72________) );
  nor2s1 _28868_inst ( .DIN1(_28999), .DIN2(_29000), .Q(_28997) );
  and2s1 _28869_inst ( .DIN1(_28922), .DIN2(_52875), .Q(_29000) );
  nor2s1 _28870_inst ( .DIN1(_29001), .DIN2(_29002), .Q(_28999) );
  nnd2s1 _28871_inst ( .DIN1(_28849), .DIN2(______[0]), .Q(_29002) );
  xor2s1 _28872_inst ( .DIN1(_52998), .DIN2(_53001), .Q(_29001) );
  nnd2s1 _28873_inst ( .DIN1(_29003), .DIN2(_28569), .Q(
        ______________________________71________) );
  nor2s1 _28874_inst ( .DIN1(_29004), .DIN2(_29005), .Q(_29003) );
  nor2s1 _28875_inst ( .DIN1(_28575), .DIN2(_29006), .Q(_29005) );
  nnd2s1 _28876_inst ( .DIN1(_29007), .DIN2(_29008), .Q(_29006) );
  nnd2s1 _28877_inst ( .DIN1(_28922), .DIN2(_26426), .Q(_29008) );
  nnd2s1 _28878_inst ( .DIN1(_29009), .DIN2(_28849), .Q(_29007) );
  xor2s1 _28879_inst ( .DIN1(_29010), .DIN2(_52995), .Q(_29009) );
  nnd2s1 _28880_inst ( .DIN1(_53095), .DIN2(_52998), .Q(_29010) );
  nor2s1 _28881_inst ( .DIN1(_28572), .DIN2(_29011), .Q(_29004) );
  nor2s1 _28882_inst ( .DIN1(_29012), .DIN2(_27082), .Q(_29011) );
  xor2s1 _28883_inst ( .DIN1(_29013), .DIN2(_29014), .Q(_29012) );
  xor2s1 _28884_inst ( .DIN1(_52999), .DIN2(_53138), .Q(_29014) );
  nnd2s1 _28885_inst ( .DIN1(_53095), .DIN2(_53018), .Q(_29013) );
  nor2s1 _28886_inst ( .DIN1(_29015), .DIN2(_27593), .Q(
        ______________________________70________) );
  nor2s1 _28887_inst ( .DIN1(_29016), .DIN2(_29017), .Q(_29015) );
  nor2s1 _28888_inst ( .DIN1(_28986), .DIN2(_26608), .Q(_29017) );
  nor2s1 _28889_inst ( .DIN1(_28985), .DIN2(_26405), .Q(_29016) );
  nnd2s1 _28890_inst ( .DIN1(_29018), .DIN2(_29019), .Q(
        ______________________________6________) );
  nnd2s1 _28891_inst ( .DIN1(_29020), .DIN2(_29021), .Q(_29019) );
  nnd2s1 _28892_inst ( .DIN1(_29022), .DIN2(_29023), .Q(_29020) );
  nor2s1 _28893_inst ( .DIN1(_28930), .DIN2(_28808), .Q(_29023) );
  nor2s1 _28894_inst ( .DIN1(_27651), .DIN2(_29024), .Q(_29022) );
  nnd2s1 _28895_inst ( .DIN1(_29025), .DIN2(_29026), .Q(_29024) );
  nnd2s1 _28896_inst ( .DIN1(_26304), .DIN2(_26568), .Q(_29026) );
  nnd2s1 _28897_inst ( .DIN1(_29027), .DIN2(_52966), .Q(_29025) );
  nnd2s1 _28898_inst ( .DIN1(_28932), .DIN2(_29028), .Q(_29018) );
  nnd2s1 _28899_inst ( .DIN1(_29029), .DIN2(_29030), .Q(_29028) );
  nnd2s1 _28900_inst ( .DIN1(_28809), .DIN2(_26568), .Q(_29030) );
  nnd2s1 _28901_inst ( .DIN1(_28935), .DIN2(_52838), .Q(_29029) );
  nnd2s1 _28902_inst ( .DIN1(_29031), .DIN2(_29032), .Q(
        ______________________________69________) );
  nnd2s1 _28903_inst ( .DIN1(_28738), .DIN2(_29033), .Q(_29032) );
  nnd2s1 _28904_inst ( .DIN1(_29034), .DIN2(_29035), .Q(_29033) );
  nnd2s1 _28905_inst ( .DIN1(_29036), .DIN2(_29037), .Q(_29035) );
  xnr2s1 _28906_inst ( .DIN1(_52998), .DIN2(_52995), .Q(_29037) );
  nor2s1 _28907_inst ( .DIN1(_27039), .DIN2(_28985), .Q(_29036) );
  nnd2s1 _28908_inst ( .DIN1(_52878), .DIN2(_28922), .Q(_29034) );
  nnd2s1 _28909_inst ( .DIN1(_29038), .DIN2(_29039), .Q(_29031) );
  xor2s1 _28910_inst ( .DIN1(_26383), .DIN2(_29040), .Q(_29038) );
  nnd2s1 _28911_inst ( .DIN1(_29041), .DIN2(_29042), .Q(
        ______________________________68________) );
  nnd2s1 _28912_inst ( .DIN1(_29043), .DIN2(_28980), .Q(_29042) );
  hi1s1 _28913_inst ( .DIN(_29044), .Q(_28980) );
  xnr2s1 _28914_inst ( .DIN1(_29045), .DIN2(_52934), .Q(_29043) );
  nnd2s1 _28915_inst ( .DIN1(_28957), .DIN2(_29046), .Q(_29041) );
  nnd2s1 _28916_inst ( .DIN1(_29047), .DIN2(_29048), .Q(_29046) );
  xnr2s1 _28917_inst ( .DIN1(_29049), .DIN2(_29050), .Q(_29048) );
  nnd2s1 _28918_inst ( .DIN1(_29051), .DIN2(_29052), .Q(_29050) );
  nor2s1 _28919_inst ( .DIN1(_29053), .DIN2(_29054), .Q(_29052) );
  nor2s1 _28920_inst ( .DIN1(_53007), .DIN2(_26359), .Q(_29054) );
  nor2s1 _28921_inst ( .DIN1(_53426), .DIN2(_29055), .Q(_29053) );
  nnd2s1 _28922_inst ( .DIN1(_53007), .DIN2(_29056), .Q(_29055) );
  nor2s1 _28923_inst ( .DIN1(_29057), .DIN2(_29058), .Q(_29051) );
  nor2s1 _28924_inst ( .DIN1(_29059), .DIN2(_29056), .Q(_29058) );
  nor2s1 _28925_inst ( .DIN1(_29060), .DIN2(_29061), .Q(_29047) );
  and2s1 _28926_inst ( .DIN1(_29057), .DIN2(_52882), .Q(_29061) );
  nnd2s1 _28927_inst ( .DIN1(_29062), .DIN2(_29063), .Q(
        ______________________________67________) );
  nnd2s1 _28928_inst ( .DIN1(_29064), .DIN2(_29065), .Q(_29063) );
  xor2s1 _28929_inst ( .DIN1(_29066), .DIN2(_29067), .Q(_29065) );
  xor2s1 _28930_inst ( .DIN1(_52943), .DIN2(_53051), .Q(_29067) );
  nor2s1 _28931_inst ( .DIN1(_53007), .DIN2(_52941), .Q(_29066) );
  nnd2s1 _28932_inst ( .DIN1(_27782), .DIN2(_29068), .Q(_29062) );
  nnd2s1 _28933_inst ( .DIN1(_29069), .DIN2(_29070), .Q(_29068) );
  nor2s1 _28934_inst ( .DIN1(_29071), .DIN2(_29072), .Q(_29069) );
  nor2s1 _28935_inst ( .DIN1(_29057), .DIN2(_29073), .Q(_29072) );
  nor2s1 _28936_inst ( .DIN1(_53006), .DIN2(_26773), .Q(_29073) );
  and2s1 _28937_inst ( .DIN1(_29057), .DIN2(_53025), .Q(_29071) );
  nnd2s1 _28938_inst ( .DIN1(_27183), .DIN2(_29074), .Q(
        ______________________________66________) );
  nnd2s1 _28939_inst ( .DIN1(_29075), .DIN2(_29070), .Q(_29074) );
  nor2s1 _28940_inst ( .DIN1(_29076), .DIN2(_29077), .Q(_29075) );
  nor2s1 _28941_inst ( .DIN1(_53007), .DIN2(_29057), .Q(_29077) );
  nor2s1 _28942_inst ( .DIN1(_52912), .DIN2(_29078), .Q(_29076) );
  nnd2s1 _28943_inst ( .DIN1(_29079), .DIN2(_29080), .Q(
        ______________________________65________) );
  nnd2s1 _28944_inst ( .DIN1(_29081), .DIN2(_29082), .Q(_29080) );
  xor2s1 _28945_inst ( .DIN1(_53427), .DIN2(_53428), .Q(_29081) );
  nnd2s1 _28946_inst ( .DIN1(_29083), .DIN2(_29084), .Q(_29079) );
  nnd2s1 _28947_inst ( .DIN1(_29085), .DIN2(_29070), .Q(_29084) );
  nor2s1 _28948_inst ( .DIN1(_29086), .DIN2(_29087), .Q(_29085) );
  nor2s1 _28949_inst ( .DIN1(_29057), .DIN2(_29088), .Q(_29087) );
  nor2s1 _28950_inst ( .DIN1(_29089), .DIN2(_29090), .Q(_29088) );
  nor2s1 _28951_inst ( .DIN1(_26359), .DIN2(_29056), .Q(_29090) );
  nnd2s1 _28952_inst ( .DIN1(_52853), .DIN2(_53007), .Q(_29056) );
  and2s1 _28953_inst ( .DIN1(_26732), .DIN2(_29059), .Q(_29089) );
  nnd2s1 _28954_inst ( .DIN1(_53007), .DIN2(_53426), .Q(_29059) );
  and2s1 _28955_inst ( .DIN1(_29057), .DIN2(_52876), .Q(_29086) );
  nnd2s1 _28956_inst ( .DIN1(_29091), .DIN2(_29092), .Q(
        ______________________________64________) );
  nnd2s1 _28957_inst ( .DIN1(_29093), .DIN2(_29094), .Q(_29092) );
  nor2s1 _28958_inst ( .DIN1(_29095), .DIN2(_28646), .Q(_29093) );
  xor2s1 _28959_inst ( .DIN1(_53119), .DIN2(_26516), .Q(_29095) );
  nnd2s1 _28960_inst ( .DIN1(_29096), .DIN2(_29097), .Q(_29091) );
  nnd2s1 _28961_inst ( .DIN1(_29098), .DIN2(_29099), .Q(_29097) );
  nnd2s1 _28962_inst ( .DIN1(_29100), .DIN2(_29101), .Q(_29099) );
  xor2s1 _28963_inst ( .DIN1(_27157), .DIN2(_29102), .Q(_29100) );
  xor2s1 _28964_inst ( .DIN1(_26618), .DIN2(_29103), .Q(_29102) );
  nnd2s1 _28965_inst ( .DIN1(_29104), .DIN2(_29105), .Q(_29103) );
  nnd2s1 _28966_inst ( .DIN1(_29106), .DIN2(_26653), .Q(_29105) );
  nnd2s1 _28967_inst ( .DIN1(_27157), .DIN2(_29107), .Q(_29106) );
  or2s1 _28968_inst ( .DIN1(_29107), .DIN2(_26796), .Q(_29104) );
  nnd2s1 _28969_inst ( .DIN1(_29108), .DIN2(_26296), .Q(_29098) );
  nnd2s1 _28970_inst ( .DIN1(_29109), .DIN2(_29110), .Q(
        ______________________________63________) );
  nor2s1 _28971_inst ( .DIN1(_29111), .DIN2(_29112), .Q(_29110) );
  nor2s1 _28972_inst ( .DIN1(_28151), .DIN2(_29113), .Q(_29112) );
  nnd2s1 _28973_inst ( .DIN1(_29114), .DIN2(_29115), .Q(_29113) );
  nnd2s1 _28974_inst ( .DIN1(_29116), .DIN2(_29101), .Q(_29115) );
  xor2s1 _28975_inst ( .DIN1(_27157), .DIN2(_29117), .Q(_29116) );
  xor2s1 _28976_inst ( .DIN1(_26653), .DIN2(_29107), .Q(_29117) );
  nnd2s1 _28977_inst ( .DIN1(_29118), .DIN2(_29119), .Q(_29107) );
  nnd2s1 _28978_inst ( .DIN1(_29120), .DIN2(_26402), .Q(_29119) );
  or2s1 _28979_inst ( .DIN1(_29121), .DIN2(_26796), .Q(_29120) );
  nnd2s1 _28980_inst ( .DIN1(_27157), .DIN2(_29121), .Q(_29118) );
  nnd2s1 _28981_inst ( .DIN1(_29122), .DIN2(_29123), .Q(_29114) );
  nnd2s1 _28982_inst ( .DIN1(_29124), .DIN2(_29125), .Q(_29123) );
  nor2s1 _28983_inst ( .DIN1(_29126), .DIN2(_29127), .Q(_29125) );
  nor2s1 _28984_inst ( .DIN1(_29128), .DIN2(_27393), .Q(_29124) );
  nor2s1 _28985_inst ( .DIN1(_53126), .DIN2(_26296), .Q(_29128) );
  nor2s1 _28986_inst ( .DIN1(_28153), .DIN2(_29129), .Q(_29111) );
  nor2s1 _28987_inst ( .DIN1(_29130), .DIN2(_27651), .Q(_29129) );
  nor2s1 _28988_inst ( .DIN1(_29131), .DIN2(_26368), .Q(_29130) );
  nor2s1 _28989_inst ( .DIN1(_29132), .DIN2(_29133), .Q(_29109) );
  nor2s1 _28990_inst ( .DIN1(_52904), .DIN2(_29134), .Q(_29133) );
  nnd2s1 _28991_inst ( .DIN1(_29135), .DIN2(_29136), .Q(
        ______________________________62________) );
  nnd2s1 _28992_inst ( .DIN1(_29137), .DIN2(_29138), .Q(_29136) );
  xor2s1 _28993_inst ( .DIN1(_52923), .DIN2(_52925), .Q(_29138) );
  nnd2s1 _28994_inst ( .DIN1(_29139), .DIN2(_29140), .Q(_29135) );
  nnd2s1 _28995_inst ( .DIN1(_29141), .DIN2(_29142), .Q(_29140) );
  nnd2s1 _28996_inst ( .DIN1(_29101), .DIN2(_29143), .Q(_29142) );
  xor2s1 _28997_inst ( .DIN1(_27175), .DIN2(_29144), .Q(_29143) );
  xor2s1 _28998_inst ( .DIN1(_26402), .DIN2(_29121), .Q(_29144) );
  nnd2s1 _28999_inst ( .DIN1(_29145), .DIN2(_29146), .Q(_29121) );
  nnd2s1 _29000_inst ( .DIN1(_53106), .DIN2(_29147), .Q(_29146) );
  or2s1 _29001_inst ( .DIN1(_29148), .DIN2(_27209), .Q(_29147) );
  nnd2s1 _29002_inst ( .DIN1(_29148), .DIN2(_27209), .Q(_29145) );
  nnd2s1 _29003_inst ( .DIN1(_29149), .DIN2(_29122), .Q(_29141) );
  nnd2s1 _29004_inst ( .DIN1(_29150), .DIN2(_29108), .Q(_29149) );
  xnr2s1 _29005_inst ( .DIN1(_53181), .DIN2(_52955), .Q(_29150) );
  nnd2s1 _29006_inst ( .DIN1(_29151), .DIN2(_27113), .Q(
        ______________________________61________) );
  nor2s1 _29007_inst ( .DIN1(_29152), .DIN2(_29153), .Q(_29151) );
  nor2s1 _29008_inst ( .DIN1(_29154), .DIN2(_29155), .Q(_29153) );
  nnd2s1 _29009_inst ( .DIN1(_29156), .DIN2(_27108), .Q(_29155) );
  nnd2s1 _29010_inst ( .DIN1(_29157), .DIN2(_29158), .Q(_27108) );
  nor2s1 _29011_inst ( .DIN1(_27058), .DIN2(_27360), .Q(_29158) );
  nor2s1 _29012_inst ( .DIN1(_29159), .DIN2(_27013), .Q(_29157) );
  nor2s1 _29013_inst ( .DIN1(_29160), .DIN2(_29161), .Q(_29156) );
  nor2s1 _29014_inst ( .DIN1(_27101), .DIN2(_29162), .Q(_29161) );
  xnr2s1 _29015_inst ( .DIN1(_29148), .DIN2(_29163), .Q(_29162) );
  xnr2s1 _29016_inst ( .DIN1(_53106), .DIN2(_27209), .Q(_29163) );
  nnd2s1 _29017_inst ( .DIN1(_27175), .DIN2(_29164), .Q(_27209) );
  nnd2s1 _29018_inst ( .DIN1(_29165), .DIN2(_29166), .Q(_29164) );
  hi1s1 _29019_inst ( .DIN(_27157), .Q(_27175) );
  xor2s1 _29020_inst ( .DIN1(_29167), .DIN2(_29168), .Q(_27157) );
  nnd2s1 _29021_inst ( .DIN1(_26836), .DIN2(_29170), .Q(_29167) );
  nnd2s1 _29022_inst ( .DIN1(_29171), .DIN2(_29172), .Q(_29148) );
  nnd2s1 _29023_inst ( .DIN1(_29173), .DIN2(_26752), .Q(_29172) );
  nnd2s1 _29024_inst ( .DIN1(_29174), .DIN2(_27223), .Q(_29173) );
  xor2s1 _29025_inst ( .DIN1(_26998), .DIN2(_29175), .Q(_29171) );
  or2s1 _29026_inst ( .DIN1(_27223), .DIN2(_29174), .Q(_29175) );
  nor2s1 _29027_inst ( .DIN1(_27058), .DIN2(_29176), .Q(_29160) );
  nor2s1 _29028_inst ( .DIN1(_27651), .DIN2(_29177), .Q(_29176) );
  xor2s1 _29029_inst ( .DIN1(_26299), .DIN2(_29178), .Q(_29177) );
  nnd2s1 _29030_inst ( .DIN1(_52859), .DIN2(_52860), .Q(_29178) );
  nor2s1 _29031_inst ( .DIN1(_27105), .DIN2(_29179), .Q(_29152) );
  nor2s1 _29032_inst ( .DIN1(_27061), .DIN2(_27048), .Q(_29179) );
  hi1s1 _29033_inst ( .DIN(_27091), .Q(_27048) );
  nnd2s1 _29034_inst ( .DIN1(_52866), .DIN2(_52872), .Q(_27091) );
  nor2s1 _29035_inst ( .DIN1(_52872), .DIN2(_52866), .Q(_27061) );
  nnd2s1 _29036_inst ( .DIN1(_29180), .DIN2(_29181), .Q(
        ______________________________60________) );
  nor2s1 _29037_inst ( .DIN1(_29182), .DIN2(_29183), .Q(_29180) );
  nor2s1 _29038_inst ( .DIN1(_29184), .DIN2(_29185), .Q(_29183) );
  nnd2s1 _29039_inst ( .DIN1(_29186), .DIN2(_29187), .Q(_29185) );
  nnd2s1 _29040_inst ( .DIN1(_27058), .DIN2(_29188), .Q(_29187) );
  xnr2s1 _29041_inst ( .DIN1(_29174), .DIN2(_29189), .Q(_29188) );
  xor2s1 _29042_inst ( .DIN1(_27223), .DIN2(_52890), .Q(_29189) );
  nnd2s1 _29043_inst ( .DIN1(_29170), .DIN2(_29190), .Q(_27223) );
  nnd2s1 _29044_inst ( .DIN1(_15544), .DIN2(_29191), .Q(_29190) );
  hi1s1 _29045_inst ( .DIN(_29165), .Q(_29170) );
  nor2s1 _29046_inst ( .DIN1(_29191), .DIN2(_15544), .Q(_29165) );
  and2s1 _29047_inst ( .DIN1(_29192), .DIN2(_29193), .Q(_29174) );
  nnd2s1 _29048_inst ( .DIN1(_29194), .DIN2(_26655), .Q(_29193) );
  nnd2s1 _29049_inst ( .DIN1(_29195), .DIN2(_29196), .Q(_29194) );
  or2s1 _29050_inst ( .DIN1(_29196), .DIN2(_29195), .Q(_29192) );
  nnd2s1 _29051_inst ( .DIN1(_29197), .DIN2(______[10]), .Q(_29186) );
  nor2s1 _29052_inst ( .DIN1(_29198), .DIN2(_27063), .Q(_29197) );
  nnd2s1 _29053_inst ( .DIN1(_29199), .DIN2(_27101), .Q(_27063) );
  hi1s1 _29054_inst ( .DIN(_27058), .Q(_27101) );
  nor2s1 _29055_inst ( .DIN1(_29200), .DIN2(_27004), .Q(_27058) );
  nnd2s1 _29056_inst ( .DIN1(_29201), .DIN2(_27412), .Q(_29199) );
  hi1s1 _29057_inst ( .DIN(_27013), .Q(_27412) );
  nnd2s1 _29058_inst ( .DIN1(_27332), .DIN2(_29202), .Q(_27013) );
  nor2s1 _29059_inst ( .DIN1(_29203), .DIN2(_29204), .Q(_29202) );
  nor2s1 _29060_inst ( .DIN1(_29205), .DIN2(_27343), .Q(_27332) );
  nor2s1 _29061_inst ( .DIN1(_27360), .DIN2(_29159), .Q(_29201) );
  xnr2s1 _29062_inst ( .DIN1(_52857), .DIN2(_52860), .Q(_29198) );
  nor2s1 _29063_inst ( .DIN1(_29206), .DIN2(_29207), .Q(_29182) );
  xor2s1 _29064_inst ( .DIN1(_29208), .DIN2(_29209), .Q(_29207) );
  xor2s1 _29065_inst ( .DIN1(_53100), .DIN2(_53180), .Q(_29209) );
  nnd2s1 _29066_inst ( .DIN1(_52859), .DIN2(_52881), .Q(_29208) );
  nnd2s1 _29067_inst ( .DIN1(_29210), .DIN2(_29211), .Q(
        ______________________________5________) );
  nnd2s1 _29068_inst ( .DIN1(_29212), .DIN2(_29213), .Q(_29211) );
  xor2s1 _29069_inst ( .DIN1(_29214), .DIN2(_53049), .Q(_29213) );
  nnd2s1 _29070_inst ( .DIN1(_53315), .DIN2(_53325), .Q(_29214) );
  nor2s1 _29071_inst ( .DIN1(_29215), .DIN2(_27651), .Q(_29212) );
  nnd2s1 _29072_inst ( .DIN1(_28542), .DIN2(_29216), .Q(_29210) );
  nnd2s1 _29073_inst ( .DIN1(_29217), .DIN2(_29218), .Q(_29216) );
  nnd2s1 _29074_inst ( .DIN1(_29219), .DIN2(_28809), .Q(_29218) );
  nor2s1 _29075_inst ( .DIN1(_28808), .DIN2(_29027), .Q(_29219) );
  nor2s1 _29076_inst ( .DIN1(_26568), .DIN2(_26301), .Q(_29027) );
  nor2s1 _29077_inst ( .DIN1(_52874), .DIN2(_52965), .Q(_28808) );
  nnd2s1 _29078_inst ( .DIN1(_28935), .DIN2(_26572), .Q(_29217) );
  nnd2s1 _29079_inst ( .DIN1(_29220), .DIN2(_29221), .Q(
        ______________________________59________) );
  nor2s1 _29080_inst ( .DIN1(_29222), .DIN2(_29223), .Q(_29220) );
  nor2s1 _29081_inst ( .DIN1(_29224), .DIN2(_29225), .Q(_29223) );
  xor2s1 _29082_inst ( .DIN1(_29195), .DIN2(_29226), .Q(_29225) );
  xor2s1 _29083_inst ( .DIN1(_26655), .DIN2(_29196), .Q(_29226) );
  nnd2s1 _29084_inst ( .DIN1(_29227), .DIN2(_29228), .Q(_29196) );
  nnd2s1 _29085_inst ( .DIN1(_52889), .DIN2(_29229), .Q(_29228) );
  or2s1 _29086_inst ( .DIN1(_27238), .DIN2(_29230), .Q(_29229) );
  nnd2s1 _29087_inst ( .DIN1(_29230), .DIN2(_27238), .Q(_29227) );
  xnr2s1 _29088_inst ( .DIN1(_27232), .DIN2(_29231), .Q(_29195) );
  nnd2s1 _29089_inst ( .DIN1(_29191), .DIN2(_29232), .Q(_27232) );
  nnd2s1 _29090_inst ( .DIN1(_359), .DIN2(_29233), .Q(_29232) );
  or2s1 _29091_inst ( .DIN1(_29233), .DIN2(_359), .Q(_29191) );
  nor2s1 _29092_inst ( .DIN1(_29234), .DIN2(_29235), .Q(_29222) );
  and2s1 _29093_inst ( .DIN1(_29236), .DIN2(_52859), .Q(_29235) );
  nnd2s1 _29094_inst ( .DIN1(_29237), .DIN2(_27050), .Q(
        ______________________________58________) );
  nor2s1 _29095_inst ( .DIN1(_29238), .DIN2(_29239), .Q(_29237) );
  nor2s1 _29096_inst ( .DIN1(_27053), .DIN2(_29240), .Q(_29239) );
  nor2s1 _29097_inst ( .DIN1(_29241), .DIN2(_29242), .Q(_29240) );
  nor2s1 _29098_inst ( .DIN1(_29224), .DIN2(_29243), .Q(_29242) );
  xor2s1 _29099_inst ( .DIN1(_29244), .DIN2(_29230), .Q(_29243) );
  and2s1 _29100_inst ( .DIN1(_29245), .DIN2(_29246), .Q(_29230) );
  nnd2s1 _29101_inst ( .DIN1(_52887), .DIN2(_29247), .Q(_29246) );
  or2s1 _29102_inst ( .DIN1(_29248), .DIN2(_27254), .Q(_29247) );
  nnd2s1 _29103_inst ( .DIN1(_27254), .DIN2(_29248), .Q(_29245) );
  xor2s1 _29104_inst ( .DIN1(_27238), .DIN2(_52889), .Q(_29244) );
  nnd2s1 _29105_inst ( .DIN1(_29233), .DIN2(_29249), .Q(_27238) );
  nnd2s1 _29106_inst ( .DIN1(_15546), .DIN2(_29250), .Q(_29249) );
  or2s1 _29107_inst ( .DIN1(_29250), .DIN2(_15546), .Q(_29233) );
  nnd2s1 _29108_inst ( .DIN1(_29251), .DIN2(_29252), .Q(_29250) );
  nor2s1 _29109_inst ( .DIN1(_29234), .DIN2(_29253), .Q(_29241) );
  nnd2s1 _29110_inst ( .DIN1(_29254), .DIN2(_29236), .Q(_29253) );
  xor2s1 _29111_inst ( .DIN1(_52859), .DIN2(_52860), .Q(_29254) );
  nor2s1 _29112_inst ( .DIN1(_52905), .DIN2(_27064), .Q(_29238) );
  nnd2s1 _29113_inst ( .DIN1(_29255), .DIN2(_29256), .Q(
        ______________________________57________) );
  nor2s1 _29114_inst ( .DIN1(_29257), .DIN2(_29258), .Q(_29256) );
  nor2s1 _29115_inst ( .DIN1(_29259), .DIN2(_29260), .Q(_29258) );
  nnd2s1 _29116_inst ( .DIN1(_29261), .DIN2(______[0]), .Q(_29260) );
  xor2s1 _29117_inst ( .DIN1(_52864), .DIN2(_29262), .Q(_29259) );
  nor2s1 _29118_inst ( .DIN1(_29263), .DIN2(_29264), .Q(_29255) );
  nnd2s1 _29119_inst ( .DIN1(_29265), .DIN2(_29266), .Q(_29264) );
  or2s1 _29120_inst ( .DIN1(_29267), .DIN2(_26293), .Q(_29266) );
  nnd2s1 _29121_inst ( .DIN1(_29268), .DIN2(_26293), .Q(_29265) );
  nnd2s1 _29122_inst ( .DIN1(_29269), .DIN2(_29270), .Q(_29268) );
  nnd2s1 _29123_inst ( .DIN1(_29271), .DIN2(_52862), .Q(_29270) );
  nor2s1 _29124_inst ( .DIN1(_29272), .DIN2(_29273), .Q(_29263) );
  xnr2s1 _29125_inst ( .DIN1(_27254), .DIN2(_29274), .Q(_29273) );
  xnr2s1 _29126_inst ( .DIN1(_52887), .DIN2(_29248), .Q(_29274) );
  nnd2s1 _29127_inst ( .DIN1(_29275), .DIN2(_29276), .Q(_29248) );
  nnd2s1 _29128_inst ( .DIN1(_29277), .DIN2(_26389), .Q(_29276) );
  or2s1 _29129_inst ( .DIN1(_29278), .DIN2(_27277), .Q(_29277) );
  nnd2s1 _29130_inst ( .DIN1(_27277), .DIN2(_29278), .Q(_29275) );
  xor2s1 _29131_inst ( .DIN1(_29251), .DIN2(_29252), .Q(_27254) );
  nor2s1 _29132_inst ( .DIN1(_29279), .DIN2(_356), .Q(_29251) );
  nnd2s1 _29133_inst ( .DIN1(_29280), .DIN2(_29281), .Q(
        ______________________________56________) );
  nor2s1 _29134_inst ( .DIN1(_29257), .DIN2(_29282), .Q(_29281) );
  nor2s1 _29135_inst ( .DIN1(_29283), .DIN2(_29284), .Q(_29282) );
  nnd2s1 _29136_inst ( .DIN1(_29261), .DIN2(______[30]), .Q(_29284) );
  and2s1 _29137_inst ( .DIN1(_29154), .DIN2(_29285), .Q(_29261) );
  nnd2s1 _29138_inst ( .DIN1(_29286), .DIN2(_29287), .Q(_29285) );
  nor2s1 _29139_inst ( .DIN1(_29288), .DIN2(_29289), .Q(_29287) );
  xor2s1 _29140_inst ( .DIN1(_52861), .DIN2(_29262), .Q(_29283) );
  nor2s1 _29141_inst ( .DIN1(_29290), .DIN2(_29291), .Q(_29280) );
  nnd2s1 _29142_inst ( .DIN1(_29292), .DIN2(_29293), .Q(_29291) );
  or2s1 _29143_inst ( .DIN1(_29269), .DIN2(_52861), .Q(_29293) );
  hi1s1 _29144_inst ( .DIN(_29294), .Q(_29269) );
  nnd2s1 _29145_inst ( .DIN1(_29295), .DIN2(_52861), .Q(_29292) );
  and2s1 _29146_inst ( .DIN1(_29271), .DIN2(_52863), .Q(_29295) );
  hi1s1 _29147_inst ( .DIN(_29296), .Q(_29271) );
  nor2s1 _29148_inst ( .DIN1(_29272), .DIN2(_29297), .Q(_29290) );
  xor2s1 _29149_inst ( .DIN1(_27277), .DIN2(_29298), .Q(_29297) );
  xor2s1 _29150_inst ( .DIN1(_26389), .DIN2(_29278), .Q(_29298) );
  nnd2s1 _29151_inst ( .DIN1(_29299), .DIN2(_29300), .Q(_29278) );
  nnd2s1 _29152_inst ( .DIN1(_29301), .DIN2(_26234), .Q(_29300) );
  or2s1 _29153_inst ( .DIN1(_29302), .DIN2(_27297), .Q(_29301) );
  nnd2s1 _29154_inst ( .DIN1(_27297), .DIN2(_29302), .Q(_29299) );
  xor2s1 _29155_inst ( .DIN1(_29279), .DIN2(_356), .Q(_27277) );
  nnd2s1 _29156_inst ( .DIN1(_29303), .DIN2(_29304), .Q(_29279) );
  nor2s1 _29157_inst ( .DIN1(_28218), .DIN2(_29305), .Q(
        ______________________________55________) );
  nnd2s1 _29158_inst ( .DIN1(_29306), .DIN2(_29307), .Q(_29305) );
  nnd2s1 _29159_inst ( .DIN1(_29308), .DIN2(_29224), .Q(_29307) );
  nnd2s1 _29160_inst ( .DIN1(_29236), .DIN2(_26666), .Q(_29308) );
  nnd2s1 _29161_inst ( .DIN1(_29309), .DIN2(_29234), .Q(_29306) );
  xnr2s1 _29162_inst ( .DIN1(_27297), .DIN2(_29310), .Q(_29309) );
  xor2s1 _29163_inst ( .DIN1(_26234), .DIN2(_29302), .Q(_29310) );
  nnd2s1 _29164_inst ( .DIN1(_29311), .DIN2(_29312), .Q(_29302) );
  nnd2s1 _29165_inst ( .DIN1(_29313), .DIN2(_26674), .Q(_29312) );
  nnd2s1 _29166_inst ( .DIN1(_29314), .DIN2(_27323), .Q(_29313) );
  or2s1 _29167_inst ( .DIN1(_27323), .DIN2(_29314), .Q(_29311) );
  xor2s1 _29168_inst ( .DIN1(_29315), .DIN2(_355), .Q(_27297) );
  nnd2s1 _29169_inst ( .DIN1(_29316), .DIN2(_29317), .Q(
        ______________________________54________) );
  nor2s1 _29170_inst ( .DIN1(_29318), .DIN2(_29319), .Q(_29317) );
  nnd2s1 _29171_inst ( .DIN1(_29320), .DIN2(_29321), .Q(_29319) );
  hi1s1 _29172_inst ( .DIN(_29257), .Q(_29321) );
  nor2s1 _29173_inst ( .DIN1(_29236), .DIN2(_29296), .Q(_29257) );
  nnd2s1 _29174_inst ( .DIN1(_29322), .DIN2(_29323), .Q(_29236) );
  hi1s1 _29175_inst ( .DIN(_27343), .Q(_29323) );
  and2s1 _29176_inst ( .DIN1(_27470), .DIN2(_27496), .Q(_29322) );
  nor2s1 _29177_inst ( .DIN1(_29324), .DIN2(_29325), .Q(_27496) );
  hi1s1 _29178_inst ( .DIN(_27360), .Q(_27470) );
  nnd2s1 _29179_inst ( .DIN1(_29326), .DIN2(_29327), .Q(_29320) );
  xor2s1 _29180_inst ( .DIN1(_29314), .DIN2(_29328), .Q(_29327) );
  xor2s1 _29181_inst ( .DIN1(_27323), .DIN2(_52918), .Q(_29328) );
  nnd2s1 _29182_inst ( .DIN1(_29315), .DIN2(_29329), .Q(_27323) );
  nnd2s1 _29183_inst ( .DIN1(_353), .DIN2(_29330), .Q(_29329) );
  hi1s1 _29184_inst ( .DIN(_29303), .Q(_29315) );
  nor2s1 _29185_inst ( .DIN1(_29330), .DIN2(_353), .Q(_29303) );
  nnd2s1 _29186_inst ( .DIN1(_29331), .DIN2(_29332), .Q(_29330) );
  nnd2s1 _29187_inst ( .DIN1(_29333), .DIN2(_29334), .Q(_29314) );
  nnd2s1 _29188_inst ( .DIN1(_52930), .DIN2(_29335), .Q(_29334) );
  nnd2s1 _29189_inst ( .DIN1(_29336), .DIN2(_29337), .Q(_29335) );
  or2s1 _29190_inst ( .DIN1(_29337), .DIN2(_29336), .Q(_29333) );
  hi1s1 _29191_inst ( .DIN(_29272), .Q(_29326) );
  nnd2s1 _29192_inst ( .DIN1(_29234), .DIN2(_27105), .Q(_29272) );
  hi1s1 _29193_inst ( .DIN(_29224), .Q(_29234) );
  nnd2s1 _29194_inst ( .DIN1(_29267), .DIN2(_27113), .Q(_29318) );
  nnd2s1 _29195_inst ( .DIN1(_29338), .DIN2(_52863), .Q(_29267) );
  nor2s1 _29196_inst ( .DIN1(_52862), .DIN2(_29296), .Q(_29338) );
  nor2s1 _29197_inst ( .DIN1(_29339), .DIN2(_29340), .Q(_29316) );
  nnd2s1 _29198_inst ( .DIN1(_29341), .DIN2(_29342), .Q(_29340) );
  nnd2s1 _29199_inst ( .DIN1(_29343), .DIN2(_29154), .Q(_29342) );
  nnd2s1 _29200_inst ( .DIN1(_52862), .DIN2(______[30]), .Q(_29343) );
  nnd2s1 _29201_inst ( .DIN1(_29294), .DIN2(_52862), .Q(_29341) );
  nor2s1 _29202_inst ( .DIN1(_29296), .DIN2(_52863), .Q(_29294) );
  nor2s1 _29203_inst ( .DIN1(______[14]), .DIN2(_29296), .Q(_29339) );
  nnd2s1 _29204_inst ( .DIN1(_27105), .DIN2(_29224), .Q(_29296) );
  nnd2s1 _29205_inst ( .DIN1(_29344), .DIN2(_29345), .Q(_29224) );
  nor2s1 _29206_inst ( .DIN1(_29346), .DIN2(_29200), .Q(_29344) );
  nnd2s1 _29207_inst ( .DIN1(_29347), .DIN2(_29348), .Q(_29200) );
  nor2s1 _29208_inst ( .DIN1(_27296), .DIN2(_29349), .Q(_29348) );
  nnd2s1 _29209_inst ( .DIN1(_27497), .DIN2(_27335), .Q(_29349) );
  nor2s1 _29210_inst ( .DIN1(_29324), .DIN2(_29350), .Q(_29347) );
  nnd2s1 _29211_inst ( .DIN1(_27471), .DIN2(_29351), .Q(_29350) );
  nnd2s1 _29212_inst ( .DIN1(_29352), .DIN2(_29353), .Q(_29324) );
  nor2s1 _29213_inst ( .DIN1(_29354), .DIN2(_29204), .Q(_29352) );
  nnd2s1 _29214_inst ( .DIN1(_29355), .DIN2(_28045), .Q(
        ______________________________53________) );
  nor2s1 _29215_inst ( .DIN1(_29356), .DIN2(_29357), .Q(_29355) );
  nor2s1 _29216_inst ( .DIN1(_29358), .DIN2(_28049), .Q(_29357) );
  nor2s1 _29217_inst ( .DIN1(_29359), .DIN2(_29360), .Q(_29358) );
  nor2s1 _29218_inst ( .DIN1(_29361), .DIN2(_29362), .Q(_29360) );
  xor2s1 _29219_inst ( .DIN1(_27337), .DIN2(_29363), .Q(_29361) );
  xnr2s1 _29220_inst ( .DIN1(_52930), .DIN2(_29337), .Q(_29363) );
  nnd2s1 _29221_inst ( .DIN1(_29364), .DIN2(_29365), .Q(_29337) );
  nnd2s1 _29222_inst ( .DIN1(_29366), .DIN2(_26637), .Q(_29365) );
  nnd2s1 _29223_inst ( .DIN1(_27368), .DIN2(_29367), .Q(_29366) );
  or2s1 _29224_inst ( .DIN1(_27368), .DIN2(_29367), .Q(_29364) );
  hi1s1 _29225_inst ( .DIN(_29336), .Q(_27337) );
  xnr2s1 _29226_inst ( .DIN1(_29368), .DIN2(_29332), .Q(_29336) );
  nor2s1 _29227_inst ( .DIN1(_29369), .DIN2(_29370), .Q(_29359) );
  xor2s1 _29228_inst ( .DIN1(_52864), .DIN2(_29371), .Q(_29370) );
  nor2s1 _29229_inst ( .DIN1(_28056), .DIN2(_26345), .Q(_29356) );
  nnd2s1 _29230_inst ( .DIN1(_29372), .DIN2(_29373), .Q(
        ______________________________52________) );
  nnd2s1 _29231_inst ( .DIN1(_28250), .DIN2(_29374), .Q(_29373) );
  nnd2s1 _29232_inst ( .DIN1(_29375), .DIN2(_29376), .Q(_29374) );
  nnd2s1 _29233_inst ( .DIN1(_29377), .DIN2(_29378), .Q(_29376) );
  xor2s1 _29234_inst ( .DIN1(_29379), .DIN2(_53413), .Q(_29377) );
  nnd2s1 _29235_inst ( .DIN1(_29380), .DIN2(_29381), .Q(_29375) );
  xor2s1 _29236_inst ( .DIN1(_29367), .DIN2(_29382), .Q(_29380) );
  xor2s1 _29237_inst ( .DIN1(_26637), .DIN2(_27368), .Q(_29382) );
  nnd2s1 _29238_inst ( .DIN1(_29368), .DIN2(_29383), .Q(_27368) );
  nnd2s1 _29239_inst ( .DIN1(_15550), .DIN2(_29384), .Q(_29383) );
  hi1s1 _29240_inst ( .DIN(_29331), .Q(_29368) );
  nor2s1 _29241_inst ( .DIN1(_29384), .DIN2(_15550), .Q(_29331) );
  or2s1 _29242_inst ( .DIN1(_29385), .DIN2(_15551), .Q(_29384) );
  nnd2s1 _29243_inst ( .DIN1(_29386), .DIN2(_29387), .Q(_29367) );
  nnd2s1 _29244_inst ( .DIN1(_29388), .DIN2(_26667), .Q(_29387) );
  nnd2s1 _29245_inst ( .DIN1(_27380), .DIN2(_29389), .Q(_29388) );
  or2s1 _29246_inst ( .DIN1(_29389), .DIN2(_27380), .Q(_29386) );
  nnd2s1 _29247_inst ( .DIN1(_29390), .DIN2(_52850), .Q(_29372) );
  nnd2s1 _29248_inst ( .DIN1(_29391), .DIN2(_29392), .Q(
        ______________________________51________) );
  nnd2s1 _29249_inst ( .DIN1(_29393), .DIN2(_29039), .Q(_29392) );
  and2s1 _29250_inst ( .DIN1(______[10]), .DIN2(_52900), .Q(_29393) );
  nnd2s1 _29251_inst ( .DIN1(_28738), .DIN2(_29394), .Q(_29391) );
  nnd2s1 _29252_inst ( .DIN1(_29395), .DIN2(_29396), .Q(_29394) );
  nnd2s1 _29253_inst ( .DIN1(_29397), .DIN2(_29378), .Q(_29396) );
  nor2s1 _29254_inst ( .DIN1(_28100), .DIN2(_26305), .Q(_29397) );
  nnd2s1 _29255_inst ( .DIN1(_29381), .DIN2(_29398), .Q(_29395) );
  xnr2s1 _29256_inst ( .DIN1(_27380), .DIN2(_29399), .Q(_29398) );
  xor2s1 _29257_inst ( .DIN1(_26667), .DIN2(_29389), .Q(_29399) );
  nnd2s1 _29258_inst ( .DIN1(_29400), .DIN2(_29401), .Q(_29389) );
  nnd2s1 _29259_inst ( .DIN1(_53162), .DIN2(_29402), .Q(_29401) );
  or2s1 _29260_inst ( .DIN1(_29403), .DIN2(_27403), .Q(_29402) );
  nnd2s1 _29261_inst ( .DIN1(_27403), .DIN2(_29403), .Q(_29400) );
  xnr2s1 _29262_inst ( .DIN1(_29385), .DIN2(_29404), .Q(_27380) );
  nnd2s1 _29263_inst ( .DIN1(_29405), .DIN2(_27113), .Q(
        ______________________________50________) );
  nnd2s1 _29264_inst ( .DIN1(_29286), .DIN2(_29406), .Q(_27113) );
  nor2s1 _29265_inst ( .DIN1(_27105), .DIN2(_29407), .Q(_29406) );
  nnd2s1 _29266_inst ( .DIN1(_27445), .DIN2(_29408), .Q(_29407) );
  nor2s1 _29267_inst ( .DIN1(_27431), .DIN2(_29409), .Q(_29286) );
  nor2s1 _29268_inst ( .DIN1(_29410), .DIN2(_29411), .Q(_29405) );
  nor2s1 _29269_inst ( .DIN1(_29154), .DIN2(_29412), .Q(_29411) );
  nnd2s1 _29270_inst ( .DIN1(_29413), .DIN2(_29414), .Q(_29412) );
  nnd2s1 _29271_inst ( .DIN1(_29415), .DIN2(_29381), .Q(_29414) );
  xnr2s1 _29272_inst ( .DIN1(_29416), .DIN2(_29403), .Q(_29415) );
  nnd2s1 _29273_inst ( .DIN1(_29417), .DIN2(_29418), .Q(_29403) );
  nnd2s1 _29274_inst ( .DIN1(_29419), .DIN2(_26486), .Q(_29418) );
  or2s1 _29275_inst ( .DIN1(_29420), .DIN2(_27420), .Q(_29419) );
  nnd2s1 _29276_inst ( .DIN1(_27420), .DIN2(_29420), .Q(_29417) );
  xnr2s1 _29277_inst ( .DIN1(_27403), .DIN2(_53162), .Q(_29416) );
  and2s1 _29278_inst ( .DIN1(_29421), .DIN2(_29385), .Q(_27403) );
  nnd2s1 _29279_inst ( .DIN1(_29422), .DIN2(_29423), .Q(_29385) );
  nor2s1 _29280_inst ( .DIN1(_398), .DIN2(_26205), .Q(_29422) );
  nnd2s1 _29281_inst ( .DIN1(_26205), .DIN2(_29424), .Q(_29421) );
  nnd2s1 _29282_inst ( .DIN1(_29423), .DIN2(_29425), .Q(_29424) );
  nnd2s1 _29283_inst ( .DIN1(_29426), .DIN2(_29427), .Q(_29413) );
  nor2s1 _29284_inst ( .DIN1(_29371), .DIN2(_29428), .Q(_29427) );
  nor2s1 _29285_inst ( .DIN1(_52898), .DIN2(_53396), .Q(_29428) );
  hi1s1 _29286_inst ( .DIN(_29379), .Q(_29371) );
  nnd2s1 _29287_inst ( .DIN1(_53396), .DIN2(_52898), .Q(_29379) );
  nor2s1 _29288_inst ( .DIN1(_26774), .DIN2(_29369), .Q(_29426) );
  nor2s1 _29289_inst ( .DIN1(_27105), .DIN2(_29429), .Q(_29410) );
  nor2s1 _29290_inst ( .DIN1(_29430), .DIN2(_29262), .Q(_29429) );
  nor2s1 _29291_inst ( .DIN1(_26293), .DIN2(_26666), .Q(_29262) );
  nor2s1 _29292_inst ( .DIN1(_52862), .DIN2(_52865), .Q(_29430) );
  hi1s1 _29293_inst ( .DIN(_29154), .Q(_27105) );
  nnd2s1 _29294_inst ( .DIN1(_29431), .DIN2(_29432), .Q(_29154) );
  nor2s1 _29295_inst ( .DIN1(_29433), .DIN2(_27310), .Q(_29432) );
  nor2s1 _29296_inst ( .DIN1(_29289), .DIN2(_29434), .Q(_29431) );
  hi1s1 _29297_inst ( .DIN(_27445), .Q(_29289) );
  nnd2s1 _29298_inst ( .DIN1(_29435), .DIN2(_29436), .Q(
        ______________________________4________) );
  nor2s1 _29299_inst ( .DIN1(_29437), .DIN2(_29438), .Q(_29436) );
  nor2s1 _29300_inst ( .DIN1(_27144), .DIN2(_29439), .Q(_29438) );
  nnd2s1 _29301_inst ( .DIN1(_29440), .DIN2(_29441), .Q(_29439) );
  nnd2s1 _29302_inst ( .DIN1(_29442), .DIN2(_28809), .Q(_29441) );
  xor2s1 _29303_inst ( .DIN1(_29443), .DIN2(_29444), .Q(_29442) );
  xor2s1 _29304_inst ( .DIN1(_52881), .DIN2(_52896), .Q(_29444) );
  nnd2s1 _29305_inst ( .DIN1(_52879), .DIN2(_26360), .Q(_29443) );
  nnd2s1 _29306_inst ( .DIN1(_28935), .DIN2(_26715), .Q(_29440) );
  nor2s1 _29307_inst ( .DIN1(______[6]), .DIN2(_27146), .Q(_29437) );
  nor2s1 _29308_inst ( .DIN1(_29445), .DIN2(_27149), .Q(_29435) );
  nnd2s1 _29309_inst ( .DIN1(_28284), .DIN2(_29446), .Q(_27149) );
  nnd2s1 _29310_inst ( .DIN1(_29447), .DIN2(_53250), .Q(_29446) );
  nor2s1 _29311_inst ( .DIN1(_53246), .DIN2(_27146), .Q(_29447) );
  hi1s1 _29312_inst ( .DIN(_27150), .Q(_29445) );
  nnd2s1 _29313_inst ( .DIN1(_29448), .DIN2(_53246), .Q(_27150) );
  nor2s1 _29314_inst ( .DIN1(_53250), .DIN2(_27146), .Q(_29448) );
  nnd2s1 _29315_inst ( .DIN1(_27723), .DIN2(_29449), .Q(
        ______________________________49________) );
  xor2s1 _29316_inst ( .DIN1(_29450), .DIN2(_29451), .Q(_29449) );
  nnd2s1 _29317_inst ( .DIN1(_29452), .DIN2(_29453), .Q(_29451) );
  nnd2s1 _29318_inst ( .DIN1(_29454), .DIN2(_29378), .Q(_29453) );
  hi1s1 _29319_inst ( .DIN(_29369), .Q(_29378) );
  nnd2s1 _29320_inst ( .DIN1(_29362), .DIN2(_29455), .Q(_29369) );
  or2s1 _29321_inst ( .DIN1(_27344), .DIN2(_29204), .Q(_29455) );
  nor2s1 _29322_inst ( .DIN1(_29456), .DIN2(_27039), .Q(_29454) );
  xnr2s1 _29323_inst ( .DIN1(_52931), .DIN2(_29457), .Q(_29456) );
  nnd2s1 _29324_inst ( .DIN1(_29381), .DIN2(_29458), .Q(_29452) );
  xor2s1 _29325_inst ( .DIN1(_27420), .DIN2(_29459), .Q(_29458) );
  xor2s1 _29326_inst ( .DIN1(_26486), .DIN2(_29420), .Q(_29459) );
  nnd2s1 _29327_inst ( .DIN1(_29460), .DIN2(_29461), .Q(_29420) );
  nnd2s1 _29328_inst ( .DIN1(_29462), .DIN2(_26475), .Q(_29461) );
  nnd2s1 _29329_inst ( .DIN1(_29463), .DIN2(_29464), .Q(_29462) );
  nnd2s1 _29330_inst ( .DIN1(_27436), .DIN2(_29465), .Q(_29460) );
  hi1s1 _29331_inst ( .DIN(_29463), .Q(_29465) );
  hi1s1 _29332_inst ( .DIN(_29464), .Q(_27436) );
  xor2s1 _29333_inst ( .DIN1(_29466), .DIN2(_398), .Q(_27420) );
  hi1s1 _29334_inst ( .DIN(_28925), .Q(_27723) );
  nnd2s1 _29335_inst ( .DIN1(_29467), .DIN2(_29468), .Q(
        ______________________________48________) );
  nnd2s1 _29336_inst ( .DIN1(_29094), .DIN2(_29469), .Q(_29468) );
  xor2s1 _29337_inst ( .DIN1(_53093), .DIN2(_53351), .Q(_29469) );
  nnd2s1 _29338_inst ( .DIN1(_29470), .DIN2(_29096), .Q(_29467) );
  nor2s1 _29339_inst ( .DIN1(_29471), .DIN2(_29472), .Q(_29470) );
  nor2s1 _29340_inst ( .DIN1(_29381), .DIN2(_29473), .Q(_29472) );
  nnd2s1 _29341_inst ( .DIN1(_29474), .DIN2(______[8]), .Q(_29473) );
  nor2s1 _29342_inst ( .DIN1(_29475), .DIN2(_29476), .Q(_29474) );
  xor2s1 _29343_inst ( .DIN1(_52867), .DIN2(_52868), .Q(_29476) );
  nor2s1 _29344_inst ( .DIN1(_29204), .DIN2(_27344), .Q(_29475) );
  nnd2s1 _29345_inst ( .DIN1(_29477), .DIN2(_29478), .Q(_27344) );
  nor2s1 _29346_inst ( .DIN1(_29479), .DIN2(_29480), .Q(_29478) );
  nnd2s1 _29347_inst ( .DIN1(_29481), .DIN2(_27492), .Q(_29480) );
  nnd2s1 _29348_inst ( .DIN1(_29482), .DIN2(_27336), .Q(_29479) );
  nor2s1 _29349_inst ( .DIN1(_29483), .DIN2(_29484), .Q(_29477) );
  or2s1 _29350_inst ( .DIN1(_29205), .DIN2(_27360), .Q(_29484) );
  nnd2s1 _29351_inst ( .DIN1(_29485), .DIN2(_27335), .Q(_27360) );
  hi1s1 _29352_inst ( .DIN(_29362), .Q(_29381) );
  nor2s1 _29353_inst ( .DIN1(_29362), .DIN2(_29486), .Q(_29471) );
  xor2s1 _29354_inst ( .DIN1(_29463), .DIN2(_29487), .Q(_29486) );
  xor2s1 _29355_inst ( .DIN1(_29464), .DIN2(_52928), .Q(_29487) );
  nnd2s1 _29356_inst ( .DIN1(_29466), .DIN2(_29488), .Q(_29464) );
  nnd2s1 _29357_inst ( .DIN1(_15553), .DIN2(_29489), .Q(_29488) );
  xor2s1 _29358_inst ( .DIN1(_29423), .DIN2(_29490), .Q(_29466) );
  nor2s1 _29359_inst ( .DIN1(_29489), .DIN2(_15553), .Q(_29423) );
  xor2s1 _29360_inst ( .DIN1(_29491), .DIN2(_29492), .Q(_29463) );
  nnd2s1 _29361_inst ( .DIN1(_29493), .DIN2(_29494), .Q(_29491) );
  nnd2s1 _29362_inst ( .DIN1(_53469), .DIN2(_29495), .Q(_29494) );
  nnd2s1 _29363_inst ( .DIN1(_29496), .DIN2(_27457), .Q(_29495) );
  or2s1 _29364_inst ( .DIN1(_29496), .DIN2(_27457), .Q(_29493) );
  nnd2s1 _29365_inst ( .DIN1(_29497), .DIN2(_29498), .Q(_29362) );
  nor2s1 _29366_inst ( .DIN1(_29499), .DIN2(_29500), .Q(_29498) );
  nnd2s1 _29367_inst ( .DIN1(_29501), .DIN2(_27493), .Q(_29500) );
  nor2s1 _29368_inst ( .DIN1(_27361), .DIN2(_29502), .Q(_29497) );
  or2s1 _29369_inst ( .DIN1(_27343), .DIN2(_27376), .Q(_29502) );
  nnd2s1 _29370_inst ( .DIN1(_29503), .DIN2(_29504), .Q(
        ______________________________47________) );
  nor2s1 _29371_inst ( .DIN1(_29505), .DIN2(_29506), .Q(_29503) );
  nor2s1 _29372_inst ( .DIN1(_29507), .DIN2(_29508), .Q(_29506) );
  nnd2s1 _29373_inst ( .DIN1(_29509), .DIN2(_29510), .Q(_29508) );
  nor2s1 _29374_inst ( .DIN1(_29511), .DIN2(_29512), .Q(_29509) );
  nor2s1 _29375_inst ( .DIN1(_29513), .DIN2(_29514), .Q(_29512) );
  xor2s1 _29376_inst ( .DIN1(_29496), .DIN2(_29515), .Q(_29514) );
  xor2s1 _29377_inst ( .DIN1(_53469), .DIN2(_27457), .Q(_29515) );
  nnd2s1 _29378_inst ( .DIN1(_29516), .DIN2(_29489), .Q(_27457) );
  or2s1 _29379_inst ( .DIN1(_29517), .DIN2(_26204), .Q(_29489) );
  xor2s1 _29380_inst ( .DIN1(_29518), .DIN2(_29519), .Q(_29516) );
  nnd2s1 _29381_inst ( .DIN1(_26204), .DIN2(_29517), .Q(_29519) );
  or2s1 _29382_inst ( .DIN1(_29520), .DIN2(_26826), .Q(_29517) );
  nnd2s1 _29383_inst ( .DIN1(_29521), .DIN2(_29522), .Q(_29496) );
  nnd2s1 _29384_inst ( .DIN1(_29523), .DIN2(_26628), .Q(_29522) );
  nnd2s1 _29385_inst ( .DIN1(_27006), .DIN2(_29524), .Q(_29523) );
  or2s1 _29386_inst ( .DIN1(_29524), .DIN2(_27006), .Q(_29521) );
  nor2s1 _29387_inst ( .DIN1(_29525), .DIN2(_29526), .Q(_29511) );
  nor2s1 _29388_inst ( .DIN1(_26774), .DIN2(_26442), .Q(_29526) );
  nor2s1 _29389_inst ( .DIN1(_29527), .DIN2(_29528), .Q(_29505) );
  nor2s1 _29390_inst ( .DIN1(_29529), .DIN2(_27039), .Q(_29528) );
  xnr2s1 _29391_inst ( .DIN1(_29530), .DIN2(_29531), .Q(_29529) );
  xor2s1 _29392_inst ( .DIN1(_52833), .DIN2(_52869), .Q(_29531) );
  nnd2s1 _29393_inst ( .DIN1(_29532), .DIN2(_27050), .Q(
        ______________________________46________) );
  nor2s1 _29394_inst ( .DIN1(_29533), .DIN2(_29534), .Q(_29532) );
  nor2s1 _29395_inst ( .DIN1(_27053), .DIN2(_29535), .Q(_29534) );
  nnd2s1 _29396_inst ( .DIN1(_29536), .DIN2(_29510), .Q(_29535) );
  nor2s1 _29397_inst ( .DIN1(_29537), .DIN2(_29538), .Q(_29536) );
  nor2s1 _29398_inst ( .DIN1(_29513), .DIN2(_29539), .Q(_29538) );
  xnr2s1 _29399_inst ( .DIN1(_27006), .DIN2(_29540), .Q(_29539) );
  xor2s1 _29400_inst ( .DIN1(_26628), .DIN2(_29524), .Q(_29540) );
  nnd2s1 _29401_inst ( .DIN1(_29541), .DIN2(_29542), .Q(_29524) );
  nnd2s1 _29402_inst ( .DIN1(_53016), .DIN2(_29543), .Q(_29542) );
  xor2s1 _29403_inst ( .DIN1(_29544), .DIN2(_29545), .Q(_29543) );
  xor2s1 _29404_inst ( .DIN1(_408), .DIN2(_29520), .Q(_27006) );
  nor2s1 _29405_inst ( .DIN1(_29525), .DIN2(_29546), .Q(_29537) );
  nor2s1 _29406_inst ( .DIN1(_29547), .DIN2(_29457), .Q(_29546) );
  nor2s1 _29407_inst ( .DIN1(_26442), .DIN2(_52868), .Q(_29457) );
  and2s1 _29408_inst ( .DIN1(_26442), .DIN2(_52868), .Q(_29547) );
  nor2s1 _29409_inst ( .DIN1(_27064), .DIN2(_29548), .Q(_29533) );
  nor2s1 _29410_inst ( .DIN1(_26855), .DIN2(_29549), .Q(_29548) );
  nnd2s1 _29411_inst ( .DIN1(_29550), .DIN2(_29551), .Q(_29549) );
  nnd2s1 _29412_inst ( .DIN1(_53054), .DIN2(_53074), .Q(_29550) );
  nnd2s1 _29413_inst ( .DIN1(_29552), .DIN2(_29553), .Q(
        ______________________________45________) );
  nnd2s1 _29414_inst ( .DIN1(_29554), .DIN2(_29555), .Q(_29553) );
  nnd2s1 _29415_inst ( .DIN1(_29556), .DIN2(_29557), .Q(_29554) );
  xor2s1 _29416_inst ( .DIN1(_26292), .DIN2(_29558), .Q(_29557) );
  nnd2s1 _29417_inst ( .DIN1(_29559), .DIN2(_29560), .Q(_29552) );
  nor2s1 _29418_inst ( .DIN1(_29561), .DIN2(_29562), .Q(_29559) );
  nnd2s1 _29419_inst ( .DIN1(_29563), .DIN2(_29564), .Q(_29562) );
  nnd2s1 _29420_inst ( .DIN1(_29565), .DIN2(_29525), .Q(_29564) );
  xor2s1 _29421_inst ( .DIN1(_26473), .DIN2(_29566), .Q(_29565) );
  and2s1 _29422_inst ( .DIN1(_29541), .DIN2(_29545), .Q(_29566) );
  nnd2s1 _29423_inst ( .DIN1(_29567), .DIN2(_29568), .Q(_29545) );
  nnd2s1 _29424_inst ( .DIN1(_27027), .DIN2(_29569), .Q(_29568) );
  nor2s1 _29425_inst ( .DIN1(_29570), .DIN2(_29571), .Q(_29567) );
  nor2s1 _29426_inst ( .DIN1(_53123), .DIN2(_29572), .Q(_29571) );
  nnd2s1 _29427_inst ( .DIN1(_29573), .DIN2(_29570), .Q(_29541) );
  hi1s1 _29428_inst ( .DIN(_27019), .Q(_29570) );
  nnd2s1 _29429_inst ( .DIN1(_29520), .DIN2(_29574), .Q(_27019) );
  nnd2s1 _29430_inst ( .DIN1(_15555), .DIN2(_29575), .Q(_29574) );
  or2s1 _29431_inst ( .DIN1(_29575), .DIN2(_15555), .Q(_29520) );
  nnd2s1 _29432_inst ( .DIN1(_29576), .DIN2(_29577), .Q(_29575) );
  xnr2s1 _29433_inst ( .DIN1(_29578), .DIN2(_29579), .Q(_29576) );
  nnd2s1 _29434_inst ( .DIN1(_29580), .DIN2(_29581), .Q(_29578) );
  nor2s1 _29435_inst ( .DIN1(_29582), .DIN2(_29572), .Q(_29573) );
  nor2s1 _29436_inst ( .DIN1(_27027), .DIN2(_29569), .Q(_29572) );
  nor2s1 _29437_inst ( .DIN1(_29583), .DIN2(_26365), .Q(_29582) );
  and2s1 _29438_inst ( .DIN1(_29569), .DIN2(_27027), .Q(_29583) );
  nnd2s1 _29439_inst ( .DIN1(_29584), .DIN2(_29513), .Q(_29563) );
  nnd2s1 _29440_inst ( .DIN1(_29585), .DIN2(_29586), .Q(_29584) );
  nnd2s1 _29441_inst ( .DIN1(_52987), .DIN2(_29587), .Q(_29586) );
  nnd2s1 _29442_inst ( .DIN1(_52870), .DIN2(______[16]), .Q(_29587) );
  nnd2s1 _29443_inst ( .DIN1(_29588), .DIN2(_26704), .Q(_29585) );
  nnd2s1 _29444_inst ( .DIN1(______[16]), .DIN2(_26588), .Q(_29588) );
  nnd2s1 _29445_inst ( .DIN1(_29589), .DIN2(_29590), .Q(
        ______________________________44________) );
  nnd2s1 _29446_inst ( .DIN1(_29591), .DIN2(_29592), .Q(_29590) );
  hi1s1 _29447_inst ( .DIN(_29593), .Q(_29592) );
  xnr2s1 _29448_inst ( .DIN1(_27027), .DIN2(_29594), .Q(_29591) );
  xor2s1 _29449_inst ( .DIN1(_26365), .DIN2(_29569), .Q(_29594) );
  nnd2s1 _29450_inst ( .DIN1(_29595), .DIN2(_29596), .Q(_29569) );
  nnd2s1 _29451_inst ( .DIN1(_29597), .DIN2(_26506), .Q(_29596) );
  or2s1 _29452_inst ( .DIN1(_29598), .DIN2(_27042), .Q(_29597) );
  xor2s1 _29453_inst ( .DIN1(_29599), .DIN2(_29600), .Q(_29595) );
  nnd2s1 _29454_inst ( .DIN1(_27042), .DIN2(_29598), .Q(_29600) );
  xnr2s1 _29455_inst ( .DIN1(_29601), .DIN2(_29580), .Q(_27027) );
  nnd2s1 _29456_inst ( .DIN1(_29577), .DIN2(_29581), .Q(_29601) );
  nor2s1 _29457_inst ( .DIN1(_29602), .DIN2(_29603), .Q(_29589) );
  nor2s1 _29458_inst ( .DIN1(_29527), .DIN2(_29604), .Q(_29603) );
  nnd2s1 _29459_inst ( .DIN1(_52868), .DIN2(_29605), .Q(_29604) );
  nor2s1 _29460_inst ( .DIN1(_29606), .DIN2(_29507), .Q(_29602) );
  nor2s1 _29461_inst ( .DIN1(_29607), .DIN2(_29608), .Q(_29606) );
  nor2s1 _29462_inst ( .DIN1(_29525), .DIN2(_29609), .Q(_29607) );
  nor2s1 _29463_inst ( .DIN1(_26853), .DIN2(_29610), .Q(_29609) );
  nnd2s1 _29464_inst ( .DIN1(_29611), .DIN2(_29612), .Q(_29610) );
  nnd2s1 _29465_inst ( .DIN1(_52869), .DIN2(_26561), .Q(_29612) );
  nnd2s1 _29466_inst ( .DIN1(_29613), .DIN2(_53128), .Q(_29611) );
  nor2s1 _29467_inst ( .DIN1(_52869), .DIN2(_52870), .Q(_29613) );
  nnd2s1 _29468_inst ( .DIN1(_29614), .DIN2(_29615), .Q(
        ______________________________43________) );
  nor2s1 _29469_inst ( .DIN1(_29616), .DIN2(_29617), .Q(_29615) );
  nor2s1 _29470_inst ( .DIN1(_29593), .DIN2(_29618), .Q(_29617) );
  xnr2s1 _29471_inst ( .DIN1(_27042), .DIN2(_29619), .Q(_29618) );
  xor2s1 _29472_inst ( .DIN1(_26506), .DIN2(_29598), .Q(_29619) );
  nnd2s1 _29473_inst ( .DIN1(_29620), .DIN2(_29621), .Q(_29598) );
  nnd2s1 _29474_inst ( .DIN1(_29622), .DIN2(_26304), .Q(_29621) );
  nnd2s1 _29475_inst ( .DIN1(_29623), .DIN2(_29624), .Q(_29622) );
  or2s1 _29476_inst ( .DIN1(_29624), .DIN2(_29623), .Q(_29620) );
  xor2s1 _29477_inst ( .DIN1(_29577), .DIN2(_29581), .Q(_27042) );
  nnd2s1 _29478_inst ( .DIN1(_29527), .DIN2(_29525), .Q(_29593) );
  nor2s1 _29479_inst ( .DIN1(_29625), .DIN2(_29626), .Q(_29614) );
  nor2s1 _29480_inst ( .DIN1(______[24]), .DIN2(_29527), .Q(_29626) );
  nor2s1 _29481_inst ( .DIN1(_52869), .DIN2(_29627), .Q(_29625) );
  nor2s1 _29482_inst ( .DIN1(_29628), .DIN2(_29507), .Q(_29627) );
  nor2s1 _29483_inst ( .DIN1(_29525), .DIN2(_29561), .Q(_29628) );
  hi1s1 _29484_inst ( .DIN(_29510), .Q(_29561) );
  nnd2s1 _29485_inst ( .DIN1(_29629), .DIN2(_29630), .Q(
        ______________________________42________) );
  nnd2s1 _29486_inst ( .DIN1(_27476), .DIN2(_29631), .Q(_29630) );
  nnd2s1 _29487_inst ( .DIN1(_29632), .DIN2(_29633), .Q(_29631) );
  hi1s1 _29488_inst ( .DIN(_29608), .Q(_29633) );
  nnd2s1 _29489_inst ( .DIN1(_29510), .DIN2(_29634), .Q(_29608) );
  nnd2s1 _29490_inst ( .DIN1(_29635), .DIN2(_52870), .Q(_29634) );
  nor2s1 _29491_inst ( .DIN1(_53128), .DIN2(_29525), .Q(_29635) );
  nnd2s1 _29492_inst ( .DIN1(_29636), .DIN2(_29637), .Q(_29510) );
  and2s1 _29493_inst ( .DIN1(_27497), .DIN2(_29513), .Q(_29637) );
  nor2s1 _29494_inst ( .DIN1(_29205), .DIN2(_29159), .Q(_29636) );
  nnd2s1 _29495_inst ( .DIN1(_29345), .DIN2(_29353), .Q(_29159) );
  nor2s1 _29496_inst ( .DIN1(_29638), .DIN2(_29639), .Q(_29632) );
  nor2s1 _29497_inst ( .DIN1(_29513), .DIN2(_29640), .Q(_29639) );
  xor2s1 _29498_inst ( .DIN1(_29624), .DIN2(_29641), .Q(_29640) );
  xor2s1 _29499_inst ( .DIN1(_26304), .DIN2(_29623), .Q(_29641) );
  hi1s1 _29500_inst ( .DIN(_27057), .Q(_29623) );
  nor2s1 _29501_inst ( .DIN1(_29577), .DIN2(_29642), .Q(_27057) );
  and2s1 _29502_inst ( .DIN1(_26829), .DIN2(_29643), .Q(_29642) );
  nor2s1 _29503_inst ( .DIN1(_29643), .DIN2(_420), .Q(_29577) );
  nnd2s1 _29504_inst ( .DIN1(_29644), .DIN2(_29645), .Q(_29624) );
  nnd2s1 _29505_inst ( .DIN1(_29646), .DIN2(_26251), .Q(_29645) );
  or2s1 _29506_inst ( .DIN1(_27081), .DIN2(_29647), .Q(_29646) );
  nnd2s1 _29507_inst ( .DIN1(_29647), .DIN2(_27081), .Q(_29644) );
  nor2s1 _29508_inst ( .DIN1(_29525), .DIN2(_29648), .Q(_29638) );
  nor2s1 _29509_inst ( .DIN1(_29649), .DIN2(_27393), .Q(_29648) );
  nor2s1 _29510_inst ( .DIN1(_52870), .DIN2(_26561), .Q(_29649) );
  hi1s1 _29511_inst ( .DIN(_29513), .Q(_29525) );
  nnd2s1 _29512_inst ( .DIN1(_29650), .DIN2(_29651), .Q(_29513) );
  nor2s1 _29513_inst ( .DIN1(_29203), .DIN2(_29652), .Q(_29651) );
  nnd2s1 _29514_inst ( .DIN1(_27348), .DIN2(_27467), .Q(_29652) );
  nor2s1 _29515_inst ( .DIN1(_27377), .DIN2(_29653), .Q(_29650) );
  nnd2s1 _29516_inst ( .DIN1(_29654), .DIN2(_29655), .Q(_29653) );
  hi1s1 _29517_inst ( .DIN(_29656), .Q(_29654) );
  nnd2s1 _29518_inst ( .DIN1(_29657), .DIN2(_29658), .Q(_29629) );
  nor2s1 _29519_inst ( .DIN1(_29659), .DIN2(_27614), .Q(_29657) );
  xor2s1 _29520_inst ( .DIN1(_29660), .DIN2(_29661), .Q(_29659) );
  nor2s1 _29521_inst ( .DIN1(_53289), .DIN2(_52987), .Q(_29661) );
  xor2s1 _29522_inst ( .DIN1(_26682), .DIN2(_53288), .Q(_29660) );
  nnd2s1 _29523_inst ( .DIN1(_29662), .DIN2(_29504), .Q(
        ______________________________41________) );
  nor2s1 _29524_inst ( .DIN1(_29663), .DIN2(_29664), .Q(_29662) );
  nor2s1 _29525_inst ( .DIN1(_29507), .DIN2(_29665), .Q(_29664) );
  nnd2s1 _29526_inst ( .DIN1(_29666), .DIN2(_29667), .Q(_29665) );
  nnd2s1 _29527_inst ( .DIN1(_29668), .DIN2(_29669), .Q(_29667) );
  xnr2s1 _29528_inst ( .DIN1(_29647), .DIN2(_29670), .Q(_29669) );
  xor2s1 _29529_inst ( .DIN1(_26251), .DIN2(_27081), .Q(_29670) );
  nnd2s1 _29530_inst ( .DIN1(_29643), .DIN2(_29671), .Q(_27081) );
  nnd2s1 _29531_inst ( .DIN1(_424), .DIN2(_29672), .Q(_29671) );
  or2s1 _29532_inst ( .DIN1(_29672), .DIN2(_424), .Q(_29643) );
  nnd2s1 _29533_inst ( .DIN1(_29673), .DIN2(_29674), .Q(_29647) );
  nnd2s1 _29534_inst ( .DIN1(_52871), .DIN2(_29675), .Q(_29674) );
  or2s1 _29535_inst ( .DIN1(_27099), .DIN2(_29676), .Q(_29675) );
  nnd2s1 _29536_inst ( .DIN1(_29676), .DIN2(_27099), .Q(_29673) );
  nnd2s1 _29537_inst ( .DIN1(_29677), .DIN2(_29678), .Q(_29666) );
  xor2s1 _29538_inst ( .DIN1(_26608), .DIN2(_29679), .Q(_29678) );
  nor2s1 _29539_inst ( .DIN1(_29527), .DIN2(_29680), .Q(_29663) );
  nor2s1 _29540_inst ( .DIN1(_27066), .DIN2(_29681), .Q(_29680) );
  nnd2s1 _29541_inst ( .DIN1(_29682), .DIN2(_29683), .Q(_29681) );
  nnd2s1 _29542_inst ( .DIN1(_29684), .DIN2(_26588), .Q(_29683) );
  nnd2s1 _29543_inst ( .DIN1(_52869), .DIN2(_52833), .Q(_29684) );
  nnd2s1 _29544_inst ( .DIN1(_29530), .DIN2(_52833), .Q(_29682) );
  and2s1 _29545_inst ( .DIN1(_52869), .DIN2(_52870), .Q(_29530) );
  nnd2s1 _29546_inst ( .DIN1(_29685), .DIN2(_29686), .Q(
        ______________________________40________) );
  nor2s1 _29547_inst ( .DIN1(_29687), .DIN2(_29688), .Q(_29685) );
  nor2s1 _29548_inst ( .DIN1(_29689), .DIN2(_29690), .Q(_29688) );
  nnd2s1 _29549_inst ( .DIN1(_29691), .DIN2(_29692), .Q(_29690) );
  nnd2s1 _29550_inst ( .DIN1(_29693), .DIN2(_29668), .Q(_29692) );
  xor2s1 _29551_inst ( .DIN1(_29676), .DIN2(_29694), .Q(_29693) );
  xnr2s1 _29552_inst ( .DIN1(_52871), .DIN2(_27099), .Q(_29694) );
  nnd2s1 _29553_inst ( .DIN1(_29672), .DIN2(_29695), .Q(_27099) );
  nnd2s1 _29554_inst ( .DIN1(_15560), .DIN2(_29696), .Q(_29695) );
  or2s1 _29555_inst ( .DIN1(_29696), .DIN2(_15560), .Q(_29672) );
  nnd2s1 _29556_inst ( .DIN1(_29697), .DIN2(_29698), .Q(_29676) );
  nnd2s1 _29557_inst ( .DIN1(_52874), .DIN2(_29699), .Q(_29698) );
  or2s1 _29558_inst ( .DIN1(_27111), .DIN2(_29700), .Q(_29699) );
  nnd2s1 _29559_inst ( .DIN1(_29700), .DIN2(_27111), .Q(_29697) );
  nnd2s1 _29560_inst ( .DIN1(_29677), .DIN2(_29701), .Q(_29691) );
  xor2s1 _29561_inst ( .DIN1(_52833), .DIN2(_29702), .Q(_29701) );
  nor2s1 _29562_inst ( .DIN1(_29703), .DIN2(_27448), .Q(_29677) );
  nor2s1 _29563_inst ( .DIN1(_27154), .DIN2(_29704), .Q(_29687) );
  xor2s1 _29564_inst ( .DIN1(_26406), .DIN2(_29705), .Q(_29704) );
  nnd2s1 _29565_inst ( .DIN1(_53093), .DIN2(_52875), .Q(_29705) );
  nnd2s1 _29566_inst ( .DIN1(_29706), .DIN2(_29707), .Q(
        ______________________________3________) );
  nnd2s1 _29567_inst ( .DIN1(_29708), .DIN2(______[2]), .Q(_29707) );
  nor2s1 _29568_inst ( .DIN1(_27522), .DIN2(_29709), .Q(_29708) );
  xor2s1 _29569_inst ( .DIN1(_26323), .DIN2(_29710), .Q(_29709) );
  nnd2s1 _29570_inst ( .DIN1(_27524), .DIN2(_29711), .Q(_29706) );
  nnd2s1 _29571_inst ( .DIN1(_29712), .DIN2(_29713), .Q(_29711) );
  nnd2s1 _29572_inst ( .DIN1(_52879), .DIN2(_28809), .Q(_29713) );
  nor2s1 _29573_inst ( .DIN1(_28935), .DIN2(_28938), .Q(_28809) );
  or2s1 _29574_inst ( .DIN1(_28804), .DIN2(_52872), .Q(_29712) );
  nnd2s1 _29575_inst ( .DIN1(_29714), .DIN2(_29504), .Q(
        ______________________________39________) );
  nor2s1 _29576_inst ( .DIN1(_29715), .DIN2(_29716), .Q(_29714) );
  nor2s1 _29577_inst ( .DIN1(_29717), .DIN2(_29507), .Q(_29716) );
  nor2s1 _29578_inst ( .DIN1(_29718), .DIN2(_29719), .Q(_29717) );
  nor2s1 _29579_inst ( .DIN1(_29720), .DIN2(_29721), .Q(_29719) );
  xor2s1 _29580_inst ( .DIN1(_29722), .DIN2(_29700), .Q(_29720) );
  and2s1 _29581_inst ( .DIN1(_29723), .DIN2(_29724), .Q(_29700) );
  nnd2s1 _29582_inst ( .DIN1(_29725), .DIN2(_26301), .Q(_29724) );
  nnd2s1 _29583_inst ( .DIN1(_27262), .DIN2(_29726), .Q(_29725) );
  xor2s1 _29584_inst ( .DIN1(_29727), .DIN2(_29728), .Q(_29723) );
  nor2s1 _29585_inst ( .DIN1(_27262), .DIN2(_29726), .Q(_29728) );
  xor2s1 _29586_inst ( .DIN1(_27111), .DIN2(_52874), .Q(_29722) );
  nnd2s1 _29587_inst ( .DIN1(_29729), .DIN2(_29696), .Q(_27111) );
  nnd2s1 _29588_inst ( .DIN1(_29730), .DIN2(_29731), .Q(_29696) );
  nor2s1 _29589_inst ( .DIN1(_29732), .DIN2(_433), .Q(_29730) );
  xor2s1 _29590_inst ( .DIN1(_26321), .DIN2(_29733), .Q(_29729) );
  and2s1 _29591_inst ( .DIN1(_29734), .DIN2(_15561), .Q(_29733) );
  nor2s1 _29592_inst ( .DIN1(_29703), .DIN2(_29735), .Q(_29718) );
  nnd2s1 _29593_inst ( .DIN1(_52875), .DIN2(______[22]), .Q(_29735) );
  nor2s1 _29594_inst ( .DIN1(_29527), .DIN2(_29736), .Q(_29715) );
  nor2s1 _29595_inst ( .DIN1(_26774), .DIN2(_29737), .Q(_29736) );
  xnr2s1 _29596_inst ( .DIN1(_52876), .DIN2(_29738), .Q(_29737) );
  nnd2s1 _29597_inst ( .DIN1(_52882), .DIN2(_52873), .Q(_29738) );
  nnd2s1 _29598_inst ( .DIN1(_29739), .DIN2(_29504), .Q(
        ______________________________38________) );
  hi1s1 _29599_inst ( .DIN(_29616), .Q(_29504) );
  nor2s1 _29600_inst ( .DIN1(_29605), .DIN2(_29527), .Q(_29616) );
  or2s1 _29601_inst ( .DIN1(_29740), .DIN2(_27317), .Q(_29605) );
  nnd2s1 _29602_inst ( .DIN1(_29741), .DIN2(_29742), .Q(_29740) );
  nor2s1 _29603_inst ( .DIN1(_29743), .DIN2(_29744), .Q(_29739) );
  nor2s1 _29604_inst ( .DIN1(_29507), .DIN2(_29745), .Q(_29744) );
  nnd2s1 _29605_inst ( .DIN1(_29746), .DIN2(_29747), .Q(_29745) );
  nnd2s1 _29606_inst ( .DIN1(_29748), .DIN2(_29668), .Q(_29747) );
  xor2s1 _29607_inst ( .DIN1(_29726), .DIN2(_29749), .Q(_29748) );
  xor2s1 _29608_inst ( .DIN1(_26301), .DIN2(_27262), .Q(_29749) );
  nnd2s1 _29609_inst ( .DIN1(_29734), .DIN2(_29750), .Q(_27262) );
  nnd2s1 _29610_inst ( .DIN1(_433), .DIN2(_29751), .Q(_29750) );
  nnd2s1 _29611_inst ( .DIN1(_29731), .DIN2(_29752), .Q(_29751) );
  nnd2s1 _29612_inst ( .DIN1(_29753), .DIN2(_29731), .Q(_29734) );
  nor2s1 _29613_inst ( .DIN1(_438), .DIN2(_433), .Q(_29753) );
  nnd2s1 _29614_inst ( .DIN1(_29754), .DIN2(_29755), .Q(_29726) );
  nnd2s1 _29615_inst ( .DIN1(_29756), .DIN2(_26635), .Q(_29755) );
  nnd2s1 _29616_inst ( .DIN1(_27486), .DIN2(_29757), .Q(_29756) );
  or2s1 _29617_inst ( .DIN1(_29757), .DIN2(_27486), .Q(_29754) );
  nnd2s1 _29618_inst ( .DIN1(_29758), .DIN2(_29759), .Q(_29746) );
  nor2s1 _29619_inst ( .DIN1(_29702), .DIN2(_29760), .Q(_29759) );
  nor2s1 _29620_inst ( .DIN1(_52875), .DIN2(_26426), .Q(_29760) );
  hi1s1 _29621_inst ( .DIN(_29679), .Q(_29702) );
  nnd2s1 _29622_inst ( .DIN1(_52875), .DIN2(_26426), .Q(_29679) );
  nor2s1 _29623_inst ( .DIN1(_28646), .DIN2(_29703), .Q(_29758) );
  nnd2s1 _29624_inst ( .DIN1(_29721), .DIN2(_29761), .Q(_29703) );
  nnd2s1 _29625_inst ( .DIN1(_29762), .DIN2(_27492), .Q(_29761) );
  nor2s1 _29626_inst ( .DIN1(_29527), .DIN2(_29763), .Q(_29743) );
  nor2s1 _29627_inst ( .DIN1(_29764), .DIN2(_27365), .Q(_29763) );
  xor2s1 _29628_inst ( .DIN1(_26426), .DIN2(_52882), .Q(_29764) );
  hi1s1 _29629_inst ( .DIN(_29507), .Q(_29527) );
  nnd2s1 _29630_inst ( .DIN1(_29765), .DIN2(_29766), .Q(_29507) );
  nor2s1 _29631_inst ( .DIN1(_27430), .DIN2(_29767), .Q(_29766) );
  nor2s1 _29632_inst ( .DIN1(_27433), .DIN2(_29768), .Q(_29765) );
  nnd2s1 _29633_inst ( .DIN1(_29769), .DIN2(_29770), .Q(
        ______________________________37________) );
  nnd2s1 _29634_inst ( .DIN1(_27129), .DIN2(_29771), .Q(_29770) );
  nnd2s1 _29635_inst ( .DIN1(_29772), .DIN2(_29773), .Q(_29771) );
  nor2s1 _29636_inst ( .DIN1(_29774), .DIN2(_29775), .Q(_29772) );
  nor2s1 _29637_inst ( .DIN1(_29721), .DIN2(_29776), .Q(_29775) );
  xnr2s1 _29638_inst ( .DIN1(_27486), .DIN2(_29777), .Q(_29776) );
  xor2s1 _29639_inst ( .DIN1(_26635), .DIN2(_29757), .Q(_29777) );
  nnd2s1 _29640_inst ( .DIN1(_29778), .DIN2(_29779), .Q(_29757) );
  nnd2s1 _29641_inst ( .DIN1(_52879), .DIN2(_29780), .Q(_29779) );
  nnd2s1 _29642_inst ( .DIN1(_29781), .DIN2(_29782), .Q(_29780) );
  or2s1 _29643_inst ( .DIN1(_29781), .DIN2(_29782), .Q(_29778) );
  xor2s1 _29644_inst ( .DIN1(_29731), .DIN2(_29752), .Q(_27486) );
  nor2s1 _29645_inst ( .DIN1(_29668), .DIN2(_29783), .Q(_29774) );
  xnr2s1 _29646_inst ( .DIN1(_52876), .DIN2(_29784), .Q(_29783) );
  nnd2s1 _29647_inst ( .DIN1(_29785), .DIN2(_29786), .Q(_29769) );
  nor2s1 _29648_inst ( .DIN1(_29787), .DIN2(_29788), .Q(_29786) );
  nor2s1 _29649_inst ( .DIN1(_52834), .DIN2(_26427), .Q(_29788) );
  nor2s1 _29650_inst ( .DIN1(_27039), .DIN2(_29789), .Q(_29785) );
  nnd2s1 _29651_inst ( .DIN1(_29790), .DIN2(_29791), .Q(
        ______________________________36________) );
  nnd2s1 _29652_inst ( .DIN1(_29792), .DIN2(_29793), .Q(_29791) );
  nnd2s1 _29653_inst ( .DIN1(_29794), .DIN2(_29773), .Q(_29793) );
  nnd2s1 _29654_inst ( .DIN1(_29795), .DIN2(_29762), .Q(_29773) );
  hi1s1 _29655_inst ( .DIN(_27377), .Q(_29762) );
  nnd2s1 _29656_inst ( .DIN1(_29796), .DIN2(_29797), .Q(_27377) );
  nor2s1 _29657_inst ( .DIN1(_29798), .DIN2(_29799), .Q(_29797) );
  nnd2s1 _29658_inst ( .DIN1(_27494), .DIN2(_27349), .Q(_29799) );
  hi1s1 _29659_inst ( .DIN(_27493), .Q(_29798) );
  nor2s1 _29660_inst ( .DIN1(_29483), .DIN2(_29800), .Q(_29796) );
  nnd2s1 _29661_inst ( .DIN1(_29353), .DIN2(_29501), .Q(_29800) );
  nor2s1 _29662_inst ( .DIN1(_29801), .DIN2(_29668), .Q(_29795) );
  nor2s1 _29663_inst ( .DIN1(_29802), .DIN2(_29803), .Q(_29794) );
  nor2s1 _29664_inst ( .DIN1(_29721), .DIN2(_29804), .Q(_29803) );
  xor2s1 _29665_inst ( .DIN1(_29782), .DIN2(_29805), .Q(_29804) );
  xor2s1 _29666_inst ( .DIN1(_29781), .DIN2(_52879), .Q(_29805) );
  nnd2s1 _29667_inst ( .DIN1(_29806), .DIN2(_29807), .Q(_29781) );
  nnd2s1 _29668_inst ( .DIN1(_52896), .DIN2(_29808), .Q(_29807) );
  or2s1 _29669_inst ( .DIN1(_29809), .DIN2(_29810), .Q(_29808) );
  nnd2s1 _29670_inst ( .DIN1(_29810), .DIN2(_29809), .Q(_29806) );
  or2s1 _29671_inst ( .DIN1(_29731), .DIN2(_29811), .Q(_29782) );
  and2s1 _29672_inst ( .DIN1(_441), .DIN2(_29812), .Q(_29811) );
  nor2s1 _29673_inst ( .DIN1(_29812), .DIN2(_441), .Q(_29731) );
  nor2s1 _29674_inst ( .DIN1(_29668), .DIN2(_29813), .Q(_29802) );
  xor2s1 _29675_inst ( .DIN1(_52878), .DIN2(_29784), .Q(_29813) );
  nor2s1 _29676_inst ( .DIN1(_52882), .DIN2(_53025), .Q(_29784) );
  hi1s1 _29677_inst ( .DIN(_29721), .Q(_29668) );
  nnd2s1 _29678_inst ( .DIN1(_29814), .DIN2(_29815), .Q(_29721) );
  nor2s1 _29679_inst ( .DIN1(_29816), .DIN2(_27376), .Q(_29815) );
  nor2s1 _29680_inst ( .DIN1(_29205), .DIN2(_27004), .Q(_29814) );
  nnd2s1 _29681_inst ( .DIN1(_29817), .DIN2(_29485), .Q(_27004) );
  nnd2s1 _29682_inst ( .DIN1(_29818), .DIN2(_29819), .Q(_29485) );
  nor2s1 _29683_inst ( .DIN1(_29820), .DIN2(_29801), .Q(_29817) );
  nnd2s1 _29684_inst ( .DIN1(_29821), .DIN2(_27493), .Q(_29205) );
  and2s1 _29685_inst ( .DIN1(_27467), .DIN2(_27373), .Q(_29821) );
  nnd2s1 _29686_inst ( .DIN1(_29822), .DIN2(_52873), .Q(_29790) );
  nnd2s1 _29687_inst ( .DIN1(_29823), .DIN2(_29824), .Q(
        ______________________________35________) );
  nor2s1 _29688_inst ( .DIN1(_29825), .DIN2(_29826), .Q(_29824) );
  nor2s1 _29689_inst ( .DIN1(_29827), .DIN2(_29828), .Q(_29826) );
  nor2s1 _29690_inst ( .DIN1(_29829), .DIN2(_29830), .Q(_29827) );
  nor2s1 _29691_inst ( .DIN1(_29831), .DIN2(_29832), .Q(_29830) );
  xor2s1 _29692_inst ( .DIN1(_29810), .DIN2(_29833), .Q(_29832) );
  xnr2s1 _29693_inst ( .DIN1(_52896), .DIN2(_29809), .Q(_29833) );
  nnd2s1 _29694_inst ( .DIN1(_29834), .DIN2(_29812), .Q(_29809) );
  nnd2s1 _29695_inst ( .DIN1(_29835), .DIN2(_29836), .Q(_29812) );
  nor2s1 _29696_inst ( .DIN1(_640), .DIN2(_29837), .Q(_29835) );
  nnd2s1 _29697_inst ( .DIN1(_14172), .DIN2(_29838), .Q(_29834) );
  nnd2s1 _29698_inst ( .DIN1(_29839), .DIN2(_29836), .Q(_29838) );
  nor2s1 _29699_inst ( .DIN1(_26827), .DIN2(_15563), .Q(_29839) );
  and2s1 _29700_inst ( .DIN1(_29840), .DIN2(_29841), .Q(_29810) );
  nnd2s1 _29701_inst ( .DIN1(_29842), .DIN2(_52881), .Q(_29841) );
  nor2s1 _29702_inst ( .DIN1(_29843), .DIN2(_29844), .Q(_29842) );
  nor2s1 _29703_inst ( .DIN1(_26360), .DIN2(_29845), .Q(_29843) );
  nnd2s1 _29704_inst ( .DIN1(_29845), .DIN2(_26360), .Q(_29840) );
  nor2s1 _29705_inst ( .DIN1(_29846), .DIN2(_29847), .Q(_29829) );
  nor2s1 _29706_inst ( .DIN1(_52882), .DIN2(_29848), .Q(_29847) );
  nor2s1 _29707_inst ( .DIN1(_29849), .DIN2(_29850), .Q(_29825) );
  nor2s1 _29708_inst ( .DIN1(_29851), .DIN2(_27448), .Q(_29850) );
  nor2s1 _29709_inst ( .DIN1(_29852), .DIN2(_26412), .Q(_29851) );
  nor2s1 _29710_inst ( .DIN1(_29853), .DIN2(_29854), .Q(_29823) );
  nor2s1 _29711_inst ( .DIN1(_53294), .DIN2(_29855), .Q(_29854) );
  nnd2s1 _29712_inst ( .DIN1(_29856), .DIN2(_29857), .Q(
        ______________________________34________) );
  nnd2s1 _29713_inst ( .DIN1(_29858), .DIN2(_27779), .Q(_29857) );
  nnd2s1 _29714_inst ( .DIN1(_29859), .DIN2(_29860), .Q(_29858) );
  nnd2s1 _29715_inst ( .DIN1(_52988), .DIN2(_26297), .Q(_29860) );
  nnd2s1 _29716_inst ( .DIN1(_29861), .DIN2(_27782), .Q(_29856) );
  nor2s1 _29717_inst ( .DIN1(_29862), .DIN2(_29863), .Q(_29861) );
  nor2s1 _29718_inst ( .DIN1(_29126), .DIN2(_29864), .Q(_29863) );
  xnr2s1 _29719_inst ( .DIN1(_52956), .DIN2(_29865), .Q(_29864) );
  nnd2s1 _29720_inst ( .DIN1(_52912), .DIN2(_52955), .Q(_29865) );
  nor2s1 _29721_inst ( .DIN1(_29866), .DIN2(_29867), .Q(_29862) );
  xnr2s1 _29722_inst ( .DIN1(_29845), .DIN2(_29868), .Q(_29867) );
  xor2s1 _29723_inst ( .DIN1(_26360), .DIN2(_29869), .Q(_29868) );
  nor2s1 _29724_inst ( .DIN1(_29844), .DIN2(_26603), .Q(_29869) );
  xnr2s1 _29725_inst ( .DIN1(_29870), .DIN2(_29871), .Q(_29845) );
  nnd2s1 _29726_inst ( .DIN1(_29836), .DIN2(_29872), .Q(_29870) );
  nnd2s1 _29727_inst ( .DIN1(_29873), .DIN2(_29874), .Q(
        ______________________________33________) );
  nnd2s1 _29728_inst ( .DIN1(_29875), .DIN2(_29876), .Q(_29874) );
  xor2s1 _29729_inst ( .DIN1(_26603), .DIN2(_29844), .Q(_29875) );
  xor2s1 _29730_inst ( .DIN1(_29836), .DIN2(_15563), .Q(_29844) );
  nor2s1 _29731_inst ( .DIN1(_29877), .DIN2(_29878), .Q(_29873) );
  nor2s1 _29732_inst ( .DIN1(_29879), .DIN2(_29880), .Q(_29878) );
  nnd2s1 _29733_inst ( .DIN1(______[0]), .DIN2(_29881), .Q(_29880) );
  xor2s1 _29734_inst ( .DIN1(_52873), .DIN2(_52882), .Q(_29881) );
  nor2s1 _29735_inst ( .DIN1(_29882), .DIN2(_29883), .Q(_29877) );
  nnd2s1 _29736_inst ( .DIN1(_29884), .DIN2(_29885), .Q(_29883) );
  xor2s1 _29737_inst ( .DIN1(_52882), .DIN2(_53025), .Q(_29884) );
  nnd2s1 _29738_inst ( .DIN1(_29886), .DIN2(_29887), .Q(
        ______________________________32________) );
  nnd2s1 _29739_inst ( .DIN1(_29888), .DIN2(_29889), .Q(_29887) );
  xor2s1 _29740_inst ( .DIN1(_53360), .DIN2(_53485), .Q(_29889) );
  hi1s1 _29741_inst ( .DIN(_27881), .Q(_29888) );
  nnd2s1 _29742_inst ( .DIN1(_27882), .DIN2(_29890), .Q(_29886) );
  nnd2s1 _29743_inst ( .DIN1(_29891), .DIN2(_28009), .Q(_29890) );
  nnd2s1 _29744_inst ( .DIN1(_29892), .DIN2(_29893), .Q(_28009) );
  nor2s1 _29745_inst ( .DIN1(_29894), .DIN2(_27963), .Q(_29893) );
  nor2s1 _29746_inst ( .DIN1(_29895), .DIN2(_29896), .Q(_29891) );
  nor2s1 _29747_inst ( .DIN1(_27963), .DIN2(_29897), .Q(_29896) );
  nor2s1 _29748_inst ( .DIN1(_26774), .DIN2(_29898), .Q(_29897) );
  nnd2s1 _29749_inst ( .DIN1(_29899), .DIN2(_28006), .Q(_29898) );
  nnd2s1 _29750_inst ( .DIN1(_52970), .DIN2(_53175), .Q(_28006) );
  nnd2s1 _29751_inst ( .DIN1(_26295), .DIN2(_26425), .Q(_29899) );
  hi1s1 _29752_inst ( .DIN(_27965), .Q(_27963) );
  nor2s1 _29753_inst ( .DIN1(_52979), .DIN2(_27965), .Q(_29895) );
  nnd2s1 _29754_inst ( .DIN1(_29900), .DIN2(_29901), .Q(_27965) );
  nor2s1 _29755_inst ( .DIN1(_29902), .DIN2(_29903), .Q(_29901) );
  nor2s1 _29756_inst ( .DIN1(_28215), .DIN2(_29904), .Q(_29900) );
  nnd2s1 _29757_inst ( .DIN1(_29905), .DIN2(_29906), .Q(
        ______________________________31________) );
  nnd2s1 _29758_inst ( .DIN1(_29907), .DIN2(______[18]), .Q(_29906) );
  nor2s1 _29759_inst ( .DIN1(_27522), .DIN2(_29908), .Q(_29907) );
  xor2s1 _29760_inst ( .DIN1(_26488), .DIN2(_53011), .Q(_29908) );
  nnd2s1 _29761_inst ( .DIN1(_27524), .DIN2(_29909), .Q(_29905) );
  nnd2s1 _29762_inst ( .DIN1(_29910), .DIN2(_29911), .Q(_29909) );
  nor2s1 _29763_inst ( .DIN1(_29912), .DIN2(_29913), .Q(_29910) );
  and2s1 _29764_inst ( .DIN1(_52842), .DIN2(_27951), .Q(_29913) );
  nor2s1 _29765_inst ( .DIN1(_27951), .DIN2(_29914), .Q(_29912) );
  xor2s1 _29766_inst ( .DIN1(_26730), .DIN2(_52886), .Q(_29914) );
  nnd2s1 _29767_inst ( .DIN1(_29915), .DIN2(_29916), .Q(
        ______________________________30________) );
  nnd2s1 _29768_inst ( .DIN1(_29917), .DIN2(_29918), .Q(_29916) );
  xnr2s1 _29769_inst ( .DIN1(_29919), .DIN2(_29920), .Q(_29917) );
  nnd2s1 _29770_inst ( .DIN1(_29921), .DIN2(_29922), .Q(_29915) );
  nnd2s1 _29771_inst ( .DIN1(_29923), .DIN2(_29911), .Q(_29922) );
  nor2s1 _29772_inst ( .DIN1(_29924), .DIN2(_29925), .Q(_29923) );
  nor2s1 _29773_inst ( .DIN1(_52885), .DIN2(_27951), .Q(_29925) );
  nor2s1 _29774_inst ( .DIN1(_53393), .DIN2(_29926), .Q(_29924) );
  nnd2s1 _29775_inst ( .DIN1(_29927), .DIN2(_29928), .Q(
        ______________________________2________) );
  nor2s1 _29776_inst ( .DIN1(_29929), .DIN2(_29930), .Q(_29928) );
  nor2s1 _29777_inst ( .DIN1(_28704), .DIN2(_29931), .Q(_29930) );
  nnd2s1 _29778_inst ( .DIN1(_28724), .DIN2(_52837), .Q(_29931) );
  hi1s1 _29779_inst ( .DIN(_28851), .Q(_28704) );
  nor2s1 _29780_inst ( .DIN1(_28851), .DIN2(_29932), .Q(_29929) );
  xor2s1 _29781_inst ( .DIN1(_29933), .DIN2(_29934), .Q(_29932) );
  xor2s1 _29782_inst ( .DIN1(_52954), .DIN2(_52974), .Q(_29934) );
  nor2s1 _29783_inst ( .DIN1(_26471), .DIN2(_26257), .Q(_29933) );
  nor2s1 _29784_inst ( .DIN1(_28891), .DIN2(_29935), .Q(_29927) );
  nor2s1 _29785_inst ( .DIN1(_52896), .DIN2(_28710), .Q(_29935) );
  nnd2s1 _29786_inst ( .DIN1(_29936), .DIN2(_28851), .Q(_28710) );
  nor2s1 _29787_inst ( .DIN1(_28724), .DIN2(_28727), .Q(_29936) );
  hi1s1 _29788_inst ( .DIN(_28837), .Q(_28891) );
  nnd2s1 _29789_inst ( .DIN1(_29937), .DIN2(_28887), .Q(_28837) );
  nor2s1 _29790_inst ( .DIN1(_28851), .DIN2(_29938), .Q(_29937) );
  nor2s1 _29791_inst ( .DIN1(_29939), .DIN2(_29940), .Q(_28851) );
  nnd2s1 _29792_inst ( .DIN1(_29941), .DIN2(_27560), .Q(
        ______________________________29________) );
  nor2s1 _29793_inst ( .DIN1(_29942), .DIN2(_29943), .Q(_29941) );
  nor2s1 _29794_inst ( .DIN1(_27563), .DIN2(_29944), .Q(_29943) );
  nnd2s1 _29795_inst ( .DIN1(_29945), .DIN2(_29946), .Q(_29944) );
  nnd2s1 _29796_inst ( .DIN1(_27951), .DIN2(_52884), .Q(_29946) );
  nnd2s1 _29797_inst ( .DIN1(_29947), .DIN2(_29948), .Q(_29945) );
  xor2s1 _29798_inst ( .DIN1(_26402), .DIN2(_52885), .Q(_29948) );
  nor2s1 _29799_inst ( .DIN1(_27066), .DIN2(_27955), .Q(_29947) );
  nnd2s1 _29800_inst ( .DIN1(_29949), .DIN2(_29926), .Q(_27955) );
  nor2s1 _29801_inst ( .DIN1(_27571), .DIN2(_29950), .Q(_29942) );
  and2s1 _29802_inst ( .DIN1(______[24]), .DIN2(_53029), .Q(_29950) );
  nnd2s1 _29803_inst ( .DIN1(_29951), .DIN2(_29952), .Q(
        ______________________________28________) );
  nor2s1 _29804_inst ( .DIN1(_29953), .DIN2(_29954), .Q(_29951) );
  nor2s1 _29805_inst ( .DIN1(_29955), .DIN2(_29956), .Q(_29954) );
  nnd2s1 _29806_inst ( .DIN1(_29957), .DIN2(_29911), .Q(_29956) );
  nor2s1 _29807_inst ( .DIN1(_29958), .DIN2(_29959), .Q(_29957) );
  nor2s1 _29808_inst ( .DIN1(_27951), .DIN2(_29960), .Q(_29959) );
  nor2s1 _29809_inst ( .DIN1(_29961), .DIN2(_27291), .Q(_29960) );
  xnr2s1 _29810_inst ( .DIN1(_52887), .DIN2(_29962), .Q(_29961) );
  nor2s1 _29811_inst ( .DIN1(_53274), .DIN2(_29926), .Q(_29958) );
  nor2s1 _29812_inst ( .DIN1(_52886), .DIN2(_29921), .Q(_29953) );
  nnd2s1 _29813_inst ( .DIN1(_29963), .DIN2(_29952), .Q(
        ______________________________27________) );
  nor2s1 _29814_inst ( .DIN1(_29964), .DIN2(_29965), .Q(_29963) );
  nor2s1 _29815_inst ( .DIN1(_29955), .DIN2(_29966), .Q(_29965) );
  nnd2s1 _29816_inst ( .DIN1(_29967), .DIN2(_29911), .Q(_29966) );
  or2s1 _29817_inst ( .DIN1(_29949), .DIN2(_27951), .Q(_29911) );
  nnd2s1 _29818_inst ( .DIN1(_29892), .DIN2(_29968), .Q(_29949) );
  nor2s1 _29819_inst ( .DIN1(_29969), .DIN2(_27977), .Q(_29968) );
  nor2s1 _29820_inst ( .DIN1(_28215), .DIN2(_29970), .Q(_29892) );
  nor2s1 _29821_inst ( .DIN1(_29971), .DIN2(_29972), .Q(_29967) );
  nor2s1 _29822_inst ( .DIN1(_27951), .DIN2(_29920), .Q(_29972) );
  xor2s1 _29823_inst ( .DIN1(_52890), .DIN2(_52889), .Q(_29920) );
  hi1s1 _29824_inst ( .DIN(_29926), .Q(_27951) );
  nor2s1 _29825_inst ( .DIN1(_26508), .DIN2(_29926), .Q(_29971) );
  nnd2s1 _29826_inst ( .DIN1(_29973), .DIN2(_29126), .Q(_29926) );
  nor2s1 _29827_inst ( .DIN1(_28215), .DIN2(_28168), .Q(_29973) );
  nnd2s1 _29828_inst ( .DIN1(_29974), .DIN2(_28938), .Q(_28168) );
  nor2s1 _29829_inst ( .DIN1(_28115), .DIN2(_28110), .Q(_29974) );
  nor2s1 _29830_inst ( .DIN1(_52890), .DIN2(_29921), .Q(_29964) );
  nnd2s1 _29831_inst ( .DIN1(_29975), .DIN2(_29976), .Q(
        ______________________________26________) );
  nor2s1 _29832_inst ( .DIN1(_29977), .DIN2(_29978), .Q(_29976) );
  nor2s1 _29833_inst ( .DIN1(_29919), .DIN2(_29979), .Q(_29978) );
  nnd2s1 _29834_inst ( .DIN1(_52889), .DIN2(_29955), .Q(_29979) );
  nnd2s1 _29835_inst ( .DIN1(_52891), .DIN2(_52890), .Q(_29919) );
  nor2s1 _29836_inst ( .DIN1(_29980), .DIN2(_29981), .Q(_29975) );
  nor2s1 _29837_inst ( .DIN1(_52888), .DIN2(_29982), .Q(_29981) );
  nor2s1 _29838_inst ( .DIN1(_52891), .DIN2(_29983), .Q(_29980) );
  nor2s1 _29839_inst ( .DIN1(_29984), .DIN2(_29985), .Q(_29983) );
  nor2s1 _29840_inst ( .DIN1(_29921), .DIN2(_29986), .Q(_29985) );
  and2s1 _29841_inst ( .DIN1(_52889), .DIN2(_52890), .Q(_29986) );
  nor2s1 _29842_inst ( .DIN1(_27774), .DIN2(_29987), .Q(_29984) );
  nnd2s1 _29843_inst ( .DIN1(_27325), .DIN2(_29988), .Q(
        ______________________________25________) );
  nnd2s1 _29844_inst ( .DIN1(_29989), .DIN2(_29990), .Q(_29988) );
  nnd2s1 _29845_inst ( .DIN1(_29991), .DIN2(_29992), .Q(_29990) );
  xnr2s1 _29846_inst ( .DIN1(_29993), .DIN2(_29994), .Q(_29992) );
  nnd2s1 _29847_inst ( .DIN1(______[20]), .DIN2(_29995), .Q(_29993) );
  nnd2s1 _29848_inst ( .DIN1(_52891), .DIN2(_52889), .Q(_29995) );
  nor2s1 _29849_inst ( .DIN1(_29962), .DIN2(_29996), .Q(_29991) );
  nor2s1 _29850_inst ( .DIN1(_29997), .DIN2(_29998), .Q(_29996) );
  nnd2s1 _29851_inst ( .DIN1(_28214), .DIN2(_29999), .Q(_29998) );
  nor2s1 _29852_inst ( .DIN1(_52889), .DIN2(_52891), .Q(_29962) );
  nnd2s1 _29853_inst ( .DIN1(_30000), .DIN2(_53311), .Q(_29989) );
  nnd2s1 _29854_inst ( .DIN1(_30001), .DIN2(_30002), .Q(
        ______________________________24________) );
  nor2s1 _29855_inst ( .DIN1(_29977), .DIN2(_30003), .Q(_30002) );
  nor2s1 _29856_inst ( .DIN1(_30004), .DIN2(_29987), .Q(_30003) );
  nnd2s1 _29857_inst ( .DIN1(_30005), .DIN2(_29921), .Q(_29987) );
  nor2s1 _29858_inst ( .DIN1(_30000), .DIN2(_30006), .Q(_30005) );
  xor2s1 _29859_inst ( .DIN1(_30007), .DIN2(_30008), .Q(_30004) );
  nor2s1 _29860_inst ( .DIN1(_52918), .DIN2(_52893), .Q(_30008) );
  xor2s1 _29861_inst ( .DIN1(_52930), .DIN2(_26234), .Q(_30007) );
  hi1s1 _29862_inst ( .DIN(_29952), .Q(_29977) );
  nnd2s1 _29863_inst ( .DIN1(_30009), .DIN2(_29955), .Q(_29952) );
  nor2s1 _29864_inst ( .DIN1(_30010), .DIN2(_30011), .Q(_30001) );
  nor2s1 _29865_inst ( .DIN1(_26494), .DIN2(_29982), .Q(_30011) );
  nnd2s1 _29866_inst ( .DIN1(_30000), .DIN2(_29921), .Q(_29982) );
  nor2s1 _29867_inst ( .DIN1(_29921), .DIN2(_30012), .Q(_30010) );
  nor2s1 _29868_inst ( .DIN1(_30013), .DIN2(_27082), .Q(_30012) );
  xor2s1 _29869_inst ( .DIN1(_26475), .DIN2(_52918), .Q(_30013) );
  nnd2s1 _29870_inst ( .DIN1(_30014), .DIN2(_30015), .Q(
        ______________________________23________) );
  nnd2s1 _29871_inst ( .DIN1(_30016), .DIN2(______[14]), .Q(_30015) );
  nor2s1 _29872_inst ( .DIN1(_30009), .DIN2(_30017), .Q(_30016) );
  xor2s1 _29873_inst ( .DIN1(_30018), .DIN2(_26389), .Q(_30017) );
  hi1s1 _29874_inst ( .DIN(_29918), .Q(_30009) );
  nnd2s1 _29875_inst ( .DIN1(_29921), .DIN2(_30019), .Q(_30014) );
  nnd2s1 _29876_inst ( .DIN1(_30020), .DIN2(_30021), .Q(_30019) );
  nor2s1 _29877_inst ( .DIN1(_30022), .DIN2(_30023), .Q(_30020) );
  and2s1 _29878_inst ( .DIN1(_53237), .DIN2(_30000), .Q(_30023) );
  nor2s1 _29879_inst ( .DIN1(_30000), .DIN2(_26389), .Q(_30022) );
  hi1s1 _29880_inst ( .DIN(_29955), .Q(_29921) );
  nnd2s1 _29881_inst ( .DIN1(_30024), .DIN2(_30025), .Q(_29955) );
  nor2s1 _29882_inst ( .DIN1(_30026), .DIN2(_29940), .Q(_30025) );
  nor2s1 _29883_inst ( .DIN1(_30027), .DIN2(_29918), .Q(_30024) );
  nnd2s1 _29884_inst ( .DIN1(_30028), .DIN2(_28887), .Q(_29918) );
  nor2s1 _29885_inst ( .DIN1(_30029), .DIN2(_30030), .Q(_30028) );
  nnd2s1 _29886_inst ( .DIN1(_30031), .DIN2(_30032), .Q(
        ______________________________22________) );
  nnd2s1 _29887_inst ( .DIN1(_30033), .DIN2(_52894), .Q(_30032) );
  nor2s1 _29888_inst ( .DIN1(_28930), .DIN2(_26987), .Q(_30033) );
  nnd2s1 _29889_inst ( .DIN1(_28932), .DIN2(_30034), .Q(_30031) );
  nnd2s1 _29890_inst ( .DIN1(_30035), .DIN2(_30021), .Q(_30034) );
  nor2s1 _29891_inst ( .DIN1(_30036), .DIN2(_30037), .Q(_30035) );
  nor2s1 _29892_inst ( .DIN1(_30000), .DIN2(_26234), .Q(_30037) );
  nor2s1 _29893_inst ( .DIN1(_53385), .DIN2(_30038), .Q(_30036) );
  nnd2s1 _29894_inst ( .DIN1(_30039), .DIN2(_30040), .Q(
        ______________________________21________) );
  nnd2s1 _29895_inst ( .DIN1(_30041), .DIN2(_28069), .Q(_30040) );
  nnd2s1 _29896_inst ( .DIN1(_30042), .DIN2(______[6]), .Q(_30041) );
  nor2s1 _29897_inst ( .DIN1(_30043), .DIN2(_26659), .Q(_30042) );
  nnd2s1 _29898_inst ( .DIN1(_30044), .DIN2(_28060), .Q(_30039) );
  nor2s1 _29899_inst ( .DIN1(_30006), .DIN2(_30045), .Q(_30044) );
  nnd2s1 _29900_inst ( .DIN1(_30046), .DIN2(_30047), .Q(_30045) );
  nnd2s1 _29901_inst ( .DIN1(_30000), .DIN2(_26502), .Q(_30047) );
  nnd2s1 _29902_inst ( .DIN1(_30048), .DIN2(_30038), .Q(_30046) );
  hi1s1 _29903_inst ( .DIN(_30000), .Q(_30038) );
  nnd2s1 _29904_inst ( .DIN1(_30049), .DIN2(______[26]), .Q(_30048) );
  nor2s1 _29905_inst ( .DIN1(_30018), .DIN2(_30050), .Q(_30049) );
  nor2s1 _29906_inst ( .DIN1(_52894), .DIN2(_52918), .Q(_30050) );
  nor2s1 _29907_inst ( .DIN1(_26674), .DIN2(_26234), .Q(_30018) );
  hi1s1 _29908_inst ( .DIN(_30021), .Q(_30006) );
  nnd2s1 _29909_inst ( .DIN1(_30051), .DIN2(_30052), .Q(_30021) );
  nor2s1 _29910_inst ( .DIN1(_29894), .DIN2(_28116), .Q(_30052) );
  nor2s1 _29911_inst ( .DIN1(_30000), .DIN2(_29997), .Q(_30051) );
  nor2s1 _29912_inst ( .DIN1(_28804), .DIN2(_29970), .Q(_30000) );
  or2s1 _29913_inst ( .DIN1(_30053), .DIN2(_29904), .Q(_29970) );
  hi1s1 _29914_inst ( .DIN(_28935), .Q(_28804) );
  nor2s1 _29915_inst ( .DIN1(_30054), .DIN2(_29902), .Q(_28935) );
  nnd2s1 _29916_inst ( .DIN1(_30055), .DIN2(_30056), .Q(
        ______________________________20________) );
  nnd2s1 _29917_inst ( .DIN1(_30057), .DIN2(_30058), .Q(_30056) );
  nnd2s1 _29918_inst ( .DIN1(_30059), .DIN2(______[30]), .Q(_30058) );
  xor2s1 _29919_inst ( .DIN1(_30060), .DIN2(_53144), .Q(_30059) );
  nor2s1 _29920_inst ( .DIN1(_30061), .DIN2(_30062), .Q(_30055) );
  nor2s1 _29921_inst ( .DIN1(_30063), .DIN2(_28329), .Q(_30062) );
  nor2s1 _29922_inst ( .DIN1(_30064), .DIN2(_30065), .Q(_30063) );
  nor2s1 _29923_inst ( .DIN1(_26544), .DIN2(_30066), .Q(_30064) );
  nor2s1 _29924_inst ( .DIN1(_30067), .DIN2(_30068), .Q(_30061) );
  xor2s1 _29925_inst ( .DIN1(_26393), .DIN2(_52851), .Q(_30067) );
  nnd2s1 _29926_inst ( .DIN1(_30069), .DIN2(_29181), .Q(
        ______________________________1________) );
  nor2s1 _29927_inst ( .DIN1(_30070), .DIN2(_30071), .Q(_30069) );
  nor2s1 _29928_inst ( .DIN1(_29184), .DIN2(_30072), .Q(_30071) );
  nor2s1 _29929_inst ( .DIN1(_30073), .DIN2(_30074), .Q(_30072) );
  nor2s1 _29930_inst ( .DIN1(_28724), .DIN2(_30075), .Q(_30074) );
  nor2s1 _29931_inst ( .DIN1(_27651), .DIN2(_30076), .Q(_30075) );
  nnd2s1 _29932_inst ( .DIN1(_30077), .DIN2(_28844), .Q(_30076) );
  xor2s1 _29933_inst ( .DIN1(_52880), .DIN2(_52896), .Q(_30077) );
  nor2s1 _29934_inst ( .DIN1(_53064), .DIN2(_28705), .Q(_30073) );
  nor2s1 _29935_inst ( .DIN1(_53180), .DIN2(_29206), .Q(_30070) );
  nor2s1 _29936_inst ( .DIN1(_30078), .DIN2(_27749), .Q(
        ______________________________19________) );
  nor2s1 _29937_inst ( .DIN1(_30079), .DIN2(_30080), .Q(_30078) );
  xor2s1 _29938_inst ( .DIN1(_30081), .DIN2(_30082), .Q(_30080) );
  nnd2s1 _29939_inst ( .DIN1(_30083), .DIN2(_30084), .Q(_30082) );
  nnd2s1 _29940_inst ( .DIN1(_30085), .DIN2(_52849), .Q(_30084) );
  nor2s1 _29941_inst ( .DIN1(_30085), .DIN2(_30086), .Q(_30079) );
  xor2s1 _29942_inst ( .DIN1(_30060), .DIN2(_52897), .Q(_30086) );
  nnd2s1 _29943_inst ( .DIN1(_52908), .DIN2(_53162), .Q(_30060) );
  nnd2s1 _29944_inst ( .DIN1(_30087), .DIN2(_30088), .Q(
        ______________________________192________) );
  nnd2s1 _29945_inst ( .DIN1(_30089), .DIN2(_29039), .Q(_30088) );
  nor2s1 _29946_inst ( .DIN1(_30090), .DIN2(_26773), .Q(_30089) );
  xor2s1 _29947_inst ( .DIN1(_30091), .DIN2(_30092), .Q(_30090) );
  xor2s1 _29948_inst ( .DIN1(_52883), .DIN2(_52898), .Q(_30092) );
  nnd2s1 _29949_inst ( .DIN1(_52899), .DIN2(_52898), .Q(_30091) );
  nnd2s1 _29950_inst ( .DIN1(_28738), .DIN2(_30093), .Q(_30087) );
  nnd2s1 _29951_inst ( .DIN1(_30094), .DIN2(_30095), .Q(_30093) );
  nnd2s1 _29952_inst ( .DIN1(_30096), .DIN2(_30097), .Q(_30095) );
  xor2s1 _29953_inst ( .DIN1(_30098), .DIN2(_52953), .Q(_30097) );
  nnd2s1 _29954_inst ( .DIN1(_53464), .DIN2(_52900), .Q(_30098) );
  nor2s1 _29955_inst ( .DIN1(_28129), .DIN2(_27448), .Q(_30096) );
  nnd2s1 _29956_inst ( .DIN1(_30099), .DIN2(_30100), .Q(_30094) );
  xor2s1 _29957_inst ( .DIN1(_30101), .DIN2(_30102), .Q(_30100) );
  xor2s1 _29958_inst ( .DIN1(_30103), .DIN2(_30104), .Q(_30102) );
  nnd2s1 _29959_inst ( .DIN1(_30105), .DIN2(_30106), .Q(_30103) );
  nnd2s1 _29960_inst ( .DIN1(_30107), .DIN2(_26472), .Q(_30106) );
  nnd2s1 _29961_inst ( .DIN1(_30108), .DIN2(_30109), .Q(_30107) );
  or2s1 _29962_inst ( .DIN1(_30109), .DIN2(_30108), .Q(_30105) );
  xor2s1 _29963_inst ( .DIN1(_26498), .DIN2(_30110), .Q(_30101) );
  nnd2s1 _29964_inst ( .DIN1(_30111), .DIN2(_30112), .Q(
        ______________________________191________) );
  nor2s1 _29965_inst ( .DIN1(_30113), .DIN2(_30114), .Q(_30111) );
  nor2s1 _29966_inst ( .DIN1(_28032), .DIN2(_30115), .Q(_30114) );
  nnd2s1 _29967_inst ( .DIN1(_30116), .DIN2(_30117), .Q(_30115) );
  nnd2s1 _29968_inst ( .DIN1(_30118), .DIN2(_30099), .Q(_30117) );
  xnr2s1 _29969_inst ( .DIN1(_30108), .DIN2(_30119), .Q(_30118) );
  xor2s1 _29970_inst ( .DIN1(_26472), .DIN2(_30109), .Q(_30119) );
  nnd2s1 _29971_inst ( .DIN1(_30120), .DIN2(_30121), .Q(_30109) );
  nnd2s1 _29972_inst ( .DIN1(_30122), .DIN2(_30123), .Q(_30121) );
  and2s1 _29973_inst ( .DIN1(_30124), .DIN2(_30110), .Q(_30108) );
  nnd2s1 _29974_inst ( .DIN1(_52900), .DIN2(_28223), .Q(_30116) );
  nor2s1 _29975_inst ( .DIN1(_53463), .DIN2(_28037), .Q(_30113) );
  nnd2s1 _29976_inst ( .DIN1(_30125), .DIN2(_30126), .Q(
        ______________________________190________) );
  nnd2s1 _29977_inst ( .DIN1(_30127), .DIN2(_28084), .Q(_30126) );
  nnd2s1 _29978_inst ( .DIN1(_30128), .DIN2(_30129), .Q(_30127) );
  xor2s1 _29979_inst ( .DIN1(_26377), .DIN2(_30130), .Q(_30128) );
  nnd2s1 _29980_inst ( .DIN1(_52902), .DIN2(_53273), .Q(_30130) );
  nnd2s1 _29981_inst ( .DIN1(_30131), .DIN2(_27183), .Q(_30125) );
  nnd2s1 _29982_inst ( .DIN1(_30132), .DIN2(_30133), .Q(_30131) );
  nnd2s1 _29983_inst ( .DIN1(_30134), .DIN2(_30135), .Q(_30133) );
  nnd2s1 _29984_inst ( .DIN1(_30136), .DIN2(______[22]), .Q(_30134) );
  nor2s1 _29985_inst ( .DIN1(_30137), .DIN2(_30138), .Q(_30136) );
  xor2s1 _29986_inst ( .DIN1(_30139), .DIN2(_53002), .Q(_30138) );
  nnd2s1 _29987_inst ( .DIN1(_52902), .DIN2(_53040), .Q(_30139) );
  nnd2s1 _29988_inst ( .DIN1(_30140), .DIN2(_30141), .Q(_30132) );
  xor2s1 _29989_inst ( .DIN1(_30142), .DIN2(_30122), .Q(_30140) );
  and2s1 _29990_inst ( .DIN1(_30143), .DIN2(_30110), .Q(_30122) );
  nnd2s1 _29991_inst ( .DIN1(_30123), .DIN2(_30120), .Q(_30142) );
  nnd2s1 _29992_inst ( .DIN1(_30144), .DIN2(_26584), .Q(_30120) );
  or2s1 _29993_inst ( .DIN1(_30144), .DIN2(_26584), .Q(_30123) );
  nnd2s1 _29994_inst ( .DIN1(_30145), .DIN2(_30146), .Q(_30144) );
  nnd2s1 _29995_inst ( .DIN1(_52927), .DIN2(_30147), .Q(_30146) );
  nnd2s1 _29996_inst ( .DIN1(_30148), .DIN2(_30149), .Q(_30147) );
  or2s1 _29997_inst ( .DIN1(_30149), .DIN2(_30148), .Q(_30145) );
  hi1s1 _29998_inst ( .DIN(_30150), .Q(_30148) );
  nnd2s1 _29999_inst ( .DIN1(_30151), .DIN2(_28782), .Q(
        ______________________________18________) );
  nor2s1 _30000_inst ( .DIN1(_30152), .DIN2(_30153), .Q(_30151) );
  nor2s1 _30001_inst ( .DIN1(_30154), .DIN2(_28786), .Q(_30153) );
  nor2s1 _30002_inst ( .DIN1(_30155), .DIN2(_30156), .Q(_30154) );
  nnd2s1 _30003_inst ( .DIN1(_30157), .DIN2(_30158), .Q(_30156) );
  nnd2s1 _30004_inst ( .DIN1(_30159), .DIN2(_28521), .Q(_30158) );
  nor2s1 _30005_inst ( .DIN1(_30160), .DIN2(_30161), .Q(_30159) );
  nnd2s1 _30006_inst ( .DIN1(_30162), .DIN2(_30066), .Q(_30161) );
  nnd2s1 _30007_inst ( .DIN1(_30163), .DIN2(_30164), .Q(_30157) );
  nnd2s1 _30008_inst ( .DIN1(_30083), .DIN2(_30165), .Q(_30164) );
  nnd2s1 _30009_inst ( .DIN1(_30160), .DIN2(_30066), .Q(_30165) );
  nnd2s1 _30010_inst ( .DIN1(_52908), .DIN2(______[22]), .Q(_30160) );
  nor2s1 _30011_inst ( .DIN1(_26264), .DIN2(_30066), .Q(_30155) );
  nor2s1 _30012_inst ( .DIN1(_28792), .DIN2(_30166), .Q(_30152) );
  nor2s1 _30013_inst ( .DIN1(_27066), .DIN2(_30167), .Q(_30166) );
  xor2s1 _30014_inst ( .DIN1(_26463), .DIN2(_30168), .Q(_30167) );
  nnd2s1 _30015_inst ( .DIN1(_30169), .DIN2(_30170), .Q(
        ______________________________189________) );
  nnd2s1 _30016_inst ( .DIN1(_30171), .DIN2(_30172), .Q(_30170) );
  xor2s1 _30017_inst ( .DIN1(_30173), .DIN2(_52901), .Q(_30172) );
  nnd2s1 _30018_inst ( .DIN1(_53072), .DIN2(_53328), .Q(_30173) );
  nor2s1 _30019_inst ( .DIN1(_26809), .DIN2(_30174), .Q(_30171) );
  nnd2s1 _30020_inst ( .DIN1(_30175), .DIN2(_30176), .Q(_30169) );
  nnd2s1 _30021_inst ( .DIN1(_30177), .DIN2(_30178), .Q(_30176) );
  nnd2s1 _30022_inst ( .DIN1(_30179), .DIN2(_52902), .Q(_30178) );
  nor2s1 _30023_inst ( .DIN1(_27614), .DIN2(_30180), .Q(_30179) );
  nnd2s1 _30024_inst ( .DIN1(_30181), .DIN2(_30141), .Q(_30177) );
  xor2s1 _30025_inst ( .DIN1(_30149), .DIN2(_30182), .Q(_30181) );
  xor2s1 _30026_inst ( .DIN1(_26583), .DIN2(_30150), .Q(_30182) );
  nnd2s1 _30027_inst ( .DIN1(_30183), .DIN2(_30184), .Q(_30150) );
  nnd2s1 _30028_inst ( .DIN1(_53019), .DIN2(_30185), .Q(_30184) );
  xor2s1 _30029_inst ( .DIN1(_30186), .DIN2(_30187), .Q(_30183) );
  nnd2s1 _30030_inst ( .DIN1(_30188), .DIN2(_30189), .Q(_30187) );
  or2s1 _30031_inst ( .DIN1(_30185), .DIN2(_53019), .Q(_30189) );
  nnd2s1 _30032_inst ( .DIN1(_30190), .DIN2(_30110), .Q(_30149) );
  nnd2s1 _30033_inst ( .DIN1(_30191), .DIN2(_30192), .Q(
        ______________________________188________) );
  nor2s1 _30034_inst ( .DIN1(_28654), .DIN2(_30193), .Q(_30192) );
  nor2s1 _30035_inst ( .DIN1(_28696), .DIN2(_30194), .Q(_30193) );
  xnr2s1 _30036_inst ( .DIN1(_30188), .DIN2(_30195), .Q(_30194) );
  xor2s1 _30037_inst ( .DIN1(_53019), .DIN2(_30185), .Q(_30195) );
  nnd2s1 _30038_inst ( .DIN1(_30196), .DIN2(_30197), .Q(_30185) );
  nnd2s1 _30039_inst ( .DIN1(_30198), .DIN2(_30199), .Q(_30197) );
  and2s1 _30040_inst ( .DIN1(_30200), .DIN2(_30110), .Q(_30188) );
  nnd2s1 _30041_inst ( .DIN1(_30141), .DIN2(_28650), .Q(_28696) );
  nor2s1 _30042_inst ( .DIN1(_30201), .DIN2(_30202), .Q(_30191) );
  nor2s1 _30043_inst ( .DIN1(_28650), .DIN2(_30203), .Q(_30202) );
  nor2s1 _30044_inst ( .DIN1(_30204), .DIN2(_26773), .Q(_30203) );
  xor2s1 _30045_inst ( .DIN1(_30205), .DIN2(_30206), .Q(_30204) );
  xor2s1 _30046_inst ( .DIN1(_52910), .DIN2(_52911), .Q(_30206) );
  nor2s1 _30047_inst ( .DIN1(_30207), .DIN2(_28694), .Q(_30201) );
  or2s1 _30048_inst ( .DIN1(_30180), .DIN2(_28657), .Q(_28694) );
  xor2s1 _30049_inst ( .DIN1(_26728), .DIN2(_53002), .Q(_30207) );
  nnd2s1 _30050_inst ( .DIN1(_30208), .DIN2(_27126), .Q(
        ______________________________187________) );
  nor2s1 _30051_inst ( .DIN1(_30209), .DIN2(_30210), .Q(_30208) );
  nor2s1 _30052_inst ( .DIN1(_27132), .DIN2(_30211), .Q(_30210) );
  nor2s1 _30053_inst ( .DIN1(_30212), .DIN2(_30213), .Q(_30211) );
  nor2s1 _30054_inst ( .DIN1(_30135), .DIN2(_30214), .Q(_30213) );
  xnr2s1 _30055_inst ( .DIN1(_30198), .DIN2(_30215), .Q(_30214) );
  nnd2s1 _30056_inst ( .DIN1(_30199), .DIN2(_30196), .Q(_30215) );
  nnd2s1 _30057_inst ( .DIN1(_30216), .DIN2(_26250), .Q(_30196) );
  or2s1 _30058_inst ( .DIN1(_30216), .DIN2(_26250), .Q(_30199) );
  nnd2s1 _30059_inst ( .DIN1(_30217), .DIN2(_30218), .Q(_30216) );
  nnd2s1 _30060_inst ( .DIN1(_30219), .DIN2(_30220), .Q(_30218) );
  and2s1 _30061_inst ( .DIN1(_30221), .DIN2(_30110), .Q(_30198) );
  nor2s1 _30062_inst ( .DIN1(_30141), .DIN2(_30222), .Q(_30212) );
  nor2s1 _30063_inst ( .DIN1(_30137), .DIN2(_30223), .Q(_30222) );
  xor2s1 _30064_inst ( .DIN1(_30224), .DIN2(_30225), .Q(_30223) );
  nor2s1 _30065_inst ( .DIN1(_52910), .DIN2(_26382), .Q(_30225) );
  xor2s1 _30066_inst ( .DIN1(_53173), .DIN2(_26382), .Q(_30224) );
  hi1s1 _30067_inst ( .DIN(_30226), .Q(_30137) );
  hi1s1 _30068_inst ( .DIN(_30135), .Q(_30141) );
  nor2s1 _30069_inst ( .DIN1(_27129), .DIN2(_26427), .Q(_30209) );
  nnd2s1 _30070_inst ( .DIN1(_30227), .DIN2(_30228), .Q(
        ______________________________186________) );
  nor2s1 _30071_inst ( .DIN1(_30229), .DIN2(_30230), .Q(_30227) );
  nor2s1 _30072_inst ( .DIN1(_29560), .DIN2(_30231), .Q(_30230) );
  nor2s1 _30073_inst ( .DIN1(_53288), .DIN2(_27614), .Q(_30231) );
  nor2s1 _30074_inst ( .DIN1(_30232), .DIN2(_29555), .Q(_30229) );
  nor2s1 _30075_inst ( .DIN1(_30233), .DIN2(_30234), .Q(_30232) );
  nor2s1 _30076_inst ( .DIN1(_30180), .DIN2(_26679), .Q(_30234) );
  nnd2s1 _30077_inst ( .DIN1(_30226), .DIN2(_30135), .Q(_30180) );
  nor2s1 _30078_inst ( .DIN1(_30235), .DIN2(_30135), .Q(_30233) );
  nnd2s1 _30079_inst ( .DIN1(_29846), .DIN2(_30236), .Q(_30135) );
  xnr2s1 _30080_inst ( .DIN1(_30219), .DIN2(_30237), .Q(_30235) );
  and2s1 _30081_inst ( .DIN1(_30220), .DIN2(_30217), .Q(_30237) );
  nnd2s1 _30082_inst ( .DIN1(_30238), .DIN2(_52934), .Q(_30217) );
  nor2s1 _30083_inst ( .DIN1(_30239), .DIN2(_30240), .Q(_30238) );
  nor2s1 _30084_inst ( .DIN1(_30241), .DIN2(_26368), .Q(_30239) );
  and2s1 _30085_inst ( .DIN1(_30242), .DIN2(_30243), .Q(_30241) );
  nnd2s1 _30086_inst ( .DIN1(_30244), .DIN2(_30245), .Q(_30220) );
  nnd2s1 _30087_inst ( .DIN1(_30243), .DIN2(_30242), .Q(_30245) );
  nor2s1 _30088_inst ( .DIN1(_52934), .DIN2(_30246), .Q(_30244) );
  nor2s1 _30089_inst ( .DIN1(_52904), .DIN2(_30240), .Q(_30246) );
  nor2s1 _30090_inst ( .DIN1(_30243), .DIN2(_30242), .Q(_30240) );
  hi1s1 _30091_inst ( .DIN(_30247), .Q(_30243) );
  and2s1 _30092_inst ( .DIN1(_30248), .DIN2(_30110), .Q(_30219) );
  nnd2s1 _30093_inst ( .DIN1(_30249), .DIN2(_30250), .Q(
        ______________________________185________) );
  hi1s1 _30094_inst ( .DIN(_28654), .Q(_30250) );
  nor2s1 _30095_inst ( .DIN1(_30251), .DIN2(_28650), .Q(_28654) );
  nor2s1 _30096_inst ( .DIN1(_30252), .DIN2(_30253), .Q(_30249) );
  nor2s1 _30097_inst ( .DIN1(_28657), .DIN2(_30254), .Q(_30253) );
  nor2s1 _30098_inst ( .DIN1(_30255), .DIN2(_30256), .Q(_30254) );
  nor2s1 _30099_inst ( .DIN1(_30257), .DIN2(_30258), .Q(_30256) );
  xor2s1 _30100_inst ( .DIN1(_30242), .DIN2(_30259), .Q(_30258) );
  xor2s1 _30101_inst ( .DIN1(_26368), .DIN2(_30247), .Q(_30259) );
  nnd2s1 _30102_inst ( .DIN1(_30110), .DIN2(_30260), .Q(_30247) );
  nnd2s1 _30103_inst ( .DIN1(_30261), .DIN2(_30262), .Q(_30260) );
  hi1s1 _30104_inst ( .DIN(_30263), .Q(_30261) );
  nnd2s1 _30105_inst ( .DIN1(_30264), .DIN2(_30263), .Q(_30110) );
  nnd2s1 _30106_inst ( .DIN1(_30265), .DIN2(_30266), .Q(_30242) );
  nnd2s1 _30107_inst ( .DIN1(_30267), .DIN2(_26511), .Q(_30266) );
  nnd2s1 _30108_inst ( .DIN1(_30268), .DIN2(_30269), .Q(_30267) );
  or2s1 _30109_inst ( .DIN1(_30268), .DIN2(_30269), .Q(_30265) );
  nor2s1 _30110_inst ( .DIN1(_30270), .DIN2(_30271), .Q(_30255) );
  nnd2s1 _30111_inst ( .DIN1(_30272), .DIN2(_53289), .Q(_30271) );
  nor2s1 _30112_inst ( .DIN1(_52903), .DIN2(_28650), .Q(_30252) );
  nnd2s1 _30113_inst ( .DIN1(_30273), .DIN2(_30274), .Q(
        ______________________________184________) );
  nnd2s1 _30114_inst ( .DIN1(_27183), .DIN2(_30275), .Q(_30274) );
  nnd2s1 _30115_inst ( .DIN1(_30276), .DIN2(_30277), .Q(_30275) );
  nnd2s1 _30116_inst ( .DIN1(_30278), .DIN2(_30270), .Q(_30277) );
  xor2s1 _30117_inst ( .DIN1(_30269), .DIN2(_30279), .Q(_30278) );
  xor2s1 _30118_inst ( .DIN1(_26511), .DIN2(_30268), .Q(_30279) );
  nnd2s1 _30119_inst ( .DIN1(_30262), .DIN2(_30280), .Q(_30268) );
  nnd2s1 _30120_inst ( .DIN1(_30281), .DIN2(_30282), .Q(_30280) );
  hi1s1 _30121_inst ( .DIN(_30264), .Q(_30262) );
  nor2s1 _30122_inst ( .DIN1(_30282), .DIN2(_30281), .Q(_30264) );
  nnd2s1 _30123_inst ( .DIN1(_30283), .DIN2(_30284), .Q(_30282) );
  nnd2s1 _30124_inst ( .DIN1(_30285), .DIN2(_30286), .Q(_30269) );
  nnd2s1 _30125_inst ( .DIN1(_52944), .DIN2(_30287), .Q(_30286) );
  nnd2s1 _30126_inst ( .DIN1(_30288), .DIN2(_30289), .Q(_30287) );
  or2s1 _30127_inst ( .DIN1(_30289), .DIN2(_30288), .Q(_30285) );
  nor2s1 _30128_inst ( .DIN1(_30290), .DIN2(_30291), .Q(_30276) );
  nor2s1 _30129_inst ( .DIN1(_26282), .DIN2(_30292), .Q(_30291) );
  nnd2s1 _30130_inst ( .DIN1(_30293), .DIN2(_53173), .Q(_30292) );
  nor2s1 _30131_inst ( .DIN1(_30294), .DIN2(_26382), .Q(_30293) );
  nor2s1 _30132_inst ( .DIN1(_52910), .DIN2(_30295), .Q(_30290) );
  nnd2s1 _30133_inst ( .DIN1(_30296), .DIN2(_30297), .Q(_30295) );
  nnd2s1 _30134_inst ( .DIN1(_53173), .DIN2(_53289), .Q(_30297) );
  nnd2s1 _30135_inst ( .DIN1(_52836), .DIN2(_30298), .Q(_30273) );
  nor2s1 _30136_inst ( .DIN1(_28925), .DIN2(_30299), .Q(
        ______________________________183________) );
  nnd2s1 _30137_inst ( .DIN1(_30300), .DIN2(_30301), .Q(_30299) );
  nnd2s1 _30138_inst ( .DIN1(_30302), .DIN2(_30270), .Q(_30301) );
  xnr2s1 _30139_inst ( .DIN1(_30303), .DIN2(_30288), .Q(_30302) );
  xor2s1 _30140_inst ( .DIN1(_30283), .DIN2(_30284), .Q(_30288) );
  xor2s1 _30141_inst ( .DIN1(_30289), .DIN2(_52944), .Q(_30303) );
  nnd2s1 _30142_inst ( .DIN1(_30304), .DIN2(_30305), .Q(_30289) );
  nnd2s1 _30143_inst ( .DIN1(_30306), .DIN2(_26522), .Q(_30305) );
  nnd2s1 _30144_inst ( .DIN1(_30307), .DIN2(_30308), .Q(_30306) );
  or2s1 _30145_inst ( .DIN1(_30307), .DIN2(_30308), .Q(_30304) );
  nnd2s1 _30146_inst ( .DIN1(_30309), .DIN2(_30257), .Q(_30300) );
  nor2s1 _30147_inst ( .DIN1(_30310), .DIN2(_30294), .Q(_30309) );
  xor2s1 _30148_inst ( .DIN1(_52905), .DIN2(_30311), .Q(_30310) );
  nnd2s1 _30149_inst ( .DIN1(_30312), .DIN2(_30313), .Q(
        ______________________________182________) );
  nnd2s1 _30150_inst ( .DIN1(_28060), .DIN2(_30314), .Q(_30313) );
  nnd2s1 _30151_inst ( .DIN1(_30315), .DIN2(_30316), .Q(_30314) );
  nnd2s1 _30152_inst ( .DIN1(_30272), .DIN2(_30317), .Q(_30316) );
  xor2s1 _30153_inst ( .DIN1(_30311), .DIN2(_26481), .Q(_30317) );
  nor2s1 _30154_inst ( .DIN1(_30294), .DIN2(_28646), .Q(_30272) );
  nnd2s1 _30155_inst ( .DIN1(_30318), .DIN2(_30270), .Q(_30315) );
  xor2s1 _30156_inst ( .DIN1(_30319), .DIN2(_30320), .Q(_30318) );
  xor2s1 _30157_inst ( .DIN1(_30307), .DIN2(_30308), .Q(_30320) );
  nnd2s1 _30158_inst ( .DIN1(_30321), .DIN2(_30322), .Q(_30308) );
  nnd2s1 _30159_inst ( .DIN1(_52906), .DIN2(_30323), .Q(_30322) );
  or2s1 _30160_inst ( .DIN1(_30324), .DIN2(_30325), .Q(_30323) );
  nnd2s1 _30161_inst ( .DIN1(_30325), .DIN2(_30324), .Q(_30321) );
  nnd2s1 _30162_inst ( .DIN1(_30326), .DIN2(_30327), .Q(_30307) );
  nnd2s1 _30163_inst ( .DIN1(_30328), .DIN2(_30329), .Q(_30327) );
  hi1s1 _30164_inst ( .DIN(_30283), .Q(_30326) );
  nor2s1 _30165_inst ( .DIN1(_30329), .DIN2(_30328), .Q(_30283) );
  xor2s1 _30166_inst ( .DIN1(_26522), .DIN2(_2064), .Q(_30319) );
  nnd2s1 _30167_inst ( .DIN1(_30330), .DIN2(_28069), .Q(_30312) );
  nor2s1 _30168_inst ( .DIN1(_28684), .DIN2(_30331), .Q(_30330) );
  nnd2s1 _30169_inst ( .DIN1(_30332), .DIN2(_28071), .Q(_30331) );
  xor2s1 _30170_inst ( .DIN1(_30333), .DIN2(_30334), .Q(_30332) );
  xor2s1 _30171_inst ( .DIN1(_52927), .DIN2(_52981), .Q(_30334) );
  nnd2s1 _30172_inst ( .DIN1(_52930), .DIN2(_52907), .Q(_30333) );
  nnd2s1 _30173_inst ( .DIN1(_30335), .DIN2(_30336), .Q(
        ______________________________181________) );
  nnd2s1 _30174_inst ( .DIN1(_30337), .DIN2(_28657), .Q(_30336) );
  nor2s1 _30175_inst ( .DIN1(_26282), .DIN2(_30338), .Q(_30337) );
  nnd2s1 _30176_inst ( .DIN1(_26856), .DIN2(_30251), .Q(_30338) );
  nnd2s1 _30177_inst ( .DIN1(_30339), .DIN2(_28650), .Q(_30335) );
  nnd2s1 _30178_inst ( .DIN1(_30340), .DIN2(_30341), .Q(_30339) );
  nnd2s1 _30179_inst ( .DIN1(_30342), .DIN2(_30257), .Q(_30341) );
  nnd2s1 _30180_inst ( .DIN1(_30343), .DIN2(_52907), .Q(_30342) );
  nor2s1 _30181_inst ( .DIN1(_30294), .DIN2(_27365), .Q(_30343) );
  nnd2s1 _30182_inst ( .DIN1(_30344), .DIN2(_30270), .Q(_30340) );
  xnr2s1 _30183_inst ( .DIN1(_30325), .DIN2(_30345), .Q(_30344) );
  xor2s1 _30184_inst ( .DIN1(_26302), .DIN2(_30324), .Q(_30345) );
  nnd2s1 _30185_inst ( .DIN1(_30346), .DIN2(_30329), .Q(_30324) );
  or2s1 _30186_inst ( .DIN1(_30347), .DIN2(_30348), .Q(_30329) );
  xor2s1 _30187_inst ( .DIN1(_30349), .DIN2(_30350), .Q(_30346) );
  nnd2s1 _30188_inst ( .DIN1(_30348), .DIN2(_30347), .Q(_30350) );
  nnd2s1 _30189_inst ( .DIN1(_30351), .DIN2(_30352), .Q(_30325) );
  nnd2s1 _30190_inst ( .DIN1(_52936), .DIN2(_30353), .Q(_30352) );
  or2s1 _30191_inst ( .DIN1(_30354), .DIN2(_30355), .Q(_30353) );
  nnd2s1 _30192_inst ( .DIN1(_30355), .DIN2(_30354), .Q(_30351) );
  nnd2s1 _30193_inst ( .DIN1(_30356), .DIN2(_27050), .Q(
        ______________________________180________) );
  nor2s1 _30194_inst ( .DIN1(_30357), .DIN2(_30358), .Q(_30356) );
  nor2s1 _30195_inst ( .DIN1(_27053), .DIN2(_30359), .Q(_30358) );
  xor2s1 _30196_inst ( .DIN1(_30360), .DIN2(_30361), .Q(_30359) );
  nnd2s1 _30197_inst ( .DIN1(_30362), .DIN2(_30363), .Q(_30361) );
  nnd2s1 _30198_inst ( .DIN1(_30364), .DIN2(_30257), .Q(_30363) );
  nnd2s1 _30199_inst ( .DIN1(_30365), .DIN2(_30296), .Q(_30364) );
  hi1s1 _30200_inst ( .DIN(_30294), .Q(_30296) );
  xor2s1 _30201_inst ( .DIN1(_30366), .DIN2(_30367), .Q(_30294) );
  or2s1 _30202_inst ( .DIN1(_30368), .DIN2(_30369), .Q(_30366) );
  nor2s1 _30203_inst ( .DIN1(_30311), .DIN2(_30370), .Q(_30365) );
  and2s1 _30204_inst ( .DIN1(_26459), .DIN2(_52832), .Q(_30370) );
  nor2s1 _30205_inst ( .DIN1(_26459), .DIN2(_52832), .Q(_30311) );
  nnd2s1 _30206_inst ( .DIN1(_30371), .DIN2(_30270), .Q(_30362) );
  hi1s1 _30207_inst ( .DIN(_30257), .Q(_30270) );
  nnd2s1 _30208_inst ( .DIN1(_30372), .DIN2(_30373), .Q(_30257) );
  nor2s1 _30209_inst ( .DIN1(_30374), .DIN2(_30375), .Q(_30373) );
  nor2s1 _30210_inst ( .DIN1(_30369), .DIN2(_30376), .Q(_30372) );
  xnr2s1 _30211_inst ( .DIN1(_30355), .DIN2(_30377), .Q(_30371) );
  xnr2s1 _30212_inst ( .DIN1(_52936), .DIN2(_30354), .Q(_30377) );
  nnd2s1 _30213_inst ( .DIN1(_30378), .DIN2(_30379), .Q(_30354) );
  nnd2s1 _30214_inst ( .DIN1(_52938), .DIN2(_30380), .Q(_30379) );
  nnd2s1 _30215_inst ( .DIN1(_30381), .DIN2(_30382), .Q(_30380) );
  or2s1 _30216_inst ( .DIN1(_30382), .DIN2(_30381), .Q(_30378) );
  nnd2s1 _30217_inst ( .DIN1(_30347), .DIN2(_30383), .Q(_30355) );
  nnd2s1 _30218_inst ( .DIN1(_30384), .DIN2(_30385), .Q(_30383) );
  nnd2s1 _30219_inst ( .DIN1(_30386), .DIN2(_30387), .Q(_30385) );
  nnd2s1 _30220_inst ( .DIN1(_30388), .DIN2(_30386), .Q(_30347) );
  nor2s1 _30221_inst ( .DIN1(_30389), .DIN2(_30384), .Q(_30388) );
  nor2s1 _30222_inst ( .DIN1(_27064), .DIN2(_30390), .Q(_30357) );
  xor2s1 _30223_inst ( .DIN1(_30391), .DIN2(_30392), .Q(_30390) );
  xor2s1 _30224_inst ( .DIN1(_26492), .DIN2(_52991), .Q(_30392) );
  nnd2s1 _30225_inst ( .DIN1(_30393), .DIN2(_30394), .Q(
        ______________________________17________) );
  nnd2s1 _30226_inst ( .DIN1(_30395), .DIN2(_30083), .Q(_30394) );
  nnd2s1 _30227_inst ( .DIN1(_30396), .DIN2(_30397), .Q(_30395) );
  nnd2s1 _30228_inst ( .DIN1(_30398), .DIN2(_30085), .Q(_30397) );
  nor2s1 _30229_inst ( .DIN1(_26599), .DIN2(_28329), .Q(_30398) );
  nnd2s1 _30230_inst ( .DIN1(_30057), .DIN2(_30399), .Q(_30396) );
  xor2s1 _30231_inst ( .DIN1(_52908), .DIN2(_53162), .Q(_30399) );
  nor2s1 _30232_inst ( .DIN1(_28329), .DIN2(_30085), .Q(_30057) );
  nor2s1 _30233_inst ( .DIN1(_30400), .DIN2(_30401), .Q(_30393) );
  nor2s1 _30234_inst ( .DIN1(_28338), .DIN2(_30402), .Q(_30401) );
  xor2s1 _30235_inst ( .DIN1(_53096), .DIN2(_53143), .Q(_30402) );
  nnd2s1 _30236_inst ( .DIN1(_30403), .DIN2(_30404), .Q(
        ______________________________179________) );
  nnd2s1 _30237_inst ( .DIN1(_30405), .DIN2(_28657), .Q(_30404) );
  hi1s1 _30238_inst ( .DIN(_28650), .Q(_28657) );
  nnd2s1 _30239_inst ( .DIN1(_30406), .DIN2(_28689), .Q(_30405) );
  and2s1 _30240_inst ( .DIN1(______[18]), .DIN2(_30251), .Q(_28689) );
  nnd2s1 _30241_inst ( .DIN1(_28888), .DIN2(_30407), .Q(_30251) );
  hi1s1 _30242_inst ( .DIN(_29938), .Q(_28888) );
  nor2s1 _30243_inst ( .DIN1(_30408), .DIN2(_30409), .Q(_30406) );
  nor2s1 _30244_inst ( .DIN1(_26670), .DIN2(_30205), .Q(_30409) );
  nnd2s1 _30245_inst ( .DIN1(_52832), .DIN2(_52910), .Q(_30205) );
  nor2s1 _30246_inst ( .DIN1(_52832), .DIN2(_30410), .Q(_30408) );
  nor2s1 _30247_inst ( .DIN1(_26282), .DIN2(_26670), .Q(_30410) );
  nnd2s1 _30248_inst ( .DIN1(_28650), .DIN2(_30411), .Q(_30403) );
  nnd2s1 _30249_inst ( .DIN1(_30412), .DIN2(_30413), .Q(_30411) );
  nnd2s1 _30250_inst ( .DIN1(_30414), .DIN2(_30415), .Q(_30413) );
  xor2s1 _30251_inst ( .DIN1(_30381), .DIN2(_30416), .Q(_30414) );
  xnr2s1 _30252_inst ( .DIN1(_52938), .DIN2(_30382), .Q(_30416) );
  nnd2s1 _30253_inst ( .DIN1(_30417), .DIN2(_30418), .Q(_30382) );
  nnd2s1 _30254_inst ( .DIN1(_30419), .DIN2(_26662), .Q(_30418) );
  nnd2s1 _30255_inst ( .DIN1(_30420), .DIN2(_30421), .Q(_30419) );
  or2s1 _30256_inst ( .DIN1(_30420), .DIN2(_30421), .Q(_30417) );
  xnr2s1 _30257_inst ( .DIN1(_30386), .DIN2(_30389), .Q(_30381) );
  hi1s1 _30258_inst ( .DIN(_30387), .Q(_30389) );
  hi1s1 _30259_inst ( .DIN(_30422), .Q(_30386) );
  nnd2s1 _30260_inst ( .DIN1(_30423), .DIN2(_30424), .Q(_30412) );
  nnd2s1 _30261_inst ( .DIN1(_30425), .DIN2(_30426), .Q(_30423) );
  nnd2s1 _30262_inst ( .DIN1(_30427), .DIN2(_52988), .Q(_30426) );
  nor2s1 _30263_inst ( .DIN1(_30428), .DIN2(_30429), .Q(_30425) );
  nor2s1 _30264_inst ( .DIN1(_53122), .DIN2(_26571), .Q(_30429) );
  nor2s1 _30265_inst ( .DIN1(_52914), .DIN2(_30430), .Q(_30428) );
  nnd2s1 _30266_inst ( .DIN1(_53122), .DIN2(_26418), .Q(_30430) );
  nor2s1 _30267_inst ( .DIN1(_30431), .DIN2(_30432), .Q(_28650) );
  nnd2s1 _30268_inst ( .DIN1(_30433), .DIN2(_30434), .Q(_30431) );
  nnd2s1 _30269_inst ( .DIN1(_28253), .DIN2(_30435), .Q(
        ______________________________178________) );
  nnd2s1 _30270_inst ( .DIN1(_30436), .DIN2(_30437), .Q(_30435) );
  nnd2s1 _30271_inst ( .DIN1(_30438), .DIN2(______[24]), .Q(_30437) );
  nor2s1 _30272_inst ( .DIN1(_52911), .DIN2(_30439), .Q(_30438) );
  nnd2s1 _30273_inst ( .DIN1(_30440), .DIN2(_30415), .Q(_30436) );
  xor2s1 _30274_inst ( .DIN1(_30421), .DIN2(_30441), .Q(_30440) );
  xor2s1 _30275_inst ( .DIN1(_26662), .DIN2(_30420), .Q(_30441) );
  nnd2s1 _30276_inst ( .DIN1(_30442), .DIN2(_30443), .Q(_30420) );
  nnd2s1 _30277_inst ( .DIN1(_53089), .DIN2(_30444), .Q(_30443) );
  or2s1 _30278_inst ( .DIN1(_30445), .DIN2(_30446), .Q(_30444) );
  nnd2s1 _30279_inst ( .DIN1(_30446), .DIN2(_30445), .Q(_30442) );
  nnd2s1 _30280_inst ( .DIN1(_30422), .DIN2(_30447), .Q(_30421) );
  nnd2s1 _30281_inst ( .DIN1(_30448), .DIN2(_30449), .Q(_30447) );
  nnd2s1 _30282_inst ( .DIN1(_30450), .DIN2(_30451), .Q(_30449) );
  nnd2s1 _30283_inst ( .DIN1(_30452), .DIN2(_30450), .Q(_30422) );
  nor2s1 _30284_inst ( .DIN1(_30453), .DIN2(_30448), .Q(_30452) );
  hi1s1 _30285_inst ( .DIN(_30454), .Q(_30448) );
  nnd2s1 _30286_inst ( .DIN1(_30455), .DIN2(_30456), .Q(
        ______________________________177________) );
  nnd2s1 _30287_inst ( .DIN1(_30457), .DIN2(_29064), .Q(_30456) );
  and2s1 _30288_inst ( .DIN1(_27780), .DIN2(_27779), .Q(_29064) );
  xor2s1 _30289_inst ( .DIN1(_26621), .DIN2(_53452), .Q(_30457) );
  nnd2s1 _30290_inst ( .DIN1(_27782), .DIN2(_30458), .Q(_30455) );
  nnd2s1 _30291_inst ( .DIN1(_30459), .DIN2(_30460), .Q(_30458) );
  nnd2s1 _30292_inst ( .DIN1(_30461), .DIN2(_30415), .Q(_30460) );
  xor2s1 _30293_inst ( .DIN1(_30446), .DIN2(_30462), .Q(_30461) );
  xnr2s1 _30294_inst ( .DIN1(_53089), .DIN2(_30445), .Q(_30462) );
  nnd2s1 _30295_inst ( .DIN1(_30463), .DIN2(_30464), .Q(_30445) );
  nnd2s1 _30296_inst ( .DIN1(_52913), .DIN2(_30465), .Q(_30464) );
  nnd2s1 _30297_inst ( .DIN1(_30466), .DIN2(_30467), .Q(_30465) );
  or2s1 _30298_inst ( .DIN1(_30467), .DIN2(_30466), .Q(_30463) );
  xor2s1 _30299_inst ( .DIN1(_30450), .DIN2(_30453), .Q(_30446) );
  nor2s1 _30300_inst ( .DIN1(_30468), .DIN2(_30469), .Q(_30450) );
  nnd2s1 _30301_inst ( .DIN1(_30424), .DIN2(_26571), .Q(_30459) );
  nnd2s1 _30302_inst ( .DIN1(_30470), .DIN2(_30471), .Q(
        ______________________________176________) );
  nnd2s1 _30303_inst ( .DIN1(_30472), .DIN2(_27546), .Q(_30471) );
  nnd2s1 _30304_inst ( .DIN1(_30473), .DIN2(_27177), .Q(_30472) );
  xnr2s1 _30305_inst ( .DIN1(_52995), .DIN2(_30474), .Q(_30473) );
  nor2s1 _30306_inst ( .DIN1(_53124), .DIN2(_53123), .Q(_30474) );
  nnd2s1 _30307_inst ( .DIN1(_27164), .DIN2(_30475), .Q(_30470) );
  nnd2s1 _30308_inst ( .DIN1(_30476), .DIN2(_30477), .Q(_30475) );
  nnd2s1 _30309_inst ( .DIN1(_30478), .DIN2(_26862), .Q(_30477) );
  nor2s1 _30310_inst ( .DIN1(_30439), .DIN2(_30479), .Q(_30478) );
  xor2s1 _30311_inst ( .DIN1(_26418), .DIN2(_30427), .Q(_30479) );
  nor2s1 _30312_inst ( .DIN1(_52914), .DIN2(_53122), .Q(_30427) );
  nnd2s1 _30313_inst ( .DIN1(_30415), .DIN2(_30480), .Q(_30476) );
  xor2s1 _30314_inst ( .DIN1(_30466), .DIN2(_30481), .Q(_30480) );
  xnr2s1 _30315_inst ( .DIN1(_52913), .DIN2(_30467), .Q(_30481) );
  nnd2s1 _30316_inst ( .DIN1(_30482), .DIN2(_30483), .Q(_30467) );
  nnd2s1 _30317_inst ( .DIN1(_30484), .DIN2(_26354), .Q(_30483) );
  or2s1 _30318_inst ( .DIN1(_30485), .DIN2(_30486), .Q(_30484) );
  nnd2s1 _30319_inst ( .DIN1(_30486), .DIN2(_30485), .Q(_30482) );
  xor2s1 _30320_inst ( .DIN1(_30468), .DIN2(_30469), .Q(_30466) );
  nnd2s1 _30321_inst ( .DIN1(_30487), .DIN2(_27198), .Q(
        ______________________________175________) );
  nor2s1 _30322_inst ( .DIN1(_30488), .DIN2(_30489), .Q(_30487) );
  nor2s1 _30323_inst ( .DIN1(_27204), .DIN2(_30490), .Q(_30489) );
  nnd2s1 _30324_inst ( .DIN1(_30491), .DIN2(_30492), .Q(_30490) );
  nnd2s1 _30325_inst ( .DIN1(_30493), .DIN2(______[30]), .Q(_30492) );
  nor2s1 _30326_inst ( .DIN1(_30439), .DIN2(_30494), .Q(_30493) );
  xor2s1 _30327_inst ( .DIN1(_30495), .DIN2(_52921), .Q(_30494) );
  nnd2s1 _30328_inst ( .DIN1(_52915), .DIN2(_26395), .Q(_30495) );
  nnd2s1 _30329_inst ( .DIN1(_30496), .DIN2(_30415), .Q(_30491) );
  xor2s1 _30330_inst ( .DIN1(_30497), .DIN2(_30485), .Q(_30496) );
  xnr2s1 _30331_inst ( .DIN1(_26321), .DIN2(_30498), .Q(_30485) );
  nor2s1 _30332_inst ( .DIN1(_30499), .DIN2(_30500), .Q(_30498) );
  hi1s1 _30333_inst ( .DIN(_30468), .Q(_30500) );
  nnd2s1 _30334_inst ( .DIN1(_30501), .DIN2(_30502), .Q(_30468) );
  and2s1 _30335_inst ( .DIN1(_30503), .DIN2(_30504), .Q(_30501) );
  nor2s1 _30336_inst ( .DIN1(_30505), .DIN2(_30503), .Q(_30499) );
  nor2s1 _30337_inst ( .DIN1(_30506), .DIN2(_30507), .Q(_30505) );
  xor2s1 _30338_inst ( .DIN1(_26354), .DIN2(_30486), .Q(_30497) );
  and2s1 _30339_inst ( .DIN1(_30508), .DIN2(_30509), .Q(_30486) );
  nnd2s1 _30340_inst ( .DIN1(_30510), .DIN2(_26548), .Q(_30509) );
  or2s1 _30341_inst ( .DIN1(_30511), .DIN2(_30512), .Q(_30510) );
  nnd2s1 _30342_inst ( .DIN1(_30512), .DIN2(_30511), .Q(_30508) );
  nor2s1 _30343_inst ( .DIN1(_53183), .DIN2(_27201), .Q(_30488) );
  nnd2s1 _30344_inst ( .DIN1(_30513), .DIN2(_28073), .Q(
        ______________________________174________) );
  nor2s1 _30345_inst ( .DIN1(_30514), .DIN2(_30515), .Q(_30513) );
  nor2s1 _30346_inst ( .DIN1(_27235), .DIN2(_30516), .Q(_30515) );
  nnd2s1 _30347_inst ( .DIN1(_30517), .DIN2(_30518), .Q(_30516) );
  nnd2s1 _30348_inst ( .DIN1(_30519), .DIN2(_30424), .Q(_30518) );
  xor2s1 _30349_inst ( .DIN1(_53182), .DIN2(_26395), .Q(_30519) );
  nnd2s1 _30350_inst ( .DIN1(_30520), .DIN2(_30415), .Q(_30517) );
  and2s1 _30351_inst ( .DIN1(_30521), .DIN2(_30439), .Q(_30415) );
  hi1s1 _30352_inst ( .DIN(_30424), .Q(_30439) );
  nnd2s1 _30353_inst ( .DIN1(_30522), .DIN2(_30523), .Q(_30424) );
  nor2s1 _30354_inst ( .DIN1(_30524), .DIN2(_30375), .Q(_30523) );
  nor2s1 _30355_inst ( .DIN1(_30369), .DIN2(_30525), .Q(_30522) );
  nor2s1 _30356_inst ( .DIN1(_30374), .DIN2(_30526), .Q(_30521) );
  xnr2s1 _30357_inst ( .DIN1(_30512), .DIN2(_30527), .Q(_30520) );
  xor2s1 _30358_inst ( .DIN1(_26548), .DIN2(_30511), .Q(_30527) );
  nnd2s1 _30359_inst ( .DIN1(_30528), .DIN2(_30529), .Q(_30511) );
  nnd2s1 _30360_inst ( .DIN1(_52942), .DIN2(_30530), .Q(_30529) );
  or2s1 _30361_inst ( .DIN1(_30531), .DIN2(_30532), .Q(_30530) );
  nnd2s1 _30362_inst ( .DIN1(_30532), .DIN2(_30531), .Q(_30528) );
  xor2s1 _30363_inst ( .DIN1(_30507), .DIN2(_30504), .Q(_30512) );
  nor2s1 _30364_inst ( .DIN1(_27325), .DIN2(_30533), .Q(_30514) );
  and2s1 _30365_inst ( .DIN1(______[26]), .DIN2(_53432), .Q(_30533) );
  nnd2s1 _30366_inst ( .DIN1(_30534), .DIN2(_30535), .Q(
        ______________________________173________) );
  nor2s1 _30367_inst ( .DIN1(_30536), .DIN2(_30537), .Q(_30535) );
  nor2s1 _30368_inst ( .DIN1(_30538), .DIN2(_30539), .Q(_30537) );
  xnr2s1 _30369_inst ( .DIN1(_30532), .DIN2(_30540), .Q(_30539) );
  xnr2s1 _30370_inst ( .DIN1(_52942), .DIN2(_30531), .Q(_30540) );
  nnd2s1 _30371_inst ( .DIN1(_30541), .DIN2(_30542), .Q(_30531) );
  nnd2s1 _30372_inst ( .DIN1(_52948), .DIN2(_30543), .Q(_30542) );
  or2s1 _30373_inst ( .DIN1(_30544), .DIN2(_30545), .Q(_30543) );
  nnd2s1 _30374_inst ( .DIN1(_30545), .DIN2(_30544), .Q(_30541) );
  nnd2s1 _30375_inst ( .DIN1(_30507), .DIN2(_30546), .Q(_30532) );
  nnd2s1 _30376_inst ( .DIN1(_30547), .DIN2(_30548), .Q(_30546) );
  hi1s1 _30377_inst ( .DIN(_30502), .Q(_30507) );
  nor2s1 _30378_inst ( .DIN1(_30548), .DIN2(_30547), .Q(_30502) );
  hi1s1 _30379_inst ( .DIN(_30549), .Q(_30547) );
  nor2s1 _30380_inst ( .DIN1(_30550), .DIN2(_30551), .Q(_30534) );
  nor2s1 _30381_inst ( .DIN1(_26672), .DIN2(_30552), .Q(_30551) );
  nor2s1 _30382_inst ( .DIN1(_28957), .DIN2(_30553), .Q(_30550) );
  nor2s1 _30383_inst ( .DIN1(_30554), .DIN2(_27393), .Q(_30553) );
  xor2s1 _30384_inst ( .DIN1(_30555), .DIN2(_30556), .Q(_30554) );
  xor2s1 _30385_inst ( .DIN1(_52921), .DIN2(_52926), .Q(_30556) );
  nnd2s1 _30386_inst ( .DIN1(_52921), .DIN2(_52831), .Q(_30555) );
  nnd2s1 _30387_inst ( .DIN1(_30557), .DIN2(_30558), .Q(
        ______________________________172________) );
  hi1s1 _30388_inst ( .DIN(_30536), .Q(_30558) );
  nor2s1 _30389_inst ( .DIN1(_30559), .DIN2(_30560), .Q(_30557) );
  nor2s1 _30390_inst ( .DIN1(_28954), .DIN2(_30561), .Q(_30560) );
  nnd2s1 _30391_inst ( .DIN1(_30562), .DIN2(_30563), .Q(_30561) );
  nnd2s1 _30392_inst ( .DIN1(_30564), .DIN2(_30565), .Q(_30563) );
  xor2s1 _30393_inst ( .DIN1(_26395), .DIN2(_52915), .Q(_30565) );
  nor2s1 _30394_inst ( .DIN1(_27393), .DIN2(_30236), .Q(_30564) );
  nnd2s1 _30395_inst ( .DIN1(_30566), .DIN2(_30567), .Q(_30562) );
  xor2s1 _30396_inst ( .DIN1(_30545), .DIN2(_30568), .Q(_30566) );
  xnr2s1 _30397_inst ( .DIN1(_52948), .DIN2(_30544), .Q(_30568) );
  nnd2s1 _30398_inst ( .DIN1(_30569), .DIN2(_30570), .Q(_30544) );
  nnd2s1 _30399_inst ( .DIN1(_52945), .DIN2(_30571), .Q(_30570) );
  nnd2s1 _30400_inst ( .DIN1(_30572), .DIN2(_30573), .Q(_30571) );
  or2s1 _30401_inst ( .DIN1(_30573), .DIN2(_30572), .Q(_30569) );
  nnd2s1 _30402_inst ( .DIN1(_30548), .DIN2(_30574), .Q(_30545) );
  nnd2s1 _30403_inst ( .DIN1(_30575), .DIN2(_30576), .Q(_30574) );
  or2s1 _30404_inst ( .DIN1(_30576), .DIN2(_30575), .Q(_30548) );
  or2s1 _30405_inst ( .DIN1(_30577), .DIN2(_30578), .Q(_30576) );
  nor2s1 _30406_inst ( .DIN1(_52916), .DIN2(_28957), .Q(_30559) );
  nnd2s1 _30407_inst ( .DIN1(_30579), .DIN2(_30580), .Q(
        ______________________________171________) );
  nor2s1 _30408_inst ( .DIN1(_30581), .DIN2(_30582), .Q(_30579) );
  nor2s1 _30409_inst ( .DIN1(_27967), .DIN2(_30583), .Q(_30582) );
  nnd2s1 _30410_inst ( .DIN1(_30584), .DIN2(_30585), .Q(_30583) );
  nnd2s1 _30411_inst ( .DIN1(_30567), .DIN2(_30586), .Q(_30585) );
  xor2s1 _30412_inst ( .DIN1(_30572), .DIN2(_30587), .Q(_30586) );
  xnr2s1 _30413_inst ( .DIN1(_52945), .DIN2(_30573), .Q(_30587) );
  nnd2s1 _30414_inst ( .DIN1(_30588), .DIN2(_30589), .Q(_30573) );
  nnd2s1 _30415_inst ( .DIN1(_53292), .DIN2(_30590), .Q(_30589) );
  nnd2s1 _30416_inst ( .DIN1(_30591), .DIN2(_30592), .Q(_30590) );
  or2s1 _30417_inst ( .DIN1(_30591), .DIN2(_30592), .Q(_30588) );
  xnr2s1 _30418_inst ( .DIN1(_30577), .DIN2(_30593), .Q(_30572) );
  nnd2s1 _30419_inst ( .DIN1(_30594), .DIN2(_30595), .Q(_30584) );
  xor2s1 _30420_inst ( .DIN1(_26614), .DIN2(_52964), .Q(_30594) );
  nor2s1 _30421_inst ( .DIN1(_28755), .DIN2(_30596), .Q(_30581) );
  nor2s1 _30422_inst ( .DIN1(_30597), .DIN2(_27448), .Q(_30596) );
  xor2s1 _30423_inst ( .DIN1(_30598), .DIN2(_30599), .Q(_30597) );
  xor2s1 _30424_inst ( .DIN1(_53136), .DIN2(_53175), .Q(_30599) );
  nnd2s1 _30425_inst ( .DIN1(_30600), .DIN2(_30601), .Q(
        ______________________________170________) );
  nor2s1 _30426_inst ( .DIN1(_30602), .DIN2(_30603), .Q(_30600) );
  nor2s1 _30427_inst ( .DIN1(_30604), .DIN2(_27392), .Q(_30603) );
  nor2s1 _30428_inst ( .DIN1(_30605), .DIN2(_30606), .Q(_30604) );
  nor2s1 _30429_inst ( .DIN1(_30607), .DIN2(_30608), .Q(_30606) );
  xnr2s1 _30430_inst ( .DIN1(_30609), .DIN2(_30592), .Q(_30607) );
  nnd2s1 _30431_inst ( .DIN1(_30610), .DIN2(_30611), .Q(_30592) );
  nnd2s1 _30432_inst ( .DIN1(_52939), .DIN2(_30612), .Q(_30611) );
  or2s1 _30433_inst ( .DIN1(_30613), .DIN2(_30614), .Q(_30612) );
  nnd2s1 _30434_inst ( .DIN1(_30614), .DIN2(_30613), .Q(_30610) );
  xor2s1 _30435_inst ( .DIN1(_30591), .DIN2(_53292), .Q(_30609) );
  nnd2s1 _30436_inst ( .DIN1(_30577), .DIN2(_30615), .Q(_30591) );
  nnd2s1 _30437_inst ( .DIN1(_30616), .DIN2(_30617), .Q(_30615) );
  nnd2s1 _30438_inst ( .DIN1(_30618), .DIN2(_30619), .Q(_30617) );
  nnd2s1 _30439_inst ( .DIN1(_30620), .DIN2(_30618), .Q(_30577) );
  nor2s1 _30440_inst ( .DIN1(_30621), .DIN2(_30616), .Q(_30620) );
  hi1s1 _30441_inst ( .DIN(_30622), .Q(_30616) );
  nor2s1 _30442_inst ( .DIN1(_30236), .DIN2(_30623), .Q(_30605) );
  nnd2s1 _30443_inst ( .DIN1(______[12]), .DIN2(_30624), .Q(_30623) );
  xnr2s1 _30444_inst ( .DIN1(_52920), .DIN2(_30625), .Q(_30624) );
  nnd2s1 _30445_inst ( .DIN1(_52964), .DIN2(_52917), .Q(_30625) );
  nor2s1 _30446_inst ( .DIN1(_27397), .DIN2(_30626), .Q(_30602) );
  nor2s1 _30447_inst ( .DIN1(_30627), .DIN2(_30628), .Q(_30626) );
  nor2s1 _30448_inst ( .DIN1(_53382), .DIN2(_26228), .Q(_30627) );
  nnd2s1 _30449_inst ( .DIN1(_30629), .DIN2(_30630), .Q(
        ______________________________16________) );
  nnd2s1 _30450_inst ( .DIN1(_28932), .DIN2(_30631), .Q(_30630) );
  nnd2s1 _30451_inst ( .DIN1(_30632), .DIN2(_30083), .Q(_30631) );
  hi1s1 _30452_inst ( .DIN(_30065), .Q(_30083) );
  nor2s1 _30453_inst ( .DIN1(_30162), .DIN2(_30085), .Q(_30065) );
  nor2s1 _30454_inst ( .DIN1(_30633), .DIN2(_30634), .Q(_30632) );
  nor2s1 _30455_inst ( .DIN1(_30085), .DIN2(_30635), .Q(_30634) );
  nor2s1 _30456_inst ( .DIN1(_30636), .DIN2(_27774), .Q(_30635) );
  xor2s1 _30457_inst ( .DIN1(_30637), .DIN2(_30638), .Q(_30636) );
  xor2s1 _30458_inst ( .DIN1(_53016), .DIN2(_53469), .Q(_30638) );
  nnd2s1 _30459_inst ( .DIN1(_53192), .DIN2(_26475), .Q(_30637) );
  nor2s1 _30460_inst ( .DIN1(_30066), .DIN2(_26693), .Q(_30633) );
  hi1s1 _30461_inst ( .DIN(_29021), .Q(_28932) );
  nnd2s1 _30462_inst ( .DIN1(_30639), .DIN2(_30640), .Q(_30629) );
  xor2s1 _30463_inst ( .DIN1(_52893), .DIN2(_52918), .Q(_30639) );
  nnd2s1 _30464_inst ( .DIN1(_30641), .DIN2(_27983), .Q(
        ______________________________169________) );
  nor2s1 _30465_inst ( .DIN1(_30642), .DIN2(_30643), .Q(_30641) );
  nor2s1 _30466_inst ( .DIN1(_27994), .DIN2(_30644), .Q(_30643) );
  nor2s1 _30467_inst ( .DIN1(_26774), .DIN2(_30645), .Q(_30644) );
  xor2s1 _30468_inst ( .DIN1(_30646), .DIN2(_30647), .Q(_30645) );
  xor2s1 _30469_inst ( .DIN1(_52968), .DIN2(_53336), .Q(_30647) );
  nor2s1 _30470_inst ( .DIN1(_52964), .DIN2(_26689), .Q(_30646) );
  nor2s1 _30471_inst ( .DIN1(_30648), .DIN2(_27500), .Q(_30642) );
  nor2s1 _30472_inst ( .DIN1(_30649), .DIN2(_30650), .Q(_30648) );
  and2s1 _30473_inst ( .DIN1(_52917), .DIN2(_30595), .Q(_30650) );
  nor2s1 _30474_inst ( .DIN1(_30236), .DIN2(_26771), .Q(_30595) );
  nor2s1 _30475_inst ( .DIN1(_30651), .DIN2(_30608), .Q(_30649) );
  xnr2s1 _30476_inst ( .DIN1(_30614), .DIN2(_30652), .Q(_30651) );
  xnr2s1 _30477_inst ( .DIN1(_52939), .DIN2(_30613), .Q(_30652) );
  nnd2s1 _30478_inst ( .DIN1(_30653), .DIN2(_30654), .Q(_30613) );
  nnd2s1 _30479_inst ( .DIN1(_53386), .DIN2(_30655), .Q(_30654) );
  nnd2s1 _30480_inst ( .DIN1(_30656), .DIN2(_30657), .Q(_30655) );
  or2s1 _30481_inst ( .DIN1(_30657), .DIN2(_30656), .Q(_30653) );
  xor2s1 _30482_inst ( .DIN1(_30618), .DIN2(_30621), .Q(_30614) );
  hi1s1 _30483_inst ( .DIN(_30619), .Q(_30621) );
  nor2s1 _30484_inst ( .DIN1(_30658), .DIN2(_30659), .Q(_30618) );
  nnd2s1 _30485_inst ( .DIN1(_30660), .DIN2(_30661), .Q(
        ______________________________168________) );
  nor2s1 _30486_inst ( .DIN1(_30536), .DIN2(_30662), .Q(_30661) );
  nor2s1 _30487_inst ( .DIN1(_30663), .DIN2(_30552), .Q(_30662) );
  nnd2s1 _30488_inst ( .DIN1(_30664), .DIN2(_30526), .Q(_30552) );
  nor2s1 _30489_inst ( .DIN1(_26853), .DIN2(_28954), .Q(_30664) );
  xnr2s1 _30490_inst ( .DIN1(_52920), .DIN2(_52964), .Q(_30663) );
  nor2s1 _30491_inst ( .DIN1(_29939), .DIN2(_28957), .Q(_30536) );
  nor2s1 _30492_inst ( .DIN1(_30665), .DIN2(_30666), .Q(_30660) );
  nor2s1 _30493_inst ( .DIN1(_52921), .DIN2(_28957), .Q(_30666) );
  nor2s1 _30494_inst ( .DIN1(_30538), .DIN2(_30667), .Q(_30665) );
  xnr2s1 _30495_inst ( .DIN1(_30656), .DIN2(_30668), .Q(_30667) );
  xor2s1 _30496_inst ( .DIN1(_26591), .DIN2(_30657), .Q(_30668) );
  nnd2s1 _30497_inst ( .DIN1(_30669), .DIN2(_30670), .Q(_30657) );
  nnd2s1 _30498_inst ( .DIN1(_53020), .DIN2(_30671), .Q(_30670) );
  nnd2s1 _30499_inst ( .DIN1(_30672), .DIN2(_30673), .Q(_30671) );
  xor2s1 _30500_inst ( .DIN1(_30674), .DIN2(_30675), .Q(_30669) );
  or2s1 _30501_inst ( .DIN1(_30672), .DIN2(_30673), .Q(_30675) );
  xor2s1 _30502_inst ( .DIN1(_30659), .DIN2(_30658), .Q(_30656) );
  nnd2s1 _30503_inst ( .DIN1(_30567), .DIN2(_28957), .Q(_30538) );
  hi1s1 _30504_inst ( .DIN(_30608), .Q(_30567) );
  nnd2s1 _30505_inst ( .DIN1(_30676), .DIN2(_30677), .Q(_30608) );
  nnd2s1 _30506_inst ( .DIN1(_30678), .DIN2(_30679), .Q(
        ______________________________167________) );
  nnd2s1 _30507_inst ( .DIN1(_30680), .DIN2(_52902), .Q(_30679) );
  nor2s1 _30508_inst ( .DIN1(_26987), .DIN2(_27182), .Q(_30680) );
  nor2s1 _30509_inst ( .DIN1(_30681), .DIN2(_30682), .Q(_30678) );
  nor2s1 _30510_inst ( .DIN1(_30683), .DIN2(_30684), .Q(_30682) );
  nnd2s1 _30511_inst ( .DIN1(_30685), .DIN2(_27183), .Q(_30684) );
  nor2s1 _30512_inst ( .DIN1(_30686), .DIN2(_30687), .Q(_30685) );
  xor2s1 _30513_inst ( .DIN1(_30688), .DIN2(_30689), .Q(_30687) );
  xor2s1 _30514_inst ( .DIN1(_52924), .DIN2(_52926), .Q(_30689) );
  and2s1 _30515_inst ( .DIN1(_26581), .DIN2(_53273), .Q(_30688) );
  nor2s1 _30516_inst ( .DIN1(_30690), .DIN2(_30691), .Q(_30681) );
  nnd2s1 _30517_inst ( .DIN1(_27183), .DIN2(_30692), .Q(_30691) );
  xnr2s1 _30518_inst ( .DIN1(_30673), .DIN2(_30693), .Q(_30692) );
  xnr2s1 _30519_inst ( .DIN1(_53020), .DIN2(_30672), .Q(_30693) );
  nnd2s1 _30520_inst ( .DIN1(_30694), .DIN2(_30695), .Q(_30672) );
  nnd2s1 _30521_inst ( .DIN1(_52947), .DIN2(_30696), .Q(_30695) );
  or2s1 _30522_inst ( .DIN1(_30697), .DIN2(_30698), .Q(_30696) );
  nnd2s1 _30523_inst ( .DIN1(_30698), .DIN2(_30697), .Q(_30694) );
  nnd2s1 _30524_inst ( .DIN1(_30658), .DIN2(_30699), .Q(_30673) );
  nnd2s1 _30525_inst ( .DIN1(_30700), .DIN2(_30701), .Q(_30699) );
  or2s1 _30526_inst ( .DIN1(_30701), .DIN2(_30700), .Q(_30658) );
  nnd2s1 _30527_inst ( .DIN1(_30702), .DIN2(_30703), .Q(
        ______________________________166________) );
  nnd2s1 _30528_inst ( .DIN1(_30704), .DIN2(_30705), .Q(_30703) );
  nnd2s1 _30529_inst ( .DIN1(_30706), .DIN2(_53273), .Q(_30705) );
  nor2s1 _30530_inst ( .DIN1(_30686), .DIN2(_26771), .Q(_30706) );
  nor2s1 _30531_inst ( .DIN1(_30707), .DIN2(_30708), .Q(_30702) );
  nor2s1 _30532_inst ( .DIN1(_30709), .DIN2(_30710), .Q(_30708) );
  xor2s1 _30533_inst ( .DIN1(_30698), .DIN2(_30711), .Q(_30709) );
  xnr2s1 _30534_inst ( .DIN1(_52947), .DIN2(_30697), .Q(_30711) );
  nnd2s1 _30535_inst ( .DIN1(_30701), .DIN2(_30712), .Q(_30697) );
  nnd2s1 _30536_inst ( .DIN1(_30713), .DIN2(_30714), .Q(_30712) );
  or2s1 _30537_inst ( .DIN1(_30714), .DIN2(_30713), .Q(_30701) );
  nnd2s1 _30538_inst ( .DIN1(_30715), .DIN2(_30716), .Q(_30714) );
  nnd2s1 _30539_inst ( .DIN1(_30717), .DIN2(_30718), .Q(_30698) );
  nnd2s1 _30540_inst ( .DIN1(_52922), .DIN2(_30719), .Q(_30718) );
  nnd2s1 _30541_inst ( .DIN1(_30720), .DIN2(_30721), .Q(_30719) );
  or2s1 _30542_inst ( .DIN1(_30721), .DIN2(_30720), .Q(_30717) );
  nor2s1 _30543_inst ( .DIN1(_30722), .DIN2(_30723), .Q(_30707) );
  xor2s1 _30544_inst ( .DIN1(_30724), .DIN2(_52831), .Q(_30722) );
  nnd2s1 _30545_inst ( .DIN1(_52921), .DIN2(_52926), .Q(_30724) );
  nnd2s1 _30546_inst ( .DIN1(_30725), .DIN2(_30726), .Q(
        ______________________________165________) );
  nnd2s1 _30547_inst ( .DIN1(_30704), .DIN2(_30727), .Q(_30726) );
  nor2s1 _30548_inst ( .DIN1(_30728), .DIN2(_30729), .Q(_30725) );
  nor2s1 _30549_inst ( .DIN1(_30710), .DIN2(_30730), .Q(_30729) );
  xor2s1 _30550_inst ( .DIN1(_30720), .DIN2(_30731), .Q(_30730) );
  xnr2s1 _30551_inst ( .DIN1(_52922), .DIN2(_30721), .Q(_30731) );
  nnd2s1 _30552_inst ( .DIN1(_30732), .DIN2(_30733), .Q(_30721) );
  nnd2s1 _30553_inst ( .DIN1(_30734), .DIN2(_26532), .Q(_30733) );
  nnd2s1 _30554_inst ( .DIN1(_30735), .DIN2(_30736), .Q(_30734) );
  or2s1 _30555_inst ( .DIN1(_30735), .DIN2(_30736), .Q(_30732) );
  xor2s1 _30556_inst ( .DIN1(_30737), .DIN2(_30738), .Q(_30720) );
  nor2s1 _30557_inst ( .DIN1(_30723), .DIN2(_30739), .Q(_30728) );
  nnd2s1 _30558_inst ( .DIN1(_26857), .DIN2(_30740), .Q(_30739) );
  xor2s1 _30559_inst ( .DIN1(_52925), .DIN2(_52956), .Q(_30740) );
  nnd2s1 _30560_inst ( .DIN1(_30741), .DIN2(_30742), .Q(
        ______________________________164________) );
  nnd2s1 _30561_inst ( .DIN1(_30743), .DIN2(_30744), .Q(_30742) );
  hi1s1 _30562_inst ( .DIN(_30710), .Q(_30744) );
  nnd2s1 _30563_inst ( .DIN1(_30683), .DIN2(_28957), .Q(_30710) );
  xor2s1 _30564_inst ( .DIN1(_30736), .DIN2(_30745), .Q(_30743) );
  xor2s1 _30565_inst ( .DIN1(_26532), .DIN2(_30735), .Q(_30745) );
  nnd2s1 _30566_inst ( .DIN1(_30746), .DIN2(_30747), .Q(_30735) );
  nnd2s1 _30567_inst ( .DIN1(_30748), .DIN2(_26392), .Q(_30747) );
  or2s1 _30568_inst ( .DIN1(_30749), .DIN2(_30750), .Q(_30748) );
  nnd2s1 _30569_inst ( .DIN1(_30750), .DIN2(_30749), .Q(_30746) );
  nnd2s1 _30570_inst ( .DIN1(_30737), .DIN2(_30751), .Q(_30736) );
  nnd2s1 _30571_inst ( .DIN1(_30752), .DIN2(_30753), .Q(_30751) );
  hi1s1 _30572_inst ( .DIN(_30715), .Q(_30737) );
  nor2s1 _30573_inst ( .DIN1(_30753), .DIN2(_30752), .Q(_30715) );
  hi1s1 _30574_inst ( .DIN(_30754), .Q(_30752) );
  nnd2s1 _30575_inst ( .DIN1(_30755), .DIN2(______[22]), .Q(_30741) );
  nor2s1 _30576_inst ( .DIN1(_30756), .DIN2(_30757), .Q(_30755) );
  nor2s1 _30577_inst ( .DIN1(_26581), .DIN2(_30758), .Q(_30757) );
  nnd2s1 _30578_inst ( .DIN1(_30759), .DIN2(_30760), .Q(_30758) );
  nnd2s1 _30579_inst ( .DIN1(_30761), .DIN2(_30762), .Q(_30760) );
  nnd2s1 _30580_inst ( .DIN1(_52924), .DIN2(_52925), .Q(_30762) );
  nnd2s1 _30581_inst ( .DIN1(_30763), .DIN2(_30704), .Q(_30759) );
  hi1s1 _30582_inst ( .DIN(_30727), .Q(_30763) );
  nnd2s1 _30583_inst ( .DIN1(_26527), .DIN2(_30376), .Q(_30727) );
  nor2s1 _30584_inst ( .DIN1(_52923), .DIN2(_30764), .Q(_30756) );
  nnd2s1 _30585_inst ( .DIN1(_30765), .DIN2(_30766), .Q(_30764) );
  nnd2s1 _30586_inst ( .DIN1(_30767), .DIN2(_30704), .Q(_30766) );
  nor2s1 _30587_inst ( .DIN1(_28954), .DIN2(_30683), .Q(_30704) );
  nor2s1 _30588_inst ( .DIN1(_30686), .DIN2(_26527), .Q(_30767) );
  nnd2s1 _30589_inst ( .DIN1(_30768), .DIN2(_30761), .Q(_30765) );
  hi1s1 _30590_inst ( .DIN(_30723), .Q(_30761) );
  nnd2s1 _30591_inst ( .DIN1(_29939), .DIN2(_28954), .Q(_30723) );
  nnd2s1 _30592_inst ( .DIN1(_30769), .DIN2(_30770), .Q(_29939) );
  nor2s1 _30593_inst ( .DIN1(_30771), .DIN2(_30772), .Q(_30770) );
  nor2s1 _30594_inst ( .DIN1(_30640), .DIN2(_29938), .Q(_30769) );
  nor2s1 _30595_inst ( .DIN1(_26296), .DIN2(_26688), .Q(_30768) );
  nnd2s1 _30596_inst ( .DIN1(_30773), .DIN2(_30774), .Q(
        ______________________________163________) );
  nor2s1 _30597_inst ( .DIN1(_30775), .DIN2(_30776), .Q(_30773) );
  nor2s1 _30598_inst ( .DIN1(_30777), .DIN2(_30778), .Q(_30776) );
  nor2s1 _30599_inst ( .DIN1(_30779), .DIN2(_30780), .Q(_30778) );
  nor2s1 _30600_inst ( .DIN1(_30683), .DIN2(_30781), .Q(_30780) );
  nnd2s1 _30601_inst ( .DIN1(_30782), .DIN2(_28195), .Q(_30781) );
  nor2s1 _30602_inst ( .DIN1(_30686), .DIN2(_30783), .Q(_30782) );
  xor2s1 _30603_inst ( .DIN1(_29518), .DIN2(_30784), .Q(_30783) );
  nnd2s1 _30604_inst ( .DIN1(______[28]), .DIN2(_30785), .Q(_30784) );
  xor2s1 _30605_inst ( .DIN1(_53058), .DIN2(_29127), .Q(_30785) );
  hi1s1 _30606_inst ( .DIN(_30376), .Q(_30686) );
  nor2s1 _30607_inst ( .DIN1(_30690), .DIN2(_30786), .Q(_30779) );
  nnd2s1 _30608_inst ( .DIN1(_30787), .DIN2(_30788), .Q(_30786) );
  xor2s1 _30609_inst ( .DIN1(_30789), .DIN2(_30790), .Q(_30788) );
  xor2s1 _30610_inst ( .DIN1(_30749), .DIN2(_30750), .Q(_30790) );
  nnd2s1 _30611_inst ( .DIN1(_30753), .DIN2(_30791), .Q(_30750) );
  nnd2s1 _30612_inst ( .DIN1(_30792), .DIN2(_30793), .Q(_30791) );
  or2s1 _30613_inst ( .DIN1(_30793), .DIN2(_30792), .Q(_30753) );
  hi1s1 _30614_inst ( .DIN(_30794), .Q(_30792) );
  nnd2s1 _30615_inst ( .DIN1(_30795), .DIN2(_30796), .Q(_30749) );
  nnd2s1 _30616_inst ( .DIN1(_52952), .DIN2(_30797), .Q(_30796) );
  or2s1 _30617_inst ( .DIN1(_30798), .DIN2(_30799), .Q(_30797) );
  nnd2s1 _30618_inst ( .DIN1(_30799), .DIN2(_30798), .Q(_30795) );
  xor2s1 _30619_inst ( .DIN1(_26392), .DIN2(_28195), .Q(_30789) );
  nor2s1 _30620_inst ( .DIN1(_27227), .DIN2(_30800), .Q(_30775) );
  xor2s1 _30621_inst ( .DIN1(_53190), .DIN2(_53237), .Q(_30800) );
  nnd2s1 _30622_inst ( .DIN1(_30801), .DIN2(_30802), .Q(
        ______________________________162________) );
  nnd2s1 _30623_inst ( .DIN1(_30803), .DIN2(_28670), .Q(_30802) );
  nnd2s1 _30624_inst ( .DIN1(_30804), .DIN2(_28672), .Q(_30803) );
  xor2s1 _30625_inst ( .DIN1(_53062), .DIN2(_26622), .Q(_30804) );
  nor2s1 _30626_inst ( .DIN1(_30805), .DIN2(_30806), .Q(_30801) );
  nor2s1 _30627_inst ( .DIN1(_28683), .DIN2(_30807), .Q(_30806) );
  xor2s1 _30628_inst ( .DIN1(_52953), .DIN2(_53464), .Q(_30807) );
  nnd2s1 _30629_inst ( .DIN1(_29139), .DIN2(_28223), .Q(_28683) );
  nor2s1 _30630_inst ( .DIN1(_28677), .DIN2(_30808), .Q(_30805) );
  xor2s1 _30631_inst ( .DIN1(_30799), .DIN2(_30809), .Q(_30808) );
  xor2s1 _30632_inst ( .DIN1(_30798), .DIN2(_52952), .Q(_30809) );
  nnd2s1 _30633_inst ( .DIN1(_30793), .DIN2(_30810), .Q(_30799) );
  nnd2s1 _30634_inst ( .DIN1(_30811), .DIN2(_30812), .Q(_30810) );
  nnd2s1 _30635_inst ( .DIN1(_30813), .DIN2(_30814), .Q(_30812) );
  nnd2s1 _30636_inst ( .DIN1(_30815), .DIN2(_30813), .Q(_30793) );
  and2s1 _30637_inst ( .DIN1(_30816), .DIN2(_30814), .Q(_30815) );
  nnd2s1 _30638_inst ( .DIN1(_29139), .DIN2(_30099), .Q(_28677) );
  hi1s1 _30639_inst ( .DIN(_28133), .Q(_30099) );
  nnd2s1 _30640_inst ( .DIN1(_30817), .DIN2(_30818), .Q(_28133) );
  nor2s1 _30641_inst ( .DIN1(_29969), .DIN2(_28110), .Q(_30818) );
  nor2s1 _30642_inst ( .DIN1(_28177), .DIN2(_30053), .Q(_30817) );
  nnd2s1 _30643_inst ( .DIN1(_30819), .DIN2(_30820), .Q(_30053) );
  nor2s1 _30644_inst ( .DIN1(_28116), .DIN2(_30821), .Q(_30819) );
  nnd2s1 _30645_inst ( .DIN1(_30822), .DIN2(_30823), .Q(
        ______________________________161________) );
  nnd2s1 _30646_inst ( .DIN1(_30824), .DIN2(_29139), .Q(_30823) );
  nor2s1 _30647_inst ( .DIN1(_30825), .DIN2(_30826), .Q(_30824) );
  nor2s1 _30648_inst ( .DIN1(_30683), .DIN2(_30827), .Q(_30826) );
  nnd2s1 _30649_inst ( .DIN1(_30828), .DIN2(_30376), .Q(_30827) );
  nnd2s1 _30650_inst ( .DIN1(_30829), .DIN2(_30830), .Q(_30376) );
  nor2s1 _30651_inst ( .DIN1(_30831), .DIN2(_30832), .Q(_30830) );
  nor2s1 _30652_inst ( .DIN1(_30526), .DIN2(_30368), .Q(_30829) );
  nnd2s1 _30653_inst ( .DIN1(_30833), .DIN2(_30834), .Q(_30368) );
  xnr2s1 _30654_inst ( .DIN1(_53238), .DIN2(_29127), .Q(_30828) );
  and2s1 _30655_inst ( .DIN1(_53126), .DIN2(_26296), .Q(_29127) );
  nor2s1 _30656_inst ( .DIN1(_30690), .DIN2(_30835), .Q(_30825) );
  nnd2s1 _30657_inst ( .DIN1(_30836), .DIN2(_30798), .Q(_30835) );
  or2s1 _30658_inst ( .DIN1(_30837), .DIN2(_52951), .Q(_30798) );
  nnd2s1 _30659_inst ( .DIN1(_30837), .DIN2(_52951), .Q(_30836) );
  xnr2s1 _30660_inst ( .DIN1(_30813), .DIN2(_30814), .Q(_30837) );
  and2s1 _30661_inst ( .DIN1(_30838), .DIN2(_30839), .Q(_30813) );
  nor2s1 _30662_inst ( .DIN1(_30840), .DIN2(_30841), .Q(_30839) );
  nor2s1 _30663_inst ( .DIN1(_30842), .DIN2(_30843), .Q(_30838) );
  hi1s1 _30664_inst ( .DIN(_30683), .Q(_30690) );
  xor2s1 _30665_inst ( .DIN1(_30844), .DIN2(_29168), .Q(_30683) );
  nnd2s1 _30666_inst ( .DIN1(_30845), .DIN2(_30846), .Q(_30844) );
  nor2s1 _30667_inst ( .DIN1(_30374), .DIN2(_30847), .Q(_30846) );
  nnd2s1 _30668_inst ( .DIN1(_30848), .DIN2(_30849), .Q(_30847) );
  nor2s1 _30669_inst ( .DIN1(_30524), .DIN2(_30525), .Q(_30845) );
  hi1s1 _30670_inst ( .DIN(_30834), .Q(_30525) );
  nnd2s1 _30671_inst ( .DIN1(_52924), .DIN2(_29137), .Q(_30822) );
  nnd2s1 _30672_inst ( .DIN1(_30850), .DIN2(_30851), .Q(
        ______________________________160________) );
  nnd2s1 _30673_inst ( .DIN1(_30852), .DIN2(_30853), .Q(_30851) );
  nnd2s1 _30674_inst ( .DIN1(_26669), .DIN2(_30854), .Q(_30852) );
  nnd2s1 _30675_inst ( .DIN1(_30855), .DIN2(_30856), .Q(_30850) );
  nor2s1 _30676_inst ( .DIN1(_29060), .DIN2(_30857), .Q(_30855) );
  nnd2s1 _30677_inst ( .DIN1(_30858), .DIN2(_30859), .Q(_30857) );
  or2s1 _30678_inst ( .DIN1(_29078), .DIN2(_52955), .Q(_30859) );
  nnd2s1 _30679_inst ( .DIN1(_30860), .DIN2(_29078), .Q(_30858) );
  xor2s1 _30680_inst ( .DIN1(_30861), .DIN2(_30862), .Q(_30860) );
  nor2s1 _30681_inst ( .DIN1(_52932), .DIN2(_26498), .Q(_30862) );
  xor2s1 _30682_inst ( .DIN1(_26583), .DIN2(_53279), .Q(_30861) );
  nnd2s1 _30683_inst ( .DIN1(_30863), .DIN2(_30864), .Q(
        ______________________________15________) );
  nnd2s1 _30684_inst ( .DIN1(_30865), .DIN2(_53468), .Q(_30864) );
  nor2s1 _30685_inst ( .DIN1(_30866), .DIN2(_28684), .Q(_30865) );
  nnd2s1 _30686_inst ( .DIN1(_30867), .DIN2(_29083), .Q(_30863) );
  nor2s1 _30687_inst ( .DIN1(_30868), .DIN2(_30869), .Q(_30867) );
  nor2s1 _30688_inst ( .DIN1(_30085), .DIN2(_30870), .Q(_30869) );
  and2s1 _30689_inst ( .DIN1(_26475), .DIN2(_30162), .Q(_30870) );
  nnd2s1 _30690_inst ( .DIN1(_30871), .DIN2(_28129), .Q(_30162) );
  and2s1 _30691_inst ( .DIN1(_30872), .DIN2(_28938), .Q(_30871) );
  nor2s1 _30692_inst ( .DIN1(_29997), .DIN2(_29902), .Q(_28938) );
  and2s1 _30693_inst ( .DIN1(_52929), .DIN2(_30085), .Q(_30868) );
  hi1s1 _30694_inst ( .DIN(_30066), .Q(_30085) );
  nnd2s1 _30695_inst ( .DIN1(_30873), .DIN2(_30874), .Q(_30066) );
  nor2s1 _30696_inst ( .DIN1(_29902), .DIN2(_29904), .Q(_30874) );
  hi1s1 _30697_inst ( .DIN(_28114), .Q(_29904) );
  nor2s1 _30698_inst ( .DIN1(_28110), .DIN2(_28223), .Q(_30873) );
  nnd2s1 _30699_inst ( .DIN1(_30872), .DIN2(_30875), .Q(_28110) );
  nnd2s1 _30700_inst ( .DIN1(_30876), .DIN2(_28811), .Q(
        ______________________________159________) );
  nor2s1 _30701_inst ( .DIN1(_30877), .DIN2(_30878), .Q(_30876) );
  nor2s1 _30702_inst ( .DIN1(_28356), .DIN2(_30879), .Q(_30878) );
  xor2s1 _30703_inst ( .DIN1(_53226), .DIN2(_53278), .Q(_30879) );
  nor2s1 _30704_inst ( .DIN1(_30880), .DIN2(_28814), .Q(_30877) );
  nor2s1 _30705_inst ( .DIN1(_29060), .DIN2(_30881), .Q(_30880) );
  nnd2s1 _30706_inst ( .DIN1(_30882), .DIN2(_30883), .Q(_30881) );
  nnd2s1 _30707_inst ( .DIN1(_53181), .DIN2(_29057), .Q(_30883) );
  nnd2s1 _30708_inst ( .DIN1(_29078), .DIN2(_26498), .Q(_30882) );
  hi1s1 _30709_inst ( .DIN(_29070), .Q(_29060) );
  nnd2s1 _30710_inst ( .DIN1(_28727), .DIN2(_29078), .Q(_29070) );
  hi1s1 _30711_inst ( .DIN(_29057), .Q(_29078) );
  nor2s1 _30712_inst ( .DIN1(_30884), .DIN2(_28909), .Q(_29057) );
  nnd2s1 _30713_inst ( .DIN1(_30885), .DIN2(_28951), .Q(
        ______________________________158________) );
  nor2s1 _30714_inst ( .DIN1(_30886), .DIN2(_30887), .Q(_30885) );
  nor2s1 _30715_inst ( .DIN1(_28954), .DIN2(_30888), .Q(_30887) );
  nnd2s1 _30716_inst ( .DIN1(_30889), .DIN2(_30890), .Q(_30888) );
  nor2s1 _30717_inst ( .DIN1(_30891), .DIN2(_30892), .Q(_30889) );
  nor2s1 _30718_inst ( .DIN1(_53279), .DIN2(_28724), .Q(_30892) );
  nor2s1 _30719_inst ( .DIN1(_28705), .DIN2(_26461), .Q(_30891) );
  nor2s1 _30720_inst ( .DIN1(_28957), .DIN2(_30893), .Q(_30886) );
  xor2s1 _30721_inst ( .DIN1(_52933), .DIN2(_53006), .Q(_30893) );
  nnd2s1 _30722_inst ( .DIN1(_30894), .DIN2(_30895), .Q(
        ______________________________157________) );
  nnd2s1 _30723_inst ( .DIN1(_30896), .DIN2(_28069), .Q(_30895) );
  nnd2s1 _30724_inst ( .DIN1(_28123), .DIN2(_30897), .Q(_30896) );
  xor2s1 _30725_inst ( .DIN1(_52930), .DIN2(_52981), .Q(_30897) );
  nor2s1 _30726_inst ( .DIN1(_27365), .DIN2(_30043), .Q(_28123) );
  nnd2s1 _30727_inst ( .DIN1(_30898), .DIN2(_28060), .Q(_30894) );
  nor2s1 _30728_inst ( .DIN1(_30899), .DIN2(_30900), .Q(_30898) );
  nnd2s1 _30729_inst ( .DIN1(_30901), .DIN2(_30902), .Q(_30900) );
  nnd2s1 _30730_inst ( .DIN1(_28724), .DIN2(_26440), .Q(_30902) );
  nnd2s1 _30731_inst ( .DIN1(_30903), .DIN2(_28705), .Q(_30901) );
  nnd2s1 _30732_inst ( .DIN1(_30904), .DIN2(______[14]), .Q(_30903) );
  xor2s1 _30733_inst ( .DIN1(_26472), .DIN2(_52932), .Q(_30904) );
  nnd2s1 _30734_inst ( .DIN1(_30905), .DIN2(_30906), .Q(
        ______________________________156________) );
  nnd2s1 _30735_inst ( .DIN1(_27868), .DIN2(_30907), .Q(_30906) );
  nnd2s1 _30736_inst ( .DIN1(_30908), .DIN2(_30909), .Q(_30907) );
  nor2s1 _30737_inst ( .DIN1(_30910), .DIN2(_30911), .Q(_30909) );
  nor2s1 _30738_inst ( .DIN1(_30912), .DIN2(_30913), .Q(_30911) );
  nor2s1 _30739_inst ( .DIN1(_28724), .DIN2(_30914), .Q(_30913) );
  xor2s1 _30740_inst ( .DIN1(_52934), .DIN2(_26368), .Q(_30914) );
  nor2s1 _30741_inst ( .DIN1(_30360), .DIN2(_30915), .Q(_30910) );
  nnd2s1 _30742_inst ( .DIN1(_30916), .DIN2(_28705), .Q(_30915) );
  xor2s1 _30743_inst ( .DIN1(_52904), .DIN2(_52934), .Q(_30916) );
  nor2s1 _30744_inst ( .DIN1(_30899), .DIN2(_30917), .Q(_30908) );
  nor2s1 _30745_inst ( .DIN1(_28705), .DIN2(_26536), .Q(_30917) );
  hi1s1 _30746_inst ( .DIN(_30890), .Q(_30899) );
  nnd2s1 _30747_inst ( .DIN1(_30918), .DIN2(_27875), .Q(_30905) );
  xor2s1 _30748_inst ( .DIN1(_52931), .DIN2(_29551), .Q(_30918) );
  or2s1 _30749_inst ( .DIN1(_53054), .DIN2(_53074), .Q(_29551) );
  nnd2s1 _30750_inst ( .DIN1(_30919), .DIN2(_30920), .Q(
        ______________________________155________) );
  nnd2s1 _30751_inst ( .DIN1(_30921), .DIN2(_52932), .Q(_30920) );
  nor2s1 _30752_inst ( .DIN1(_27066), .DIN2(_29044), .Q(_30921) );
  nnd2s1 _30753_inst ( .DIN1(_28954), .DIN2(_30922), .Q(_29044) );
  nnd2s1 _30754_inst ( .DIN1(_30923), .DIN2(_30924), .Q(_30922) );
  nor2s1 _30755_inst ( .DIN1(_30030), .DIN2(_30925), .Q(_30924) );
  nnd2s1 _30756_inst ( .DIN1(_28957), .DIN2(_30926), .Q(_30919) );
  nnd2s1 _30757_inst ( .DIN1(_30927), .DIN2(_30928), .Q(_30926) );
  nor2s1 _30758_inst ( .DIN1(_30929), .DIN2(_30930), .Q(_30928) );
  nor2s1 _30759_inst ( .DIN1(_28724), .DIN2(_30931), .Q(_30930) );
  nor2s1 _30760_inst ( .DIN1(_30932), .DIN2(_27082), .Q(_30931) );
  nor2s1 _30761_inst ( .DIN1(_53019), .DIN2(_26250), .Q(_30932) );
  and2s1 _30762_inst ( .DIN1(_28724), .DIN2(_52961), .Q(_30929) );
  nor2s1 _30763_inst ( .DIN1(_30933), .DIN2(_30934), .Q(_30927) );
  nor2s1 _30764_inst ( .DIN1(_52933), .DIN2(_30935), .Q(_30933) );
  nnd2s1 _30765_inst ( .DIN1(_30936), .DIN2(_28951), .Q(
        ______________________________154________) );
  nnd2s1 _30766_inst ( .DIN1(_30923), .DIN2(_30937), .Q(_28951) );
  nor2s1 _30767_inst ( .DIN1(_30925), .DIN2(_30938), .Q(_30937) );
  nnd2s1 _30768_inst ( .DIN1(_30939), .DIN2(_28954), .Q(_30938) );
  nor2s1 _30769_inst ( .DIN1(_30772), .DIN2(_29938), .Q(_30923) );
  nnd2s1 _30770_inst ( .DIN1(_30434), .DIN2(_30940), .Q(_29938) );
  nor2s1 _30771_inst ( .DIN1(_30941), .DIN2(_30942), .Q(_30936) );
  nor2s1 _30772_inst ( .DIN1(_28954), .DIN2(_30943), .Q(_30942) );
  nnd2s1 _30773_inst ( .DIN1(_30944), .DIN2(_30890), .Q(_30943) );
  nor2s1 _30774_inst ( .DIN1(_30945), .DIN2(_30946), .Q(_30944) );
  nor2s1 _30775_inst ( .DIN1(_28724), .DIN2(_26250), .Q(_30946) );
  nor2s1 _30776_inst ( .DIN1(_52963), .DIN2(_28705), .Q(_30945) );
  nor2s1 _30777_inst ( .DIN1(_28957), .DIN2(_30947), .Q(_30941) );
  nor2s1 _30778_inst ( .DIN1(_30948), .DIN2(_29045), .Q(_30947) );
  nor2s1 _30779_inst ( .DIN1(_26584), .DIN2(_26250), .Q(_29045) );
  nor2s1 _30780_inst ( .DIN1(_52932), .DIN2(_52933), .Q(_30948) );
  hi1s1 _30781_inst ( .DIN(_28954), .Q(_28957) );
  nnd2s1 _30782_inst ( .DIN1(_30949), .DIN2(_30939), .Q(_28954) );
  nnd2s1 _30783_inst ( .DIN1(_30950), .DIN2(_30951), .Q(
        ______________________________153________) );
  nor2s1 _30784_inst ( .DIN1(_30952), .DIN2(_30953), .Q(_30951) );
  nor2s1 _30785_inst ( .DIN1(_28153), .DIN2(_30954), .Q(_30953) );
  nor2s1 _30786_inst ( .DIN1(_30955), .DIN2(_27448), .Q(_30954) );
  nor2s1 _30787_inst ( .DIN1(_53059), .DIN2(_53060), .Q(_30955) );
  nor2s1 _30788_inst ( .DIN1(_30956), .DIN2(_28151), .Q(_30952) );
  nor2s1 _30789_inst ( .DIN1(_30934), .DIN2(_30957), .Q(_30956) );
  nnd2s1 _30790_inst ( .DIN1(_30958), .DIN2(_30935), .Q(_30957) );
  nnd2s1 _30791_inst ( .DIN1(_30959), .DIN2(_53019), .Q(_30935) );
  and2s1 _30792_inst ( .DIN1(_28705), .DIN2(_52934), .Q(_30959) );
  nnd2s1 _30793_inst ( .DIN1(_28724), .DIN2(_26685), .Q(_30958) );
  nnd2s1 _30794_inst ( .DIN1(_30890), .DIN2(_30960), .Q(_30934) );
  nnd2s1 _30795_inst ( .DIN1(_30961), .DIN2(_28705), .Q(_30960) );
  nor2s1 _30796_inst ( .DIN1(_52934), .DIN2(_53019), .Q(_30961) );
  nnd2s1 _30797_inst ( .DIN1(_30962), .DIN2(_28727), .Q(_30890) );
  hi1s1 _30798_inst ( .DIN(_28844), .Q(_28727) );
  nnd2s1 _30799_inst ( .DIN1(_30963), .DIN2(_30964), .Q(_28844) );
  nor2s1 _30800_inst ( .DIN1(_30965), .DIN2(_28724), .Q(_30962) );
  hi1s1 _30801_inst ( .DIN(_28705), .Q(_28724) );
  nnd2s1 _30802_inst ( .DIN1(_28922), .DIN2(_30964), .Q(_28705) );
  and2s1 _30803_inst ( .DIN1(_28148), .DIN2(_29134), .Q(_30950) );
  nnd2s1 _30804_inst ( .DIN1(_30966), .DIN2(_30967), .Q(
        ______________________________152________) );
  nnd2s1 _30805_inst ( .DIN1(_30968), .DIN2(_30969), .Q(_30967) );
  nnd2s1 _30806_inst ( .DIN1(_30970), .DIN2(_52968), .Q(_30969) );
  nnd2s1 _30807_inst ( .DIN1(_30971), .DIN2(_30972), .Q(_30966) );
  nor2s1 _30808_inst ( .DIN1(_30973), .DIN2(_30974), .Q(_30971) );
  xor2s1 _30809_inst ( .DIN1(_30975), .DIN2(_30976), .Q(_30974) );
  xor2s1 _30810_inst ( .DIN1(_52935), .DIN2(_52937), .Q(_30976) );
  nnd2s1 _30811_inst ( .DIN1(_52935), .DIN2(_52936), .Q(_30975) );
  nnd2s1 _30812_inst ( .DIN1(_30977), .DIN2(_28941), .Q(
        ______________________________151________) );
  nor2s1 _30813_inst ( .DIN1(_30978), .DIN2(_30979), .Q(_30977) );
  nor2s1 _30814_inst ( .DIN1(_30980), .DIN2(_28949), .Q(_30979) );
  and2s1 _30815_inst ( .DIN1(_30970), .DIN2(_52962), .Q(_30980) );
  and2s1 _30816_inst ( .DIN1(_28949), .DIN2(_52983), .Q(_30978) );
  nnd2s1 _30817_inst ( .DIN1(_30981), .DIN2(_30982), .Q(
        ______________________________150________) );
  nor2s1 _30818_inst ( .DIN1(_30983), .DIN2(_30984), .Q(_30981) );
  nor2s1 _30819_inst ( .DIN1(_30972), .DIN2(_30985), .Q(_30984) );
  nnd2s1 _30820_inst ( .DIN1(_30970), .DIN2(_26705), .Q(_30985) );
  nor2s1 _30821_inst ( .DIN1(_30968), .DIN2(_30986), .Q(_30983) );
  nor2s1 _30822_inst ( .DIN1(_26987), .DIN2(_26511), .Q(_30986) );
  nnd2s1 _30823_inst ( .DIN1(_30987), .DIN2(_30988), .Q(
        ______________________________14________) );
  nnd2s1 _30824_inst ( .DIN1(_27968), .DIN2(_30989), .Q(_30988) );
  xor2s1 _30825_inst ( .DIN1(_30990), .DIN2(_30991), .Q(_30989) );
  xor2s1 _30826_inst ( .DIN1(_52844), .DIN2(_53150), .Q(_30991) );
  nor2s1 _30827_inst ( .DIN1(_26261), .DIN2(_26391), .Q(_30990) );
  nor2s1 _30828_inst ( .DIN1(_28755), .DIN2(_30992), .Q(_27968) );
  nnd2s1 _30829_inst ( .DIN1(_28755), .DIN2(_30993), .Q(_30987) );
  nnd2s1 _30830_inst ( .DIN1(_30994), .DIN2(_30995), .Q(_30993) );
  nnd2s1 _30831_inst ( .DIN1(_30996), .DIN2(_53469), .Q(_30995) );
  nor2s1 _30832_inst ( .DIN1(_27873), .DIN2(_27039), .Q(_30996) );
  nnd2s1 _30833_inst ( .DIN1(_28642), .DIN2(_53183), .Q(_30994) );
  nnd2s1 _30834_inst ( .DIN1(_30997), .DIN2(_30998), .Q(
        ______________________________149________) );
  nnd2s1 _30835_inst ( .DIN1(_30999), .DIN2(_28949), .Q(_30998) );
  nor2s1 _30836_inst ( .DIN1(_28100), .DIN2(_31000), .Q(_30999) );
  nnd2s1 _30837_inst ( .DIN1(_31001), .DIN2(_26710), .Q(_31000) );
  nnd2s1 _30838_inst ( .DIN1(_31002), .DIN2(_28944), .Q(_30997) );
  nor2s1 _30839_inst ( .DIN1(_52975), .DIN2(_31003), .Q(_31002) );
  nnd2s1 _30840_inst ( .DIN1(_31004), .DIN2(_31005), .Q(
        ______________________________148________) );
  nnd2s1 _30841_inst ( .DIN1(_30968), .DIN2(_31006), .Q(_31005) );
  nnd2s1 _30842_inst ( .DIN1(_30970), .DIN2(_26687), .Q(_31006) );
  nnd2s1 _30843_inst ( .DIN1(_31007), .DIN2(_30972), .Q(_31004) );
  nor2s1 _30844_inst ( .DIN1(_26522), .DIN2(_31008), .Q(_31007) );
  nnd2s1 _30845_inst ( .DIN1(______[20]), .DIN2(_31009), .Q(_31008) );
  nor2s1 _30846_inst ( .DIN1(_31003), .DIN2(_31010), .Q(
        ______________________________147________) );
  nnd2s1 _30847_inst ( .DIN1(_28010), .DIN2(_26718), .Q(_31010) );
  nnd2s1 _30848_inst ( .DIN1(_31011), .DIN2(_31012), .Q(
        ______________________________146________) );
  nnd2s1 _30849_inst ( .DIN1(_31013), .DIN2(_30972), .Q(_31012) );
  xor2s1 _30850_inst ( .DIN1(_31014), .DIN2(_52936), .Q(_31013) );
  nnd2s1 _30851_inst ( .DIN1(_52937), .DIN2(_52935), .Q(_31014) );
  nor2s1 _30852_inst ( .DIN1(_31015), .DIN2(_31016), .Q(_31011) );
  nor2s1 _30853_inst ( .DIN1(_31017), .DIN2(_31018), .Q(_31016) );
  nnd2s1 _30854_inst ( .DIN1(_31019), .DIN2(_31020), .Q(_31018) );
  nnd2s1 _30855_inst ( .DIN1(_31021), .DIN2(_26711), .Q(_31020) );
  nnd2s1 _30856_inst ( .DIN1(_52938), .DIN2(_31022), .Q(_31019) );
  nnd2s1 _30857_inst ( .DIN1(_31023), .DIN2(_31024), .Q(
        ______________________________145________) );
  nnd2s1 _30858_inst ( .DIN1(_31025), .DIN2(_31026), .Q(_31024) );
  nnd2s1 _30859_inst ( .DIN1(_26403), .DIN2(_31027), .Q(_31025) );
  nnd2s1 _30860_inst ( .DIN1(_27247), .DIN2(_31028), .Q(_31023) );
  nnd2s1 _30861_inst ( .DIN1(_31029), .DIN2(_31030), .Q(_31028) );
  nor2s1 _30862_inst ( .DIN1(_31031), .DIN2(_31032), .Q(_31029) );
  nor2s1 _30863_inst ( .DIN1(_31021), .DIN2(_31033), .Q(_31032) );
  nor2s1 _30864_inst ( .DIN1(_28684), .DIN2(_31034), .Q(_31033) );
  xor2s1 _30865_inst ( .DIN1(_52937), .DIN2(_31035), .Q(_31034) );
  nor2s1 _30866_inst ( .DIN1(_53089), .DIN2(_52938), .Q(_31035) );
  nor2s1 _30867_inst ( .DIN1(_53332), .DIN2(_31022), .Q(_31031) );
  nor2s1 _30868_inst ( .DIN1(_31036), .DIN2(_31037), .Q(
        ______________________________144________) );
  nor2s1 _30869_inst ( .DIN1(_31038), .DIN2(_31039), .Q(_31036) );
  nnd2s1 _30870_inst ( .DIN1(_31040), .DIN2(_31041), .Q(_31039) );
  or2s1 _30871_inst ( .DIN1(_31022), .DIN2(_52836), .Q(_31041) );
  nnd2s1 _30872_inst ( .DIN1(_31042), .DIN2(_31022), .Q(_31040) );
  xnr2s1 _30873_inst ( .DIN1(_52942), .DIN2(_31043), .Q(_31042) );
  hi1s1 _30874_inst ( .DIN(_31030), .Q(_31038) );
  nnd2s1 _30875_inst ( .DIN1(_31044), .DIN2(_31045), .Q(
        ______________________________143________) );
  nnd2s1 _30876_inst ( .DIN1(_31046), .DIN2(_30972), .Q(_31045) );
  xor2s1 _30877_inst ( .DIN1(_31047), .DIN2(_31048), .Q(_31046) );
  xor2s1 _30878_inst ( .DIN1(_52948), .DIN2(_52949), .Q(_31048) );
  nnd2s1 _30879_inst ( .DIN1(_52948), .DIN2(_52939), .Q(_31047) );
  nor2s1 _30880_inst ( .DIN1(_31015), .DIN2(_31049), .Q(_31044) );
  nor2s1 _30881_inst ( .DIN1(_31017), .DIN2(_31050), .Q(_31049) );
  nnd2s1 _30882_inst ( .DIN1(_31051), .DIN2(_31052), .Q(_31050) );
  nnd2s1 _30883_inst ( .DIN1(_31021), .DIN2(_26270), .Q(_31052) );
  nnd2s1 _30884_inst ( .DIN1(_31053), .DIN2(_31022), .Q(_31051) );
  xor2s1 _30885_inst ( .DIN1(_52913), .DIN2(_52943), .Q(_31053) );
  nnd2s1 _30886_inst ( .DIN1(_30968), .DIN2(_31030), .Q(_31017) );
  hi1s1 _30887_inst ( .DIN(_30982), .Q(_31015) );
  nnd2s1 _30888_inst ( .DIN1(_31054), .DIN2(_31055), .Q(
        ______________________________142________) );
  nnd2s1 _30889_inst ( .DIN1(_31056), .DIN2(_31057), .Q(_31055) );
  xor2s1 _30890_inst ( .DIN1(_52941), .DIN2(_53051), .Q(_31057) );
  nnd2s1 _30891_inst ( .DIN1(_30856), .DIN2(_31058), .Q(_31054) );
  nnd2s1 _30892_inst ( .DIN1(_31059), .DIN2(_31030), .Q(_31058) );
  nor2s1 _30893_inst ( .DIN1(_31060), .DIN2(_31061), .Q(_31059) );
  nor2s1 _30894_inst ( .DIN1(_31021), .DIN2(_26354), .Q(_31061) );
  nor2s1 _30895_inst ( .DIN1(_53000), .DIN2(_31022), .Q(_31060) );
  nnd2s1 _30896_inst ( .DIN1(_31062), .DIN2(_31063), .Q(
        ______________________________141________) );
  nnd2s1 _30897_inst ( .DIN1(_31064), .DIN2(_31065), .Q(_31063) );
  hi1s1 _30898_inst ( .DIN(_30068), .Q(_31065) );
  nor2s1 _30899_inst ( .DIN1(_31066), .DIN2(_26773), .Q(_31064) );
  xor2s1 _30900_inst ( .DIN1(_31067), .DIN2(_53144), .Q(_31066) );
  nnd2s1 _30901_inst ( .DIN1(_52942), .DIN2(_53096), .Q(_31067) );
  nnd2s1 _30902_inst ( .DIN1(_28338), .DIN2(_31068), .Q(_31062) );
  nnd2s1 _30903_inst ( .DIN1(_31069), .DIN2(_31030), .Q(_31068) );
  nnd2s1 _30904_inst ( .DIN1(_28843), .DIN2(_31022), .Q(_31030) );
  nor2s1 _30905_inst ( .DIN1(_31070), .DIN2(_31071), .Q(_31069) );
  nor2s1 _30906_inst ( .DIN1(_31021), .DIN2(_31072), .Q(_31071) );
  nor2s1 _30907_inst ( .DIN1(_27614), .DIN2(_31073), .Q(_31072) );
  nnd2s1 _30908_inst ( .DIN1(_31074), .DIN2(_31043), .Q(_31073) );
  nnd2s1 _30909_inst ( .DIN1(_52943), .DIN2(_26354), .Q(_31043) );
  nnd2s1 _30910_inst ( .DIN1(_52940), .DIN2(_26548), .Q(_31074) );
  hi1s1 _30911_inst ( .DIN(_31022), .Q(_31021) );
  nor2s1 _30912_inst ( .DIN1(_53288), .DIN2(_31022), .Q(_31070) );
  nnd2s1 _30913_inst ( .DIN1(_28956), .DIN2(_28864), .Q(_31022) );
  nnd2s1 _30914_inst ( .DIN1(_31075), .DIN2(_30982), .Q(
        ______________________________140________) );
  nnd2s1 _30915_inst ( .DIN1(_30973), .DIN2(_30972), .Q(_30982) );
  hi1s1 _30916_inst ( .DIN(_31009), .Q(_30973) );
  nnd2s1 _30917_inst ( .DIN1(_31076), .DIN2(_28887), .Q(_31009) );
  nor2s1 _30918_inst ( .DIN1(_30771), .DIN2(_31077), .Q(_31076) );
  nor2s1 _30919_inst ( .DIN1(_31078), .DIN2(_31079), .Q(_31075) );
  nor2s1 _30920_inst ( .DIN1(_30972), .DIN2(_31080), .Q(_31079) );
  or2s1 _30921_inst ( .DIN1(_26634), .DIN2(_30884), .Q(_31080) );
  hi1s1 _30922_inst ( .DIN(_30968), .Q(_30972) );
  nor2s1 _30923_inst ( .DIN1(_30968), .DIN2(_31081), .Q(_31078) );
  nor2s1 _30924_inst ( .DIN1(_26855), .DIN2(_26354), .Q(_31081) );
  nor2s1 _30925_inst ( .DIN1(_31082), .DIN2(_31083), .Q(_30968) );
  or2s1 _30926_inst ( .DIN1(_30925), .DIN2(_31084), .Q(_31082) );
  nnd2s1 _30927_inst ( .DIN1(_31085), .DIN2(_31086), .Q(
        ______________________________13________) );
  nnd2s1 _30928_inst ( .DIN1(_27146), .DIN2(_31087), .Q(_31086) );
  nnd2s1 _30929_inst ( .DIN1(_31088), .DIN2(_31089), .Q(_31087) );
  nnd2s1 _30930_inst ( .DIN1(_28209), .DIN2(_31090), .Q(_31089) );
  xor2s1 _30931_inst ( .DIN1(_53192), .DIN2(_53469), .Q(_31090) );
  or2s1 _30932_inst ( .DIN1(_31091), .DIN2(_53046), .Q(_31088) );
  nnd2s1 _30933_inst ( .DIN1(_31092), .DIN2(_27144), .Q(_31085) );
  nor2s1 _30934_inst ( .DIN1(_27606), .DIN2(_31093), .Q(_31092) );
  xor2s1 _30935_inst ( .DIN1(_53508), .DIN2(_28296), .Q(_31093) );
  nnd2s1 _30936_inst ( .DIN1(_31094), .DIN2(_28941), .Q(
        ______________________________139________) );
  nor2s1 _30937_inst ( .DIN1(_31095), .DIN2(_31096), .Q(_31094) );
  nor2s1 _30938_inst ( .DIN1(_31097), .DIN2(_28949), .Q(_31096) );
  nor2s1 _30939_inst ( .DIN1(_53434), .DIN2(_30884), .Q(_31097) );
  nor2s1 _30940_inst ( .DIN1(_28944), .DIN2(_31098), .Q(_31095) );
  nor2s1 _30941_inst ( .DIN1(_31099), .DIN2(_31100), .Q(_31098) );
  nor2s1 _30942_inst ( .DIN1(_52945), .DIN2(_28946), .Q(_31100) );
  nnd2s1 _30943_inst ( .DIN1(_26302), .DIN2(_26710), .Q(_28946) );
  nor2s1 _30944_inst ( .DIN1(_31101), .DIN2(_26302), .Q(_31099) );
  nor2s1 _30945_inst ( .DIN1(_52945), .DIN2(_52944), .Q(_31101) );
  nnd2s1 _30946_inst ( .DIN1(_31102), .DIN2(_52993), .Q(
        ______________________________138________) );
  nor2s1 _30947_inst ( .DIN1(_28925), .DIN2(_30884), .Q(_31102) );
  nnd2s1 _30948_inst ( .DIN1(_27201), .DIN2(_31103), .Q(_28925) );
  nnd2s1 _30949_inst ( .DIN1(_31104), .DIN2(_31105), .Q(
        ______________________________137________) );
  nnd2s1 _30950_inst ( .DIN1(_31106), .DIN2(_31107), .Q(_31105) );
  nnd2s1 _30951_inst ( .DIN1(_31108), .DIN2(_52948), .Q(_31106) );
  nor2s1 _30952_inst ( .DIN1(_31109), .DIN2(_27241), .Q(_31108) );
  nnd2s1 _30953_inst ( .DIN1(_31110), .DIN2(_27806), .Q(_31104) );
  nor2s1 _30954_inst ( .DIN1(_26391), .DIN2(_30884), .Q(_31110) );
  nnd2s1 _30955_inst ( .DIN1(_31111), .DIN2(_31112), .Q(
        ______________________________136________) );
  nnd2s1 _30956_inst ( .DIN1(_31113), .DIN2(_28923), .Q(_31112) );
  nor2s1 _30957_inst ( .DIN1(_31114), .DIN2(_28646), .Q(_31113) );
  xor2s1 _30958_inst ( .DIN1(_53388), .DIN2(_26470), .Q(_31114) );
  nnd2s1 _30959_inst ( .DIN1(_31115), .DIN2(_52996), .Q(_31111) );
  nor2s1 _30960_inst ( .DIN1(_28302), .DIN2(_30884), .Q(_31115) );
  nnd2s1 _30961_inst ( .DIN1(_31116), .DIN2(_31117), .Q(
        ______________________________135________) );
  nor2s1 _30962_inst ( .DIN1(_31118), .DIN2(_31119), .Q(_31117) );
  nor2s1 _30963_inst ( .DIN1(_31120), .DIN2(_28733), .Q(_31119) );
  nor2s1 _30964_inst ( .DIN1(_53382), .DIN2(_30884), .Q(_31120) );
  nnd2s1 _30965_inst ( .DIN1(_30963), .DIN2(_31121), .Q(_30884) );
  nor2s1 _30966_inst ( .DIN1(_28738), .DIN2(_31122), .Q(_31118) );
  nor2s1 _30967_inst ( .DIN1(_26772), .DIN2(_31123), .Q(_31122) );
  nnd2s1 _30968_inst ( .DIN1(_31124), .DIN2(_31125), .Q(_31123) );
  nnd2s1 _30969_inst ( .DIN1(_29040), .DIN2(_52958), .Q(_31125) );
  nor2s1 _30970_inst ( .DIN1(_26617), .DIN2(_53001), .Q(_29040) );
  nnd2s1 _30971_inst ( .DIN1(_53001), .DIN2(_26383), .Q(_31124) );
  nor2s1 _30972_inst ( .DIN1(_28740), .DIN2(_31126), .Q(_31116) );
  and2s1 _30973_inst ( .DIN1(_53001), .DIN2(_28739), .Q(_31126) );
  nor2s1 _30974_inst ( .DIN1(_28738), .DIN2(_53021), .Q(_28739) );
  hi1s1 _30975_inst ( .DIN(_31127), .Q(_28740) );
  nnd2s1 _30976_inst ( .DIN1(_31128), .DIN2(_28941), .Q(
        ______________________________134________) );
  nor2s1 _30977_inst ( .DIN1(_31129), .DIN2(_31130), .Q(_31128) );
  nor2s1 _30978_inst ( .DIN1(_28949), .DIN2(_31131), .Q(_31130) );
  nnd2s1 _30979_inst ( .DIN1(_31132), .DIN2(_31133), .Q(_31131) );
  nnd2s1 _30980_inst ( .DIN1(_30970), .DIN2(_52946), .Q(_31133) );
  nnd2s1 _30981_inst ( .DIN1(_31134), .DIN2(_53020), .Q(_31132) );
  nor2s1 _30982_inst ( .DIN1(_28843), .DIN2(_28100), .Q(_31134) );
  nor2s1 _30983_inst ( .DIN1(_28944), .DIN2(_31135), .Q(_31129) );
  xnr2s1 _30984_inst ( .DIN1(_53082), .DIN2(_31136), .Q(_31135) );
  nnd2s1 _30985_inst ( .DIN1(_31137), .DIN2(_31138), .Q(
        ______________________________133________) );
  nnd2s1 _30986_inst ( .DIN1(_27875), .DIN2(_31139), .Q(_31138) );
  xor2s1 _30987_inst ( .DIN1(_52843), .DIN2(_53497), .Q(_31139) );
  nnd2s1 _30988_inst ( .DIN1(_27868), .DIN2(_31140), .Q(_31137) );
  nnd2s1 _30989_inst ( .DIN1(_31141), .DIN2(_31142), .Q(_31140) );
  nnd2s1 _30990_inst ( .DIN1(_31143), .DIN2(_31144), .Q(_31142) );
  xor2s1 _30991_inst ( .DIN1(_52947), .DIN2(_53386), .Q(_31143) );
  or2s1 _30992_inst ( .DIN1(_31003), .DIN2(_53004), .Q(_31141) );
  nnd2s1 _30993_inst ( .DIN1(_31145), .DIN2(_31146), .Q(
        ______________________________132________) );
  nnd2s1 _30994_inst ( .DIN1(_31147), .DIN2(_53003), .Q(_31146) );
  nor2s1 _30995_inst ( .DIN1(_31148), .DIN2(_31149), .Q(_31145) );
  nor2s1 _30996_inst ( .DIN1(_31150), .DIN2(_31151), .Q(_31149) );
  nor2s1 _30997_inst ( .DIN1(_28843), .DIN2(_31152), .Q(_31150) );
  xor2s1 _30998_inst ( .DIN1(_31153), .DIN2(_31154), .Q(_31152) );
  xor2s1 _30999_inst ( .DIN1(_52950), .DIN2(_52951), .Q(_31154) );
  nor2s1 _31000_inst ( .DIN1(_52952), .DIN2(_52949), .Q(_31153) );
  nor2s1 _31001_inst ( .DIN1(_27804), .DIN2(_31155), .Q(_31148) );
  nnd2s1 _31002_inst ( .DIN1(______[16]), .DIN2(_31156), .Q(_31155) );
  xnr2s1 _31003_inst ( .DIN1(_52939), .DIN2(_31157), .Q(_31156) );
  nnd2s1 _31004_inst ( .DIN1(_52949), .DIN2(_52948), .Q(_31157) );
  nnd2s1 _31005_inst ( .DIN1(_31158), .DIN2(_31159), .Q(
        ______________________________131________) );
  nnd2s1 _31006_inst ( .DIN1(_31147), .DIN2(_53005), .Q(_31159) );
  hi1s1 _31007_inst ( .DIN(_31160), .Q(_31147) );
  nor2s1 _31008_inst ( .DIN1(_31161), .DIN2(_31162), .Q(_31158) );
  nor2s1 _31009_inst ( .DIN1(_31163), .DIN2(_31151), .Q(_31162) );
  nor2s1 _31010_inst ( .DIN1(_27039), .DIN2(_31164), .Q(_31163) );
  nnd2s1 _31011_inst ( .DIN1(_31144), .DIN2(_26532), .Q(_31164) );
  nor2s1 _31012_inst ( .DIN1(_31165), .DIN2(_27804), .Q(_31161) );
  xor2s1 _31013_inst ( .DIN1(_31166), .DIN2(_53052), .Q(_31165) );
  nnd2s1 _31014_inst ( .DIN1(_31167), .DIN2(_31168), .Q(
        ______________________________130________) );
  or2s1 _31015_inst ( .DIN1(_31151), .DIN2(_31169), .Q(_31168) );
  nor2s1 _31016_inst ( .DIN1(_31170), .DIN2(_31171), .Q(_31167) );
  nor2s1 _31017_inst ( .DIN1(_26622), .DIN2(_31160), .Q(_31171) );
  nor2s1 _31018_inst ( .DIN1(_27804), .DIN2(_31172), .Q(_31170) );
  xor2s1 _31019_inst ( .DIN1(_26392), .DIN2(_31166), .Q(_31172) );
  nnd2s1 _31020_inst ( .DIN1(_52952), .DIN2(_52951), .Q(_31166) );
  nnd2s1 _31021_inst ( .DIN1(_31173), .DIN2(_31107), .Q(_27804) );
  nor2s1 _31022_inst ( .DIN1(_31174), .DIN2(_28998), .Q(
        ______________________________12________) );
  nor2s1 _31023_inst ( .DIN1(_31175), .DIN2(_31176), .Q(_31174) );
  nor2s1 _31024_inst ( .DIN1(_52839), .DIN2(_31091), .Q(_31176) );
  nor2s1 _31025_inst ( .DIN1(_27651), .DIN2(_31177), .Q(_31175) );
  nnd2s1 _31026_inst ( .DIN1(_31178), .DIN2(_31179), .Q(_31177) );
  or2s1 _31027_inst ( .DIN1(_26251), .DIN2(_28643), .Q(_31179) );
  nor2s1 _31028_inst ( .DIN1(_27873), .DIN2(_31180), .Q(_28643) );
  nnd2s1 _31029_inst ( .DIN1(_31181), .DIN2(_26251), .Q(_31178) );
  nnd2s1 _31030_inst ( .DIN1(_31180), .DIN2(_28177), .Q(_31181) );
  nnd2s1 _31031_inst ( .DIN1(_31182), .DIN2(_31183), .Q(
        ______________________________129________) );
  nor2s1 _31032_inst ( .DIN1(_31184), .DIN2(_31185), .Q(_31183) );
  nor2s1 _31033_inst ( .DIN1(_26733), .DIN2(_31186), .Q(_31185) );
  nnd2s1 _31034_inst ( .DIN1(_31169), .DIN2(_31187), .Q(_31186) );
  hi1s1 _31035_inst ( .DIN(_31151), .Q(_31187) );
  nnd2s1 _31036_inst ( .DIN1(_27806), .DIN2(_31003), .Q(_31151) );
  nor2s1 _31037_inst ( .DIN1(_26392), .DIN2(_28843), .Q(_31169) );
  nor2s1 _31038_inst ( .DIN1(_52952), .DIN2(_31188), .Q(_31184) );
  nor2s1 _31039_inst ( .DIN1(_31189), .DIN2(_31107), .Q(_31188) );
  nor2s1 _31040_inst ( .DIN1(_52950), .DIN2(_28843), .Q(_31189) );
  hi1s1 _31041_inst ( .DIN(_31144), .Q(_28843) );
  nnd2s1 _31042_inst ( .DIN1(_28985), .DIN2(_31190), .Q(_31144) );
  nor2s1 _31043_inst ( .DIN1(_31191), .DIN2(_31192), .Q(_31182) );
  nor2s1 _31044_inst ( .DIN1(_27806), .DIN2(_31173), .Q(_31192) );
  nor2s1 _31045_inst ( .DIN1(_26736), .DIN2(_31160), .Q(_31191) );
  nnd2s1 _31046_inst ( .DIN1(_30970), .DIN2(_27806), .Q(_31160) );
  hi1s1 _31047_inst ( .DIN(_31107), .Q(_27806) );
  nnd2s1 _31048_inst ( .DIN1(_31193), .DIN2(_31194), .Q(_31107) );
  nor2s1 _31049_inst ( .DIN1(_31195), .DIN2(_31196), .Q(_31194) );
  hi1s1 _31050_inst ( .DIN(_31003), .Q(_30970) );
  nnd2s1 _31051_inst ( .DIN1(_28922), .DIN2(_30963), .Q(_31003) );
  hi1s1 _31052_inst ( .DIN(_28986), .Q(_28922) );
  nnd2s1 _31053_inst ( .DIN1(_28956), .DIN2(_28985), .Q(_28986) );
  hi1s1 _31054_inst ( .DIN(_28926), .Q(_28956) );
  nnd2s1 _31055_inst ( .DIN1(_31121), .DIN2(_31190), .Q(_28926) );
  nor2s1 _31056_inst ( .DIN1(_28218), .DIN2(_31197), .Q(
        ______________________________128________) );
  nor2s1 _31057_inst ( .DIN1(_31198), .DIN2(_31199), .Q(_31197) );
  nor2s1 _31058_inst ( .DIN1(_31200), .DIN2(_29866), .Q(_31199) );
  hi1s1 _31059_inst ( .DIN(_29101), .Q(_29866) );
  xor2s1 _31060_inst ( .DIN1(_31201), .DIN2(_31202), .Q(_31200) );
  xor2s1 _31061_inst ( .DIN1(_31203), .DIN2(_31204), .Q(_31202) );
  nnd2s1 _31062_inst ( .DIN1(_26836), .DIN2(_31205), .Q(_31204) );
  nnd2s1 _31063_inst ( .DIN1(_31206), .DIN2(_31207), .Q(_31203) );
  nnd2s1 _31064_inst ( .DIN1(_52957), .DIN2(_31208), .Q(_31207) );
  nnd2s1 _31065_inst ( .DIN1(_31209), .DIN2(_31210), .Q(_31208) );
  or2s1 _31066_inst ( .DIN1(_31210), .DIN2(_31209), .Q(_31206) );
  xor2s1 _31067_inst ( .DIN1(_27346), .DIN2(_52954), .Q(_31201) );
  nor2s1 _31068_inst ( .DIN1(_26621), .DIN2(_31211), .Q(_31198) );
  nnd2s1 _31069_inst ( .DIN1(______[0]), .DIN2(_29108), .Q(_31211) );
  nnd2s1 _31070_inst ( .DIN1(_31212), .DIN2(_31213), .Q(
        ______________________________127________) );
  nnd2s1 _31071_inst ( .DIN1(_31214), .DIN2(_28992), .Q(_31213) );
  nor2s1 _31072_inst ( .DIN1(_31215), .DIN2(_26771), .Q(_31214) );
  xnr2s1 _31073_inst ( .DIN1(_53182), .DIN2(_53183), .Q(_31215) );
  nnd2s1 _31074_inst ( .DIN1(_27201), .DIN2(_31216), .Q(_31212) );
  nnd2s1 _31075_inst ( .DIN1(_31217), .DIN2(_31218), .Q(_31216) );
  nnd2s1 _31076_inst ( .DIN1(_31219), .DIN2(_31220), .Q(_31218) );
  xnr2s1 _31077_inst ( .DIN1(_52956), .DIN2(_52955), .Q(_31220) );
  nor2s1 _31078_inst ( .DIN1(_29126), .DIN2(_27614), .Q(_31219) );
  hi1s1 _31079_inst ( .DIN(_29108), .Q(_29126) );
  nnd2s1 _31080_inst ( .DIN1(_31221), .DIN2(_29101), .Q(_31217) );
  xnr2s1 _31081_inst ( .DIN1(_31222), .DIN2(_29122), .Q(_29101) );
  nnd2s1 _31082_inst ( .DIN1(_31223), .DIN2(_31224), .Q(_29122) );
  nor2s1 _31083_inst ( .DIN1(_30821), .DIN2(_29903), .Q(_31224) );
  nnd2s1 _31084_inst ( .DIN1(_29999), .DIN2(_30875), .Q(_29903) );
  nor2s1 _31085_inst ( .DIN1(_29997), .DIN2(_29108), .Q(_31223) );
  nnd2s1 _31086_inst ( .DIN1(_28114), .DIN2(_28169), .Q(_29108) );
  xnr2s1 _31087_inst ( .DIN1(_31209), .DIN2(_31225), .Q(_31221) );
  xor2s1 _31088_inst ( .DIN1(_26349), .DIN2(_31210), .Q(_31225) );
  nnd2s1 _31089_inst ( .DIN1(_31226), .DIN2(_31227), .Q(_31210) );
  nnd2s1 _31090_inst ( .DIN1(_52958), .DIN2(_31228), .Q(_31227) );
  nnd2s1 _31091_inst ( .DIN1(_31229), .DIN2(_31230), .Q(_31228) );
  or2s1 _31092_inst ( .DIN1(_31230), .DIN2(_31229), .Q(_31226) );
  nnd2s1 _31093_inst ( .DIN1(_31231), .DIN2(_31232), .Q(_31209) );
  nnd2s1 _31094_inst ( .DIN1(_31233), .DIN2(_31234), .Q(_31232) );
  nnd2s1 _31095_inst ( .DIN1(_31205), .DIN2(_31235), .Q(_31234) );
  nnd2s1 _31096_inst ( .DIN1(_30104), .DIN2(_31236), .Q(_31235) );
  or2s1 _31097_inst ( .DIN1(_31236), .DIN2(_30104), .Q(_31205) );
  nnd2s1 _31098_inst ( .DIN1(_31237), .DIN2(_922), .Q(_31231) );
  hi1s1 _31099_inst ( .DIN(_31233), .Q(_922) );
  xor2s1 _31100_inst ( .DIN1(_31236), .DIN2(_30104), .Q(_31237) );
  xnr2s1 _31101_inst ( .DIN1(_31238), .DIN2(_31239), .Q(_30104) );
  xor2s1 _31102_inst ( .DIN1(_31240), .DIN2(_31233), .Q(_31239) );
  nnd2s1 _31103_inst ( .DIN1(_31241), .DIN2(_31242), .Q(_31240) );
  nnd2s1 _31104_inst ( .DIN1(_26836), .DIN2(_31243), .Q(_31242) );
  nnd2s1 _31105_inst ( .DIN1(_31244), .DIN2(_31245), .Q(_31243) );
  nnd2s1 _31106_inst ( .DIN1(_31246), .DIN2(_31247), .Q(_31241) );
  nnd2s1 _31107_inst ( .DIN1(_31248), .DIN2(_31249), .Q(_31236) );
  nnd2s1 _31108_inst ( .DIN1(_26836), .DIN2(_31250), .Q(_31249) );
  nnd2s1 _31109_inst ( .DIN1(_30124), .DIN2(_31251), .Q(_31250) );
  or2s1 _31110_inst ( .DIN1(_30124), .DIN2(_31251), .Q(_31248) );
  nnd2s1 _31111_inst ( .DIN1(_31252), .DIN2(_31253), .Q(
        ______________________________126________) );
  nnd2s1 _31112_inst ( .DIN1(_31254), .DIN2(_31255), .Q(_31253) );
  nnd2s1 _31113_inst ( .DIN1(_31256), .DIN2(_31257), .Q(_31254) );
  xor2s1 _31114_inst ( .DIN1(_31258), .DIN2(_52963), .Q(_31256) );
  nnd2s1 _31115_inst ( .DIN1(_52961), .DIN2(_52959), .Q(_31258) );
  nor2s1 _31116_inst ( .DIN1(_31259), .DIN2(_31260), .Q(_31252) );
  nor2s1 _31117_inst ( .DIN1(_31261), .DIN2(_31262), .Q(_31260) );
  xnr2s1 _31118_inst ( .DIN1(_31229), .DIN2(_31263), .Q(_31261) );
  xor2s1 _31119_inst ( .DIN1(_26383), .DIN2(_31230), .Q(_31263) );
  nnd2s1 _31120_inst ( .DIN1(_31264), .DIN2(_31265), .Q(_31230) );
  nnd2s1 _31121_inst ( .DIN1(_53107), .DIN2(_31266), .Q(_31265) );
  nnd2s1 _31122_inst ( .DIN1(_31267), .DIN2(_31268), .Q(_31266) );
  xor2s1 _31123_inst ( .DIN1(_31269), .DIN2(_31270), .Q(_31264) );
  nor2s1 _31124_inst ( .DIN1(_31267), .DIN2(_31268), .Q(_31270) );
  xor2s1 _31125_inst ( .DIN1(_30124), .DIN2(_31271), .Q(_31229) );
  xor2s1 _31126_inst ( .DIN1(_31251), .DIN2(_29166), .Q(_31271) );
  nnd2s1 _31127_inst ( .DIN1(_31272), .DIN2(_31273), .Q(_31251) );
  nnd2s1 _31128_inst ( .DIN1(_29166), .DIN2(_31274), .Q(_31273) );
  nnd2s1 _31129_inst ( .DIN1(_31275), .DIN2(_31276), .Q(_31274) );
  or2s1 _31130_inst ( .DIN1(_31276), .DIN2(_31275), .Q(_31272) );
  hi1s1 _31131_inst ( .DIN(_30143), .Q(_31275) );
  xnr2s1 _31132_inst ( .DIN1(_31277), .DIN2(_31246), .Q(_30124) );
  hi1s1 _31133_inst ( .DIN(_31245), .Q(_31246) );
  xor2s1 _31134_inst ( .DIN1(_29166), .DIN2(_31244), .Q(_31277) );
  hi1s1 _31135_inst ( .DIN(_31247), .Q(_31244) );
  nnd2s1 _31136_inst ( .DIN1(_31278), .DIN2(_31279), .Q(_31247) );
  nnd2s1 _31137_inst ( .DIN1(_31280), .DIN2(_31281), .Q(_31279) );
  xor2s1 _31138_inst ( .DIN1(_31282), .DIN2(_31283), .Q(_31278) );
  or2s1 _31139_inst ( .DIN1(_29166), .DIN2(_31284), .Q(_31283) );
  nor2s1 _31140_inst ( .DIN1(_29882), .DIN2(_31285), .Q(_31259) );
  nnd2s1 _31141_inst ( .DIN1(_31286), .DIN2(_29885), .Q(_31285) );
  nnd2s1 _31142_inst ( .DIN1(_31287), .DIN2(_31288), .Q(
        ______________________________125________) );
  nnd2s1 _31143_inst ( .DIN1(_31289), .DIN2(______[14]), .Q(_31288) );
  nor2s1 _31144_inst ( .DIN1(_31290), .DIN2(_31291), .Q(_31289) );
  xor2s1 _31145_inst ( .DIN1(_31292), .DIN2(_26564), .Q(_31290) );
  nnd2s1 _31146_inst ( .DIN1(_31293), .DIN2(_27154), .Q(_31287) );
  nor2s1 _31147_inst ( .DIN1(_31294), .DIN2(_31295), .Q(_31293) );
  nor2s1 _31148_inst ( .DIN1(_29831), .DIN2(_31296), .Q(_31295) );
  xnr2s1 _31149_inst ( .DIN1(_31267), .DIN2(_31297), .Q(_31296) );
  xor2s1 _31150_inst ( .DIN1(_26731), .DIN2(_31268), .Q(_31297) );
  nnd2s1 _31151_inst ( .DIN1(_31298), .DIN2(_31299), .Q(_31268) );
  nnd2s1 _31152_inst ( .DIN1(_53174), .DIN2(_31300), .Q(_31299) );
  nnd2s1 _31153_inst ( .DIN1(_31301), .DIN2(_31302), .Q(_31300) );
  or2s1 _31154_inst ( .DIN1(_31302), .DIN2(_31301), .Q(_31298) );
  xnr2s1 _31155_inst ( .DIN1(_26836), .DIN2(_31303), .Q(_31267) );
  xor2s1 _31156_inst ( .DIN1(_30143), .DIN2(_31276), .Q(_31303) );
  nnd2s1 _31157_inst ( .DIN1(_31304), .DIN2(_31305), .Q(_31276) );
  nnd2s1 _31158_inst ( .DIN1(_31306), .DIN2(_26836), .Q(_31305) );
  xor2s1 _31159_inst ( .DIN1(_31307), .DIN2(_31308), .Q(_31306) );
  nnd2s1 _31160_inst ( .DIN1(_31309), .DIN2(_31310), .Q(_30143) );
  nnd2s1 _31161_inst ( .DIN1(_31284), .DIN2(_29166), .Q(_31310) );
  nor2s1 _31162_inst ( .DIN1(_31281), .DIN2(_31280), .Q(_31284) );
  nor2s1 _31163_inst ( .DIN1(_31311), .DIN2(_31312), .Q(_31309) );
  nor2s1 _31164_inst ( .DIN1(_31313), .DIN2(_31314), .Q(_31312) );
  xor2s1 _31165_inst ( .DIN1(_31280), .DIN2(_29166), .Q(_31314) );
  nor2s1 _31166_inst ( .DIN1(_31281), .DIN2(_31315), .Q(_31311) );
  nnd2s1 _31167_inst ( .DIN1(_31280), .DIN2(_26836), .Q(_31315) );
  and2s1 _31168_inst ( .DIN1(_31316), .DIN2(_31317), .Q(_31280) );
  nnd2s1 _31169_inst ( .DIN1(_31318), .DIN2(_31319), .Q(_31317) );
  nnd2s1 _31170_inst ( .DIN1(_26836), .DIN2(_31320), .Q(_31319) );
  or2s1 _31171_inst ( .DIN1(_31320), .DIN2(_26836), .Q(_31316) );
  nor2s1 _31172_inst ( .DIN1(_29846), .DIN2(_31321), .Q(_31294) );
  nor2s1 _31173_inst ( .DIN1(_29848), .DIN2(_31322), .Q(_31321) );
  xor2s1 _31174_inst ( .DIN1(_26461), .DIN2(_31323), .Q(_31322) );
  nnd2s1 _31175_inst ( .DIN1(_53395), .DIN2(_26536), .Q(_31323) );
  nnd2s1 _31176_inst ( .DIN1(_31324), .DIN2(_31325), .Q(
        ______________________________124________) );
  nnd2s1 _31177_inst ( .DIN1(_31326), .DIN2(_29876), .Q(_31325) );
  hi1s1 _31178_inst ( .DIN(_31262), .Q(_29876) );
  xnr2s1 _31179_inst ( .DIN1(_31301), .DIN2(_31327), .Q(_31326) );
  xnr2s1 _31180_inst ( .DIN1(_53174), .DIN2(_31302), .Q(_31327) );
  nnd2s1 _31181_inst ( .DIN1(_31328), .DIN2(_31329), .Q(_31302) );
  nnd2s1 _31182_inst ( .DIN1(_52855), .DIN2(_31330), .Q(_31329) );
  nnd2s1 _31183_inst ( .DIN1(_31331), .DIN2(_31332), .Q(_31330) );
  or2s1 _31184_inst ( .DIN1(_31332), .DIN2(_31331), .Q(_31328) );
  nnd2s1 _31185_inst ( .DIN1(_31333), .DIN2(_31334), .Q(_31301) );
  nnd2s1 _31186_inst ( .DIN1(_29166), .DIN2(_31335), .Q(_31334) );
  nnd2s1 _31187_inst ( .DIN1(_31308), .DIN2(_31304), .Q(_31335) );
  nnd2s1 _31188_inst ( .DIN1(_31336), .DIN2(_31337), .Q(_31304) );
  hi1s1 _31189_inst ( .DIN(_30190), .Q(_31337) );
  hi1s1 _31190_inst ( .DIN(_31338), .Q(_31336) );
  nnd2s1 _31191_inst ( .DIN1(_30190), .DIN2(_31338), .Q(_31308) );
  nnd2s1 _31192_inst ( .DIN1(_31339), .DIN2(_26836), .Q(_31333) );
  xor2s1 _31193_inst ( .DIN1(_31338), .DIN2(_30190), .Q(_31339) );
  xnr2s1 _31194_inst ( .DIN1(_31318), .DIN2(_31340), .Q(_30190) );
  xor2s1 _31195_inst ( .DIN1(_31320), .DIN2(_29166), .Q(_31340) );
  nnd2s1 _31196_inst ( .DIN1(_31341), .DIN2(_31342), .Q(_31320) );
  nnd2s1 _31197_inst ( .DIN1(_31343), .DIN2(_31344), .Q(_31342) );
  or2s1 _31198_inst ( .DIN1(_31345), .DIN2(_26836), .Q(_31344) );
  nnd2s1 _31199_inst ( .DIN1(_26836), .DIN2(_31345), .Q(_31341) );
  nnd2s1 _31200_inst ( .DIN1(_31346), .DIN2(_31347), .Q(_31338) );
  nnd2s1 _31201_inst ( .DIN1(_30200), .DIN2(_31348), .Q(_31347) );
  or2s1 _31202_inst ( .DIN1(_31349), .DIN2(_31350), .Q(_31348) );
  nnd2s1 _31203_inst ( .DIN1(_31349), .DIN2(_31350), .Q(_31346) );
  nor2s1 _31204_inst ( .DIN1(_31351), .DIN2(_31352), .Q(_31324) );
  nor2s1 _31205_inst ( .DIN1(_31353), .DIN2(_29882), .Q(_31352) );
  nor2s1 _31206_inst ( .DIN1(_29848), .DIN2(_26440), .Q(_31353) );
  nor2s1 _31207_inst ( .DIN1(_29879), .DIN2(_31354), .Q(_31351) );
  nnd2s1 _31208_inst ( .DIN1(______[0]), .DIN2(_31355), .Q(_31354) );
  xor2s1 _31209_inst ( .DIN1(_52960), .DIN2(_52961), .Q(_31355) );
  nnd2s1 _31210_inst ( .DIN1(_31356), .DIN2(_31357), .Q(
        ______________________________123________) );
  nnd2s1 _31211_inst ( .DIN1(_31358), .DIN2(_31359), .Q(_31357) );
  nnd2s1 _31212_inst ( .DIN1(_31360), .DIN2(______[0]), .Q(_31359) );
  nor2s1 _31213_inst ( .DIN1(_29848), .DIN2(_31361), .Q(_31360) );
  xor2s1 _31214_inst ( .DIN1(_26461), .DIN2(_52959), .Q(_31361) );
  hi1s1 _31215_inst ( .DIN(_29885), .Q(_29848) );
  hi1s1 _31216_inst ( .DIN(_29882), .Q(_31358) );
  nnd2s1 _31217_inst ( .DIN1(_29792), .DIN2(_29831), .Q(_29882) );
  nor2s1 _31218_inst ( .DIN1(_31362), .DIN2(_31363), .Q(_31356) );
  nor2s1 _31219_inst ( .DIN1(_31364), .DIN2(_31262), .Q(_31363) );
  nnd2s1 _31220_inst ( .DIN1(_29792), .DIN2(_29846), .Q(_31262) );
  hi1s1 _31221_inst ( .DIN(_29831), .Q(_29846) );
  nnd2s1 _31222_inst ( .DIN1(_31365), .DIN2(_31366), .Q(_29831) );
  nor2s1 _31223_inst ( .DIN1(_30524), .DIN2(_31367), .Q(_31365) );
  xnr2s1 _31224_inst ( .DIN1(_31331), .DIN2(_31368), .Q(_31364) );
  xor2s1 _31225_inst ( .DIN1(_26496), .DIN2(_31332), .Q(_31368) );
  nnd2s1 _31226_inst ( .DIN1(_31369), .DIN2(_31370), .Q(_31332) );
  nnd2s1 _31227_inst ( .DIN1(_31371), .DIN2(_26235), .Q(_31370) );
  nnd2s1 _31228_inst ( .DIN1(_31372), .DIN2(_31373), .Q(_31371) );
  or2s1 _31229_inst ( .DIN1(_31373), .DIN2(_31372), .Q(_31369) );
  xnr2s1 _31230_inst ( .DIN1(_30200), .DIN2(_31374), .Q(_31331) );
  xor2s1 _31231_inst ( .DIN1(_31350), .DIN2(_31349), .Q(_31374) );
  nnd2s1 _31232_inst ( .DIN1(_31375), .DIN2(_31376), .Q(_31349) );
  nnd2s1 _31233_inst ( .DIN1(_15544), .DIN2(_31377), .Q(_31376) );
  or2s1 _31234_inst ( .DIN1(_31378), .DIN2(_29166), .Q(_31377) );
  nnd2s1 _31235_inst ( .DIN1(_29166), .DIN2(_31378), .Q(_31375) );
  nnd2s1 _31236_inst ( .DIN1(_31379), .DIN2(_31380), .Q(_31350) );
  nnd2s1 _31237_inst ( .DIN1(_31381), .DIN2(_31382), .Q(_31380) );
  or2s1 _31238_inst ( .DIN1(_31383), .DIN2(_30221), .Q(_31382) );
  nnd2s1 _31239_inst ( .DIN1(_30221), .DIN2(_31383), .Q(_31379) );
  xor2s1 _31240_inst ( .DIN1(_31343), .DIN2(_31384), .Q(_30200) );
  xor2s1 _31241_inst ( .DIN1(_31345), .DIN2(_29166), .Q(_31384) );
  nnd2s1 _31242_inst ( .DIN1(_31385), .DIN2(_31386), .Q(_31345) );
  nnd2s1 _31243_inst ( .DIN1(_31387), .DIN2(_31388), .Q(_31386) );
  or2s1 _31244_inst ( .DIN1(_31389), .DIN2(_26836), .Q(_31388) );
  nnd2s1 _31245_inst ( .DIN1(_26836), .DIN2(_31389), .Q(_31385) );
  nor2s1 _31246_inst ( .DIN1(_26536), .DIN2(_31390), .Q(_31362) );
  nnd2s1 _31247_inst ( .DIN1(_29822), .DIN2(______[22]), .Q(_31390) );
  nnd2s1 _31248_inst ( .DIN1(_31391), .DIN2(_31392), .Q(
        ______________________________122________) );
  nnd2s1 _31249_inst ( .DIN1(_31393), .DIN2(_29822), .Q(_31392) );
  hi1s1 _31250_inst ( .DIN(_29879), .Q(_29822) );
  nnd2s1 _31251_inst ( .DIN1(_31255), .DIN2(_31257), .Q(_29879) );
  nnd2s1 _31252_inst ( .DIN1(_31394), .DIN2(_31395), .Q(_31257) );
  nor2s1 _31253_inst ( .DIN1(_29433), .DIN2(_31396), .Q(_31395) );
  nor2s1 _31254_inst ( .DIN1(_31397), .DIN2(_29409), .Q(_31394) );
  nnd2s1 _31255_inst ( .DIN1(_31398), .DIN2(_31399), .Q(_29409) );
  nor2s1 _31256_inst ( .DIN1(_31400), .DIN2(_27310), .Q(_31398) );
  and2s1 _31257_inst ( .DIN1(_31286), .DIN2(______[22]), .Q(_31393) );
  xor2s1 _31258_inst ( .DIN1(_52961), .DIN2(_52959), .Q(_31286) );
  nnd2s1 _31259_inst ( .DIN1(_31401), .DIN2(_29792), .Q(_31391) );
  hi1s1 _31260_inst ( .DIN(_31255), .Q(_29792) );
  nnd2s1 _31261_inst ( .DIN1(_31402), .DIN2(_31403), .Q(_31255) );
  nor2s1 _31262_inst ( .DIN1(_29288), .DIN2(_31404), .Q(_31403) );
  nor2s1 _31263_inst ( .DIN1(_29768), .DIN2(_31405), .Q(_31402) );
  nnd2s1 _31264_inst ( .DIN1(_31406), .DIN2(_29742), .Q(_29768) );
  nor2s1 _31265_inst ( .DIN1(_27316), .DIN2(_27310), .Q(_31406) );
  nor2s1 _31266_inst ( .DIN1(_31407), .DIN2(_31408), .Q(_31401) );
  nor2s1 _31267_inst ( .DIN1(_31409), .DIN2(_31410), .Q(_31408) );
  nnd2s1 _31268_inst ( .DIN1(_31411), .DIN2(______[16]), .Q(_31410) );
  nor2s1 _31269_inst ( .DIN1(_31412), .DIN2(_31413), .Q(_31411) );
  xor2s1 _31270_inst ( .DIN1(_31414), .DIN2(_52962), .Q(_31413) );
  nnd2s1 _31271_inst ( .DIN1(_52968), .DIN2(_52967), .Q(_31414) );
  nor2s1 _31272_inst ( .DIN1(_31415), .DIN2(_31416), .Q(_31407) );
  xor2s1 _31273_inst ( .DIN1(_31372), .DIN2(_31417), .Q(_31416) );
  xor2s1 _31274_inst ( .DIN1(_26235), .DIN2(_31373), .Q(_31417) );
  nnd2s1 _31275_inst ( .DIN1(_31418), .DIN2(_31419), .Q(_31373) );
  nnd2s1 _31276_inst ( .DIN1(_31420), .DIN2(_26512), .Q(_31419) );
  or2s1 _31277_inst ( .DIN1(_31421), .DIN2(_31422), .Q(_31420) );
  nnd2s1 _31278_inst ( .DIN1(_31422), .DIN2(_31421), .Q(_31418) );
  xor2s1 _31279_inst ( .DIN1(_31381), .DIN2(_31423), .Q(_31372) );
  xor2s1 _31280_inst ( .DIN1(_31383), .DIN2(_30221), .Q(_31423) );
  xor2s1 _31281_inst ( .DIN1(_31387), .DIN2(_31424), .Q(_30221) );
  xor2s1 _31282_inst ( .DIN1(_31389), .DIN2(_29166), .Q(_31424) );
  nnd2s1 _31283_inst ( .DIN1(_31425), .DIN2(_31426), .Q(_31389) );
  nnd2s1 _31284_inst ( .DIN1(_31427), .DIN2(_31428), .Q(_31426) );
  or2s1 _31285_inst ( .DIN1(_31429), .DIN2(_31238), .Q(_31428) );
  nnd2s1 _31286_inst ( .DIN1(_31238), .DIN2(_31429), .Q(_31425) );
  nnd2s1 _31287_inst ( .DIN1(_31430), .DIN2(_31431), .Q(_31383) );
  nnd2s1 _31288_inst ( .DIN1(_31432), .DIN2(_31433), .Q(_31431) );
  xnr2s1 _31289_inst ( .DIN1(_29492), .DIN2(_31434), .Q(_31432) );
  nnd2s1 _31290_inst ( .DIN1(_31435), .DIN2(_31436), .Q(_31434) );
  or2s1 _31291_inst ( .DIN1(_31435), .DIN2(_31436), .Q(_31430) );
  hi1s1 _31292_inst ( .DIN(_30248), .Q(_31436) );
  xnr2s1 _31293_inst ( .DIN1(_31378), .DIN2(_31437), .Q(_31381) );
  nnd2s1 _31294_inst ( .DIN1(_31438), .DIN2(_31439), .Q(_31378) );
  nnd2s1 _31295_inst ( .DIN1(_359), .DIN2(_31440), .Q(_31439) );
  or2s1 _31296_inst ( .DIN1(_31441), .DIN2(_29166), .Q(_31440) );
  nnd2s1 _31297_inst ( .DIN1(_29166), .DIN2(_31441), .Q(_31438) );
  nnd2s1 _31298_inst ( .DIN1(_31442), .DIN2(_26993), .Q(
        ______________________________121________) );
  nor2s1 _31299_inst ( .DIN1(_31443), .DIN2(_31444), .Q(_31442) );
  nor2s1 _31300_inst ( .DIN1(_26996), .DIN2(_31445), .Q(_31444) );
  nor2s1 _31301_inst ( .DIN1(_31446), .DIN2(_31447), .Q(_31445) );
  nor2s1 _31302_inst ( .DIN1(_31415), .DIN2(_31448), .Q(_31447) );
  xor2s1 _31303_inst ( .DIN1(_31449), .DIN2(_31450), .Q(_31448) );
  xor2s1 _31304_inst ( .DIN1(_26512), .DIN2(_31421), .Q(_31450) );
  nnd2s1 _31305_inst ( .DIN1(_31451), .DIN2(_31452), .Q(_31421) );
  nnd2s1 _31306_inst ( .DIN1(_26401), .DIN2(_31453), .Q(_31452) );
  nnd2s1 _31307_inst ( .DIN1(_31454), .DIN2(_31455), .Q(_31453) );
  xor2s1 _31308_inst ( .DIN1(_31456), .DIN2(_31457), .Q(_31451) );
  xor2s1 _31309_inst ( .DIN1(_31458), .DIN2(_28195), .Q(_31457) );
  xor2s1 _31310_inst ( .DIN1(_31459), .DIN2(_31422), .Q(_31449) );
  xnr2s1 _31311_inst ( .DIN1(_30248), .DIN2(_31460), .Q(_31422) );
  xnr2s1 _31312_inst ( .DIN1(_31433), .DIN2(_31461), .Q(_31460) );
  nor2s1 _31313_inst ( .DIN1(_31462), .DIN2(_31435), .Q(_31461) );
  xnr2s1 _31314_inst ( .DIN1(_31441), .DIN2(_31463), .Q(_31435) );
  nnd2s1 _31315_inst ( .DIN1(_31464), .DIN2(_31465), .Q(_31441) );
  nnd2s1 _31316_inst ( .DIN1(_15546), .DIN2(_31466), .Q(_31465) );
  or2s1 _31317_inst ( .DIN1(_31467), .DIN2(_15544), .Q(_31466) );
  nnd2s1 _31318_inst ( .DIN1(_15544), .DIN2(_31467), .Q(_31464) );
  nnd2s1 _31319_inst ( .DIN1(_31468), .DIN2(_31469), .Q(_31433) );
  nnd2s1 _31320_inst ( .DIN1(_31470), .DIN2(_31471), .Q(_31469) );
  or2s1 _31321_inst ( .DIN1(_31472), .DIN2(_30263), .Q(_31471) );
  nnd2s1 _31322_inst ( .DIN1(_30263), .DIN2(_31472), .Q(_31468) );
  xnr2s1 _31323_inst ( .DIN1(_31238), .DIN2(_31473), .Q(_30248) );
  xor2s1 _31324_inst ( .DIN1(_31429), .DIN2(_31427), .Q(_31473) );
  nnd2s1 _31325_inst ( .DIN1(_31474), .DIN2(_31475), .Q(_31429) );
  nnd2s1 _31326_inst ( .DIN1(_31476), .DIN2(_31477), .Q(_31475) );
  or2s1 _31327_inst ( .DIN1(_31478), .DIN2(_31245), .Q(_31477) );
  nnd2s1 _31328_inst ( .DIN1(_31245), .DIN2(_31478), .Q(_31474) );
  xnr2s1 _31329_inst ( .DIN1(_31437), .DIN2(_31479), .Q(_31238) );
  xor2s1 _31330_inst ( .DIN1(_15544), .DIN2(_26836), .Q(_31437) );
  xnr2s1 _31331_inst ( .DIN1(_31480), .DIN2(_29994), .Q(_31479) );
  nnd2s1 _31332_inst ( .DIN1(_31481), .DIN2(_31482), .Q(_31480) );
  nnd2s1 _31333_inst ( .DIN1(_31483), .DIN2(_31484), .Q(_31482) );
  nnd2s1 _31334_inst ( .DIN1(_26836), .DIN2(_31485), .Q(_31484) );
  or2s1 _31335_inst ( .DIN1(_31485), .DIN2(_26836), .Q(_31481) );
  nor2s1 _31336_inst ( .DIN1(_31409), .DIN2(_31486), .Q(_31446) );
  nnd2s1 _31337_inst ( .DIN1(_31487), .DIN2(______[20]), .Q(_31486) );
  nor2s1 _31338_inst ( .DIN1(_31412), .DIN2(_31488), .Q(_31487) );
  xnr2s1 _31339_inst ( .DIN1(_52963), .DIN2(_52968), .Q(_31488) );
  nor2s1 _31340_inst ( .DIN1(_27007), .DIN2(_26447), .Q(_31443) );
  nnd2s1 _31341_inst ( .DIN1(_31489), .DIN2(_27983), .Q(
        ______________________________120________) );
  nor2s1 _31342_inst ( .DIN1(_31490), .DIN2(_31491), .Q(_31489) );
  nor2s1 _31343_inst ( .DIN1(_31492), .DIN2(_27500), .Q(_31491) );
  nor2s1 _31344_inst ( .DIN1(_31493), .DIN2(_31494), .Q(_31492) );
  nnd2s1 _31345_inst ( .DIN1(_31495), .DIN2(_31496), .Q(_31494) );
  nnd2s1 _31346_inst ( .DIN1(_31497), .DIN2(_26401), .Q(_31496) );
  nor2s1 _31347_inst ( .DIN1(_31498), .DIN2(_31415), .Q(_31497) );
  xnr2s1 _31348_inst ( .DIN1(_31455), .DIN2(_31454), .Q(_31498) );
  nnd2s1 _31349_inst ( .DIN1(_31499), .DIN2(_53339), .Q(_31495) );
  nor2s1 _31350_inst ( .DIN1(_31500), .DIN2(_31415), .Q(_31499) );
  nor2s1 _31351_inst ( .DIN1(_31501), .DIN2(_31458), .Q(_31500) );
  nor2s1 _31352_inst ( .DIN1(_31455), .DIN2(_31454), .Q(_31458) );
  and2s1 _31353_inst ( .DIN1(_31455), .DIN2(_31454), .Q(_31501) );
  xnr2s1 _31354_inst ( .DIN1(_31470), .DIN2(_31502), .Q(_31454) );
  xor2s1 _31355_inst ( .DIN1(_31472), .DIN2(_30263), .Q(_31502) );
  xor2s1 _31356_inst ( .DIN1(_31503), .DIN2(_31504), .Q(_30263) );
  xor2s1 _31357_inst ( .DIN1(_31478), .DIN2(_31245), .Q(_31504) );
  xor2s1 _31358_inst ( .DIN1(_31485), .DIN2(_31463), .Q(_31245) );
  xor2s1 _31359_inst ( .DIN1(_31483), .DIN2(_26836), .Q(_31463) );
  xor2s1 _31360_inst ( .DIN1(_31505), .DIN2(_31506), .Q(_31233) );
  xor2s1 _31361_inst ( .DIN1(_52883), .DIN2(_53378), .Q(_31506) );
  nnd2s1 _31362_inst ( .DIN1(_31507), .DIN2(_31508), .Q(_31505) );
  nnd2s1 _31363_inst ( .DIN1(_52851), .DIN2(_31509), .Q(_31508) );
  nnd2s1 _31364_inst ( .DIN1(_26295), .DIN2(_31510), .Q(_31509) );
  or2s1 _31365_inst ( .DIN1(_26295), .DIN2(_31510), .Q(_31507) );
  nnd2s1 _31366_inst ( .DIN1(_31511), .DIN2(_31512), .Q(_31485) );
  nnd2s1 _31367_inst ( .DIN1(_15546), .DIN2(_31513), .Q(_31512) );
  or2s1 _31368_inst ( .DIN1(_31514), .DIN2(_31515), .Q(_31513) );
  nnd2s1 _31369_inst ( .DIN1(_31515), .DIN2(_31514), .Q(_31511) );
  nnd2s1 _31370_inst ( .DIN1(_31516), .DIN2(_31517), .Q(_31478) );
  nnd2s1 _31371_inst ( .DIN1(_31518), .DIN2(_31519), .Q(_31517) );
  or2s1 _31372_inst ( .DIN1(_31313), .DIN2(_31520), .Q(_31519) );
  nnd2s1 _31373_inst ( .DIN1(_31313), .DIN2(_31520), .Q(_31516) );
  nnd2s1 _31374_inst ( .DIN1(_31521), .DIN2(_31522), .Q(_31472) );
  nnd2s1 _31375_inst ( .DIN1(_31523), .DIN2(_31524), .Q(_31522) );
  nnd2s1 _31376_inst ( .DIN1(_31525), .DIN2(_30281), .Q(_31524) );
  or2s1 _31377_inst ( .DIN1(_31525), .DIN2(_30281), .Q(_31521) );
  xnr2s1 _31378_inst ( .DIN1(_31467), .DIN2(_31526), .Q(_31470) );
  nnd2s1 _31379_inst ( .DIN1(_31527), .DIN2(_31528), .Q(_31467) );
  nnd2s1 _31380_inst ( .DIN1(_15547), .DIN2(_31529), .Q(_31528) );
  or2s1 _31381_inst ( .DIN1(_31530), .DIN2(_359), .Q(_31529) );
  nnd2s1 _31382_inst ( .DIN1(_359), .DIN2(_31530), .Q(_31527) );
  nnd2s1 _31383_inst ( .DIN1(_31531), .DIN2(_31532), .Q(_31455) );
  nnd2s1 _31384_inst ( .DIN1(_52969), .DIN2(_31533), .Q(_31532) );
  nnd2s1 _31385_inst ( .DIN1(_31534), .DIN2(_31535), .Q(_31533) );
  or2s1 _31386_inst ( .DIN1(_31535), .DIN2(_31534), .Q(_31531) );
  nor2s1 _31387_inst ( .DIN1(_31409), .DIN2(_31536), .Q(_31493) );
  nor2s1 _31388_inst ( .DIN1(_26685), .DIN2(_31537), .Q(_31536) );
  nnd2s1 _31389_inst ( .DIN1(______[2]), .DIN2(_31538), .Q(_31537) );
  nor2s1 _31390_inst ( .DIN1(_27994), .DIN2(_31539), .Q(_31490) );
  nor2s1 _31391_inst ( .DIN1(_52964), .DIN2(_26991), .Q(_31539) );
  nnd2s1 _31392_inst ( .DIN1(_31540), .DIN2(_31541), .Q(
        ______________________________11________) );
  nnd2s1 _31393_inst ( .DIN1(_31542), .DIN2(_31543), .Q(_31541) );
  nnd2s1 _31394_inst ( .DIN1(_31544), .DIN2(_28209), .Q(_31543) );
  nor2s1 _31395_inst ( .DIN1(_26774), .DIN2(_27873), .Q(_28209) );
  xor2s1 _31396_inst ( .DIN1(_26365), .DIN2(_31180), .Q(_31544) );
  nor2s1 _31397_inst ( .DIN1(_52966), .DIN2(_52986), .Q(_31180) );
  nor2s1 _31398_inst ( .DIN1(_31545), .DIN2(_31546), .Q(_31540) );
  nor2s1 _31399_inst ( .DIN1(_28930), .DIN2(_31547), .Q(_31546) );
  xor2s1 _31400_inst ( .DIN1(_31548), .DIN2(_31549), .Q(_31547) );
  xor2s1 _31401_inst ( .DIN1(_52965), .DIN2(_52966), .Q(_31549) );
  nnd2s1 _31402_inst ( .DIN1(_52874), .DIN2(_52966), .Q(_31548) );
  nor2s1 _31403_inst ( .DIN1(_29021), .DIN2(_31550), .Q(_31545) );
  or2s1 _31404_inst ( .DIN1(_31091), .DIN2(_53199), .Q(_31550) );
  nnd2s1 _31405_inst ( .DIN1(_31551), .DIN2(_31552), .Q(
        ______________________________119________) );
  nnd2s1 _31406_inst ( .DIN1(_31553), .DIN2(_31554), .Q(_31552) );
  nor2s1 _31407_inst ( .DIN1(_31555), .DIN2(_31556), .Q(_31553) );
  nor2s1 _31408_inst ( .DIN1(_31415), .DIN2(_31557), .Q(_31556) );
  xor2s1 _31409_inst ( .DIN1(_31534), .DIN2(_31558), .Q(_31557) );
  xor2s1 _31410_inst ( .DIN1(_26257), .DIN2(_31535), .Q(_31558) );
  nnd2s1 _31411_inst ( .DIN1(_31559), .DIN2(_31560), .Q(_31535) );
  nnd2s1 _31412_inst ( .DIN1(_53468), .DIN2(_31561), .Q(_31560) );
  nnd2s1 _31413_inst ( .DIN1(_31562), .DIN2(_31563), .Q(_31561) );
  nnd2s1 _31414_inst ( .DIN1(_31564), .DIN2(_31565), .Q(_31559) );
  xnr2s1 _31415_inst ( .DIN1(_31525), .DIN2(_31566), .Q(_31534) );
  xnr2s1 _31416_inst ( .DIN1(_30281), .DIN2(_31523), .Q(_31566) );
  xor2s1 _31417_inst ( .DIN1(_31567), .DIN2(_31568), .Q(_30281) );
  xor2s1 _31418_inst ( .DIN1(_31569), .DIN2(_31520), .Q(_31568) );
  nnd2s1 _31419_inst ( .DIN1(_31570), .DIN2(_31571), .Q(_31520) );
  nnd2s1 _31420_inst ( .DIN1(_31572), .DIN2(_31573), .Q(_31571) );
  or2s1 _31421_inst ( .DIN1(_31574), .DIN2(_31318), .Q(_31573) );
  nnd2s1 _31422_inst ( .DIN1(_31318), .DIN2(_31574), .Q(_31570) );
  xor2s1 _31423_inst ( .DIN1(_31518), .DIN2(_31313), .Q(_31567) );
  hi1s1 _31424_inst ( .DIN(_31281), .Q(_31313) );
  xor2s1 _31425_inst ( .DIN1(_31526), .DIN2(_31514), .Q(_31281) );
  nnd2s1 _31426_inst ( .DIN1(_31575), .DIN2(_31576), .Q(_31514) );
  nnd2s1 _31427_inst ( .DIN1(_15547), .DIN2(_31577), .Q(_31576) );
  or2s1 _31428_inst ( .DIN1(_31578), .DIN2(_31483), .Q(_31577) );
  nnd2s1 _31429_inst ( .DIN1(_31483), .DIN2(_31578), .Q(_31575) );
  xnr2s1 _31430_inst ( .DIN1(_31579), .DIN2(_15544), .Q(_31526) );
  xor2s1 _31431_inst ( .DIN1(_31510), .DIN2(_31580), .Q(_31515) );
  xor2s1 _31432_inst ( .DIN1(_52851), .DIN2(_53175), .Q(_31580) );
  nnd2s1 _31433_inst ( .DIN1(_31581), .DIN2(_31582), .Q(_31510) );
  nnd2s1 _31434_inst ( .DIN1(_31583), .DIN2(_26425), .Q(_31582) );
  or2s1 _31435_inst ( .DIN1(_31584), .DIN2(_52971), .Q(_31583) );
  nnd2s1 _31436_inst ( .DIN1(_52971), .DIN2(_31584), .Q(_31581) );
  xor2s1 _31437_inst ( .DIN1(_31585), .DIN2(_15546), .Q(_31579) );
  and2s1 _31438_inst ( .DIN1(_31586), .DIN2(_31587), .Q(_31523) );
  nnd2s1 _31439_inst ( .DIN1(_31588), .DIN2(_31589), .Q(_31587) );
  nnd2s1 _31440_inst ( .DIN1(_30284), .DIN2(_31590), .Q(_31589) );
  or2s1 _31441_inst ( .DIN1(_31590), .DIN2(_30284), .Q(_31586) );
  xor2s1 _31442_inst ( .DIN1(_31530), .DIN2(_31591), .Q(_31525) );
  nnd2s1 _31443_inst ( .DIN1(_31592), .DIN2(_31593), .Q(_31530) );
  nnd2s1 _31444_inst ( .DIN1(_15546), .DIN2(_31594), .Q(_31593) );
  or2s1 _31445_inst ( .DIN1(_31595), .DIN2(_26830), .Q(_31594) );
  nnd2s1 _31446_inst ( .DIN1(_356), .DIN2(_31595), .Q(_31592) );
  nor2s1 _31447_inst ( .DIN1(_31409), .DIN2(_31596), .Q(_31555) );
  nor2s1 _31448_inst ( .DIN1(_27651), .DIN2(_31597), .Q(_31596) );
  nnd2s1 _31449_inst ( .DIN1(_31598), .DIN2(_31538), .Q(_31597) );
  xor2s1 _31450_inst ( .DIN1(_52967), .DIN2(_52968), .Q(_31598) );
  nnd2s1 _31451_inst ( .DIN1(_31599), .DIN2(_31600), .Q(_31551) );
  xor2s1 _31452_inst ( .DIN1(_31601), .DIN2(_31602), .Q(_31600) );
  nor2s1 _31453_inst ( .DIN1(_26271), .DIN2(_26705), .Q(_31601) );
  nnd2s1 _31454_inst ( .DIN1(_31603), .DIN2(_31604), .Q(
        ______________________________118________) );
  nnd2s1 _31455_inst ( .DIN1(_31605), .DIN2(_31606), .Q(_31604) );
  nnd2s1 _31456_inst ( .DIN1(_52962), .DIN2(_31405), .Q(_31605) );
  nnd2s1 _31457_inst ( .DIN1(_31607), .DIN2(_31554), .Q(_31603) );
  nnd2s1 _31458_inst ( .DIN1(_31608), .DIN2(_31609), .Q(_31607) );
  nnd2s1 _31459_inst ( .DIN1(_31610), .DIN2(_31415), .Q(_31609) );
  nor2s1 _31460_inst ( .DIN1(_31412), .DIN2(_31611), .Q(_31610) );
  xor2s1 _31461_inst ( .DIN1(_53211), .DIN2(_31612), .Q(_31611) );
  hi1s1 _31462_inst ( .DIN(_31538), .Q(_31412) );
  nnd2s1 _31463_inst ( .DIN1(_31613), .DIN2(_31409), .Q(_31608) );
  nnd2s1 _31464_inst ( .DIN1(_31614), .DIN2(_31615), .Q(_31613) );
  nnd2s1 _31465_inst ( .DIN1(_31616), .DIN2(_26745), .Q(_31615) );
  xor2s1 _31466_inst ( .DIN1(_31564), .DIN2(_31565), .Q(_31616) );
  hi1s1 _31467_inst ( .DIN(_31562), .Q(_31565) );
  nnd2s1 _31468_inst ( .DIN1(_31617), .DIN2(_53468), .Q(_31614) );
  xor2s1 _31469_inst ( .DIN1(_31562), .DIN2(_31564), .Q(_31617) );
  hi1s1 _31470_inst ( .DIN(_31563), .Q(_31564) );
  nnd2s1 _31471_inst ( .DIN1(_31618), .DIN2(_31619), .Q(_31563) );
  nnd2s1 _31472_inst ( .DIN1(_53027), .DIN2(_31620), .Q(_31619) );
  or2s1 _31473_inst ( .DIN1(_31621), .DIN2(_31622), .Q(_31620) );
  nnd2s1 _31474_inst ( .DIN1(_31622), .DIN2(_31621), .Q(_31618) );
  xnr2s1 _31475_inst ( .DIN1(_31623), .DIN2(_31588), .Q(_31562) );
  xor2s1 _31476_inst ( .DIN1(_31595), .DIN2(_31624), .Q(_31588) );
  nnd2s1 _31477_inst ( .DIN1(_31625), .DIN2(_31626), .Q(_31595) );
  nnd2s1 _31478_inst ( .DIN1(_15547), .DIN2(_31627), .Q(_31626) );
  or2s1 _31479_inst ( .DIN1(_31628), .DIN2(_355), .Q(_31627) );
  nnd2s1 _31480_inst ( .DIN1(_355), .DIN2(_31628), .Q(_31625) );
  xnr2s1 _31481_inst ( .DIN1(_30284), .DIN2(_31590), .Q(_31623) );
  xor2s1 _31482_inst ( .DIN1(_31572), .DIN2(_31629), .Q(_30284) );
  xnr2s1 _31483_inst ( .DIN1(_31574), .DIN2(_31318), .Q(_31629) );
  xnr2s1 _31484_inst ( .DIN1(_31591), .DIN2(_31578), .Q(_31318) );
  xor2s1 _31485_inst ( .DIN1(_15547), .DIN2(_31483), .Q(_31591) );
  xnr2s1 _31486_inst ( .DIN1(_31630), .DIN2(_31584), .Q(_359) );
  nnd2s1 _31487_inst ( .DIN1(_31631), .DIN2(_31632), .Q(_31584) );
  nnd2s1 _31488_inst ( .DIN1(_31633), .DIN2(_26756), .Q(_31632) );
  or2s1 _31489_inst ( .DIN1(_26434), .DIN2(_31634), .Q(_31633) );
  nnd2s1 _31490_inst ( .DIN1(_31634), .DIN2(_26434), .Q(_31631) );
  xor2s1 _31491_inst ( .DIN1(_52971), .DIN2(_26425), .Q(_31630) );
  nnd2s1 _31492_inst ( .DIN1(_31635), .DIN2(_31636), .Q(_31578) );
  nnd2s1 _31493_inst ( .DIN1(_31637), .DIN2(_31638), .Q(_31636) );
  or2s1 _31494_inst ( .DIN1(_31639), .DIN2(_26830), .Q(_31638) );
  nnd2s1 _31495_inst ( .DIN1(_26830), .DIN2(_31639), .Q(_31635) );
  nnd2s1 _31496_inst ( .DIN1(_31640), .DIN2(_31641), .Q(_31574) );
  nnd2s1 _31497_inst ( .DIN1(_31642), .DIN2(_31643), .Q(_31641) );
  or2s1 _31498_inst ( .DIN1(_31644), .DIN2(_31645), .Q(_31643) );
  nnd2s1 _31499_inst ( .DIN1(_31645), .DIN2(_31644), .Q(_31640) );
  hi1s1 _31500_inst ( .DIN(_31343), .Q(_31645) );
  nnd2s1 _31501_inst ( .DIN1(_31646), .DIN2(_31647), .Q(_31590) );
  nnd2s1 _31502_inst ( .DIN1(_31648), .DIN2(_31649), .Q(_31647) );
  nnd2s1 _31503_inst ( .DIN1(_30328), .DIN2(_31650), .Q(_31649) );
  or2s1 _31504_inst ( .DIN1(_31650), .DIN2(_30328), .Q(_31646) );
  nnd2s1 _31505_inst ( .DIN1(_31651), .DIN2(_31652), .Q(
        ______________________________117________) );
  nnd2s1 _31506_inst ( .DIN1(_31653), .DIN2(_31606), .Q(_31652) );
  nnd2s1 _31507_inst ( .DIN1(_52973), .DIN2(_31405), .Q(_31653) );
  nnd2s1 _31508_inst ( .DIN1(_31654), .DIN2(_31554), .Q(_31651) );
  nor2s1 _31509_inst ( .DIN1(_31655), .DIN2(_31656), .Q(_31654) );
  xor2s1 _31510_inst ( .DIN1(_31657), .DIN2(_31658), .Q(_31656) );
  nnd2s1 _31511_inst ( .DIN1(_31659), .DIN2(_31409), .Q(_31657) );
  xnr2s1 _31512_inst ( .DIN1(_31622), .DIN2(_31660), .Q(_31659) );
  xor2s1 _31513_inst ( .DIN1(_26729), .DIN2(_31621), .Q(_31660) );
  nnd2s1 _31514_inst ( .DIN1(_31661), .DIN2(_31662), .Q(_31621) );
  nnd2s1 _31515_inst ( .DIN1(_52974), .DIN2(_31663), .Q(_31662) );
  nnd2s1 _31516_inst ( .DIN1(_31664), .DIN2(_31665), .Q(_31663) );
  nnd2s1 _31517_inst ( .DIN1(_31666), .DIN2(_31667), .Q(_31661) );
  hi1s1 _31518_inst ( .DIN(_31664), .Q(_31667) );
  hi1s1 _31519_inst ( .DIN(_31665), .Q(_31666) );
  xor2s1 _31520_inst ( .DIN1(_31648), .DIN2(_31668), .Q(_31622) );
  xnr2s1 _31521_inst ( .DIN1(_31650), .DIN2(_30328), .Q(_31668) );
  xnr2s1 _31522_inst ( .DIN1(_31642), .DIN2(_31669), .Q(_30328) );
  xor2s1 _31523_inst ( .DIN1(_31644), .DIN2(_31343), .Q(_31669) );
  xor2s1 _31524_inst ( .DIN1(_31639), .DIN2(_31624), .Q(_31343) );
  xor2s1 _31525_inst ( .DIN1(_31670), .DIN2(_15546), .Q(_31624) );
  hi1s1 _31526_inst ( .DIN(_31637), .Q(_15546) );
  xor2s1 _31527_inst ( .DIN1(_31634), .DIN2(_31671), .Q(_31637) );
  xor2s1 _31528_inst ( .DIN1(_52972), .DIN2(_53188), .Q(_31671) );
  nnd2s1 _31529_inst ( .DIN1(_31672), .DIN2(_31673), .Q(_31634) );
  nnd2s1 _31530_inst ( .DIN1(_52852), .DIN2(_31674), .Q(_31673) );
  nnd2s1 _31531_inst ( .DIN1(_53099), .DIN2(_31675), .Q(_31674) );
  or2s1 _31532_inst ( .DIN1(_31675), .DIN2(_53099), .Q(_31672) );
  nnd2s1 _31533_inst ( .DIN1(_31676), .DIN2(_31677), .Q(_31639) );
  nnd2s1 _31534_inst ( .DIN1(_29252), .DIN2(_31678), .Q(_31677) );
  or2s1 _31535_inst ( .DIN1(_31679), .DIN2(_355), .Q(_31678) );
  nnd2s1 _31536_inst ( .DIN1(_355), .DIN2(_31679), .Q(_31676) );
  nnd2s1 _31537_inst ( .DIN1(_31680), .DIN2(_31681), .Q(_31644) );
  xnr2s1 _31538_inst ( .DIN1(_29994), .DIN2(_31682), .Q(_31680) );
  nor2s1 _31539_inst ( .DIN1(_31683), .DIN2(_31684), .Q(_31682) );
  nnd2s1 _31540_inst ( .DIN1(_31685), .DIN2(_31686), .Q(_31650) );
  nnd2s1 _31541_inst ( .DIN1(_31687), .DIN2(_31688), .Q(_31686) );
  nnd2s1 _31542_inst ( .DIN1(_31689), .DIN2(_31690), .Q(_31688) );
  or2s1 _31543_inst ( .DIN1(_31690), .DIN2(_31689), .Q(_31685) );
  hi1s1 _31544_inst ( .DIN(_30348), .Q(_31689) );
  xnr2s1 _31545_inst ( .DIN1(_31628), .DIN2(_31691), .Q(_31648) );
  nnd2s1 _31546_inst ( .DIN1(_31692), .DIN2(_31693), .Q(_31628) );
  nnd2s1 _31547_inst ( .DIN1(_353), .DIN2(_31694), .Q(_31693) );
  or2s1 _31548_inst ( .DIN1(_31695), .DIN2(_26830), .Q(_31694) );
  nnd2s1 _31549_inst ( .DIN1(_26830), .DIN2(_31695), .Q(_31692) );
  nor2s1 _31550_inst ( .DIN1(_31696), .DIN2(_31409), .Q(_31655) );
  hi1s1 _31551_inst ( .DIN(_31415), .Q(_31409) );
  nnd2s1 _31552_inst ( .DIN1(_31697), .DIN2(_31698), .Q(_31415) );
  nor2s1 _31553_inst ( .DIN1(_31699), .DIN2(_31700), .Q(_31698) );
  nnd2s1 _31554_inst ( .DIN1(_30677), .DIN2(_30849), .Q(_31700) );
  nor2s1 _31555_inst ( .DIN1(_30832), .DIN2(_30226), .Q(_31697) );
  nnd2s1 _31556_inst ( .DIN1(_31701), .DIN2(_31702), .Q(_30226) );
  nor2s1 _31557_inst ( .DIN1(_27066), .DIN2(_31703), .Q(_31696) );
  nnd2s1 _31558_inst ( .DIN1(_31602), .DIN2(_31538), .Q(_31703) );
  xor2s1 _31559_inst ( .DIN1(_52976), .DIN2(_52973), .Q(_31602) );
  nnd2s1 _31560_inst ( .DIN1(_31704), .DIN2(_31705), .Q(
        ______________________________116________) );
  nnd2s1 _31561_inst ( .DIN1(_31599), .DIN2(_31706), .Q(_31705) );
  xor2s1 _31562_inst ( .DIN1(_26271), .DIN2(_31707), .Q(_31706) );
  nnd2s1 _31563_inst ( .DIN1(_52976), .DIN2(_52973), .Q(_31707) );
  hi1s1 _31564_inst ( .DIN(_31708), .Q(_31599) );
  nnd2s1 _31565_inst ( .DIN1(_31709), .DIN2(_31554), .Q(_31704) );
  nor2s1 _31566_inst ( .DIN1(_31710), .DIN2(_31711), .Q(_31709) );
  nor2s1 _31567_inst ( .DIN1(_28684), .DIN2(_31712), .Q(_31711) );
  nnd2s1 _31568_inst ( .DIN1(_31713), .DIN2(_26271), .Q(_31712) );
  nor2s1 _31569_inst ( .DIN1(_31714), .DIN2(_31715), .Q(_31710) );
  xor2s1 _31570_inst ( .DIN1(_31664), .DIN2(_31716), .Q(_31714) );
  xor2s1 _31571_inst ( .DIN1(_31665), .DIN2(_52974), .Q(_31716) );
  xor2s1 _31572_inst ( .DIN1(_30348), .DIN2(_31717), .Q(_31665) );
  xor2s1 _31573_inst ( .DIN1(_31690), .DIN2(_31687), .Q(_31717) );
  xor2s1 _31574_inst ( .DIN1(_31695), .DIN2(_26789), .Q(_31687) );
  nnd2s1 _31575_inst ( .DIN1(_31719), .DIN2(_31720), .Q(_31695) );
  nnd2s1 _31576_inst ( .DIN1(_355), .DIN2(_31721), .Q(_31720) );
  xor2s1 _31577_inst ( .DIN1(_30787), .DIN2(_31722), .Q(_31721) );
  nor2s1 _31578_inst ( .DIN1(_382), .DIN2(_26777), .Q(_31722) );
  nnd2s1 _31579_inst ( .DIN1(_382), .DIN2(_26777), .Q(_31719) );
  nnd2s1 _31580_inst ( .DIN1(_31724), .DIN2(_31725), .Q(_31690) );
  nnd2s1 _31581_inst ( .DIN1(_31726), .DIN2(_31727), .Q(_31725) );
  nnd2s1 _31582_inst ( .DIN1(_30384), .DIN2(_31728), .Q(_31727) );
  or2s1 _31583_inst ( .DIN1(_31728), .DIN2(_30384), .Q(_31724) );
  nnd2s1 _31584_inst ( .DIN1(_31729), .DIN2(_31730), .Q(_30348) );
  nnd2s1 _31585_inst ( .DIN1(_31731), .DIN2(_31732), .Q(_31730) );
  nnd2s1 _31586_inst ( .DIN1(_31733), .DIN2(_31681), .Q(_31732) );
  nnd2s1 _31587_inst ( .DIN1(_31734), .DIN2(_31735), .Q(_31681) );
  hi1s1 _31588_inst ( .DIN(_31683), .Q(_31733) );
  nor2s1 _31589_inst ( .DIN1(_31735), .DIN2(_31734), .Q(_31683) );
  hi1s1 _31590_inst ( .DIN(_31684), .Q(_31731) );
  nnd2s1 _31591_inst ( .DIN1(_31736), .DIN2(_31684), .Q(_31729) );
  xor2s1 _31592_inst ( .DIN1(_31735), .DIN2(_31734), .Q(_31736) );
  hi1s1 _31593_inst ( .DIN(_31387), .Q(_31734) );
  xor2s1 _31594_inst ( .DIN1(_31679), .DIN2(_31691), .Q(_31387) );
  xor2s1 _31595_inst ( .DIN1(_29304), .DIN2(_15547), .Q(_31691) );
  hi1s1 _31596_inst ( .DIN(_29252), .Q(_15547) );
  xor2s1 _31597_inst ( .DIN1(_31675), .DIN2(_31737), .Q(_29252) );
  xor2s1 _31598_inst ( .DIN1(_52852), .DIN2(_53099), .Q(_31737) );
  nnd2s1 _31599_inst ( .DIN1(_31738), .DIN2(_31739), .Q(_31675) );
  nnd2s1 _31600_inst ( .DIN1(_53176), .DIN2(_31740), .Q(_31739) );
  nnd2s1 _31601_inst ( .DIN1(_53463), .DIN2(_31741), .Q(_31740) );
  or2s1 _31602_inst ( .DIN1(_31741), .DIN2(_53463), .Q(_31738) );
  nnd2s1 _31603_inst ( .DIN1(_31742), .DIN2(_31743), .Q(_31679) );
  nnd2s1 _31604_inst ( .DIN1(_353), .DIN2(_31744), .Q(_31743) );
  or2s1 _31605_inst ( .DIN1(_31745), .DIN2(_31670), .Q(_31744) );
  nnd2s1 _31606_inst ( .DIN1(_31670), .DIN2(_31745), .Q(_31742) );
  nnd2s1 _31607_inst ( .DIN1(_31746), .DIN2(_31747), .Q(_31735) );
  nnd2s1 _31608_inst ( .DIN1(_31748), .DIN2(_31749), .Q(_31747) );
  nnd2s1 _31609_inst ( .DIN1(_31427), .DIN2(_31750), .Q(_31749) );
  or2s1 _31610_inst ( .DIN1(_31750), .DIN2(_31427), .Q(_31746) );
  xor2s1 _31611_inst ( .DIN1(_31751), .DIN2(_31752), .Q(_31664) );
  nnd2s1 _31612_inst ( .DIN1(_31753), .DIN2(_31754), .Q(_31751) );
  nnd2s1 _31613_inst ( .DIN1(_52977), .DIN2(_31755), .Q(_31754) );
  nnd2s1 _31614_inst ( .DIN1(_31756), .DIN2(_31757), .Q(_31755) );
  or2s1 _31615_inst ( .DIN1(_31757), .DIN2(_31756), .Q(_31753) );
  nnd2s1 _31616_inst ( .DIN1(_31758), .DIN2(_31759), .Q(
        ______________________________115________) );
  nnd2s1 _31617_inst ( .DIN1(_31760), .DIN2(_30175), .Q(_31759) );
  nor2s1 _31618_inst ( .DIN1(_31761), .DIN2(_31762), .Q(_31760) );
  nor2s1 _31619_inst ( .DIN1(_31763), .DIN2(_31764), .Q(_31762) );
  nnd2s1 _31620_inst ( .DIN1(_31765), .DIN2(______[24]), .Q(_31764) );
  nor2s1 _31621_inst ( .DIN1(_31766), .DIN2(_31767), .Q(_31765) );
  xor2s1 _31622_inst ( .DIN1(_31768), .DIN2(_31769), .Q(_31767) );
  or2s1 _31623_inst ( .DIN1(_31770), .DIN2(_31612), .Q(_31769) );
  nor2s1 _31624_inst ( .DIN1(_52975), .DIN2(_52976), .Q(_31612) );
  nor2s1 _31625_inst ( .DIN1(_26271), .DIN2(_26687), .Q(_31766) );
  nor2s1 _31626_inst ( .DIN1(_31715), .DIN2(_31771), .Q(_31761) );
  xnr2s1 _31627_inst ( .DIN1(_31756), .DIN2(_31772), .Q(_31771) );
  xor2s1 _31628_inst ( .DIN1(_26388), .DIN2(_31757), .Q(_31772) );
  nnd2s1 _31629_inst ( .DIN1(_31773), .DIN2(_31774), .Q(_31757) );
  nnd2s1 _31630_inst ( .DIN1(_31775), .DIN2(_26226), .Q(_31774) );
  nnd2s1 _31631_inst ( .DIN1(_31776), .DIN2(_31777), .Q(_31775) );
  or2s1 _31632_inst ( .DIN1(_31777), .DIN2(_31776), .Q(_31773) );
  xnr2s1 _31633_inst ( .DIN1(_31726), .DIN2(_31778), .Q(_31756) );
  xnr2s1 _31634_inst ( .DIN1(_31728), .DIN2(_30384), .Q(_31778) );
  xnr2s1 _31635_inst ( .DIN1(_31779), .DIN2(_31780), .Q(_30384) );
  hi1s1 _31636_inst ( .DIN(_31427), .Q(_31780) );
  xor2s1 _31637_inst ( .DIN1(_31745), .DIN2(_26789), .Q(_31427) );
  xor2s1 _31638_inst ( .DIN1(_353), .DIN2(_31670), .Q(_31718) );
  hi1s1 _31639_inst ( .DIN(_356), .Q(_31670) );
  xor2s1 _31640_inst ( .DIN1(_31741), .DIN2(_31781), .Q(_356) );
  xor2s1 _31641_inst ( .DIN1(_53176), .DIN2(_53463), .Q(_31781) );
  nnd2s1 _31642_inst ( .DIN1(_31782), .DIN2(_31783), .Q(_31741) );
  nnd2s1 _31643_inst ( .DIN1(_52978), .DIN2(_31784), .Q(_31783) );
  nnd2s1 _31644_inst ( .DIN1(_26429), .DIN2(_31785), .Q(_31784) );
  or2s1 _31645_inst ( .DIN1(_26429), .DIN2(_31785), .Q(_31782) );
  nnd2s1 _31646_inst ( .DIN1(_31786), .DIN2(_31787), .Q(_31745) );
  nnd2s1 _31647_inst ( .DIN1(_382), .DIN2(_31788), .Q(_31787) );
  or2s1 _31648_inst ( .DIN1(_31789), .DIN2(_29304), .Q(_31788) );
  nnd2s1 _31649_inst ( .DIN1(_29304), .DIN2(_31789), .Q(_31786) );
  xor2s1 _31650_inst ( .DIN1(_31750), .DIN2(_31748), .Q(_31779) );
  hi1s1 _31651_inst ( .DIN(_31790), .Q(_31748) );
  nnd2s1 _31652_inst ( .DIN1(_31791), .DIN2(_31792), .Q(_31750) );
  nnd2s1 _31653_inst ( .DIN1(_31793), .DIN2(_31794), .Q(_31792) );
  nnd2s1 _31654_inst ( .DIN1(_31503), .DIN2(_31795), .Q(_31794) );
  or2s1 _31655_inst ( .DIN1(_31795), .DIN2(_31503), .Q(_31791) );
  nnd2s1 _31656_inst ( .DIN1(_31796), .DIN2(_31797), .Q(_31728) );
  nnd2s1 _31657_inst ( .DIN1(_31798), .DIN2(_31799), .Q(_31797) );
  nnd2s1 _31658_inst ( .DIN1(_30387), .DIN2(_31800), .Q(_31799) );
  or2s1 _31659_inst ( .DIN1(_31800), .DIN2(_30387), .Q(_31796) );
  xor2s1 _31660_inst ( .DIN1(_31801), .DIN2(_26777), .Q(_31726) );
  nor2s1 _31661_inst ( .DIN1(_31804), .DIN2(_31805), .Q(_31803) );
  and2s1 _31662_inst ( .DIN1(_31806), .DIN2(_353), .Q(_31805) );
  nor2s1 _31663_inst ( .DIN1(_31807), .DIN2(_31808), .Q(_31804) );
  nor2s1 _31664_inst ( .DIN1(_353), .DIN2(_31806), .Q(_31807) );
  nnd2s1 _31665_inst ( .DIN1(_53256), .DIN2(_31809), .Q(_31758) );
  nnd2s1 _31666_inst ( .DIN1(_31810), .DIN2(_27126), .Q(
        ______________________________114________) );
  nor2s1 _31667_inst ( .DIN1(_31811), .DIN2(_31812), .Q(_31810) );
  nor2s1 _31668_inst ( .DIN1(_27132), .DIN2(_31813), .Q(_31812) );
  nnd2s1 _31669_inst ( .DIN1(_31814), .DIN2(_31815), .Q(_31813) );
  nnd2s1 _31670_inst ( .DIN1(_31816), .DIN2(_31763), .Q(_31815) );
  xor2s1 _31671_inst ( .DIN1(_31776), .DIN2(_31817), .Q(_31816) );
  xor2s1 _31672_inst ( .DIN1(_26226), .DIN2(_31777), .Q(_31817) );
  nnd2s1 _31673_inst ( .DIN1(_31818), .DIN2(_31819), .Q(_31777) );
  nnd2s1 _31674_inst ( .DIN1(_53388), .DIN2(_31820), .Q(_31819) );
  nnd2s1 _31675_inst ( .DIN1(_31821), .DIN2(_31822), .Q(_31820) );
  or2s1 _31676_inst ( .DIN1(_31822), .DIN2(_31821), .Q(_31818) );
  xor2s1 _31677_inst ( .DIN1(_31798), .DIN2(_31823), .Q(_31776) );
  xor2s1 _31678_inst ( .DIN1(_31800), .DIN2(_30387), .Q(_31823) );
  xor2s1 _31679_inst ( .DIN1(_31793), .DIN2(_31824), .Q(_30387) );
  xor2s1 _31680_inst ( .DIN1(_31795), .DIN2(_31503), .Q(_31824) );
  hi1s1 _31681_inst ( .DIN(_31476), .Q(_31503) );
  xnr2s1 _31682_inst ( .DIN1(_31789), .DIN2(_31801), .Q(_31476) );
  xnr2s1 _31683_inst ( .DIN1(_382), .DIN2(_29304), .Q(_31801) );
  xor2s1 _31684_inst ( .DIN1(_31785), .DIN2(_31825), .Q(_355) );
  xor2s1 _31685_inst ( .DIN1(_52978), .DIN2(_53045), .Q(_31825) );
  nnd2s1 _31686_inst ( .DIN1(_31826), .DIN2(_31827), .Q(_31785) );
  nnd2s1 _31687_inst ( .DIN1(_52980), .DIN2(_31828), .Q(_31827) );
  nnd2s1 _31688_inst ( .DIN1(_31829), .DIN2(_26659), .Q(_31828) );
  nnd2s1 _31689_inst ( .DIN1(_52981), .DIN2(_31830), .Q(_31826) );
  hi1s1 _31690_inst ( .DIN(_31829), .Q(_31830) );
  nnd2s1 _31691_inst ( .DIN1(_31831), .DIN2(_31832), .Q(_31789) );
  nnd2s1 _31692_inst ( .DIN1(_15550), .DIN2(_31833), .Q(_31832) );
  or2s1 _31693_inst ( .DIN1(_31834), .DIN2(_31835), .Q(_31833) );
  nnd2s1 _31694_inst ( .DIN1(_31835), .DIN2(_31834), .Q(_31831) );
  nnd2s1 _31695_inst ( .DIN1(_31836), .DIN2(_31837), .Q(_31795) );
  nnd2s1 _31696_inst ( .DIN1(_31838), .DIN2(_31839), .Q(_31837) );
  or2s1 _31697_inst ( .DIN1(_31840), .DIN2(_31841), .Q(_31839) );
  hi1s1 _31698_inst ( .DIN(_31518), .Q(_31838) );
  nnd2s1 _31699_inst ( .DIN1(_31840), .DIN2(_31841), .Q(_31836) );
  xor2s1 _31700_inst ( .DIN1(_31842), .DIN2(_31843), .Q(_31840) );
  nnd2s1 _31701_inst ( .DIN1(_31844), .DIN2(_31845), .Q(_31800) );
  nnd2s1 _31702_inst ( .DIN1(_31846), .DIN2(_31847), .Q(_31845) );
  or2s1 _31703_inst ( .DIN1(_31848), .DIN2(_30454), .Q(_31847) );
  nnd2s1 _31704_inst ( .DIN1(_30454), .DIN2(_31848), .Q(_31844) );
  xor2s1 _31705_inst ( .DIN1(_31806), .DIN2(_26764), .Q(_31798) );
  nnd2s1 _31706_inst ( .DIN1(_31849), .DIN2(_31850), .Q(_31806) );
  nnd2s1 _31707_inst ( .DIN1(_15551), .DIN2(_31851), .Q(_31850) );
  xor2s1 _31708_inst ( .DIN1(_31456), .DIN2(_31852), .Q(_31849) );
  xor2s1 _31709_inst ( .DIN1(_28088), .DIN2(_31853), .Q(_31852) );
  nor2s1 _31710_inst ( .DIN1(_31854), .DIN2(_29332), .Q(_31853) );
  nor2s1 _31711_inst ( .DIN1(_15551), .DIN2(_31851), .Q(_31854) );
  nnd2s1 _31712_inst ( .DIN1(_31855), .DIN2(_31713), .Q(_31814) );
  xor2s1 _31713_inst ( .DIN1(_31856), .DIN2(_31857), .Q(_31855) );
  xor2s1 _31714_inst ( .DIN1(_53055), .DIN2(_53332), .Q(_31857) );
  nor2s1 _31715_inst ( .DIN1(_27129), .DIN2(_31858), .Q(_31811) );
  xnr2s1 _31716_inst ( .DIN1(_52979), .DIN2(_31859), .Q(_31858) );
  nnd2s1 _31717_inst ( .DIN1(_52984), .DIN2(_53000), .Q(_31859) );
  nnd2s1 _31718_inst ( .DIN1(_31860), .DIN2(_31861), .Q(
        ______________________________113________) );
  nor2s1 _31719_inst ( .DIN1(_31862), .DIN2(_31863), .Q(_31860) );
  nor2s1 _31720_inst ( .DIN1(_31864), .DIN2(_31865), .Q(_31863) );
  nnd2s1 _31721_inst ( .DIN1(_31866), .DIN2(_31867), .Q(_31865) );
  nnd2s1 _31722_inst ( .DIN1(_52984), .DIN2(_31713), .Q(_31867) );
  nnd2s1 _31723_inst ( .DIN1(_31763), .DIN2(_31868), .Q(_31866) );
  xor2s1 _31724_inst ( .DIN1(_31821), .DIN2(_31869), .Q(_31868) );
  xnr2s1 _31725_inst ( .DIN1(_53388), .DIN2(_31822), .Q(_31869) );
  nnd2s1 _31726_inst ( .DIN1(_31870), .DIN2(_31871), .Q(_31822) );
  nnd2s1 _31727_inst ( .DIN1(_52982), .DIN2(_31872), .Q(_31871) );
  nnd2s1 _31728_inst ( .DIN1(_31873), .DIN2(_31874), .Q(_31872) );
  or2s1 _31729_inst ( .DIN1(_31874), .DIN2(_31873), .Q(_31870) );
  xor2s1 _31730_inst ( .DIN1(_31846), .DIN2(_31875), .Q(_31821) );
  xor2s1 _31731_inst ( .DIN1(_31848), .DIN2(_30454), .Q(_31875) );
  xor2s1 _31732_inst ( .DIN1(_31518), .DIN2(_31876), .Q(_30454) );
  xor2s1 _31733_inst ( .DIN1(_31841), .DIN2(_31843), .Q(_31876) );
  nnd2s1 _31734_inst ( .DIN1(_31877), .DIN2(_31878), .Q(_31841) );
  nnd2s1 _31735_inst ( .DIN1(_31879), .DIN2(_31880), .Q(_31878) );
  or2s1 _31736_inst ( .DIN1(_31881), .DIN2(_31882), .Q(_31880) );
  hi1s1 _31737_inst ( .DIN(_31883), .Q(_31879) );
  nnd2s1 _31738_inst ( .DIN1(_31882), .DIN2(_31881), .Q(_31877) );
  xor2s1 _31739_inst ( .DIN1(_31834), .DIN2(_26764), .Q(_31518) );
  xor2s1 _31740_inst ( .DIN1(_31885), .DIN2(_353), .Q(_31884) );
  hi1s1 _31741_inst ( .DIN(_31835), .Q(_353) );
  xor2s1 _31742_inst ( .DIN1(_31829), .DIN2(_31886), .Q(_31835) );
  xor2s1 _31743_inst ( .DIN1(_52980), .DIN2(_52981), .Q(_31886) );
  xor2s1 _31744_inst ( .DIN1(_31887), .DIN2(_31888), .Q(_31829) );
  nnd2s1 _31745_inst ( .DIN1(_31889), .DIN2(_31890), .Q(_31887) );
  nnd2s1 _31746_inst ( .DIN1(_31891), .DIN2(_26477), .Q(_31890) );
  nnd2s1 _31747_inst ( .DIN1(_26560), .DIN2(_31892), .Q(_31891) );
  or2s1 _31748_inst ( .DIN1(_26560), .DIN2(_31892), .Q(_31889) );
  nnd2s1 _31749_inst ( .DIN1(_31893), .DIN2(_31894), .Q(_31834) );
  nnd2s1 _31750_inst ( .DIN1(_15551), .DIN2(_31895), .Q(_31894) );
  or2s1 _31751_inst ( .DIN1(_31896), .DIN2(_29332), .Q(_31895) );
  nnd2s1 _31752_inst ( .DIN1(_29332), .DIN2(_31896), .Q(_31893) );
  nnd2s1 _31753_inst ( .DIN1(_31897), .DIN2(_31898), .Q(_31848) );
  nnd2s1 _31754_inst ( .DIN1(_31899), .DIN2(_31900), .Q(_31898) );
  or2s1 _31755_inst ( .DIN1(_31901), .DIN2(_30451), .Q(_31900) );
  nnd2s1 _31756_inst ( .DIN1(_30451), .DIN2(_31901), .Q(_31897) );
  hi1s1 _31757_inst ( .DIN(_30453), .Q(_30451) );
  xnr2s1 _31758_inst ( .DIN1(_31902), .DIN2(_31851), .Q(_31846) );
  nnd2s1 _31759_inst ( .DIN1(_31903), .DIN2(_31904), .Q(_31851) );
  nnd2s1 _31760_inst ( .DIN1(_26205), .DIN2(_31905), .Q(_31904) );
  or2s1 _31761_inst ( .DIN1(_31906), .DIN2(_15550), .Q(_31905) );
  nnd2s1 _31762_inst ( .DIN1(_15550), .DIN2(_31906), .Q(_31903) );
  hi1s1 _31763_inst ( .DIN(_31808), .Q(_15550) );
  nor2s1 _31764_inst ( .DIN1(_31907), .DIN2(_31908), .Q(_31862) );
  xor2s1 _31765_inst ( .DIN1(_31909), .DIN2(_31910), .Q(_31908) );
  xor2s1 _31766_inst ( .DIN1(_53329), .DIN2(_53488), .Q(_31910) );
  nor2s1 _31767_inst ( .DIN1(_52967), .DIN2(_26645), .Q(_31909) );
  nnd2s1 _31768_inst ( .DIN1(_27183), .DIN2(_31911), .Q(
        ______________________________112________) );
  nnd2s1 _31769_inst ( .DIN1(_31912), .DIN2(_31913), .Q(_31911) );
  nnd2s1 _31770_inst ( .DIN1(_31914), .DIN2(_31763), .Q(_31913) );
  xnr2s1 _31771_inst ( .DIN1(_31873), .DIN2(_31915), .Q(_31914) );
  xnr2s1 _31772_inst ( .DIN1(_52982), .DIN2(_31874), .Q(_31915) );
  nnd2s1 _31773_inst ( .DIN1(_31916), .DIN2(_31917), .Q(_31874) );
  nnd2s1 _31774_inst ( .DIN1(_52983), .DIN2(_31918), .Q(_31917) );
  nnd2s1 _31775_inst ( .DIN1(_31919), .DIN2(_31920), .Q(_31918) );
  or2s1 _31776_inst ( .DIN1(_31920), .DIN2(_31919), .Q(_31916) );
  xor2s1 _31777_inst ( .DIN1(_31899), .DIN2(_31921), .Q(_31873) );
  xor2s1 _31778_inst ( .DIN1(_31901), .DIN2(_30453), .Q(_31921) );
  xor2s1 _31779_inst ( .DIN1(_31883), .DIN2(_31922), .Q(_30453) );
  xor2s1 _31780_inst ( .DIN1(_31881), .DIN2(_31572), .Q(_31922) );
  hi1s1 _31781_inst ( .DIN(_31882), .Q(_31572) );
  xnr2s1 _31782_inst ( .DIN1(_31896), .DIN2(_31902), .Q(_31882) );
  xnr2s1 _31783_inst ( .DIN1(_29404), .DIN2(_29332), .Q(_31902) );
  xor2s1 _31784_inst ( .DIN1(_31923), .DIN2(_31924), .Q(_382) );
  xor2s1 _31785_inst ( .DIN1(_31925), .DIN2(_31892), .Q(_31924) );
  nnd2s1 _31786_inst ( .DIN1(_31926), .DIN2(_31927), .Q(_31892) );
  nnd2s1 _31787_inst ( .DIN1(_53184), .DIN2(_31928), .Q(_31927) );
  nnd2s1 _31788_inst ( .DIN1(_26435), .DIN2(_31929), .Q(_31928) );
  or2s1 _31789_inst ( .DIN1(_26435), .DIN2(_31929), .Q(_31926) );
  xor2s1 _31790_inst ( .DIN1(_26560), .DIN2(_53504), .Q(_31923) );
  nnd2s1 _31791_inst ( .DIN1(_31930), .DIN2(_31931), .Q(_31896) );
  nnd2s1 _31792_inst ( .DIN1(_26205), .DIN2(_31932), .Q(_31931) );
  or2s1 _31793_inst ( .DIN1(_31933), .DIN2(_31808), .Q(_31932) );
  nnd2s1 _31794_inst ( .DIN1(_31808), .DIN2(_31933), .Q(_31930) );
  nnd2s1 _31795_inst ( .DIN1(_31934), .DIN2(_31935), .Q(_31881) );
  nnd2s1 _31796_inst ( .DIN1(_31936), .DIN2(_31937), .Q(_31935) );
  or2s1 _31797_inst ( .DIN1(_31938), .DIN2(_31939), .Q(_31937) );
  hi1s1 _31798_inst ( .DIN(_31940), .Q(_31936) );
  nnd2s1 _31799_inst ( .DIN1(_31939), .DIN2(_31938), .Q(_31934) );
  hi1s1 _31800_inst ( .DIN(_31642), .Q(_31939) );
  nnd2s1 _31801_inst ( .DIN1(_31941), .DIN2(_31942), .Q(_31901) );
  nnd2s1 _31802_inst ( .DIN1(_31943), .DIN2(_31944), .Q(_31942) );
  nnd2s1 _31803_inst ( .DIN1(_30469), .DIN2(_31945), .Q(_31943) );
  hi1s1 _31804_inst ( .DIN(_31946), .Q(_31945) );
  xor2s1 _31805_inst ( .DIN1(_31947), .DIN2(_31948), .Q(_31941) );
  nnd2s1 _31806_inst ( .DIN1(_31946), .DIN2(_31949), .Q(_31948) );
  hi1s1 _31807_inst ( .DIN(_30469), .Q(_31949) );
  xnr2s1 _31808_inst ( .DIN1(_31906), .DIN2(_31950), .Q(_31899) );
  nnd2s1 _31809_inst ( .DIN1(_31951), .DIN2(_31952), .Q(_31906) );
  nnd2s1 _31810_inst ( .DIN1(_15551), .DIN2(_31953), .Q(_31952) );
  or2s1 _31811_inst ( .DIN1(_31954), .DIN2(_398), .Q(_31953) );
  nnd2s1 _31812_inst ( .DIN1(_398), .DIN2(_31954), .Q(_31951) );
  nnd2s1 _31813_inst ( .DIN1(_53332), .DIN2(_31713), .Q(_31912) );
  nnd2s1 _31814_inst ( .DIN1(_31955), .DIN2(_27256), .Q(
        ______________________________111________) );
  nor2s1 _31815_inst ( .DIN1(_31956), .DIN2(_31957), .Q(_31955) );
  nor2s1 _31816_inst ( .DIN1(_27122), .DIN2(_31958), .Q(_31957) );
  nnd2s1 _31817_inst ( .DIN1(_31959), .DIN2(_31960), .Q(_31958) );
  nnd2s1 _31818_inst ( .DIN1(_31961), .DIN2(_31763), .Q(_31960) );
  hi1s1 _31819_inst ( .DIN(_31715), .Q(_31763) );
  nnd2s1 _31820_inst ( .DIN1(_31962), .DIN2(_31963), .Q(_31715) );
  nor2s1 _31821_inst ( .DIN1(_31964), .DIN2(_30374), .Q(_31963) );
  nor2s1 _31822_inst ( .DIN1(_31367), .DIN2(_31713), .Q(_31962) );
  xor2s1 _31823_inst ( .DIN1(_31965), .DIN2(_31966), .Q(_31961) );
  xnr2s1 _31824_inst ( .DIN1(_31920), .DIN2(_31919), .Q(_31966) );
  xnr2s1 _31825_inst ( .DIN1(_31946), .DIN2(_31967), .Q(_31919) );
  xor2s1 _31826_inst ( .DIN1(_31944), .DIN2(_30469), .Q(_31967) );
  xor2s1 _31827_inst ( .DIN1(_31940), .DIN2(_31968), .Q(_30469) );
  xor2s1 _31828_inst ( .DIN1(_31938), .DIN2(_31642), .Q(_31968) );
  xor2s1 _31829_inst ( .DIN1(_31950), .DIN2(_31933), .Q(_31642) );
  nnd2s1 _31830_inst ( .DIN1(_31969), .DIN2(_31970), .Q(_31933) );
  nnd2s1 _31831_inst ( .DIN1(_29404), .DIN2(_31971), .Q(_31970) );
  or2s1 _31832_inst ( .DIN1(_31972), .DIN2(_398), .Q(_31971) );
  xnr2s1 _31833_inst ( .DIN1(_29049), .DIN2(_31973), .Q(_31969) );
  nnd2s1 _31834_inst ( .DIN1(_398), .DIN2(_31972), .Q(_31973) );
  xnr2s1 _31835_inst ( .DIN1(_31808), .DIN2(_31974), .Q(_31950) );
  xor2s1 _31836_inst ( .DIN1(_31975), .DIN2(_31976), .Q(_31974) );
  xor2s1 _31837_inst ( .DIN1(_31929), .DIN2(_31977), .Q(_31808) );
  xor2s1 _31838_inst ( .DIN1(_53184), .DIN2(_53480), .Q(_31977) );
  nnd2s1 _31839_inst ( .DIN1(_31978), .DIN2(_31979), .Q(_31929) );
  nnd2s1 _31840_inst ( .DIN1(_31980), .DIN2(_26703), .Q(_31979) );
  nnd2s1 _31841_inst ( .DIN1(_26457), .DIN2(_31981), .Q(_31980) );
  or2s1 _31842_inst ( .DIN1(_26457), .DIN2(_31981), .Q(_31978) );
  nnd2s1 _31843_inst ( .DIN1(_31982), .DIN2(_31983), .Q(_31938) );
  xor2s1 _31844_inst ( .DIN1(_31984), .DIN2(_31985), .Q(_31982) );
  nor2s1 _31845_inst ( .DIN1(_31986), .DIN2(_31987), .Q(_31985) );
  hi1s1 _31846_inst ( .DIN(_31947), .Q(_31984) );
  nnd2s1 _31847_inst ( .DIN1(_31988), .DIN2(_31989), .Q(_31944) );
  nnd2s1 _31848_inst ( .DIN1(_31990), .DIN2(_31991), .Q(_31989) );
  or2s1 _31849_inst ( .DIN1(_31992), .DIN2(_30503), .Q(_31991) );
  nnd2s1 _31850_inst ( .DIN1(_30503), .DIN2(_31992), .Q(_31988) );
  xor2s1 _31851_inst ( .DIN1(_31954), .DIN2(_26817), .Q(_31946) );
  nnd2s1 _31852_inst ( .DIN1(_31994), .DIN2(_31995), .Q(_31954) );
  nnd2s1 _31853_inst ( .DIN1(_26205), .DIN2(_31996), .Q(_31995) );
  or2s1 _31854_inst ( .DIN1(_31997), .DIN2(_15553), .Q(_31996) );
  nnd2s1 _31855_inst ( .DIN1(_15553), .DIN2(_31997), .Q(_31994) );
  nnd2s1 _31856_inst ( .DIN1(_31998), .DIN2(_31999), .Q(_31920) );
  nnd2s1 _31857_inst ( .DIN1(_32000), .DIN2(_26700), .Q(_31999) );
  nnd2s1 _31858_inst ( .DIN1(_32001), .DIN2(_32002), .Q(_32000) );
  hi1s1 _31859_inst ( .DIN(_32003), .Q(_32002) );
  nnd2s1 _31860_inst ( .DIN1(_32003), .DIN2(_32004), .Q(_31998) );
  xnr2s1 _31861_inst ( .DIN1(_52983), .DIN2(_32005), .Q(_31965) );
  nnd2s1 _31862_inst ( .DIN1(_32006), .DIN2(_32007), .Q(_31959) );
  nnd2s1 _31863_inst ( .DIN1(_31856), .DIN2(_53055), .Q(_32007) );
  and2s1 _31864_inst ( .DIN1(_53332), .DIN2(_52836), .Q(_31856) );
  nor2s1 _31865_inst ( .DIN1(_31770), .DIN2(_32008), .Q(_32006) );
  nor2s1 _31866_inst ( .DIN1(_52836), .DIN2(_32009), .Q(_32008) );
  nor2s1 _31867_inst ( .DIN1(_26270), .DIN2(_26645), .Q(_32009) );
  hi1s1 _31868_inst ( .DIN(_31713), .Q(_31770) );
  nnd2s1 _31869_inst ( .DIN1(_31701), .DIN2(_32010), .Q(_31713) );
  and2s1 _31870_inst ( .DIN1(_32011), .DIN2(_32012), .Q(_31701) );
  nor2s1 _31871_inst ( .DIN1(_30831), .DIN2(_30526), .Q(_32011) );
  nor2s1 _31872_inst ( .DIN1(_27116), .DIN2(_32013), .Q(_31956) );
  xor2s1 _31873_inst ( .DIN1(_52837), .DIN2(_53022), .Q(_32013) );
  nnd2s1 _31874_inst ( .DIN1(_32014), .DIN2(_27281), .Q(
        ______________________________110________) );
  nnd2s1 _31875_inst ( .DIN1(_27284), .DIN2(_32015), .Q(_27281) );
  nor2s1 _31876_inst ( .DIN1(_32016), .DIN2(_32017), .Q(_32014) );
  nor2s1 _31877_inst ( .DIN1(_27284), .DIN2(_32018), .Q(_32017) );
  nor2s1 _31878_inst ( .DIN1(_32019), .DIN2(_32020), .Q(_32018) );
  nor2s1 _31879_inst ( .DIN1(_32021), .DIN2(_32022), .Q(_32020) );
  xor2s1 _31880_inst ( .DIN1(_32003), .DIN2(_32023), .Q(_32021) );
  xor2s1 _31881_inst ( .DIN1(_52985), .DIN2(_32001), .Q(_32023) );
  hi1s1 _31882_inst ( .DIN(_32004), .Q(_32001) );
  nnd2s1 _31883_inst ( .DIN1(_32024), .DIN2(_32025), .Q(_32004) );
  nnd2s1 _31884_inst ( .DIN1(_32026), .DIN2(_26525), .Q(_32025) );
  nnd2s1 _31885_inst ( .DIN1(_32027), .DIN2(_32028), .Q(_32026) );
  or2s1 _31886_inst ( .DIN1(_32028), .DIN2(_32027), .Q(_32024) );
  hi1s1 _31887_inst ( .DIN(_32029), .Q(_32027) );
  xor2s1 _31888_inst ( .DIN1(_30503), .DIN2(_32030), .Q(_32003) );
  xor2s1 _31889_inst ( .DIN1(_31992), .DIN2(_31990), .Q(_32030) );
  xor2s1 _31890_inst ( .DIN1(_31997), .DIN2(_32031), .Q(_31990) );
  nnd2s1 _31891_inst ( .DIN1(_32032), .DIN2(_32033), .Q(_31997) );
  nnd2s1 _31892_inst ( .DIN1(_26204), .DIN2(_32034), .Q(_32033) );
  or2s1 _31893_inst ( .DIN1(_32035), .DIN2(_398), .Q(_32034) );
  nnd2s1 _31894_inst ( .DIN1(_398), .DIN2(_32035), .Q(_32032) );
  nnd2s1 _31895_inst ( .DIN1(_32036), .DIN2(_32037), .Q(_31992) );
  nnd2s1 _31896_inst ( .DIN1(_32038), .DIN2(_32039), .Q(_32037) );
  nnd2s1 _31897_inst ( .DIN1(_32040), .DIN2(_32041), .Q(_32038) );
  hi1s1 _31898_inst ( .DIN(_32042), .Q(_32041) );
  xor2s1 _31899_inst ( .DIN1(_31282), .DIN2(_30506), .Q(_32040) );
  hi1s1 _31900_inst ( .DIN(_30504), .Q(_30506) );
  nnd2s1 _31901_inst ( .DIN1(_32042), .DIN2(_30504), .Q(_32036) );
  nnd2s1 _31902_inst ( .DIN1(_32043), .DIN2(_32044), .Q(_30503) );
  nnd2s1 _31903_inst ( .DIN1(_31987), .DIN2(_32045), .Q(_32044) );
  nnd2s1 _31904_inst ( .DIN1(_32046), .DIN2(_31983), .Q(_32045) );
  nnd2s1 _31905_inst ( .DIN1(_31684), .DIN2(_32047), .Q(_31983) );
  hi1s1 _31906_inst ( .DIN(_31986), .Q(_32046) );
  nor2s1 _31907_inst ( .DIN1(_32047), .DIN2(_31684), .Q(_31986) );
  nnd2s1 _31908_inst ( .DIN1(_32048), .DIN2(_32049), .Q(_32043) );
  hi1s1 _31909_inst ( .DIN(_31987), .Q(_32049) );
  xor2s1 _31910_inst ( .DIN1(_32047), .DIN2(_31684), .Q(_32048) );
  xor2s1 _31911_inst ( .DIN1(_31972), .DIN2(_26817), .Q(_31684) );
  hi1s1 _31912_inst ( .DIN(_29404), .Q(_15551) );
  xor2s1 _31913_inst ( .DIN1(_31981), .DIN2(_32050), .Q(_29404) );
  xor2s1 _31914_inst ( .DIN1(_53481), .DIN2(_53482), .Q(_32050) );
  nnd2s1 _31915_inst ( .DIN1(_32051), .DIN2(_32052), .Q(_31981) );
  nnd2s1 _31916_inst ( .DIN1(_32053), .DIN2(_26702), .Q(_32052) );
  nnd2s1 _31917_inst ( .DIN1(_53483), .DIN2(_32054), .Q(_32053) );
  or2s1 _31918_inst ( .DIN1(_32054), .DIN2(_53483), .Q(_32051) );
  nnd2s1 _31919_inst ( .DIN1(_32055), .DIN2(_32056), .Q(_31972) );
  nnd2s1 _31920_inst ( .DIN1(_31976), .DIN2(_32057), .Q(_32056) );
  or2s1 _31921_inst ( .DIN1(_32058), .DIN2(_15553), .Q(_32057) );
  nnd2s1 _31922_inst ( .DIN1(_15553), .DIN2(_32058), .Q(_32055) );
  nnd2s1 _31923_inst ( .DIN1(_32059), .DIN2(_32060), .Q(_32047) );
  nnd2s1 _31924_inst ( .DIN1(_32061), .DIN2(_32062), .Q(_32060) );
  or2s1 _31925_inst ( .DIN1(_32063), .DIN2(_31790), .Q(_32062) );
  hi1s1 _31926_inst ( .DIN(_32064), .Q(_32061) );
  nnd2s1 _31927_inst ( .DIN1(_31790), .DIN2(_32063), .Q(_32059) );
  nor2s1 _31928_inst ( .DIN1(_32065), .DIN2(_32066), .Q(_32019) );
  nor2s1 _31929_inst ( .DIN1(_32067), .DIN2(_32068), .Q(_32066) );
  nnd2s1 _31930_inst ( .DIN1(_32069), .DIN2(______[20]), .Q(_32068) );
  nor2s1 _31931_inst ( .DIN1(_32070), .DIN2(_32071), .Q(_32069) );
  and2s1 _31932_inst ( .DIN1(_53433), .DIN2(_53434), .Q(_32071) );
  and2s1 _31933_inst ( .DIN1(_26634), .DIN2(_32072), .Q(_32070) );
  nnd2s1 _31934_inst ( .DIN1(_32073), .DIN2(_32074), .Q(_32067) );
  nnd2s1 _31935_inst ( .DIN1(_53434), .DIN2(_26497), .Q(_32073) );
  nor2s1 _31936_inst ( .DIN1(_27298), .DIN2(_32075), .Q(_32016) );
  nor2s1 _31937_inst ( .DIN1(_27082), .DIN2(_26711), .Q(_32075) );
  nnd2s1 _31938_inst ( .DIN1(_32076), .DIN2(_32077), .Q(
        ______________________________10________) );
  nnd2s1 _31939_inst ( .DIN1(_31542), .DIN2(_32078), .Q(_32077) );
  nnd2s1 _31940_inst ( .DIN1(_32079), .DIN2(______[18]), .Q(_32078) );
  nor2s1 _31941_inst ( .DIN1(_52986), .DIN2(_27873), .Q(_32079) );
  hi1s1 _31942_inst ( .DIN(_28177), .Q(_27873) );
  nnd2s1 _31943_inst ( .DIN1(_32080), .DIN2(_32081), .Q(_28177) );
  nor2s1 _31944_inst ( .DIN1(_29021), .DIN2(_28642), .Q(_31542) );
  nor2s1 _31945_inst ( .DIN1(_32082), .DIN2(_32083), .Q(_32076) );
  nor2s1 _31946_inst ( .DIN1(_26506), .DIN2(_32084), .Q(_32083) );
  nnd2s1 _31947_inst ( .DIN1(______[6]), .DIN2(_30640), .Q(_32084) );
  nor2s1 _31948_inst ( .DIN1(_29021), .DIN2(_32085), .Q(_32082) );
  nnd2s1 _31949_inst ( .DIN1(_28642), .DIN2(_26640), .Q(_32085) );
  hi1s1 _31950_inst ( .DIN(_31091), .Q(_28642) );
  nnd2s1 _31951_inst ( .DIN1(_32086), .DIN2(_28129), .Q(_31091) );
  hi1s1 _31952_inst ( .DIN(_28223), .Q(_28129) );
  nnd2s1 _31953_inst ( .DIN1(_32081), .DIN2(_28170), .Q(_28223) );
  nor2s1 _31954_inst ( .DIN1(_28215), .DIN2(_30054), .Q(_32086) );
  nnd2s1 _31955_inst ( .DIN1(_32087), .DIN2(_29999), .Q(_30054) );
  nor2s1 _31956_inst ( .DIN1(_28115), .DIN2(_32088), .Q(_32087) );
  nnd2s1 _31957_inst ( .DIN1(_32089), .DIN2(_28887), .Q(_29021) );
  nor2s1 _31958_inst ( .DIN1(_32090), .DIN2(_31084), .Q(_32089) );
  hi1s1 _31959_inst ( .DIN(_32091), .Q(_32090) );
  nnd2s1 _31960_inst ( .DIN1(_32092), .DIN2(_27450), .Q(
        ______________________________109________) );
  nor2s1 _31961_inst ( .DIN1(_32093), .DIN2(_32094), .Q(_32092) );
  nor2s1 _31962_inst ( .DIN1(_27453), .DIN2(_32095), .Q(_32094) );
  nor2s1 _31963_inst ( .DIN1(_32096), .DIN2(_32097), .Q(_32095) );
  nor2s1 _31964_inst ( .DIN1(_32065), .DIN2(_32098), .Q(_32097) );
  nnd2s1 _31965_inst ( .DIN1(_53000), .DIN2(_32074), .Q(_32098) );
  nor2s1 _31966_inst ( .DIN1(_32099), .DIN2(_32022), .Q(_32096) );
  xor2s1 _31967_inst ( .DIN1(_32028), .DIN2(_32100), .Q(_32099) );
  xor2s1 _31968_inst ( .DIN1(_26525), .DIN2(_32029), .Q(_32100) );
  nnd2s1 _31969_inst ( .DIN1(_32101), .DIN2(_32102), .Q(_32029) );
  nnd2s1 _31970_inst ( .DIN1(_52989), .DIN2(_32103), .Q(_32102) );
  nnd2s1 _31971_inst ( .DIN1(_32104), .DIN2(_32105), .Q(_32103) );
  or2s1 _31972_inst ( .DIN1(_32105), .DIN2(_32104), .Q(_32101) );
  xnr2s1 _31973_inst ( .DIN1(_32042), .DIN2(_32106), .Q(_32028) );
  xor2s1 _31974_inst ( .DIN1(_32039), .DIN2(_30504), .Q(_32106) );
  xor2s1 _31975_inst ( .DIN1(_32064), .DIN2(_32107), .Q(_30504) );
  xor2s1 _31976_inst ( .DIN1(_32063), .DIN2(_31790), .Q(_32107) );
  xor2s1 _31977_inst ( .DIN1(_32058), .DIN2(_32031), .Q(_31790) );
  xor2s1 _31978_inst ( .DIN1(_26205), .DIN2(_15553), .Q(_32031) );
  xor2s1 _31979_inst ( .DIN1(_32054), .DIN2(_32108), .Q(_31976) );
  xor2s1 _31980_inst ( .DIN1(_52846), .DIN2(_53483), .Q(_32108) );
  nnd2s1 _31981_inst ( .DIN1(_32109), .DIN2(_32110), .Q(_32054) );
  nnd2s1 _31982_inst ( .DIN1(_32111), .DIN2(_26393), .Q(_32110) );
  nnd2s1 _31983_inst ( .DIN1(_26726), .DIN2(_32112), .Q(_32111) );
  or2s1 _31984_inst ( .DIN1(_26726), .DIN2(_32112), .Q(_32109) );
  nnd2s1 _31985_inst ( .DIN1(_32113), .DIN2(_32114), .Q(_32058) );
  nnd2s1 _31986_inst ( .DIN1(_26204), .DIN2(_32115), .Q(_32114) );
  or2s1 _31987_inst ( .DIN1(_32116), .DIN2(_29425), .Q(_32115) );
  nnd2s1 _31988_inst ( .DIN1(_29425), .DIN2(_32116), .Q(_32113) );
  nnd2s1 _31989_inst ( .DIN1(_32117), .DIN2(_32118), .Q(_32063) );
  nnd2s1 _31990_inst ( .DIN1(_32119), .DIN2(_32120), .Q(_32118) );
  or2s1 _31991_inst ( .DIN1(_32121), .DIN2(_31793), .Q(_32120) );
  nnd2s1 _31992_inst ( .DIN1(_31793), .DIN2(_32121), .Q(_32117) );
  nnd2s1 _31993_inst ( .DIN1(_32122), .DIN2(_32123), .Q(_32039) );
  nnd2s1 _31994_inst ( .DIN1(_32124), .DIN2(_32125), .Q(_32123) );
  or2s1 _31995_inst ( .DIN1(_32126), .DIN2(_30549), .Q(_32125) );
  nnd2s1 _31996_inst ( .DIN1(_30549), .DIN2(_32126), .Q(_32122) );
  xor2s1 _31997_inst ( .DIN1(_32035), .DIN2(_32127), .Q(_32042) );
  nnd2s1 _31998_inst ( .DIN1(_32128), .DIN2(_32129), .Q(_32035) );
  nnd2s1 _31999_inst ( .DIN1(_15553), .DIN2(_32130), .Q(_32129) );
  or2s1 _32000_inst ( .DIN1(_32131), .DIN2(_26826), .Q(_32130) );
  nnd2s1 _32001_inst ( .DIN1(_408), .DIN2(_32131), .Q(_32128) );
  nor2s1 _32002_inst ( .DIN1(_27476), .DIN2(_32132), .Q(_32093) );
  nor2s1 _32003_inst ( .DIN1(_52987), .DIN2(_27291), .Q(_32132) );
  nnd2s1 _32004_inst ( .DIN1(_32133), .DIN2(_32134), .Q(
        ______________________________108________) );
  nnd2s1 _32005_inst ( .DIN1(_32135), .DIN2(_27779), .Q(_32134) );
  nnd2s1 _32006_inst ( .DIN1(_32136), .DIN2(_29859), .Q(_32135) );
  and2s1 _32007_inst ( .DIN1(_27780), .DIN2(_32137), .Q(_29859) );
  nnd2s1 _32008_inst ( .DIN1(_53452), .DIN2(_26418), .Q(_32137) );
  nor2s1 _32009_inst ( .DIN1(_32138), .DIN2(_32139), .Q(_32136) );
  nor2s1 _32010_inst ( .DIN1(_26418), .DIN2(_32140), .Q(_32139) );
  nnd2s1 _32011_inst ( .DIN1(_53433), .DIN2(_26297), .Q(_32140) );
  nor2s1 _32012_inst ( .DIN1(_52988), .DIN2(_53433), .Q(_32138) );
  nnd2s1 _32013_inst ( .DIN1(_32141), .DIN2(_27782), .Q(_32133) );
  nnd2s1 _32014_inst ( .DIN1(_32142), .DIN2(_32143), .Q(_32141) );
  nnd2s1 _32015_inst ( .DIN1(_32144), .DIN2(_32022), .Q(_32143) );
  nnd2s1 _32016_inst ( .DIN1(_32065), .DIN2(_32145), .Q(_32142) );
  xor2s1 _32017_inst ( .DIN1(_32104), .DIN2(_32146), .Q(_32145) );
  xnr2s1 _32018_inst ( .DIN1(_52989), .DIN2(_32105), .Q(_32146) );
  nnd2s1 _32019_inst ( .DIN1(_32147), .DIN2(_32148), .Q(_32105) );
  nnd2s1 _32020_inst ( .DIN1(_53432), .DIN2(_32149), .Q(_32148) );
  nnd2s1 _32021_inst ( .DIN1(_32150), .DIN2(_32151), .Q(_32149) );
  or2s1 _32022_inst ( .DIN1(_32151), .DIN2(_32150), .Q(_32147) );
  xnr2s1 _32023_inst ( .DIN1(_32124), .DIN2(_32152), .Q(_32104) );
  xor2s1 _32024_inst ( .DIN1(_32126), .DIN2(_30549), .Q(_32152) );
  xor2s1 _32025_inst ( .DIN1(_32153), .DIN2(_32154), .Q(_30549) );
  xor2s1 _32026_inst ( .DIN1(_30674), .DIN2(_32121), .Q(_32154) );
  nnd2s1 _32027_inst ( .DIN1(_32155), .DIN2(_32156), .Q(_32121) );
  nnd2s1 _32028_inst ( .DIN1(_32157), .DIN2(_32158), .Q(_32156) );
  or2s1 _32029_inst ( .DIN1(_32159), .DIN2(_32160), .Q(_32158) );
  nnd2s1 _32030_inst ( .DIN1(_32160), .DIN2(_32159), .Q(_32155) );
  hi1s1 _32031_inst ( .DIN(_31843), .Q(_32160) );
  xor2s1 _32032_inst ( .DIN1(_32161), .DIN2(_31793), .Q(_32153) );
  xor2s1 _32033_inst ( .DIN1(_32116), .DIN2(_32127), .Q(_31793) );
  xor2s1 _32034_inst ( .DIN1(_26204), .DIN2(_398), .Q(_32127) );
  hi1s1 _32035_inst ( .DIN(_29425), .Q(_398) );
  xor2s1 _32036_inst ( .DIN1(_32112), .DIN2(_32162), .Q(_29425) );
  xor2s1 _32037_inst ( .DIN1(_53484), .DIN2(_53485), .Q(_32162) );
  nnd2s1 _32038_inst ( .DIN1(_32163), .DIN2(_32164), .Q(_32112) );
  nnd2s1 _32039_inst ( .DIN1(_32165), .DIN2(_26680), .Q(_32164) );
  nnd2s1 _32040_inst ( .DIN1(_53461), .DIN2(_32166), .Q(_32165) );
  or2s1 _32041_inst ( .DIN1(_32166), .DIN2(_53461), .Q(_32163) );
  nnd2s1 _32042_inst ( .DIN1(_32167), .DIN2(_32168), .Q(_32116) );
  nnd2s1 _32043_inst ( .DIN1(_32169), .DIN2(_32170), .Q(_32168) );
  or2s1 _32044_inst ( .DIN1(_32171), .DIN2(_26826), .Q(_32170) );
  nnd2s1 _32045_inst ( .DIN1(_26826), .DIN2(_32171), .Q(_32167) );
  nnd2s1 _32046_inst ( .DIN1(_32172), .DIN2(_32173), .Q(_32126) );
  nnd2s1 _32047_inst ( .DIN1(_32174), .DIN2(_32175), .Q(_32173) );
  nnd2s1 _32048_inst ( .DIN1(_30575), .DIN2(_32176), .Q(_32175) );
  or2s1 _32049_inst ( .DIN1(_32176), .DIN2(_30575), .Q(_32172) );
  xnr2s1 _32050_inst ( .DIN1(_32131), .DIN2(_32177), .Q(_32124) );
  nnd2s1 _32051_inst ( .DIN1(_32178), .DIN2(_32179), .Q(_32131) );
  nnd2s1 _32052_inst ( .DIN1(_26204), .DIN2(_32180), .Q(_32179) );
  or2s1 _32053_inst ( .DIN1(_32181), .DIN2(_15555), .Q(_32180) );
  nnd2s1 _32054_inst ( .DIN1(_15555), .DIN2(_32181), .Q(_32178) );
  nnd2s1 _32055_inst ( .DIN1(_32182), .DIN2(_28045), .Q(
        ______________________________107________) );
  nnd2s1 _32056_inst ( .DIN1(_32183), .DIN2(_28049), .Q(_28045) );
  nor2s1 _32057_inst ( .DIN1(_32184), .DIN2(_32185), .Q(_32182) );
  nor2s1 _32058_inst ( .DIN1(_28049), .DIN2(_32186), .Q(_32185) );
  nor2s1 _32059_inst ( .DIN1(_32187), .DIN2(_32188), .Q(_32186) );
  nor2s1 _32060_inst ( .DIN1(_32065), .DIN2(_32189), .Q(_32188) );
  nnd2s1 _32061_inst ( .DIN1(______[0]), .DIN2(_32190), .Q(_32189) );
  nor2s1 _32062_inst ( .DIN1(_32191), .DIN2(_32192), .Q(_32190) );
  nor2s1 _32063_inst ( .DIN1(_32193), .DIN2(_26634), .Q(_32192) );
  nor2s1 _32064_inst ( .DIN1(_30676), .DIN2(_32072), .Q(_32193) );
  nor2s1 _32065_inst ( .DIN1(_26497), .DIN2(_53434), .Q(_32072) );
  hi1s1 _32066_inst ( .DIN(_32074), .Q(_30676) );
  nor2s1 _32067_inst ( .DIN1(_53433), .DIN2(_32194), .Q(_32191) );
  nor2s1 _32068_inst ( .DIN1(_53434), .DIN2(_32144), .Q(_32194) );
  nnd2s1 _32069_inst ( .DIN1(_53288), .DIN2(_32074), .Q(_32144) );
  nor2s1 _32070_inst ( .DIN1(_32195), .DIN2(_32022), .Q(_32187) );
  xnr2s1 _32071_inst ( .DIN1(_32150), .DIN2(_32196), .Q(_32195) );
  xnr2s1 _32072_inst ( .DIN1(_53432), .DIN2(_32151), .Q(_32196) );
  nnd2s1 _32073_inst ( .DIN1(_32197), .DIN2(_32198), .Q(_32151) );
  nnd2s1 _32074_inst ( .DIN1(_32199), .DIN2(_26478), .Q(_32198) );
  nnd2s1 _32075_inst ( .DIN1(_32200), .DIN2(_32201), .Q(_32199) );
  or2s1 _32076_inst ( .DIN1(_32201), .DIN2(_32200), .Q(_32197) );
  xor2s1 _32077_inst ( .DIN1(_32202), .DIN2(_32203), .Q(_32150) );
  xnr2s1 _32078_inst ( .DIN1(_30575), .DIN2(_32176), .Q(_32203) );
  xnr2s1 _32079_inst ( .DIN1(_32181), .DIN2(_26819), .Q(_32176) );
  nnd2s1 _32080_inst ( .DIN1(_32205), .DIN2(_32206), .Q(_32181) );
  nnd2s1 _32081_inst ( .DIN1(_26826), .DIN2(_32207), .Q(_32206) );
  xnr2s1 _32082_inst ( .DIN1(_29492), .DIN2(_32208), .Q(_32207) );
  or2s1 _32083_inst ( .DIN1(_32209), .DIN2(_414), .Q(_32208) );
  nnd2s1 _32084_inst ( .DIN1(_414), .DIN2(_32209), .Q(_32205) );
  xnr2s1 _32085_inst ( .DIN1(_32157), .DIN2(_32210), .Q(_30575) );
  xor2s1 _32086_inst ( .DIN1(_32159), .DIN2(_31843), .Q(_32210) );
  xor2s1 _32087_inst ( .DIN1(_32171), .DIN2(_32177), .Q(_31843) );
  xor2s1 _32088_inst ( .DIN1(_15553), .DIN2(_32211), .Q(_32177) );
  xor2s1 _32089_inst ( .DIN1(_32166), .DIN2(_32212), .Q(_32169) );
  xor2s1 _32090_inst ( .DIN1(_52990), .DIN2(_53461), .Q(_32212) );
  nnd2s1 _32091_inst ( .DIN1(_32213), .DIN2(_32214), .Q(_32166) );
  nnd2s1 _32092_inst ( .DIN1(_32215), .DIN2(_26314), .Q(_32214) );
  nnd2s1 _32093_inst ( .DIN1(_26291), .DIN2(_32216), .Q(_32215) );
  or2s1 _32094_inst ( .DIN1(_26291), .DIN2(_32216), .Q(_32213) );
  nnd2s1 _32095_inst ( .DIN1(_32217), .DIN2(_32218), .Q(_32171) );
  nnd2s1 _32096_inst ( .DIN1(_32219), .DIN2(_32220), .Q(_32218) );
  or2s1 _32097_inst ( .DIN1(_32221), .DIN2(_15555), .Q(_32220) );
  nnd2s1 _32098_inst ( .DIN1(_15555), .DIN2(_32221), .Q(_32217) );
  nnd2s1 _32099_inst ( .DIN1(_32222), .DIN2(_32223), .Q(_32159) );
  nnd2s1 _32100_inst ( .DIN1(_32224), .DIN2(_32225), .Q(_32223) );
  or2s1 _32101_inst ( .DIN1(_32226), .DIN2(_31883), .Q(_32225) );
  nnd2s1 _32102_inst ( .DIN1(_31883), .DIN2(_32226), .Q(_32222) );
  xnr2s1 _32103_inst ( .DIN1(_32174), .DIN2(_32227), .Q(_32202) );
  xor2s1 _32104_inst ( .DIN1(_32228), .DIN2(_29492), .Q(_32227) );
  and2s1 _32105_inst ( .DIN1(_32229), .DIN2(_32230), .Q(_32174) );
  nnd2s1 _32106_inst ( .DIN1(_32231), .DIN2(_32232), .Q(_32230) );
  nnd2s1 _32107_inst ( .DIN1(_30593), .DIN2(_32233), .Q(_32232) );
  or2s1 _32108_inst ( .DIN1(_32233), .DIN2(_30593), .Q(_32229) );
  hi1s1 _32109_inst ( .DIN(_30578), .Q(_30593) );
  hi1s1 _32110_inst ( .DIN(_28056), .Q(_28049) );
  nor2s1 _32111_inst ( .DIN1(_28056), .DIN2(_32234), .Q(_32184) );
  nor2s1 _32112_inst ( .DIN1(_32235), .DIN2(_27365), .Q(_32234) );
  xor2s1 _32113_inst ( .DIN1(_32236), .DIN2(_32237), .Q(_32235) );
  xor2s1 _32114_inst ( .DIN1(_53423), .DIN2(_53450), .Q(_32237) );
  nnd2s1 _32115_inst ( .DIN1(_53434), .DIN2(_53413), .Q(_32236) );
  nnd2s1 _32116_inst ( .DIN1(_32238), .DIN2(_27050), .Q(
        ______________________________106________) );
  nnd2s1 _32117_inst ( .DIN1(_32239), .DIN2(_27053), .Q(_27050) );
  nor2s1 _32118_inst ( .DIN1(_32240), .DIN2(_32241), .Q(_32238) );
  nor2s1 _32119_inst ( .DIN1(_27053), .DIN2(_32242), .Q(_32241) );
  nor2s1 _32120_inst ( .DIN1(_32243), .DIN2(_32244), .Q(_32242) );
  nor2s1 _32121_inst ( .DIN1(_32022), .DIN2(_32245), .Q(_32244) );
  xor2s1 _32122_inst ( .DIN1(_32200), .DIN2(_32246), .Q(_32245) );
  xor2s1 _32123_inst ( .DIN1(_26478), .DIN2(_32201), .Q(_32246) );
  nnd2s1 _32124_inst ( .DIN1(_32247), .DIN2(_32248), .Q(_32201) );
  nnd2s1 _32125_inst ( .DIN1(_52994), .DIN2(_32249), .Q(_32248) );
  or2s1 _32126_inst ( .DIN1(_32250), .DIN2(_32251), .Q(_32249) );
  nnd2s1 _32127_inst ( .DIN1(_32251), .DIN2(_32250), .Q(_32247) );
  xnr2s1 _32128_inst ( .DIN1(_32231), .DIN2(_32252), .Q(_32200) );
  xor2s1 _32129_inst ( .DIN1(_32233), .DIN2(_30578), .Q(_32252) );
  xor2s1 _32130_inst ( .DIN1(_32224), .DIN2(_32253), .Q(_30578) );
  xor2s1 _32131_inst ( .DIN1(_32226), .DIN2(_31883), .Q(_32253) );
  xor2s1 _32132_inst ( .DIN1(_32221), .DIN2(_26819), .Q(_31883) );
  xor2s1 _32133_inst ( .DIN1(_32216), .DIN2(_32254), .Q(_32219) );
  xor2s1 _32134_inst ( .DIN1(_53486), .DIN2(_53487), .Q(_32254) );
  nnd2s1 _32135_inst ( .DIN1(_32255), .DIN2(_32256), .Q(_32216) );
  nnd2s1 _32136_inst ( .DIN1(_52845), .DIN2(_32257), .Q(_32256) );
  nnd2s1 _32137_inst ( .DIN1(_53387), .DIN2(_32258), .Q(_32257) );
  or2s1 _32138_inst ( .DIN1(_32258), .DIN2(_53387), .Q(_32255) );
  nnd2s1 _32139_inst ( .DIN1(_32259), .DIN2(_32260), .Q(_32221) );
  nnd2s1 _32140_inst ( .DIN1(_414), .DIN2(_32261), .Q(_32260) );
  or2s1 _32141_inst ( .DIN1(_32262), .DIN2(_32211), .Q(_32261) );
  nnd2s1 _32142_inst ( .DIN1(_32211), .DIN2(_32262), .Q(_32259) );
  nnd2s1 _32143_inst ( .DIN1(_32263), .DIN2(_32264), .Q(_32226) );
  nnd2s1 _32144_inst ( .DIN1(_32265), .DIN2(_32266), .Q(_32264) );
  or2s1 _32145_inst ( .DIN1(_32267), .DIN2(_31940), .Q(_32266) );
  hi1s1 _32146_inst ( .DIN(_32268), .Q(_32265) );
  nnd2s1 _32147_inst ( .DIN1(_31940), .DIN2(_32267), .Q(_32263) );
  nnd2s1 _32148_inst ( .DIN1(_32269), .DIN2(_32270), .Q(_32233) );
  nnd2s1 _32149_inst ( .DIN1(_32271), .DIN2(_32272), .Q(_32270) );
  or2s1 _32150_inst ( .DIN1(_32273), .DIN2(_30622), .Q(_32272) );
  nnd2s1 _32151_inst ( .DIN1(_30622), .DIN2(_32273), .Q(_32269) );
  xnr2s1 _32152_inst ( .DIN1(_32209), .DIN2(_32274), .Q(_32231) );
  nnd2s1 _32153_inst ( .DIN1(_32275), .DIN2(_32276), .Q(_32209) );
  nnd2s1 _32154_inst ( .DIN1(_26206), .DIN2(_32277), .Q(_32276) );
  or2s1 _32155_inst ( .DIN1(_32278), .DIN2(_15555), .Q(_32277) );
  nnd2s1 _32156_inst ( .DIN1(_15555), .DIN2(_32278), .Q(_32275) );
  nor2s1 _32157_inst ( .DIN1(_32065), .DIN2(_32279), .Q(_32243) );
  nor2s1 _32158_inst ( .DIN1(_32280), .DIN2(_32281), .Q(_32279) );
  nnd2s1 _32159_inst ( .DIN1(______[30]), .DIN2(_32074), .Q(_32281) );
  xor2s1 _32160_inst ( .DIN1(_26493), .DIN2(_32282), .Q(_32280) );
  nnd2s1 _32161_inst ( .DIN1(_52996), .DIN2(_52997), .Q(_32282) );
  nor2s1 _32162_inst ( .DIN1(_27064), .DIN2(_32283), .Q(_32240) );
  nor2s1 _32163_inst ( .DIN1(_32284), .DIN2(_32285), .Q(_32283) );
  nor2s1 _32164_inst ( .DIN1(_26492), .DIN2(_30391), .Q(_32285) );
  nnd2s1 _32165_inst ( .DIN1(_52838), .DIN2(_52991), .Q(_30391) );
  nor2s1 _32166_inst ( .DIN1(_52838), .DIN2(_32286), .Q(_32284) );
  nor2s1 _32167_inst ( .DIN1(_26299), .DIN2(_26492), .Q(_32286) );
  nnd2s1 _32168_inst ( .DIN1(_32287), .DIN2(_32288), .Q(
        ______________________________105________) );
  nnd2s1 _32169_inst ( .DIN1(_32289), .DIN2(_28069), .Q(_32288) );
  nor2s1 _32170_inst ( .DIN1(_26261), .DIN2(_32290), .Q(_32289) );
  nnd2s1 _32171_inst ( .DIN1(______[6]), .DIN2(_28071), .Q(_32290) );
  nnd2s1 _32172_inst ( .DIN1(_32291), .DIN2(_28060), .Q(_32287) );
  hi1s1 _32173_inst ( .DIN(_28069), .Q(_28060) );
  nnd2s1 _32174_inst ( .DIN1(_32292), .DIN2(_28144), .Q(_28069) );
  nnd2s1 _32175_inst ( .DIN1(_32293), .DIN2(_32294), .Q(_32291) );
  nnd2s1 _32176_inst ( .DIN1(_32065), .DIN2(_32295), .Q(_32294) );
  xor2s1 _32177_inst ( .DIN1(_32296), .DIN2(_32297), .Q(_32295) );
  xnr2s1 _32178_inst ( .DIN1(_32250), .DIN2(_32251), .Q(_32297) );
  xnr2s1 _32179_inst ( .DIN1(_32271), .DIN2(_32298), .Q(_32251) );
  xor2s1 _32180_inst ( .DIN1(_32273), .DIN2(_30622), .Q(_32298) );
  xor2s1 _32181_inst ( .DIN1(_31940), .DIN2(_32299), .Q(_30622) );
  xor2s1 _32182_inst ( .DIN1(_32267), .DIN2(_32268), .Q(_32299) );
  nnd2s1 _32183_inst ( .DIN1(_32300), .DIN2(_32301), .Q(_32267) );
  nnd2s1 _32184_inst ( .DIN1(_32302), .DIN2(_32303), .Q(_32301) );
  or2s1 _32185_inst ( .DIN1(_32304), .DIN2(_31987), .Q(_32303) );
  nnd2s1 _32186_inst ( .DIN1(_31987), .DIN2(_32304), .Q(_32300) );
  xor2s1 _32187_inst ( .DIN1(_32262), .DIN2(_32274), .Q(_31940) );
  xor2s1 _32188_inst ( .DIN1(_32211), .DIN2(_29580), .Q(_32274) );
  xor2s1 _32189_inst ( .DIN1(_32258), .DIN2(_32305), .Q(_408) );
  xor2s1 _32190_inst ( .DIN1(_52845), .DIN2(_53387), .Q(_32305) );
  nnd2s1 _32191_inst ( .DIN1(_32306), .DIN2(_32307), .Q(_32258) );
  nnd2s1 _32192_inst ( .DIN1(_32308), .DIN2(_26742), .Q(_32307) );
  nnd2s1 _32193_inst ( .DIN1(_26464), .DIN2(_32309), .Q(_32308) );
  or2s1 _32194_inst ( .DIN1(_26464), .DIN2(_32309), .Q(_32306) );
  nnd2s1 _32195_inst ( .DIN1(_32310), .DIN2(_32311), .Q(_32262) );
  nnd2s1 _32196_inst ( .DIN1(_26206), .DIN2(_32312), .Q(_32311) );
  or2s1 _32197_inst ( .DIN1(_32313), .DIN2(_32314), .Q(_32312) );
  nnd2s1 _32198_inst ( .DIN1(_32314), .DIN2(_32313), .Q(_32310) );
  nnd2s1 _32199_inst ( .DIN1(_32315), .DIN2(_32316), .Q(_32273) );
  nnd2s1 _32200_inst ( .DIN1(_32317), .DIN2(_32318), .Q(_32316) );
  or2s1 _32201_inst ( .DIN1(_32319), .DIN2(_30619), .Q(_32318) );
  nnd2s1 _32202_inst ( .DIN1(_30619), .DIN2(_32319), .Q(_32315) );
  xor2s1 _32203_inst ( .DIN1(_32278), .DIN2(_32320), .Q(_32271) );
  nnd2s1 _32204_inst ( .DIN1(_32321), .DIN2(_32322), .Q(_32278) );
  nnd2s1 _32205_inst ( .DIN1(_26829), .DIN2(_32323), .Q(_32322) );
  or2s1 _32206_inst ( .DIN1(_32324), .DIN2(_414), .Q(_32323) );
  nnd2s1 _32207_inst ( .DIN1(_414), .DIN2(_32324), .Q(_32321) );
  nnd2s1 _32208_inst ( .DIN1(_32325), .DIN2(_32326), .Q(_32250) );
  nnd2s1 _32209_inst ( .DIN1(_52995), .DIN2(_32327), .Q(_32326) );
  or2s1 _32210_inst ( .DIN1(_32328), .DIN2(_32329), .Q(_32327) );
  nnd2s1 _32211_inst ( .DIN1(_32329), .DIN2(_32328), .Q(_32325) );
  xor2s1 _32212_inst ( .DIN1(_52994), .DIN2(_32330), .Q(_32296) );
  hi1s1 _32213_inst ( .DIN(_32022), .Q(_32065) );
  nnd2s1 _32214_inst ( .DIN1(_32331), .DIN2(_32022), .Q(_32293) );
  nnd2s1 _32215_inst ( .DIN1(_32332), .DIN2(_32333), .Q(_32022) );
  nor2s1 _32216_inst ( .DIN1(_31367), .DIN2(_30375), .Q(_32332) );
  nor2s1 _32217_inst ( .DIN1(_27774), .DIN2(_32334), .Q(_32331) );
  nnd2s1 _32218_inst ( .DIN1(_32335), .DIN2(_32074), .Q(_32334) );
  nnd2s1 _32219_inst ( .DIN1(_32336), .DIN2(_32337), .Q(_32074) );
  nor2s1 _32220_inst ( .DIN1(_30832), .DIN2(_32338), .Q(_32337) );
  nnd2s1 _32221_inst ( .DIN1(_32339), .DIN2(_32340), .Q(_32338) );
  hi1s1 _32222_inst ( .DIN(_32341), .Q(_30832) );
  nor2s1 _32223_inst ( .DIN1(_30526), .DIN2(_30369), .Q(_32336) );
  xor2s1 _32224_inst ( .DIN1(_52993), .DIN2(_52996), .Q(_32335) );
  nor2s1 _32225_inst ( .DIN1(_27500), .DIN2(_32342), .Q(
        ______________________________104________) );
  nnd2s1 _32226_inst ( .DIN1(_32343), .DIN2(_32344), .Q(_32342) );
  nnd2s1 _32227_inst ( .DIN1(_32345), .DIN2(_28660), .Q(_32344) );
  nor2s1 _32228_inst ( .DIN1(_26391), .DIN2(_32346), .Q(_32345) );
  nnd2s1 _32229_inst ( .DIN1(______[4]), .DIN2(_29885), .Q(_32346) );
  nnd2s1 _32230_inst ( .DIN1(_32347), .DIN2(_32348), .Q(_32343) );
  xor2s1 _32231_inst ( .DIN1(_32329), .DIN2(_32349), .Q(_32347) );
  xnr2s1 _32232_inst ( .DIN1(_52995), .DIN2(_32328), .Q(_32349) );
  nnd2s1 _32233_inst ( .DIN1(_32350), .DIN2(_32351), .Q(_32328) );
  nnd2s1 _32234_inst ( .DIN1(_32352), .DIN2(_26405), .Q(_32351) );
  nnd2s1 _32235_inst ( .DIN1(_32353), .DIN2(_32354), .Q(_32352) );
  or2s1 _32236_inst ( .DIN1(_32354), .DIN2(_32353), .Q(_32350) );
  xnr2s1 _32237_inst ( .DIN1(_32317), .DIN2(_32355), .Q(_32329) );
  xor2s1 _32238_inst ( .DIN1(_32319), .DIN2(_30619), .Q(_32355) );
  xor2s1 _32239_inst ( .DIN1(_31987), .DIN2(_32356), .Q(_30619) );
  xor2s1 _32240_inst ( .DIN1(_32304), .DIN2(_32357), .Q(_32356) );
  nnd2s1 _32241_inst ( .DIN1(_32358), .DIN2(_32359), .Q(_32304) );
  nnd2s1 _32242_inst ( .DIN1(_32360), .DIN2(_32361), .Q(_32359) );
  xor2s1 _32243_inst ( .DIN1(_32362), .DIN2(_32363), .Q(_32361) );
  xor2s1 _32244_inst ( .DIN1(_32313), .DIN2(_32320), .Q(_31987) );
  xor2s1 _32245_inst ( .DIN1(_26206), .DIN2(_15555), .Q(_32320) );
  hi1s1 _32246_inst ( .DIN(_32314), .Q(_15555) );
  xor2s1 _32247_inst ( .DIN1(_32309), .DIN2(_32364), .Q(_32314) );
  xor2s1 _32248_inst ( .DIN1(_53488), .DIN2(_53489), .Q(_32364) );
  nnd2s1 _32249_inst ( .DIN1(_32365), .DIN2(_32366), .Q(_32309) );
  nnd2s1 _32250_inst ( .DIN1(_32367), .DIN2(_26758), .Q(_32366) );
  nnd2s1 _32251_inst ( .DIN1(_26721), .DIN2(_32368), .Q(_32367) );
  or2s1 _32252_inst ( .DIN1(_26721), .DIN2(_32368), .Q(_32365) );
  nnd2s1 _32253_inst ( .DIN1(_32369), .DIN2(_32370), .Q(_32313) );
  nnd2s1 _32254_inst ( .DIN1(_26829), .DIN2(_32371), .Q(_32370) );
  or2s1 _32255_inst ( .DIN1(_32372), .DIN2(_29580), .Q(_32371) );
  nnd2s1 _32256_inst ( .DIN1(_29580), .DIN2(_32372), .Q(_32369) );
  nnd2s1 _32257_inst ( .DIN1(_32373), .DIN2(_32374), .Q(_32319) );
  nnd2s1 _32258_inst ( .DIN1(_32375), .DIN2(_32376), .Q(_32374) );
  nnd2s1 _32259_inst ( .DIN1(_32377), .DIN2(_30659), .Q(_32375) );
  xor2s1 _32260_inst ( .DIN1(_32228), .DIN2(_32378), .Q(_32373) );
  nor2s1 _32261_inst ( .DIN1(_30659), .DIN2(_32377), .Q(_32378) );
  hi1s1 _32262_inst ( .DIN(_31925), .Q(_32228) );
  xor2s1 _32263_inst ( .DIN1(_32379), .DIN2(_32324), .Q(_32317) );
  nnd2s1 _32264_inst ( .DIN1(_32380), .DIN2(_32381), .Q(_32324) );
  nnd2s1 _32265_inst ( .DIN1(_26206), .DIN2(_32382), .Q(_32381) );
  or2s1 _32266_inst ( .DIN1(_32383), .DIN2(_424), .Q(_32382) );
  nnd2s1 _32267_inst ( .DIN1(_424), .DIN2(_32383), .Q(_32380) );
  nnd2s1 _32268_inst ( .DIN1(_32384), .DIN2(_30601), .Q(
        ______________________________103________) );
  nor2s1 _32269_inst ( .DIN1(_32385), .DIN2(_32386), .Q(_32384) );
  nor2s1 _32270_inst ( .DIN1(_32387), .DIN2(_27392), .Q(_32386) );
  nor2s1 _32271_inst ( .DIN1(_32388), .DIN2(_32389), .Q(_32387) );
  nor2s1 _32272_inst ( .DIN1(_32390), .DIN2(_28660), .Q(_32389) );
  xor2s1 _32273_inst ( .DIN1(_32353), .DIN2(_32391), .Q(_32390) );
  xor2s1 _32274_inst ( .DIN1(_26405), .DIN2(_32354), .Q(_32391) );
  nnd2s1 _32275_inst ( .DIN1(_32392), .DIN2(_32393), .Q(_32354) );
  nnd2s1 _32276_inst ( .DIN1(_52998), .DIN2(_32394), .Q(_32393) );
  nnd2s1 _32277_inst ( .DIN1(_32395), .DIN2(_32396), .Q(_32394) );
  or2s1 _32278_inst ( .DIN1(_32396), .DIN2(_32395), .Q(_32392) );
  xnr2s1 _32279_inst ( .DIN1(_30659), .DIN2(_32397), .Q(_32353) );
  xnr2s1 _32280_inst ( .DIN1(_32376), .DIN2(_32377), .Q(_32397) );
  xnr2s1 _32281_inst ( .DIN1(_32383), .DIN2(_32398), .Q(_32377) );
  nnd2s1 _32282_inst ( .DIN1(_32399), .DIN2(_32400), .Q(_32383) );
  nnd2s1 _32283_inst ( .DIN1(_15560), .DIN2(_32401), .Q(_32400) );
  or2s1 _32284_inst ( .DIN1(_32402), .DIN2(_26829), .Q(_32401) );
  nnd2s1 _32285_inst ( .DIN1(_26829), .DIN2(_32402), .Q(_32399) );
  nnd2s1 _32286_inst ( .DIN1(_32403), .DIN2(_32404), .Q(_32376) );
  nnd2s1 _32287_inst ( .DIN1(_32405), .DIN2(_32406), .Q(_32404) );
  nnd2s1 _32288_inst ( .DIN1(_32407), .DIN2(_30700), .Q(_32406) );
  or2s1 _32289_inst ( .DIN1(_30700), .DIN2(_32407), .Q(_32403) );
  nnd2s1 _32290_inst ( .DIN1(_32408), .DIN2(_32409), .Q(_30659) );
  nnd2s1 _32291_inst ( .DIN1(_32360), .DIN2(_32410), .Q(_32409) );
  nnd2s1 _32292_inst ( .DIN1(_32363), .DIN2(_32358), .Q(_32410) );
  nnd2s1 _32293_inst ( .DIN1(_32064), .DIN2(_32411), .Q(_32358) );
  or2s1 _32294_inst ( .DIN1(_32411), .DIN2(_32064), .Q(_32363) );
  nnd2s1 _32295_inst ( .DIN1(_32412), .DIN2(_32413), .Q(_32408) );
  xor2s1 _32296_inst ( .DIN1(_32411), .DIN2(_32064), .Q(_32412) );
  xor2s1 _32297_inst ( .DIN1(_32372), .DIN2(_32379), .Q(_32064) );
  xnr2s1 _32298_inst ( .DIN1(_420), .DIN2(_29580), .Q(_32379) );
  xor2s1 _32299_inst ( .DIN1(_32368), .DIN2(_32414), .Q(_414) );
  xor2s1 _32300_inst ( .DIN1(_53490), .DIN2(_53491), .Q(_32414) );
  nnd2s1 _32301_inst ( .DIN1(_32415), .DIN2(_32416), .Q(_32368) );
  nnd2s1 _32302_inst ( .DIN1(_52847), .DIN2(_32417), .Q(_32416) );
  nnd2s1 _32303_inst ( .DIN1(_52999), .DIN2(_32418), .Q(_32417) );
  or2s1 _32304_inst ( .DIN1(_32418), .DIN2(_52999), .Q(_32415) );
  nnd2s1 _32305_inst ( .DIN1(_32419), .DIN2(_32420), .Q(_32372) );
  nnd2s1 _32306_inst ( .DIN1(_32421), .DIN2(_424), .Q(_32420) );
  xor2s1 _32307_inst ( .DIN1(_32422), .DIN2(_2064), .Q(_32421) );
  nnd2s1 _32308_inst ( .DIN1(_32423), .DIN2(_26206), .Q(_32422) );
  hi1s1 _32309_inst ( .DIN(_29581), .Q(_26206) );
  nnd2s1 _32310_inst ( .DIN1(_32424), .DIN2(_29581), .Q(_32419) );
  hi1s1 _32311_inst ( .DIN(_32423), .Q(_32424) );
  nnd2s1 _32312_inst ( .DIN1(_32425), .DIN2(_32426), .Q(_32411) );
  xor2s1 _32313_inst ( .DIN1(_32427), .DIN2(_32428), .Q(_32425) );
  nnd2s1 _32314_inst ( .DIN1(_32429), .DIN2(_32430), .Q(_32428) );
  nor2s1 _32315_inst ( .DIN1(_28652), .DIN2(_32431), .Q(_32388) );
  nnd2s1 _32316_inst ( .DIN1(______[24]), .DIN2(_32432), .Q(_32431) );
  xor2s1 _32317_inst ( .DIN1(_52996), .DIN2(_52997), .Q(_32432) );
  nnd2s1 _32318_inst ( .DIN1(_29885), .DIN2(_28660), .Q(_28652) );
  nor2s1 _32319_inst ( .DIN1(_27397), .DIN2(_32433), .Q(_32385) );
  nor2s1 _32320_inst ( .DIN1(_32434), .DIN2(_26773), .Q(_32433) );
  xor2s1 _32321_inst ( .DIN1(_26513), .DIN2(_53441), .Q(_32434) );
  nnd2s1 _32322_inst ( .DIN1(_32435), .DIN2(_32436), .Q(
        ______________________________102________) );
  nnd2s1 _32323_inst ( .DIN1(_32437), .DIN2(_27903), .Q(_32436) );
  nor2s1 _32324_inst ( .DIN1(_32438), .DIN2(_27082), .Q(_32437) );
  xnr2s1 _32325_inst ( .DIN1(_53000), .DIN2(_52979), .Q(_32438) );
  nnd2s1 _32326_inst ( .DIN1(_32439), .DIN2(_27298), .Q(_32435) );
  nor2s1 _32327_inst ( .DIN1(_32440), .DIN2(_32441), .Q(_32439) );
  nor2s1 _32328_inst ( .DIN1(_28660), .DIN2(_32442), .Q(_32441) );
  xnr2s1 _32329_inst ( .DIN1(_32395), .DIN2(_32443), .Q(_32442) );
  xnr2s1 _32330_inst ( .DIN1(_52998), .DIN2(_32396), .Q(_32443) );
  nnd2s1 _32331_inst ( .DIN1(_32444), .DIN2(_32445), .Q(_32396) );
  nnd2s1 _32332_inst ( .DIN1(_53001), .DIN2(_32446), .Q(_32445) );
  nnd2s1 _32333_inst ( .DIN1(_32447), .DIN2(_32448), .Q(_32446) );
  or2s1 _32334_inst ( .DIN1(_32448), .DIN2(_32447), .Q(_32444) );
  xnr2s1 _32335_inst ( .DIN1(_30700), .DIN2(_32449), .Q(_32395) );
  xor2s1 _32336_inst ( .DIN1(_32407), .DIN2(_32405), .Q(_32449) );
  xnr2s1 _32337_inst ( .DIN1(_32402), .DIN2(_32450), .Q(_32405) );
  nnd2s1 _32338_inst ( .DIN1(_32451), .DIN2(_32452), .Q(_32402) );
  nnd2s1 _32339_inst ( .DIN1(_32453), .DIN2(_15561), .Q(_32452) );
  xor2s1 _32340_inst ( .DIN1(_29544), .DIN2(_32454), .Q(_32453) );
  or2s1 _32341_inst ( .DIN1(_32455), .DIN2(_424), .Q(_32454) );
  nnd2s1 _32342_inst ( .DIN1(_424), .DIN2(_32455), .Q(_32451) );
  and2s1 _32343_inst ( .DIN1(_32456), .DIN2(_32457), .Q(_32407) );
  nnd2s1 _32344_inst ( .DIN1(_32458), .DIN2(_32459), .Q(_32457) );
  nnd2s1 _32345_inst ( .DIN1(_30713), .DIN2(_32460), .Q(_32459) );
  or2s1 _32346_inst ( .DIN1(_32460), .DIN2(_30713), .Q(_32456) );
  nnd2s1 _32347_inst ( .DIN1(_32461), .DIN2(_32462), .Q(_30700) );
  nnd2s1 _32348_inst ( .DIN1(_32429), .DIN2(_32463), .Q(_32462) );
  nnd2s1 _32349_inst ( .DIN1(_32430), .DIN2(_32426), .Q(_32463) );
  nnd2s1 _32350_inst ( .DIN1(_32161), .DIN2(_32464), .Q(_32426) );
  or2s1 _32351_inst ( .DIN1(_32464), .DIN2(_32161), .Q(_32430) );
  nnd2s1 _32352_inst ( .DIN1(_32465), .DIN2(_32466), .Q(_32461) );
  xor2s1 _32353_inst ( .DIN1(_32464), .DIN2(_32161), .Q(_32465) );
  hi1s1 _32354_inst ( .DIN(_32119), .Q(_32161) );
  xor2s1 _32355_inst ( .DIN1(_32423), .DIN2(_32398), .Q(_32119) );
  xor2s1 _32356_inst ( .DIN1(_32467), .DIN2(_29581), .Q(_32398) );
  xor2s1 _32357_inst ( .DIN1(_32418), .DIN2(_32468), .Q(_29581) );
  xor2s1 _32358_inst ( .DIN1(_52847), .DIN2(_52999), .Q(_32468) );
  nnd2s1 _32359_inst ( .DIN1(_32469), .DIN2(_32470), .Q(_32418) );
  nnd2s1 _32360_inst ( .DIN1(_32471), .DIN2(_26749), .Q(_32470) );
  nnd2s1 _32361_inst ( .DIN1(_26611), .DIN2(_32472), .Q(_32471) );
  or2s1 _32362_inst ( .DIN1(_26611), .DIN2(_32472), .Q(_32469) );
  xor2s1 _32363_inst ( .DIN1(_31569), .DIN2(_32473), .Q(_32467) );
  xor2s1 _32364_inst ( .DIN1(_32474), .DIN2(_31269), .Q(_32423) );
  nnd2s1 _32365_inst ( .DIN1(_32475), .DIN2(_32476), .Q(_32474) );
  nnd2s1 _32366_inst ( .DIN1(_15560), .DIN2(_32477), .Q(_32476) );
  or2s1 _32367_inst ( .DIN1(_32478), .DIN2(_32479), .Q(_32477) );
  nnd2s1 _32368_inst ( .DIN1(_32478), .DIN2(_32479), .Q(_32475) );
  hi1s1 _32369_inst ( .DIN(_420), .Q(_32479) );
  nnd2s1 _32370_inst ( .DIN1(_32480), .DIN2(_32481), .Q(_32464) );
  nnd2s1 _32371_inst ( .DIN1(_32482), .DIN2(_32483), .Q(_32481) );
  or2s1 _32372_inst ( .DIN1(_32484), .DIN2(_32485), .Q(_32483) );
  nnd2s1 _32373_inst ( .DIN1(_32485), .DIN2(_32484), .Q(_32480) );
  nor2s1 _32374_inst ( .DIN1(_32348), .DIN2(_32486), .Q(_32440) );
  nor2s1 _32375_inst ( .DIN1(_27241), .DIN2(_32487), .Q(_32486) );
  nnd2s1 _32376_inst ( .DIN1(_32488), .DIN2(_32489), .Q(_32487) );
  xor2s1 _32377_inst ( .DIN1(_32490), .DIN2(_32491), .Q(_32488) );
  nor2s1 _32378_inst ( .DIN1(_53004), .DIN2(_53003), .Q(_32490) );
  nnd2s1 _32379_inst ( .DIN1(_32492), .DIN2(_32493), .Q(
        ______________________________101________) );
  nnd2s1 _32380_inst ( .DIN1(_32494), .DIN2(_32495), .Q(_32493) );
  hi1s1 _32381_inst ( .DIN(_32496), .Q(_32495) );
  xnr2s1 _32382_inst ( .DIN1(_32447), .DIN2(_32497), .Q(_32494) );
  xnr2s1 _32383_inst ( .DIN1(_53001), .DIN2(_32448), .Q(_32497) );
  nnd2s1 _32384_inst ( .DIN1(_32498), .DIN2(_32499), .Q(_32448) );
  nnd2s1 _32385_inst ( .DIN1(_32500), .DIN2(_26744), .Q(_32499) );
  nnd2s1 _32386_inst ( .DIN1(_32501), .DIN2(_32502), .Q(_32500) );
  nnd2s1 _32387_inst ( .DIN1(_32503), .DIN2(_32504), .Q(_32498) );
  hi1s1 _32388_inst ( .DIN(_32501), .Q(_32504) );
  xnr2s1 _32389_inst ( .DIN1(_32505), .DIN2(_32458), .Q(_32447) );
  xnr2s1 _32390_inst ( .DIN1(_32506), .DIN2(_32455), .Q(_32458) );
  nnd2s1 _32391_inst ( .DIN1(_32507), .DIN2(_32508), .Q(_32455) );
  nnd2s1 _32392_inst ( .DIN1(_15560), .DIN2(_32509), .Q(_32508) );
  or2s1 _32393_inst ( .DIN1(_32510), .DIN2(_433), .Q(_32509) );
  nnd2s1 _32394_inst ( .DIN1(_433), .DIN2(_32510), .Q(_32507) );
  xnr2s1 _32395_inst ( .DIN1(_32460), .DIN2(_30713), .Q(_32505) );
  xnr2s1 _32396_inst ( .DIN1(_32157), .DIN2(_32511), .Q(_30713) );
  xor2s1 _32397_inst ( .DIN1(_32484), .DIN2(_32482), .Q(_32511) );
  nnd2s1 _32398_inst ( .DIN1(_32512), .DIN2(_32513), .Q(_32484) );
  nnd2s1 _32399_inst ( .DIN1(_32514), .DIN2(_32515), .Q(_32513) );
  or2s1 _32400_inst ( .DIN1(_32516), .DIN2(_32517), .Q(_32515) );
  hi1s1 _32401_inst ( .DIN(_32518), .Q(_32514) );
  xor2s1 _32402_inst ( .DIN1(_31585), .DIN2(_32519), .Q(_32512) );
  nnd2s1 _32403_inst ( .DIN1(_32516), .DIN2(_32517), .Q(_32519) );
  hi1s1 _32404_inst ( .DIN(_32224), .Q(_32516) );
  hi1s1 _32405_inst ( .DIN(_32485), .Q(_32157) );
  xnr2s1 _32406_inst ( .DIN1(_32450), .DIN2(_32478), .Q(_32485) );
  xnr2s1 _32407_inst ( .DIN1(_32520), .DIN2(_27093), .Q(_32478) );
  nnd2s1 _32408_inst ( .DIN1(_32521), .DIN2(_32522), .Q(_32520) );
  nnd2s1 _32409_inst ( .DIN1(_15561), .DIN2(_32523), .Q(_32522) );
  or2s1 _32410_inst ( .DIN1(_32524), .DIN2(_32473), .Q(_32523) );
  nnd2s1 _32411_inst ( .DIN1(_32473), .DIN2(_32524), .Q(_32521) );
  xor2s1 _32412_inst ( .DIN1(_32525), .DIN2(_420), .Q(_32450) );
  xor2s1 _32413_inst ( .DIN1(_32472), .DIN2(_32526), .Q(_420) );
  xor2s1 _32414_inst ( .DIN1(_53492), .DIN2(_53493), .Q(_32526) );
  nnd2s1 _32415_inst ( .DIN1(_32527), .DIN2(_32528), .Q(_32472) );
  nnd2s1 _32416_inst ( .DIN1(_32529), .DIN2(_26755), .Q(_32528) );
  nnd2s1 _32417_inst ( .DIN1(_53494), .DIN2(_32530), .Q(_32529) );
  or2s1 _32418_inst ( .DIN1(_32530), .DIN2(_53494), .Q(_32527) );
  nnd2s1 _32419_inst ( .DIN1(_32531), .DIN2(_32532), .Q(_32460) );
  nnd2s1 _32420_inst ( .DIN1(_32533), .DIN2(_32534), .Q(_32532) );
  nnd2s1 _32421_inst ( .DIN1(_30716), .DIN2(_32535), .Q(_32534) );
  or2s1 _32422_inst ( .DIN1(_32535), .DIN2(_30716), .Q(_32531) );
  hi1s1 _32423_inst ( .DIN(_30738), .Q(_30716) );
  nor2s1 _32424_inst ( .DIN1(_32536), .DIN2(_32537), .Q(_32492) );
  nor2s1 _32425_inst ( .DIN1(_31708), .DIN2(_32538), .Q(_32537) );
  xor2s1 _32426_inst ( .DIN1(_53002), .DIN2(_28690), .Q(_32538) );
  and2s1 _32427_inst ( .DIN1(_53005), .DIN2(_53003), .Q(_28690) );
  nor2s1 _32428_inst ( .DIN1(_32539), .DIN2(_32540), .Q(_32536) );
  and2s1 _32429_inst ( .DIN1(_29885), .DIN2(_52946), .Q(_32539) );
  nnd2s1 _32430_inst ( .DIN1(_32541), .DIN2(_32542), .Q(
        ______________________________100________) );
  nnd2s1 _32431_inst ( .DIN1(_32543), .DIN2(_32544), .Q(_32542) );
  nnd2s1 _32432_inst ( .DIN1(_32545), .DIN2(_29885), .Q(_32544) );
  xor2s1 _32433_inst ( .DIN1(_31842), .DIN2(_32489), .Q(_29885) );
  nnd2s1 _32434_inst ( .DIN1(_32546), .DIN2(_30833), .Q(_32489) );
  nor2s1 _32435_inst ( .DIN1(_31964), .DIN2(_31699), .Q(_30833) );
  nor2s1 _32436_inst ( .DIN1(_30524), .DIN2(_31538), .Q(_32546) );
  nnd2s1 _32437_inst ( .DIN1(_32547), .DIN2(_32341), .Q(_31538) );
  nor2s1 _32438_inst ( .DIN1(_30831), .DIN2(_31367), .Q(_32547) );
  hi1s1 _32439_inst ( .DIN(_32339), .Q(_31367) );
  hi1s1 _32440_inst ( .DIN(_31702), .Q(_30524) );
  xor2s1 _32441_inst ( .DIN1(_53004), .DIN2(_32548), .Q(_32545) );
  hi1s1 _32442_inst ( .DIN(_32540), .Q(_32543) );
  nnd2s1 _32443_inst ( .DIN1(_31554), .DIN2(_28660), .Q(_32540) );
  nor2s1 _32444_inst ( .DIN1(_32549), .DIN2(_32550), .Q(_32541) );
  nor2s1 _32445_inst ( .DIN1(_32496), .DIN2(_32551), .Q(_32550) );
  xor2s1 _32446_inst ( .DIN1(_32552), .DIN2(_32553), .Q(_32551) );
  xor2s1 _32447_inst ( .DIN1(_32501), .DIN2(_32503), .Q(_32553) );
  hi1s1 _32448_inst ( .DIN(_32502), .Q(_32503) );
  nnd2s1 _32449_inst ( .DIN1(_32554), .DIN2(_32555), .Q(_32502) );
  nnd2s1 _32450_inst ( .DIN1(_32556), .DIN2(_26537), .Q(_32555) );
  or2s1 _32451_inst ( .DIN1(_28662), .DIN2(_28664), .Q(_32556) );
  nnd2s1 _32452_inst ( .DIN1(_28662), .DIN2(_28664), .Q(_32554) );
  nnd2s1 _32453_inst ( .DIN1(_32557), .DIN2(_32558), .Q(_28664) );
  nnd2s1 _32454_inst ( .DIN1(_32559), .DIN2(_26732), .Q(_32558) );
  nnd2s1 _32455_inst ( .DIN1(_28699), .DIN2(_28679), .Q(_32559) );
  or2s1 _32456_inst ( .DIN1(_28679), .DIN2(_28699), .Q(_32557) );
  nor2s1 _32457_inst ( .DIN1(_26359), .DIN2(_28700), .Q(_28699) );
  xor2s1 _32458_inst ( .DIN1(_32560), .DIN2(_32561), .Q(_28700) );
  xor2s1 _32459_inst ( .DIN1(_32562), .DIN2(_30811), .Q(_32560) );
  hi1s1 _32460_inst ( .DIN(_30816), .Q(_30811) );
  xor2s1 _32461_inst ( .DIN1(_32563), .DIN2(_32564), .Q(_28679) );
  xor2s1 _32462_inst ( .DIN1(_32565), .DIN2(_30794), .Q(_32564) );
  xnr2s1 _32463_inst ( .DIN1(_32566), .DIN2(_32567), .Q(_28662) );
  xor2s1 _32464_inst ( .DIN1(_32568), .DIN2(_30754), .Q(_32567) );
  xnr2s1 _32465_inst ( .DIN1(_32533), .DIN2(_32569), .Q(_32501) );
  xor2s1 _32466_inst ( .DIN1(_32535), .DIN2(_30738), .Q(_32569) );
  xor2s1 _32467_inst ( .DIN1(_32224), .DIN2(_32570), .Q(_30738) );
  xor2s1 _32468_inst ( .DIN1(_32517), .DIN2(_32518), .Q(_32570) );
  nnd2s1 _32469_inst ( .DIN1(_32571), .DIN2(_32572), .Q(_32517) );
  nnd2s1 _32470_inst ( .DIN1(_32573), .DIN2(_32574), .Q(_32572) );
  or2s1 _32471_inst ( .DIN1(_32575), .DIN2(_32268), .Q(_32574) );
  nnd2s1 _32472_inst ( .DIN1(_32268), .DIN2(_32575), .Q(_32571) );
  xor2s1 _32473_inst ( .DIN1(_32524), .DIN2(_32506), .Q(_32224) );
  xor2s1 _32474_inst ( .DIN1(_15561), .DIN2(_32473), .Q(_32506) );
  hi1s1 _32475_inst ( .DIN(_424), .Q(_32473) );
  xor2s1 _32476_inst ( .DIN1(_32530), .DIN2(_32576), .Q(_424) );
  xor2s1 _32477_inst ( .DIN1(_52843), .DIN2(_53494), .Q(_32576) );
  nnd2s1 _32478_inst ( .DIN1(_32577), .DIN2(_32578), .Q(_32530) );
  nnd2s1 _32479_inst ( .DIN1(_52848), .DIN2(_32579), .Q(_32578) );
  or2s1 _32480_inst ( .DIN1(_26577), .DIN2(_32580), .Q(_32579) );
  nnd2s1 _32481_inst ( .DIN1(_32580), .DIN2(_26577), .Q(_32577) );
  nnd2s1 _32482_inst ( .DIN1(_32581), .DIN2(_32582), .Q(_32524) );
  nnd2s1 _32483_inst ( .DIN1(_32525), .DIN2(_32583), .Q(_32582) );
  or2s1 _32484_inst ( .DIN1(_32584), .DIN2(_433), .Q(_32583) );
  nnd2s1 _32485_inst ( .DIN1(_433), .DIN2(_32584), .Q(_32581) );
  nnd2s1 _32486_inst ( .DIN1(_32585), .DIN2(_32586), .Q(_32535) );
  nnd2s1 _32487_inst ( .DIN1(_32566), .DIN2(_32587), .Q(_32586) );
  or2s1 _32488_inst ( .DIN1(_32568), .DIN2(_30754), .Q(_32587) );
  xor2s1 _32489_inst ( .DIN1(_32588), .DIN2(_32589), .Q(_32566) );
  nnd2s1 _32490_inst ( .DIN1(_30754), .DIN2(_32568), .Q(_32585) );
  nnd2s1 _32491_inst ( .DIN1(_32590), .DIN2(_32591), .Q(_32568) );
  nnd2s1 _32492_inst ( .DIN1(_32563), .DIN2(_32592), .Q(_32591) );
  or2s1 _32493_inst ( .DIN1(_32565), .DIN2(_30794), .Q(_32592) );
  xnr2s1 _32494_inst ( .DIN1(_32593), .DIN2(_32594), .Q(_32563) );
  nnd2s1 _32495_inst ( .DIN1(_30794), .DIN2(_32565), .Q(_32590) );
  nnd2s1 _32496_inst ( .DIN1(_32595), .DIN2(_32596), .Q(_32565) );
  nnd2s1 _32497_inst ( .DIN1(_32597), .DIN2(_30816), .Q(_32596) );
  nnd2s1 _32498_inst ( .DIN1(_32598), .DIN2(_32599), .Q(_30816) );
  nnd2s1 _32499_inst ( .DIN1(_32600), .DIN2(_32601), .Q(_32599) );
  nor2s1 _32500_inst ( .DIN1(_32602), .DIN2(_32603), .Q(_32598) );
  nor2s1 _32501_inst ( .DIN1(_32360), .DIN2(_32604), .Q(_32603) );
  xor2s1 _32502_inst ( .DIN1(_32605), .DIN2(_32601), .Q(_32604) );
  nor2s1 _32503_inst ( .DIN1(_32413), .DIN2(_32606), .Q(_32602) );
  nnd2s1 _32504_inst ( .DIN1(_32605), .DIN2(_32607), .Q(_32606) );
  or2s1 _32505_inst ( .DIN1(_32562), .DIN2(_32561), .Q(_32597) );
  nnd2s1 _32506_inst ( .DIN1(_32561), .DIN2(_32562), .Q(_32595) );
  nnd2s1 _32507_inst ( .DIN1(_32608), .DIN2(_32609), .Q(_32562) );
  nnd2s1 _32508_inst ( .DIN1(_32610), .DIN2(_30814), .Q(_32609) );
  xor2s1 _32509_inst ( .DIN1(_32611), .DIN2(_32612), .Q(_32608) );
  nnd2s1 _32510_inst ( .DIN1(_32613), .DIN2(_32614), .Q(_32611) );
  xnr2s1 _32511_inst ( .DIN1(_32615), .DIN2(_32616), .Q(_32614) );
  or2s1 _32512_inst ( .DIN1(_32617), .DIN2(_30841), .Q(_32616) );
  nor2s1 _32513_inst ( .DIN1(_32618), .DIN2(_32619), .Q(_32613) );
  nor2s1 _32514_inst ( .DIN1(_32617), .DIN2(_32620), .Q(_32619) );
  nnd2s1 _32515_inst ( .DIN1(_32621), .DIN2(_32622), .Q(_32617) );
  nnd2s1 _32516_inst ( .DIN1(_30842), .DIN2(_32623), .Q(_32622) );
  nnd2s1 _32517_inst ( .DIN1(_32624), .DIN2(_32625), .Q(_32623) );
  xor2s1 _32518_inst ( .DIN1(_32626), .DIN2(_32518), .Q(_30842) );
  nor2s1 _32519_inst ( .DIN1(_32627), .DIN2(_32628), .Q(_32621) );
  nor2s1 _32520_inst ( .DIN1(_32624), .DIN2(_32625), .Q(_32628) );
  nnd2s1 _32521_inst ( .DIN1(_32629), .DIN2(_32630), .Q(_32625) );
  nnd2s1 _32522_inst ( .DIN1(_32631), .DIN2(_32632), .Q(_32630) );
  nor2s1 _32523_inst ( .DIN1(_32633), .DIN2(_30840), .Q(_32631) );
  xor2s1 _32524_inst ( .DIN1(_31768), .DIN2(_32634), .Q(_32629) );
  nnd2s1 _32525_inst ( .DIN1(_32635), .DIN2(_32636), .Q(_32634) );
  nnd2s1 _32526_inst ( .DIN1(_32637), .DIN2(_30840), .Q(_32636) );
  nor2s1 _32527_inst ( .DIN1(_32638), .DIN2(_32626), .Q(_30840) );
  and2s1 _32528_inst ( .DIN1(_32573), .DIN2(_30843), .Q(_32638) );
  nor2s1 _32529_inst ( .DIN1(_32633), .DIN2(_32632), .Q(_32637) );
  nnd2s1 _32530_inst ( .DIN1(_32639), .DIN2(_30843), .Q(_32635) );
  nnd2s1 _32531_inst ( .DIN1(_32640), .DIN2(_32641), .Q(_32639) );
  nnd2s1 _32532_inst ( .DIN1(_32642), .DIN2(_32601), .Q(_32641) );
  hi1s1 _32533_inst ( .DIN(_32607), .Q(_32601) );
  xor2s1 _32534_inst ( .DIN1(_32643), .DIN2(_32644), .Q(_32624) );
  nor2s1 _32535_inst ( .DIN1(_32620), .DIN2(_32645), .Q(_32618) );
  or2s1 _32536_inst ( .DIN1(_30841), .DIN2(_32627), .Q(_32645) );
  nor2s1 _32537_inst ( .DIN1(_30814), .DIN2(_32610), .Q(_32627) );
  xor2s1 _32538_inst ( .DIN1(_32646), .DIN2(_32647), .Q(_32610) );
  xnr2s1 _32539_inst ( .DIN1(_32648), .DIN2(_32466), .Q(_30814) );
  xor2s1 _32540_inst ( .DIN1(_32649), .DIN2(_32650), .Q(_32648) );
  and2s1 _32541_inst ( .DIN1(_32649), .DIN2(_32651), .Q(_30841) );
  nnd2s1 _32542_inst ( .DIN1(_32652), .DIN2(_32482), .Q(_32651) );
  xnr2s1 _32543_inst ( .DIN1(_32653), .DIN2(_26818), .Q(_32620) );
  xor2s1 _32544_inst ( .DIN1(_32655), .DIN2(_32656), .Q(_32561) );
  xor2s1 _32545_inst ( .DIN1(_32657), .DIN2(_32658), .Q(_30794) );
  nor2s1 _32546_inst ( .DIN1(_32659), .DIN2(_32660), .Q(_32658) );
  nnd2s1 _32547_inst ( .DIN1(_32661), .DIN2(_32662), .Q(_32660) );
  nnd2s1 _32548_inst ( .DIN1(_32663), .DIN2(_32302), .Q(_32662) );
  nor2s1 _32549_inst ( .DIN1(_32664), .DIN2(_32640), .Q(_32663) );
  nnd2s1 _32550_inst ( .DIN1(_32665), .DIN2(_32357), .Q(_32661) );
  xor2s1 _32551_inst ( .DIN1(_32666), .DIN2(_32667), .Q(_32665) );
  nor2s1 _32552_inst ( .DIN1(_32667), .DIN2(_32668), .Q(_32659) );
  hi1s1 _32553_inst ( .DIN(_32640), .Q(_32667) );
  xnr2s1 _32554_inst ( .DIN1(_32573), .DIN2(_32669), .Q(_30754) );
  xor2s1 _32555_inst ( .DIN1(_32575), .DIN2(_32268), .Q(_32669) );
  xor2s1 _32556_inst ( .DIN1(_32584), .DIN2(_26821), .Q(_32268) );
  nnd2s1 _32557_inst ( .DIN1(_32671), .DIN2(_32672), .Q(_32584) );
  nnd2s1 _32558_inst ( .DIN1(_32673), .DIN2(_32674), .Q(_32672) );
  or2s1 _32559_inst ( .DIN1(_32675), .DIN2(_26798), .Q(_32674) );
  nnd2s1 _32560_inst ( .DIN1(_438), .DIN2(_32675), .Q(_32671) );
  nnd2s1 _32561_inst ( .DIN1(_32676), .DIN2(_32677), .Q(_32575) );
  nnd2s1 _32562_inst ( .DIN1(_32357), .DIN2(_32666), .Q(_32677) );
  xnr2s1 _32563_inst ( .DIN1(_32615), .DIN2(_32678), .Q(_32676) );
  nnd2s1 _32564_inst ( .DIN1(_32640), .DIN2(_32668), .Q(_32678) );
  nnd2s1 _32565_inst ( .DIN1(_32664), .DIN2(_32302), .Q(_32668) );
  hi1s1 _32566_inst ( .DIN(_32357), .Q(_32302) );
  xor2s1 _32567_inst ( .DIN1(_32675), .DIN2(_32589), .Q(_32357) );
  and2s1 _32568_inst ( .DIN1(_32679), .DIN2(_32680), .Q(_32589) );
  or2s1 _32569_inst ( .DIN1(_29732), .DIN2(_32681), .Q(_32680) );
  nor2s1 _32570_inst ( .DIN1(_32682), .DIN2(_32683), .Q(_32679) );
  nor2s1 _32571_inst ( .DIN1(_32673), .DIN2(_32684), .Q(_32683) );
  xor2s1 _32572_inst ( .DIN1(_32681), .DIN2(_29752), .Q(_32684) );
  nor2s1 _32573_inst ( .DIN1(_15561), .DIN2(_32685), .Q(_32682) );
  nnd2s1 _32574_inst ( .DIN1(_32681), .DIN2(_26798), .Q(_32685) );
  nnd2s1 _32575_inst ( .DIN1(_32686), .DIN2(_32687), .Q(_32675) );
  nnd2s1 _32576_inst ( .DIN1(_32688), .DIN2(_32689), .Q(_32687) );
  or2s1 _32577_inst ( .DIN1(_32690), .DIN2(_441), .Q(_32689) );
  xor2s1 _32578_inst ( .DIN1(_32691), .DIN2(_32681), .Q(_32686) );
  nnd2s1 _32579_inst ( .DIN1(_441), .DIN2(_32690), .Q(_32691) );
  hi1s1 _32580_inst ( .DIN(_32666), .Q(_32664) );
  nnd2s1 _32581_inst ( .DIN1(_32692), .DIN2(_32693), .Q(_32666) );
  nnd2s1 _32582_inst ( .DIN1(_32694), .DIN2(_32607), .Q(_32693) );
  xor2s1 _32583_inst ( .DIN1(_32600), .DIN2(_32612), .Q(_32694) );
  nor2s1 _32584_inst ( .DIN1(_32605), .DIN2(_32413), .Q(_32600) );
  nnd2s1 _32585_inst ( .DIN1(_32413), .DIN2(_32605), .Q(_32692) );
  nnd2s1 _32586_inst ( .DIN1(_32695), .DIN2(_32696), .Q(_32605) );
  nnd2s1 _32587_inst ( .DIN1(_32697), .DIN2(_32698), .Q(_32696) );
  xnr2s1 _32588_inst ( .DIN1(_32615), .DIN2(_32699), .Q(_32698) );
  nnd2s1 _32589_inst ( .DIN1(_32429), .DIN2(_32649), .Q(_32699) );
  hi1s1 _32590_inst ( .DIN(_32700), .Q(_32649) );
  nnd2s1 _32591_inst ( .DIN1(_32700), .DIN2(_32466), .Q(_32695) );
  hi1s1 _32592_inst ( .DIN(_32429), .Q(_32466) );
  xnr2s1 _32593_inst ( .DIN1(_32655), .DIN2(_32701), .Q(_32429) );
  xor2s1 _32594_inst ( .DIN1(_32702), .DIN2(_29752), .Q(_32655) );
  nor2s1 _32595_inst ( .DIN1(_32482), .DIN2(_32652), .Q(_32700) );
  and2s1 _32596_inst ( .DIN1(_32703), .DIN2(_32704), .Q(_32652) );
  nnd2s1 _32597_inst ( .DIN1(_32626), .DIN2(_32518), .Q(_32704) );
  xor2s1 _32598_inst ( .DIN1(_32705), .DIN2(_26818), .Q(_32518) );
  nor2s1 _32599_inst ( .DIN1(_30843), .DIN2(_32573), .Q(_32626) );
  nnd2s1 _32600_inst ( .DIN1(_32706), .DIN2(_32642), .Q(_30843) );
  nor2s1 _32601_inst ( .DIN1(_654), .DIN2(_32697), .Q(_32642) );
  hi1s1 _32602_inst ( .DIN(_32650), .Q(_32697) );
  xnr2s1 _32603_inst ( .DIN1(_32703), .DIN2(_32707), .Q(_32650) );
  nor2s1 _32604_inst ( .DIN1(_32607), .DIN2(_32640), .Q(_32706) );
  nnd2s1 _32605_inst ( .DIN1(_32708), .DIN2(_32709), .Q(_32607) );
  nnd2s1 _32606_inst ( .DIN1(_32710), .DIN2(_32711), .Q(_32709) );
  nnd2s1 _32607_inst ( .DIN1(_648), .DIN2(_652), .Q(_32711) );
  nor2s1 _32608_inst ( .DIN1(_29836), .DIN2(_654), .Q(_32710) );
  and2s1 _32609_inst ( .DIN1(_32712), .DIN2(_32713), .Q(_29836) );
  nor2s1 _32610_inst ( .DIN1(_654), .DIN2(_652), .Q(_32712) );
  xor2s1 _32611_inst ( .DIN1(_32714), .DIN2(_32647), .Q(_32482) );
  xor2s1 _32612_inst ( .DIN1(_29871), .DIN2(_32715), .Q(_32647) );
  xor2s1 _32613_inst ( .DIN1(_32716), .DIN2(_32717), .Q(_32714) );
  hi1s1 _32614_inst ( .DIN(_32360), .Q(_32413) );
  xor2s1 _32615_inst ( .DIN1(_32690), .DIN2(_32594), .Q(_32360) );
  xor2s1 _32616_inst ( .DIN1(_32715), .DIN2(_433), .Q(_32594) );
  nnd2s1 _32617_inst ( .DIN1(_32718), .DIN2(_32719), .Q(_32690) );
  nnd2s1 _32618_inst ( .DIN1(_14172), .DIN2(_32720), .Q(_32719) );
  or2s1 _32619_inst ( .DIN1(_32701), .DIN2(_29752), .Q(_32720) );
  nnd2s1 _32620_inst ( .DIN1(_29752), .DIN2(_32701), .Q(_32718) );
  nnd2s1 _32621_inst ( .DIN1(_32721), .DIN2(_32722), .Q(_32701) );
  nnd2s1 _32622_inst ( .DIN1(_32715), .DIN2(_32723), .Q(_32722) );
  nnd2s1 _32623_inst ( .DIN1(_32717), .DIN2(_29871), .Q(_32723) );
  hi1s1 _32624_inst ( .DIN(_32724), .Q(_32717) );
  nnd2s1 _32625_inst ( .DIN1(_26827), .DIN2(_32724), .Q(_32721) );
  nnd2s1 _32626_inst ( .DIN1(_32725), .DIN2(_32726), .Q(_32724) );
  nnd2s1 _32627_inst ( .DIN1(_15563), .DIN2(_32727), .Q(_32726) );
  or2s1 _32628_inst ( .DIN1(_32705), .DIN2(_32702), .Q(_32727) );
  nnd2s1 _32629_inst ( .DIN1(_32702), .DIN2(_32705), .Q(_32725) );
  nnd2s1 _32630_inst ( .DIN1(_32728), .DIN2(_32729), .Q(_32705) );
  nnd2s1 _32631_inst ( .DIN1(_648), .DIN2(_32730), .Q(_32729) );
  or2s1 _32632_inst ( .DIN1(_32731), .DIN2(_29871), .Q(_32730) );
  nnd2s1 _32633_inst ( .DIN1(_29871), .DIN2(_32731), .Q(_32728) );
  xor2s1 _32634_inst ( .DIN1(_32732), .DIN2(_32632), .Q(_32640) );
  xor2s1 _32635_inst ( .DIN1(_32707), .DIN2(_29872), .Q(_32632) );
  xnr2s1 _32636_inst ( .DIN1(_32644), .DIN2(_32731), .Q(_32573) );
  nnd2s1 _32637_inst ( .DIN1(_32733), .DIN2(_32734), .Q(_32731) );
  or2s1 _32638_inst ( .DIN1(_32732), .DIN2(_32707), .Q(_32734) );
  nor2s1 _32639_inst ( .DIN1(_32735), .DIN2(_32736), .Q(_32733) );
  nor2s1 _32640_inst ( .DIN1(_32737), .DIN2(_15563), .Q(_32736) );
  nor2s1 _32641_inst ( .DIN1(_32738), .DIN2(_652), .Q(_32737) );
  nor2s1 _32642_inst ( .DIN1(_27329), .DIN2(_32732), .Q(_32738) );
  nor2s1 _32643_inst ( .DIN1(_27338), .DIN2(_32739), .Q(_32735) );
  nor2s1 _32644_inst ( .DIN1(_15563), .DIN2(_32732), .Q(_32739) );
  nnd2s1 _32645_inst ( .DIN1(_32713), .DIN2(_32740), .Q(_32732) );
  nnd2s1 _32646_inst ( .DIN1(_652), .DIN2(_32703), .Q(_32740) );
  hi1s1 _32647_inst ( .DIN(_648), .Q(_32713) );
  xor2s1 _32648_inst ( .DIN1(_648), .DIN2(_640), .Q(_32644) );
  xnr2s1 _32649_inst ( .DIN1(_32510), .DIN2(_26821), .Q(_32533) );
  hi1s1 _32650_inst ( .DIN(_32525), .Q(_15560) );
  xor2s1 _32651_inst ( .DIN1(_32580), .DIN2(_32741), .Q(_32525) );
  xor2s1 _32652_inst ( .DIN1(_52848), .DIN2(_53495), .Q(_32741) );
  nnd2s1 _32653_inst ( .DIN1(_32742), .DIN2(_32743), .Q(_32580) );
  nnd2s1 _32654_inst ( .DIN1(_53125), .DIN2(_32744), .Q(_32743) );
  or2s1 _32655_inst ( .DIN1(_26431), .DIN2(_32745), .Q(_32744) );
  nnd2s1 _32656_inst ( .DIN1(_32745), .DIN2(_26431), .Q(_32742) );
  nnd2s1 _32657_inst ( .DIN1(_32746), .DIN2(_32747), .Q(_32510) );
  nnd2s1 _32658_inst ( .DIN1(_32588), .DIN2(_29732), .Q(_32747) );
  nnd2s1 _32659_inst ( .DIN1(_29752), .DIN2(_32673), .Q(_29732) );
  hi1s1 _32660_inst ( .DIN(_438), .Q(_29752) );
  nnd2s1 _32661_inst ( .DIN1(_32748), .DIN2(_32749), .Q(_32588) );
  nnd2s1 _32662_inst ( .DIN1(_441), .DIN2(_32750), .Q(_32749) );
  or2s1 _32663_inst ( .DIN1(_32593), .DIN2(_433), .Q(_32750) );
  nnd2s1 _32664_inst ( .DIN1(_433), .DIN2(_32593), .Q(_32748) );
  nnd2s1 _32665_inst ( .DIN1(_32751), .DIN2(_32752), .Q(_32593) );
  nnd2s1 _32666_inst ( .DIN1(_438), .DIN2(_32656), .Q(_32752) );
  xor2s1 _32667_inst ( .DIN1(_32753), .DIN2(_32754), .Q(_32751) );
  nnd2s1 _32668_inst ( .DIN1(_14172), .DIN2(_32755), .Q(_32754) );
  or2s1 _32669_inst ( .DIN1(_32656), .DIN2(_26798), .Q(_32755) );
  nnd2s1 _32670_inst ( .DIN1(_32756), .DIN2(_32757), .Q(_32656) );
  nnd2s1 _32671_inst ( .DIN1(_441), .DIN2(_32758), .Q(_32757) );
  or2s1 _32672_inst ( .DIN1(_32646), .DIN2(_26827), .Q(_32758) );
  xor2s1 _32673_inst ( .DIN1(_32759), .DIN2(_32760), .Q(_441) );
  xor2s1 _32674_inst ( .DIN1(_53156), .DIN2(_53498), .Q(_32760) );
  xor2s1 _32675_inst ( .DIN1(_32761), .DIN2(_32762), .Q(_32759) );
  nnd2s1 _32676_inst ( .DIN1(_26827), .DIN2(_32646), .Q(_32756) );
  nnd2s1 _32677_inst ( .DIN1(_32763), .DIN2(_32764), .Q(_32646) );
  nnd2s1 _32678_inst ( .DIN1(_32653), .DIN2(_29837), .Q(_32764) );
  nnd2s1 _32679_inst ( .DIN1(_32702), .DIN2(_29872), .Q(_29837) );
  nnd2s1 _32680_inst ( .DIN1(_32765), .DIN2(_32766), .Q(_32653) );
  nnd2s1 _32681_inst ( .DIN1(_26827), .DIN2(_32767), .Q(_32766) );
  or2s1 _32682_inst ( .DIN1(_32643), .DIN2(_648), .Q(_32767) );
  xor2s1 _32683_inst ( .DIN1(_30674), .DIN2(_32768), .Q(_32765) );
  nnd2s1 _32684_inst ( .DIN1(_648), .DIN2(_32643), .Q(_32768) );
  nnd2s1 _32685_inst ( .DIN1(_32769), .DIN2(_32770), .Q(_32643) );
  nnd2s1 _32686_inst ( .DIN1(_15563), .DIN2(_32771), .Q(_32770) );
  nnd2s1 _32687_inst ( .DIN1(_32707), .DIN2(_32708), .Q(_32771) );
  nnd2s1 _32688_inst ( .DIN1(_32633), .DIN2(_652), .Q(_32769) );
  xor2s1 _32689_inst ( .DIN1(_32772), .DIN2(_32773), .Q(_652) );
  xor2s1 _32690_inst ( .DIN1(_52844), .DIN2(_53511), .Q(_32773) );
  hi1s1 _32691_inst ( .DIN(_32708), .Q(_32633) );
  nnd2s1 _32692_inst ( .DIN1(_654), .DIN2(_648), .Q(_32708) );
  hi1s1 _32693_inst ( .DIN(_32703), .Q(_654) );
  nnd2s1 _32694_inst ( .DIN1(_32772), .DIN2(_32774), .Q(_32703) );
  nnd2s1 _32695_inst ( .DIN1(_53135), .DIN2(_26562), .Q(_32774) );
  xor2s1 _32696_inst ( .DIN1(_32775), .DIN2(_32776), .Q(_648) );
  xor2s1 _32697_inst ( .DIN1(_53134), .DIN2(_53506), .Q(_32776) );
  nnd2s1 _32698_inst ( .DIN1(_14172), .DIN2(_15563), .Q(_32763) );
  hi1s1 _32699_inst ( .DIN(_29872), .Q(_15563) );
  xnr2s1 _32700_inst ( .DIN1(_32777), .DIN2(_32778), .Q(_29872) );
  xor2s1 _32701_inst ( .DIN1(_26542), .DIN2(_53510), .Q(_32777) );
  xor2s1 _32702_inst ( .DIN1(_32779), .DIN2(_32780), .Q(_640) );
  xor2s1 _32703_inst ( .DIN1(_53507), .DIN2(_53508), .Q(_32780) );
  hi1s1 _32704_inst ( .DIN(_32688), .Q(_433) );
  xnr2s1 _32705_inst ( .DIN1(_32781), .DIN2(_32782), .Q(_32688) );
  xor2s1 _32706_inst ( .DIN1(_26411), .DIN2(_52850), .Q(_32781) );
  nnd2s1 _32707_inst ( .DIN1(_26798), .DIN2(_15561), .Q(_32746) );
  hi1s1 _32708_inst ( .DIN(_32673), .Q(_15561) );
  xor2s1 _32709_inst ( .DIN1(_32745), .DIN2(_32783), .Q(_32673) );
  xor2s1 _32710_inst ( .DIN1(_53125), .DIN2(_53496), .Q(_32783) );
  nnd2s1 _32711_inst ( .DIN1(_32784), .DIN2(_32785), .Q(_32745) );
  nnd2s1 _32712_inst ( .DIN1(_52850), .DIN2(_32786), .Q(_32785) );
  nnd2s1 _32713_inst ( .DIN1(_26411), .DIN2(_32782), .Q(_32786) );
  or2s1 _32714_inst ( .DIN1(_26411), .DIN2(_32782), .Q(_32784) );
  nnd2s1 _32715_inst ( .DIN1(_32787), .DIN2(_32788), .Q(_32782) );
  nnd2s1 _32716_inst ( .DIN1(_32789), .DIN2(_26739), .Q(_32788) );
  or2s1 _32717_inst ( .DIN1(_32790), .DIN2(_53360), .Q(_32789) );
  nnd2s1 _32718_inst ( .DIN1(_53360), .DIN2(_32790), .Q(_32787) );
  xor2s1 _32719_inst ( .DIN1(_32790), .DIN2(_32791), .Q(_438) );
  xor2s1 _32720_inst ( .DIN1(_53057), .DIN2(_53360), .Q(_32791) );
  nnd2s1 _32721_inst ( .DIN1(_32792), .DIN2(_32793), .Q(_32790) );
  nnd2s1 _32722_inst ( .DIN1(_53156), .DIN2(_32794), .Q(_32793) );
  nnd2s1 _32723_inst ( .DIN1(_53498), .DIN2(_32761), .Q(_32794) );
  or2s1 _32724_inst ( .DIN1(_32761), .DIN2(_53498), .Q(_32792) );
  xor2s1 _32725_inst ( .DIN1(_32795), .DIN2(_32681), .Q(_32761) );
  nnd2s1 _32726_inst ( .DIN1(_32796), .DIN2(_32797), .Q(_32795) );
  nnd2s1 _32727_inst ( .DIN1(_53513), .DIN2(_32798), .Q(_32797) );
  nnd2s1 _32728_inst ( .DIN1(_26559), .DIN2(_32799), .Q(_32798) );
  or2s1 _32729_inst ( .DIN1(_26559), .DIN2(_32799), .Q(_32796) );
  xor2s1 _32730_inst ( .DIN1(_27413), .DIN2(_53006), .Q(_32552) );
  nnd2s1 _32731_inst ( .DIN1(_31554), .DIN2(_32348), .Q(_32496) );
  hi1s1 _32732_inst ( .DIN(_28660), .Q(_32348) );
  nnd2s1 _32733_inst ( .DIN1(_32800), .DIN2(_32333), .Q(_28660) );
  and2s1 _32734_inst ( .DIN1(_31366), .DIN2(_32340), .Q(_32333) );
  nor2s1 _32735_inst ( .DIN1(_30831), .DIN2(_30374), .Q(_31366) );
  hi1s1 _32736_inst ( .DIN(_30677), .Q(_30374) );
  nor2s1 _32737_inst ( .DIN1(_32801), .DIN2(_31964), .Q(_32800) );
  hi1s1 _32738_inst ( .DIN(_30848), .Q(_31964) );
  hi1s1 _32739_inst ( .DIN(_31606), .Q(_31554) );
  nor2s1 _32740_inst ( .DIN1(_31708), .DIN2(_32802), .Q(_32549) );
  nnd2s1 _32741_inst ( .DIN1(______[14]), .DIN2(_32491), .Q(_32802) );
  xor2s1 _32742_inst ( .DIN1(_53005), .DIN2(_53004), .Q(_32491) );
  nnd2s1 _32743_inst ( .DIN1(_31606), .DIN2(_31405), .Q(_31708) );
  nnd2s1 _32744_inst ( .DIN1(_32803), .DIN2(_32804), .Q(_31405) );
  hi1s1 _32745_inst ( .DIN(_27318), .Q(_32804) );
  nnd2s1 _32746_inst ( .DIN1(_32805), .DIN2(_32806), .Q(_27318) );
  nor2s1 _32747_inst ( .DIN1(_32807), .DIN2(_32808), .Q(_32806) );
  nnd2s1 _32748_inst ( .DIN1(_27441), .DIN2(_32809), .Q(_32808) );
  nor2s1 _32749_inst ( .DIN1(_27309), .DIN2(_27431), .Q(_32805) );
  nor2s1 _32750_inst ( .DIN1(_32810), .DIN2(_31397), .Q(_32803) );
  nnd2s1 _32751_inst ( .DIN1(_32811), .DIN2(_32812), .Q(_31606) );
  nor2s1 _32752_inst ( .DIN1(_32813), .DIN2(_32814), .Q(_32812) );
  nnd2s1 _32753_inst ( .DIN1(_32809), .DIN2(_29741), .Q(_32814) );
  nor2s1 _32754_inst ( .DIN1(_32815), .DIN2(_29434), .Q(_32811) );
  nnd2s1 _32755_inst ( .DIN1(_32816), .DIN2(_32817), .Q(_29434) );
  nor2s1 _32756_inst ( .DIN1(_32818), .DIN2(_32819), .Q(_32817) );
  nnd2s1 _32757_inst ( .DIN1(_27442), .DIN2(_32820), .Q(_32819) );
  nnd2s1 _32758_inst ( .DIN1(_32821), .DIN2(_29408), .Q(_32818) );
  nor2s1 _32759_inst ( .DIN1(_32822), .DIN2(_32823), .Q(_32816) );
  nnd2s1 _32760_inst ( .DIN1(_32824), .DIN2(_32825), .Q(_32823) );
  nnd2s1 _32761_inst ( .DIN1(_27446), .DIN2(_32826), .Q(_32822) );
  nnd2s1 _32762_inst ( .DIN1(_32827), .DIN2(_32828), .Q(
        _____________________________9________) );
  nnd2s1 _32763_inst ( .DIN1(_32829), .DIN2(_32830), .Q(_32828) );
  nnd2s1 _32764_inst ( .DIN1(_32831), .DIN2(_32832), .Q(_32829) );
  nor2s1 _32765_inst ( .DIN1(_32833), .DIN2(_32834), .Q(_32832) );
  nor2s1 _32766_inst ( .DIN1(_32835), .DIN2(_27365), .Q(_32831) );
  nor2s1 _32767_inst ( .DIN1(_53252), .DIN2(_53253), .Q(_32835) );
  nnd2s1 _32768_inst ( .DIN1(_32836), .DIN2(_32837), .Q(_32827) );
  nor2s1 _32769_inst ( .DIN1(_32838), .DIN2(_32839), .Q(_32836) );
  xor2s1 _32770_inst ( .DIN1(_32840), .DIN2(_32841), .Q(_32838) );
  xnr2s1 _32771_inst ( .DIN1(_53008), .DIN2(_32842), .Q(_32841) );
  nnd2s1 _32772_inst ( .DIN1(_32843), .DIN2(_32844), .Q(
        _____________________________99________) );
  nor2s1 _32773_inst ( .DIN1(_32845), .DIN2(_32846), .Q(_32843) );
  nor2s1 _32774_inst ( .DIN1(_32847), .DIN2(_32848), .Q(_32846) );
  nnd2s1 _32775_inst ( .DIN1(_32849), .DIN2(_32850), .Q(_32848) );
  xor2s1 _32776_inst ( .DIN1(_30163), .DIN2(_32851), .Q(_32850) );
  nor2s1 _32777_inst ( .DIN1(_32852), .DIN2(_32853), .Q(_32851) );
  nnd2s1 _32778_inst ( .DIN1(_32854), .DIN2(_32855), .Q(_32853) );
  nnd2s1 _32779_inst ( .DIN1(_32856), .DIN2(_32857), .Q(_32854) );
  nnd2s1 _32780_inst ( .DIN1(_32858), .DIN2(_32859), .Q(_32852) );
  nnd2s1 _32781_inst ( .DIN1(_53215), .DIN2(_53344), .Q(_32859) );
  nnd2s1 _32782_inst ( .DIN1(_32860), .DIN2(_26613), .Q(_32858) );
  nor2s1 _32783_inst ( .DIN1(_53215), .DIN2(_32856), .Q(_32860) );
  nor2s1 _32784_inst ( .DIN1(_32861), .DIN2(_32862), .Q(_32849) );
  nor2s1 _32785_inst ( .DIN1(_32855), .DIN2(_32863), .Q(_32862) );
  xor2s1 _32786_inst ( .DIN1(_32864), .DIN2(_32865), .Q(_32863) );
  xor2s1 _32787_inst ( .DIN1(_26220), .DIN2(_32866), .Q(_32865) );
  hi1s1 _32788_inst ( .DIN(_32867), .Q(_32864) );
  nor2s1 _32789_inst ( .DIN1(_32868), .DIN2(_32869), .Q(_32845) );
  nor2s1 _32790_inst ( .DIN1(_27291), .DIN2(_32870), .Q(_32869) );
  xnr2s1 _32791_inst ( .DIN1(_53340), .DIN2(_32871), .Q(_32870) );
  nor2s1 _32792_inst ( .DIN1(_32872), .DIN2(_32873), .Q(
        _____________________________98________) );
  nor2s1 _32793_inst ( .DIN1(_32861), .DIN2(_32874), .Q(_32872) );
  nnd2s1 _32794_inst ( .DIN1(_32875), .DIN2(_32876), .Q(_32874) );
  nnd2s1 _32795_inst ( .DIN1(_53343), .DIN2(_32855), .Q(_32876) );
  nnd2s1 _32796_inst ( .DIN1(_32877), .DIN2(_32878), .Q(_32875) );
  xor2s1 _32797_inst ( .DIN1(_32879), .DIN2(_32880), .Q(_32877) );
  xor2s1 _32798_inst ( .DIN1(_32881), .DIN2(_53015), .Q(_32879) );
  nnd2s1 _32799_inst ( .DIN1(_32882), .DIN2(_28569), .Q(
        _____________________________97________) );
  nor2s1 _32800_inst ( .DIN1(_32883), .DIN2(_32884), .Q(_32882) );
  nor2s1 _32801_inst ( .DIN1(_32885), .DIN2(_28575), .Q(_32884) );
  nor2s1 _32802_inst ( .DIN1(_32861), .DIN2(_32886), .Q(_32885) );
  nnd2s1 _32803_inst ( .DIN1(_32887), .DIN2(_32888), .Q(_32886) );
  nnd2s1 _32804_inst ( .DIN1(_53344), .DIN2(_32855), .Q(_32888) );
  nnd2s1 _32805_inst ( .DIN1(_32878), .DIN2(_32889), .Q(_32887) );
  nnd2s1 _32806_inst ( .DIN1(_32881), .DIN2(_32890), .Q(_32889) );
  nnd2s1 _32807_inst ( .DIN1(_32891), .DIN2(_53014), .Q(_32890) );
  nor2s1 _32808_inst ( .DIN1(_28572), .DIN2(_32892), .Q(_32883) );
  nor2s1 _32809_inst ( .DIN1(_32893), .DIN2(_26771), .Q(_32892) );
  xor2s1 _32810_inst ( .DIN1(_32894), .DIN2(_32895), .Q(_32893) );
  xor2s1 _32811_inst ( .DIN1(_53009), .DIN2(_53224), .Q(_32895) );
  nnd2s1 _32812_inst ( .DIN1(_53050), .DIN2(_53224), .Q(_32894) );
  nor2s1 _32813_inst ( .DIN1(_32896), .DIN2(_27235), .Q(
        _____________________________96________) );
  nor2s1 _32814_inst ( .DIN1(_32897), .DIN2(_32898), .Q(_32896) );
  nnd2s1 _32815_inst ( .DIN1(_32899), .DIN2(_32900), .Q(_32898) );
  nnd2s1 _32816_inst ( .DIN1(_32901), .DIN2(_26487), .Q(_32900) );
  nnd2s1 _32817_inst ( .DIN1(_32902), .DIN2(_32903), .Q(_32901) );
  nnd2s1 _32818_inst ( .DIN1(_32904), .DIN2(_32905), .Q(_32903) );
  nnd2s1 _32819_inst ( .DIN1(_32906), .DIN2(_32907), .Q(_32902) );
  nnd2s1 _32820_inst ( .DIN1(_32908), .DIN2(_53050), .Q(_32899) );
  nnd2s1 _32821_inst ( .DIN1(_32909), .DIN2(_32910), .Q(_32908) );
  nnd2s1 _32822_inst ( .DIN1(_32907), .DIN2(_32905), .Q(_32910) );
  nnd2s1 _32823_inst ( .DIN1(_32906), .DIN2(_32904), .Q(_32909) );
  hi1s1 _32824_inst ( .DIN(_32905), .Q(_32906) );
  nnd2s1 _32825_inst ( .DIN1(_32911), .DIN2(_32912), .Q(_32905) );
  nnd2s1 _32826_inst ( .DIN1(_53069), .DIN2(_32913), .Q(_32912) );
  nnd2s1 _32827_inst ( .DIN1(_32914), .DIN2(_32915), .Q(_32913) );
  or2s1 _32828_inst ( .DIN1(_32914), .DIN2(_32915), .Q(_32911) );
  nor2s1 _32829_inst ( .DIN1(_32916), .DIN2(_32917), .Q(_32897) );
  nor2s1 _32830_inst ( .DIN1(_26772), .DIN2(_32918), .Q(_32917) );
  nnd2s1 _32831_inst ( .DIN1(_32919), .DIN2(_32920), .Q(_32918) );
  xor2s1 _32832_inst ( .DIN1(_26300), .DIN2(_32921), .Q(_32919) );
  nnd2s1 _32833_inst ( .DIN1(_53276), .DIN2(_53277), .Q(_32921) );
  nnd2s1 _32834_inst ( .DIN1(_32922), .DIN2(_28445), .Q(
        _____________________________95________) );
  nor2s1 _32835_inst ( .DIN1(_32923), .DIN2(_32924), .Q(_32922) );
  nor2s1 _32836_inst ( .DIN1(_27845), .DIN2(_32925), .Q(_32924) );
  nnd2s1 _32837_inst ( .DIN1(_32926), .DIN2(_32927), .Q(_32925) );
  nnd2s1 _32838_inst ( .DIN1(_32928), .DIN2(_32929), .Q(_32927) );
  xor2s1 _32839_inst ( .DIN1(_32915), .DIN2(_32930), .Q(_32928) );
  xor2s1 _32840_inst ( .DIN1(_26339), .DIN2(_32914), .Q(_32930) );
  nnd2s1 _32841_inst ( .DIN1(_32931), .DIN2(_32932), .Q(_32915) );
  nnd2s1 _32842_inst ( .DIN1(_53054), .DIN2(_32933), .Q(_32932) );
  or2s1 _32843_inst ( .DIN1(_32934), .DIN2(_32935), .Q(_32933) );
  nnd2s1 _32844_inst ( .DIN1(_32935), .DIN2(_32934), .Q(_32931) );
  nnd2s1 _32845_inst ( .DIN1(_32936), .DIN2(_26554), .Q(_32926) );
  nor2s1 _32846_inst ( .DIN1(_53186), .DIN2(_27836), .Q(_32923) );
  nnd2s1 _32847_inst ( .DIN1(_32937), .DIN2(_32938), .Q(
        _____________________________94________) );
  nor2s1 _32848_inst ( .DIN1(_32939), .DIN2(_32940), .Q(_32938) );
  nor2s1 _32849_inst ( .DIN1(_28032), .DIN2(_32941), .Q(_32940) );
  nnd2s1 _32850_inst ( .DIN1(_32942), .DIN2(_32943), .Q(_32941) );
  nnd2s1 _32851_inst ( .DIN1(_32929), .DIN2(_32944), .Q(_32942) );
  xor2s1 _32852_inst ( .DIN1(_32945), .DIN2(_32946), .Q(_32944) );
  xnr2s1 _32853_inst ( .DIN1(_53054), .DIN2(_32934), .Q(_32946) );
  nnd2s1 _32854_inst ( .DIN1(_32947), .DIN2(_32948), .Q(_32934) );
  nnd2s1 _32855_inst ( .DIN1(_53021), .DIN2(_32949), .Q(_32948) );
  or2s1 _32856_inst ( .DIN1(_32950), .DIN2(_32951), .Q(_32949) );
  nnd2s1 _32857_inst ( .DIN1(_32951), .DIN2(_32950), .Q(_32947) );
  nor2s1 _32858_inst ( .DIN1(_28037), .DIN2(_32952), .Q(_32939) );
  nor2s1 _32859_inst ( .DIN1(_32953), .DIN2(_27365), .Q(_32952) );
  nor2s1 _32860_inst ( .DIN1(_53463), .DIN2(_53464), .Q(_32953) );
  nor2s1 _32861_inst ( .DIN1(_28041), .DIN2(_32954), .Q(_32937) );
  nnd2s1 _32862_inst ( .DIN1(_32955), .DIN2(_32956), .Q(
        _____________________________93________) );
  nnd2s1 _32863_inst ( .DIN1(_32957), .DIN2(_32958), .Q(_32956) );
  xor2s1 _32864_inst ( .DIN1(_32959), .DIN2(_32960), .Q(_32958) );
  xor2s1 _32865_inst ( .DIN1(_53290), .DIN2(_53299), .Q(_32960) );
  nor2s1 _32866_inst ( .DIN1(_32961), .DIN2(_32962), .Q(_32955) );
  nor2s1 _32867_inst ( .DIN1(_32963), .DIN2(_32964), .Q(_32962) );
  nor2s1 _32868_inst ( .DIN1(_32965), .DIN2(_32966), .Q(_32963) );
  nnd2s1 _32869_inst ( .DIN1(______[0]), .DIN2(_32967), .Q(_32966) );
  nnd2s1 _32870_inst ( .DIN1(_32968), .DIN2(_26420), .Q(_32967) );
  nnd2s1 _32871_inst ( .DIN1(_32969), .DIN2(_32936), .Q(_32965) );
  nnd2s1 _32872_inst ( .DIN1(_53462), .DIN2(_32970), .Q(_32969) );
  nnd2s1 _32873_inst ( .DIN1(_53280), .DIN2(_26420), .Q(_32970) );
  nor2s1 _32874_inst ( .DIN1(_32971), .DIN2(_32972), .Q(_32961) );
  xor2s1 _32875_inst ( .DIN1(_32973), .DIN2(_32974), .Q(_32972) );
  xor2s1 _32876_inst ( .DIN1(_26617), .DIN2(_32950), .Q(_32974) );
  nnd2s1 _32877_inst ( .DIN1(_32975), .DIN2(_32976), .Q(_32950) );
  nnd2s1 _32878_inst ( .DIN1(_32977), .DIN2(_26346), .Q(_32976) );
  or2s1 _32879_inst ( .DIN1(_32978), .DIN2(_32979), .Q(_32977) );
  nnd2s1 _32880_inst ( .DIN1(_32979), .DIN2(_32978), .Q(_32975) );
  nnd2s1 _32881_inst ( .DIN1(_32980), .DIN2(_32981), .Q(
        _____________________________92________) );
  nnd2s1 _32882_inst ( .DIN1(_32982), .DIN2(_28801), .Q(_32981) );
  nor2s1 _32883_inst ( .DIN1(_27614), .DIN2(_32983), .Q(_32982) );
  nnd2s1 _32884_inst ( .DIN1(_32984), .DIN2(_32985), .Q(_32983) );
  xor2s1 _32885_inst ( .DIN1(_53140), .DIN2(_53281), .Q(_32984) );
  nnd2s1 _32886_inst ( .DIN1(_32986), .DIN2(_28797), .Q(_32980) );
  nnd2s1 _32887_inst ( .DIN1(_32987), .DIN2(_32988), .Q(_32986) );
  nnd2s1 _32888_inst ( .DIN1(_32989), .DIN2(_32990), .Q(_32988) );
  nnd2s1 _32889_inst ( .DIN1(_32991), .DIN2(_32936), .Q(_32989) );
  xor2s1 _32890_inst ( .DIN1(_53293), .DIN2(_32992), .Q(_32991) );
  nnd2s1 _32891_inst ( .DIN1(_32993), .DIN2(_32929), .Q(_32987) );
  xor2s1 _32892_inst ( .DIN1(_32994), .DIN2(_32995), .Q(_32993) );
  xor2s1 _32893_inst ( .DIN1(_26346), .DIN2(_32978), .Q(_32995) );
  nnd2s1 _32894_inst ( .DIN1(_32996), .DIN2(_32997), .Q(_32978) );
  nnd2s1 _32895_inst ( .DIN1(_53223), .DIN2(_32998), .Q(_32997) );
  or2s1 _32896_inst ( .DIN1(_32999), .DIN2(_33000), .Q(_32998) );
  nnd2s1 _32897_inst ( .DIN1(_33000), .DIN2(_32999), .Q(_32996) );
  nnd2s1 _32898_inst ( .DIN1(_33001), .DIN2(_33002), .Q(
        _____________________________91________) );
  nnd2s1 _32899_inst ( .DIN1(_33003), .DIN2(_33004), .Q(_33002) );
  nnd2s1 _32900_inst ( .DIN1(_33005), .DIN2(_33006), .Q(_33004) );
  xor2s1 _32901_inst ( .DIN1(_26224), .DIN2(_32992), .Q(_33006) );
  nor2s1 _32902_inst ( .DIN1(_33007), .DIN2(_27066), .Q(_33005) );
  hi1s1 _32903_inst ( .DIN(_32964), .Q(_33003) );
  nnd2s1 _32904_inst ( .DIN1(_33008), .DIN2(_32990), .Q(_32964) );
  hi1s1 _32905_inst ( .DIN(_32929), .Q(_32990) );
  nor2s1 _32906_inst ( .DIN1(_33009), .DIN2(_33010), .Q(_33001) );
  nor2s1 _32907_inst ( .DIN1(_33011), .DIN2(_32971), .Q(_33010) );
  nnd2s1 _32908_inst ( .DIN1(_33008), .DIN2(_32929), .Q(_32971) );
  xnr2s1 _32909_inst ( .DIN1(_33000), .DIN2(_33012), .Q(_33011) );
  xnr2s1 _32910_inst ( .DIN1(_53223), .DIN2(_32999), .Q(_33012) );
  nnd2s1 _32911_inst ( .DIN1(_33013), .DIN2(_33014), .Q(_32999) );
  nnd2s1 _32912_inst ( .DIN1(_33015), .DIN2(_26376), .Q(_33014) );
  or2s1 _32913_inst ( .DIN1(_33016), .DIN2(_26828), .Q(_33015) );
  xor2s1 _32914_inst ( .DIN1(_33018), .DIN2(_31888), .Q(_33013) );
  nnd2s1 _32915_inst ( .DIN1(_26828), .DIN2(_33016), .Q(_33018) );
  nor2s1 _32916_inst ( .DIN1(_26420), .DIN2(_33019), .Q(_33009) );
  or2s1 _32917_inst ( .DIN1(_33008), .DIN2(_33020), .Q(_33019) );
  nnd2s1 _32918_inst ( .DIN1(_33021), .DIN2(_33022), .Q(
        _____________________________90________) );
  nnd2s1 _32919_inst ( .DIN1(_33023), .DIN2(_26281), .Q(_33022) );
  nnd2s1 _32920_inst ( .DIN1(_33008), .DIN2(_33024), .Q(_33023) );
  nor2s1 _32921_inst ( .DIN1(_33025), .DIN2(_33026), .Q(_33021) );
  nor2s1 _32922_inst ( .DIN1(_33027), .DIN2(_33028), .Q(_33026) );
  xor2s1 _32923_inst ( .DIN1(_33029), .DIN2(_33030), .Q(_33028) );
  xor2s1 _32924_inst ( .DIN1(_26376), .DIN2(_33016), .Q(_33030) );
  nnd2s1 _32925_inst ( .DIN1(_33031), .DIN2(_33032), .Q(_33016) );
  nnd2s1 _32926_inst ( .DIN1(_53149), .DIN2(_33033), .Q(_33032) );
  or2s1 _32927_inst ( .DIN1(_33034), .DIN2(_33035), .Q(_33033) );
  nnd2s1 _32928_inst ( .DIN1(_33035), .DIN2(_33034), .Q(_33031) );
  nnd2s1 _32929_inst ( .DIN1(_33036), .DIN2(_33037), .Q(
        _____________________________8________) );
  nnd2s1 _32930_inst ( .DIN1(_33038), .DIN2(_33039), .Q(_33037) );
  xor2s1 _32931_inst ( .DIN1(_33040), .DIN2(_33041), .Q(_33038) );
  xor2s1 _32932_inst ( .DIN1(_53032), .DIN2(_53042), .Q(_33041) );
  nnd2s1 _32933_inst ( .DIN1(_53031), .DIN2(_53038), .Q(_33040) );
  nnd2s1 _32934_inst ( .DIN1(_32837), .DIN2(_33042), .Q(_33036) );
  nnd2s1 _32935_inst ( .DIN1(_33043), .DIN2(_33044), .Q(_33042) );
  xor2s1 _32936_inst ( .DIN1(_33045), .DIN2(_53465), .Q(_33043) );
  nnd2s1 _32937_inst ( .DIN1(_33046), .DIN2(_33047), .Q(_33045) );
  nnd2s1 _32938_inst ( .DIN1(_33048), .DIN2(_33049), .Q(
        _____________________________89________) );
  or2s1 _32939_inst ( .DIN1(_33050), .DIN2(_26570), .Q(_33049) );
  nor2s1 _32940_inst ( .DIN1(_33051), .DIN2(_33052), .Q(_33048) );
  nor2s1 _32941_inst ( .DIN1(_33053), .DIN2(_33054), .Q(_33052) );
  nnd2s1 _32942_inst ( .DIN1(_33055), .DIN2(_33056), .Q(_33054) );
  nnd2s1 _32943_inst ( .DIN1(_33057), .DIN2(_33058), .Q(_33056) );
  xor2s1 _32944_inst ( .DIN1(_33059), .DIN2(_33060), .Q(_33057) );
  xor2s1 _32945_inst ( .DIN1(_33034), .DIN2(_33035), .Q(_33060) );
  nnd2s1 _32946_inst ( .DIN1(_33061), .DIN2(_33062), .Q(_33034) );
  nnd2s1 _32947_inst ( .DIN1(_53243), .DIN2(_33063), .Q(_33062) );
  or2s1 _32948_inst ( .DIN1(_33064), .DIN2(_26800), .Q(_33063) );
  xor2s1 _32949_inst ( .DIN1(_33066), .DIN2(_31888), .Q(_33061) );
  nnd2s1 _32950_inst ( .DIN1(_26800), .DIN2(_33064), .Q(_33066) );
  xor2s1 _32951_inst ( .DIN1(_26485), .DIN2(_31802), .Q(_33059) );
  nnd2s1 _32952_inst ( .DIN1(_33067), .DIN2(_33068), .Q(_33055) );
  nor2s1 _32953_inst ( .DIN1(_32992), .DIN2(_32959), .Q(_33067) );
  nor2s1 _32954_inst ( .DIN1(_33069), .DIN2(_33070), .Q(_33051) );
  nor2s1 _32955_inst ( .DIN1(_33071), .DIN2(_33072), .Q(_33070) );
  nnd2s1 _32956_inst ( .DIN1(______[0]), .DIN2(_33073), .Q(_33072) );
  nnd2s1 _32957_inst ( .DIN1(_26570), .DIN2(_26287), .Q(_33073) );
  nnd2s1 _32958_inst ( .DIN1(_33074), .DIN2(_33075), .Q(
        _____________________________88________) );
  nor2s1 _32959_inst ( .DIN1(_33076), .DIN2(_33077), .Q(_33075) );
  nor2s1 _32960_inst ( .DIN1(_29828), .DIN2(_33078), .Q(_33077) );
  nnd2s1 _32961_inst ( .DIN1(_33079), .DIN2(_33080), .Q(_33078) );
  nnd2s1 _32962_inst ( .DIN1(_33058), .DIN2(_33081), .Q(_33080) );
  xor2s1 _32963_inst ( .DIN1(_33082), .DIN2(_33083), .Q(_33081) );
  xor2s1 _32964_inst ( .DIN1(_26366), .DIN2(_33064), .Q(_33083) );
  nnd2s1 _32965_inst ( .DIN1(_33084), .DIN2(_33085), .Q(_33064) );
  nnd2s1 _32966_inst ( .DIN1(_53028), .DIN2(_33086), .Q(_33085) );
  or2s1 _32967_inst ( .DIN1(_33087), .DIN2(_33088), .Q(_33086) );
  nnd2s1 _32968_inst ( .DIN1(_33088), .DIN2(_33087), .Q(_33084) );
  nnd2s1 _32969_inst ( .DIN1(_33068), .DIN2(_33089), .Q(_33079) );
  xor2s1 _32970_inst ( .DIN1(_33090), .DIN2(_33091), .Q(_33089) );
  xor2s1 _32971_inst ( .DIN1(_53221), .DIN2(_53296), .Q(_33091) );
  nor2s1 _32972_inst ( .DIN1(_53299), .DIN2(_53294), .Q(_33090) );
  hi1s1 _32973_inst ( .DIN(_33024), .Q(_33068) );
  nor2s1 _32974_inst ( .DIN1(_29849), .DIN2(_33092), .Q(_33076) );
  nor2s1 _32975_inst ( .DIN1(_33093), .DIN2(_27241), .Q(_33092) );
  nor2s1 _32976_inst ( .DIN1(_53147), .DIN2(_53149), .Q(_33093) );
  and2s1 _32977_inst ( .DIN1(_33094), .DIN2(_29855), .Q(_33074) );
  nor2s1 _32978_inst ( .DIN1(_33095), .DIN2(_27500), .Q(
        _____________________________87________) );
  xor2s1 _32979_inst ( .DIN1(_31222), .DIN2(_33096), .Q(_33095) );
  nor2s1 _32980_inst ( .DIN1(_33097), .DIN2(_33098), .Q(_33096) );
  nor2s1 _32981_inst ( .DIN1(_33099), .DIN2(_33100), .Q(_33098) );
  xor2s1 _32982_inst ( .DIN1(_33101), .DIN2(_33102), .Q(_33099) );
  xor2s1 _32983_inst ( .DIN1(_33087), .DIN2(_33103), .Q(_33102) );
  nnd2s1 _32984_inst ( .DIN1(_33104), .DIN2(_33105), .Q(_33087) );
  nnd2s1 _32985_inst ( .DIN1(_33106), .DIN2(_26505), .Q(_33105) );
  or2s1 _32986_inst ( .DIN1(_33107), .DIN2(_26797), .Q(_33106) );
  nnd2s1 _32987_inst ( .DIN1(_33108), .DIN2(_33107), .Q(_33104) );
  xnr2s1 _32988_inst ( .DIN1(_29492), .DIN2(_53028), .Q(_33101) );
  nor2s1 _32989_inst ( .DIN1(_33024), .DIN2(_33109), .Q(_33097) );
  nnd2s1 _32990_inst ( .DIN1(______[16]), .DIN2(_26412), .Q(_33109) );
  nnd2s1 _32991_inst ( .DIN1(_33110), .DIN2(_33111), .Q(
        _____________________________86________) );
  nor2s1 _32992_inst ( .DIN1(_33112), .DIN2(_33113), .Q(_33111) );
  nor2s1 _32993_inst ( .DIN1(_33114), .DIN2(_33115), .Q(_33113) );
  nnd2s1 _32994_inst ( .DIN1(_33116), .DIN2(_53296), .Q(_33115) );
  nor2s1 _32995_inst ( .DIN1(_26772), .DIN2(_33024), .Q(_33116) );
  nor2s1 _32996_inst ( .DIN1(_33008), .DIN2(_33117), .Q(_33112) );
  nor2s1 _32997_inst ( .DIN1(_32992), .DIN2(_33118), .Q(_33117) );
  nnd2s1 _32998_inst ( .DIN1(_33119), .DIN2(_33120), .Q(_33118) );
  nnd2s1 _32999_inst ( .DIN1(_26269), .DIN2(_26423), .Q(_33120) );
  nnd2s1 _33000_inst ( .DIN1(_32959), .DIN2(_53299), .Q(_33119) );
  nor2s1 _33001_inst ( .DIN1(_26281), .DIN2(_26423), .Q(_32959) );
  nor2s1 _33002_inst ( .DIN1(_53291), .DIN2(_53290), .Q(_32992) );
  nor2s1 _33003_inst ( .DIN1(_33025), .DIN2(_33121), .Q(_33110) );
  nor2s1 _33004_inst ( .DIN1(_33027), .DIN2(_33122), .Q(_33121) );
  xor2s1 _33005_inst ( .DIN1(_33123), .DIN2(_33124), .Q(_33122) );
  xor2s1 _33006_inst ( .DIN1(_26505), .DIN2(_33107), .Q(_33124) );
  nnd2s1 _33007_inst ( .DIN1(_33125), .DIN2(_33126), .Q(_33107) );
  nnd2s1 _33008_inst ( .DIN1(_53029), .DIN2(_33127), .Q(_33126) );
  or2s1 _33009_inst ( .DIN1(_33128), .DIN2(_33129), .Q(_33127) );
  nnd2s1 _33010_inst ( .DIN1(_33129), .DIN2(_33128), .Q(_33125) );
  nnd2s1 _33011_inst ( .DIN1(_33058), .DIN2(_33008), .Q(_33027) );
  nnd2s1 _33012_inst ( .DIN1(_33130), .DIN2(_33131), .Q(
        _____________________________85________) );
  nnd2s1 _33013_inst ( .DIN1(_33132), .DIN2(_33133), .Q(_33131) );
  nnd2s1 _33014_inst ( .DIN1(_33134), .DIN2(_33135), .Q(_33133) );
  nnd2s1 _33015_inst ( .DIN1(_33136), .DIN2(_33137), .Q(_33135) );
  xor2s1 _33016_inst ( .DIN1(_53296), .DIN2(_26269), .Q(_33137) );
  nor2s1 _33017_inst ( .DIN1(_28646), .DIN2(_33024), .Q(_33136) );
  nnd2s1 _33018_inst ( .DIN1(_33100), .DIN2(_33138), .Q(_33024) );
  nnd2s1 _33019_inst ( .DIN1(_33007), .DIN2(_33139), .Q(_33138) );
  hi1s1 _33020_inst ( .DIN(_32936), .Q(_33007) );
  nnd2s1 _33021_inst ( .DIN1(_33140), .DIN2(_33058), .Q(_33134) );
  hi1s1 _33022_inst ( .DIN(_33100), .Q(_33058) );
  xor2s1 _33023_inst ( .DIN1(_33141), .DIN2(_33142), .Q(_33140) );
  xnr2s1 _33024_inst ( .DIN1(_53029), .DIN2(_33128), .Q(_33142) );
  nnd2s1 _33025_inst ( .DIN1(_33143), .DIN2(_33144), .Q(_33128) );
  nnd2s1 _33026_inst ( .DIN1(_33145), .DIN2(_26352), .Q(_33144) );
  or2s1 _33027_inst ( .DIN1(_33146), .DIN2(_26832), .Q(_33145) );
  nnd2s1 _33028_inst ( .DIN1(_26832), .DIN2(_33146), .Q(_33143) );
  nnd2s1 _33029_inst ( .DIN1(_33148), .DIN2(_33149), .Q(_33130) );
  nor2s1 _33030_inst ( .DIN1(_27774), .DIN2(_33150), .Q(_33148) );
  nnd2s1 _33031_inst ( .DIN1(_33151), .DIN2(_33152), .Q(_33150) );
  xor2s1 _33032_inst ( .DIN1(_53151), .DIN2(_53223), .Q(_33151) );
  nnd2s1 _33033_inst ( .DIN1(_33153), .DIN2(_33154), .Q(
        _____________________________84________) );
  nnd2s1 _33034_inst ( .DIN1(_33155), .DIN2(_31026), .Q(_33154) );
  nnd2s1 _33035_inst ( .DIN1(_33156), .DIN2(_33157), .Q(_33155) );
  nor2s1 _33036_inst ( .DIN1(_33158), .DIN2(_33159), .Q(_33157) );
  nor2s1 _33037_inst ( .DIN1(_33160), .DIN2(_27066), .Q(_33156) );
  and2s1 _33038_inst ( .DIN1(_53089), .DIN2(_53306), .Q(_33160) );
  nnd2s1 _33039_inst ( .DIN1(_33161), .DIN2(_27247), .Q(_33153) );
  nor2s1 _33040_inst ( .DIN1(_33162), .DIN2(_33163), .Q(_33161) );
  nor2s1 _33041_inst ( .DIN1(_33164), .DIN2(_33165), .Q(_33163) );
  xor2s1 _33042_inst ( .DIN1(_33166), .DIN2(_33167), .Q(_33164) );
  nor2s1 _33043_inst ( .DIN1(_53306), .DIN2(_53305), .Q(_33167) );
  nnd2s1 _33044_inst ( .DIN1(_33168), .DIN2(_33169), .Q(_33166) );
  nnd2s1 _33045_inst ( .DIN1(_53305), .DIN2(_26689), .Q(_33169) );
  nor2s1 _33046_inst ( .DIN1(_33170), .DIN2(_33171), .Q(_33162) );
  xor2s1 _33047_inst ( .DIN1(_33172), .DIN2(_33173), .Q(_33171) );
  xor2s1 _33048_inst ( .DIN1(_26352), .DIN2(_33146), .Q(_33173) );
  nnd2s1 _33049_inst ( .DIN1(_33174), .DIN2(_33175), .Q(_33146) );
  nnd2s1 _33050_inst ( .DIN1(_53427), .DIN2(_33176), .Q(_33175) );
  or2s1 _33051_inst ( .DIN1(_33177), .DIN2(_33178), .Q(_33176) );
  nnd2s1 _33052_inst ( .DIN1(_33178), .DIN2(_33177), .Q(_33174) );
  hi1s1 _33053_inst ( .DIN(_33147), .Q(_33172) );
  nnd2s1 _33054_inst ( .DIN1(_33179), .DIN2(_27405), .Q(
        _____________________________83________) );
  nnd2s1 _33055_inst ( .DIN1(_33180), .DIN2(_27408), .Q(_27405) );
  nor2s1 _33056_inst ( .DIN1(_33181), .DIN2(_33182), .Q(_33180) );
  nor2s1 _33057_inst ( .DIN1(_33183), .DIN2(_33184), .Q(_33179) );
  nor2s1 _33058_inst ( .DIN1(_27408), .DIN2(_33185), .Q(_33184) );
  nnd2s1 _33059_inst ( .DIN1(_33186), .DIN2(_33187), .Q(_33185) );
  or2s1 _33060_inst ( .DIN1(_33165), .DIN2(_53302), .Q(_33187) );
  nnd2s1 _33061_inst ( .DIN1(_33188), .DIN2(_33189), .Q(_33186) );
  xor2s1 _33062_inst ( .DIN1(_33190), .DIN2(_33191), .Q(_33188) );
  xnr2s1 _33063_inst ( .DIN1(_53427), .DIN2(_33177), .Q(_33191) );
  nnd2s1 _33064_inst ( .DIN1(_33192), .DIN2(_33193), .Q(_33177) );
  nnd2s1 _33065_inst ( .DIN1(_33194), .DIN2(_26380), .Q(_33193) );
  or2s1 _33066_inst ( .DIN1(_33195), .DIN2(_33196), .Q(_33194) );
  nnd2s1 _33067_inst ( .DIN1(_33196), .DIN2(_33195), .Q(_33192) );
  nor2s1 _33068_inst ( .DIN1(_27421), .DIN2(_33197), .Q(_33183) );
  nor2s1 _33069_inst ( .DIN1(_33198), .DIN2(_27291), .Q(_33197) );
  xor2s1 _33070_inst ( .DIN1(_33199), .DIN2(_33200), .Q(_33198) );
  xor2s1 _33071_inst ( .DIN1(_53064), .DIN2(_53065), .Q(_33200) );
  nnd2s1 _33072_inst ( .DIN1(_53515), .DIN2(_53064), .Q(_33199) );
  nnd2s1 _33073_inst ( .DIN1(_33201), .DIN2(_33202), .Q(
        _____________________________82________) );
  nnd2s1 _33074_inst ( .DIN1(_33203), .DIN2(_27246), .Q(_33202) );
  xor2s1 _33075_inst ( .DIN1(_26480), .DIN2(_33159), .Q(_33203) );
  nnd2s1 _33076_inst ( .DIN1(_27247), .DIN2(_33204), .Q(_33201) );
  nnd2s1 _33077_inst ( .DIN1(_33205), .DIN2(_33206), .Q(_33204) );
  nnd2s1 _33078_inst ( .DIN1(_33189), .DIN2(_33207), .Q(_33206) );
  xor2s1 _33079_inst ( .DIN1(_33196), .DIN2(_33208), .Q(_33207) );
  xor2s1 _33080_inst ( .DIN1(_26380), .DIN2(_33195), .Q(_33208) );
  nnd2s1 _33081_inst ( .DIN1(_33209), .DIN2(_33210), .Q(_33195) );
  nnd2s1 _33082_inst ( .DIN1(_53010), .DIN2(_33211), .Q(_33210) );
  or2s1 _33083_inst ( .DIN1(_33212), .DIN2(_33213), .Q(_33211) );
  xor2s1 _33084_inst ( .DIN1(_33214), .DIN2(_33215), .Q(_33209) );
  nnd2s1 _33085_inst ( .DIN1(_33213), .DIN2(_33212), .Q(_33215) );
  nnd2s1 _33086_inst ( .DIN1(_33216), .DIN2(_26378), .Q(_33205) );
  nor2s1 _33087_inst ( .DIN1(_33217), .DIN2(_27500), .Q(
        _____________________________81________) );
  nor2s1 _33088_inst ( .DIN1(_33218), .DIN2(_33219), .Q(_33217) );
  nor2s1 _33089_inst ( .DIN1(_33220), .DIN2(_33170), .Q(_33219) );
  xor2s1 _33090_inst ( .DIN1(_33213), .DIN2(_33221), .Q(_33220) );
  xnr2s1 _33091_inst ( .DIN1(_53010), .DIN2(_33212), .Q(_33221) );
  nnd2s1 _33092_inst ( .DIN1(_33222), .DIN2(_33223), .Q(_33212) );
  nnd2s1 _33093_inst ( .DIN1(_53032), .DIN2(_33224), .Q(_33223) );
  nnd2s1 _33094_inst ( .DIN1(_33225), .DIN2(_33226), .Q(_33224) );
  or2s1 _33095_inst ( .DIN1(_33226), .DIN2(_33225), .Q(_33222) );
  nor2s1 _33096_inst ( .DIN1(_33165), .DIN2(_33227), .Q(_33218) );
  xor2s1 _33097_inst ( .DIN1(_26403), .DIN2(_33168), .Q(_33227) );
  nnd2s1 _33098_inst ( .DIN1(_53308), .DIN2(_26378), .Q(_33168) );
  nnd2s1 _33099_inst ( .DIN1(_33228), .DIN2(_33229), .Q(
        _____________________________80________) );
  nor2s1 _33100_inst ( .DIN1(_33230), .DIN2(_33231), .Q(_33228) );
  nor2s1 _33101_inst ( .DIN1(_27509), .DIN2(_33232), .Q(_33231) );
  nnd2s1 _33102_inst ( .DIN1(_33233), .DIN2(_33234), .Q(_33232) );
  nnd2s1 _33103_inst ( .DIN1(_33235), .DIN2(_33216), .Q(_33234) );
  hi1s1 _33104_inst ( .DIN(_33165), .Q(_33216) );
  nnd2s1 _33105_inst ( .DIN1(_33236), .DIN2(_33170), .Q(_33165) );
  nor2s1 _33106_inst ( .DIN1(_33237), .DIN2(_27774), .Q(_33235) );
  xor2s1 _33107_inst ( .DIN1(_33238), .DIN2(_33239), .Q(_33237) );
  xor2s1 _33108_inst ( .DIN1(_53312), .DIN2(_53320), .Q(_33239) );
  nnd2s1 _33109_inst ( .DIN1(_53331), .DIN2(_26545), .Q(_33238) );
  nnd2s1 _33110_inst ( .DIN1(_33189), .DIN2(_33240), .Q(_33233) );
  xor2s1 _33111_inst ( .DIN1(_33225), .DIN2(_33241), .Q(_33240) );
  xor2s1 _33112_inst ( .DIN1(_53032), .DIN2(_33226), .Q(_33241) );
  xnr2s1 _33113_inst ( .DIN1(_33242), .DIN2(_29231), .Q(_33226) );
  nnd2s1 _33114_inst ( .DIN1(_33243), .DIN2(_33244), .Q(_33242) );
  nnd2s1 _33115_inst ( .DIN1(_33245), .DIN2(_26307), .Q(_33244) );
  nnd2s1 _33116_inst ( .DIN1(_26834), .DIN2(_33247), .Q(_33245) );
  or2s1 _33117_inst ( .DIN1(_33247), .DIN2(_26834), .Q(_33243) );
  nor2s1 _33118_inst ( .DIN1(_53330), .DIN2(_27512), .Q(_33230) );
  nnd2s1 _33119_inst ( .DIN1(_33248), .DIN2(_28794), .Q(
        _____________________________7________) );
  nor2s1 _33120_inst ( .DIN1(_33249), .DIN2(_33250), .Q(_33248) );
  nor2s1 _33121_inst ( .DIN1(_28801), .DIN2(_33251), .Q(_33250) );
  nnd2s1 _33122_inst ( .DIN1(_33044), .DIN2(_33252), .Q(_33251) );
  xnr2s1 _33123_inst ( .DIN1(_33253), .DIN2(_33254), .Q(_33252) );
  xnr2s1 _33124_inst ( .DIN1(_53011), .DIN2(_33255), .Q(_33254) );
  nor2s1 _33125_inst ( .DIN1(_53030), .DIN2(_28797), .Q(_33249) );
  nnd2s1 _33126_inst ( .DIN1(_33256), .DIN2(_33257), .Q(
        _____________________________79________) );
  nnd2s1 _33127_inst ( .DIN1(_33258), .DIN2(_32957), .Q(_33257) );
  and2s1 _33128_inst ( .DIN1(_33259), .DIN2(______[30]), .Q(_32957) );
  nor2s1 _33129_inst ( .DIN1(_33020), .DIN2(_33008), .Q(_33259) );
  xor2s1 _33130_inst ( .DIN1(_33260), .DIN2(_33261), .Q(_33258) );
  xor2s1 _33131_inst ( .DIN1(_53313), .DIN2(_53337), .Q(_33261) );
  nnd2s1 _33132_inst ( .DIN1(_53333), .DIN2(_53312), .Q(_33260) );
  nnd2s1 _33133_inst ( .DIN1(_33262), .DIN2(_33008), .Q(_33256) );
  nor2s1 _33134_inst ( .DIN1(_33263), .DIN2(_33264), .Q(_33262) );
  nor2s1 _33135_inst ( .DIN1(_33170), .DIN2(_33265), .Q(_33264) );
  xor2s1 _33136_inst ( .DIN1(_26834), .DIN2(_33266), .Q(_33265) );
  xor2s1 _33137_inst ( .DIN1(_26307), .DIN2(_33247), .Q(_33266) );
  nnd2s1 _33138_inst ( .DIN1(_33267), .DIN2(_33268), .Q(_33247) );
  nnd2s1 _33139_inst ( .DIN1(_53113), .DIN2(_33269), .Q(_33268) );
  or2s1 _33140_inst ( .DIN1(_33270), .DIN2(_33271), .Q(_33269) );
  nnd2s1 _33141_inst ( .DIN1(_33271), .DIN2(_33270), .Q(_33267) );
  nor2s1 _33142_inst ( .DIN1(_33189), .DIN2(_33272), .Q(_33263) );
  nnd2s1 _33143_inst ( .DIN1(_53331), .DIN2(_33236), .Q(_33272) );
  hi1s1 _33144_inst ( .DIN(_33170), .Q(_33189) );
  nnd2s1 _33145_inst ( .DIN1(_33273), .DIN2(_33274), .Q(_33170) );
  nor2s1 _33146_inst ( .DIN1(_33275), .DIN2(_33276), .Q(_33273) );
  nnd2s1 _33147_inst ( .DIN1(_33277), .DIN2(_33278), .Q(
        _____________________________78________) );
  nnd2s1 _33148_inst ( .DIN1(_33279), .DIN2(_26531), .Q(_33278) );
  nnd2s1 _33149_inst ( .DIN1(_33008), .DIN2(_33280), .Q(_33279) );
  nnd2s1 _33150_inst ( .DIN1(______[28]), .DIN2(_33281), .Q(_33280) );
  nor2s1 _33151_inst ( .DIN1(_33025), .DIN2(_33282), .Q(_33277) );
  nor2s1 _33152_inst ( .DIN1(_33283), .DIN2(_33284), .Q(_33282) );
  nnd2s1 _33153_inst ( .DIN1(_33285), .DIN2(_33008), .Q(_33284) );
  hi1s1 _33154_inst ( .DIN(_33114), .Q(_33008) );
  xnr2s1 _33155_inst ( .DIN1(_33271), .DIN2(_33286), .Q(_33283) );
  xor2s1 _33156_inst ( .DIN1(_53113), .DIN2(_33270), .Q(_33286) );
  nnd2s1 _33157_inst ( .DIN1(_33287), .DIN2(_33288), .Q(_33270) );
  nnd2s1 _33158_inst ( .DIN1(_33289), .DIN2(_26374), .Q(_33288) );
  or2s1 _33159_inst ( .DIN1(_33290), .DIN2(_33291), .Q(_33289) );
  nnd2s1 _33160_inst ( .DIN1(_33291), .DIN2(_33290), .Q(_33287) );
  and2s1 _33161_inst ( .DIN1(_33020), .DIN2(_33114), .Q(_33025) );
  nnd2s1 _33162_inst ( .DIN1(_33292), .DIN2(_33293), .Q(_33114) );
  nor2s1 _33163_inst ( .DIN1(_33294), .DIN2(_33295), .Q(_33020) );
  nnd2s1 _33164_inst ( .DIN1(_33296), .DIN2(_33297), .Q(
        _____________________________77________) );
  nor2s1 _33165_inst ( .DIN1(_33298), .DIN2(_33299), .Q(_33297) );
  nor2s1 _33166_inst ( .DIN1(_33300), .DIN2(_33301), .Q(_33299) );
  nnd2s1 _33167_inst ( .DIN1(______[0]), .DIN2(_33302), .Q(_33301) );
  xor2s1 _33168_inst ( .DIN1(_53312), .DIN2(_53313), .Q(_33302) );
  nor2s1 _33169_inst ( .DIN1(_33303), .DIN2(_33304), .Q(_33296) );
  nor2s1 _33170_inst ( .DIN1(_33305), .DIN2(_33306), .Q(_33304) );
  nor2s1 _33171_inst ( .DIN1(_33307), .DIN2(_28100), .Q(_33306) );
  xor2s1 _33172_inst ( .DIN1(_26380), .DIN2(_53327), .Q(_33307) );
  nor2s1 _33173_inst ( .DIN1(_33308), .DIN2(_33309), .Q(_33303) );
  xor2s1 _33174_inst ( .DIN1(_33310), .DIN2(_33311), .Q(_33308) );
  xor2s1 _33175_inst ( .DIN1(_26374), .DIN2(_33290), .Q(_33311) );
  nnd2s1 _33176_inst ( .DIN1(_33312), .DIN2(_33313), .Q(_33290) );
  nnd2s1 _33177_inst ( .DIN1(_33314), .DIN2(_26590), .Q(_33313) );
  nnd2s1 _33178_inst ( .DIN1(_33315), .DIN2(_33316), .Q(_33314) );
  or2s1 _33179_inst ( .DIN1(_33316), .DIN2(_33315), .Q(_33312) );
  nnd2s1 _33180_inst ( .DIN1(_33317), .DIN2(_33318), .Q(
        _____________________________76________) );
  nor2s1 _33181_inst ( .DIN1(_33298), .DIN2(_33319), .Q(_33318) );
  nor2s1 _33182_inst ( .DIN1(_33320), .DIN2(_33300), .Q(_33319) );
  xor2s1 _33183_inst ( .DIN1(_26582), .DIN2(_33321), .Q(_33320) );
  nor2s1 _33184_inst ( .DIN1(_33322), .DIN2(_33323), .Q(_33317) );
  nor2s1 _33185_inst ( .DIN1(_33305), .DIN2(_33324), .Q(_33323) );
  nor2s1 _33186_inst ( .DIN1(_26774), .DIN2(_26267), .Q(_33324) );
  nor2s1 _33187_inst ( .DIN1(_33309), .DIN2(_33325), .Q(_33322) );
  xor2s1 _33188_inst ( .DIN1(_33315), .DIN2(_33326), .Q(_33325) );
  xor2s1 _33189_inst ( .DIN1(_53037), .DIN2(_33316), .Q(_33326) );
  xnr2s1 _33190_inst ( .DIN1(_33327), .DIN2(_29727), .Q(_33316) );
  hi1s1 _33191_inst ( .DIN(_33328), .Q(_29727) );
  nnd2s1 _33192_inst ( .DIN1(_33329), .DIN2(_33330), .Q(_33327) );
  nnd2s1 _33193_inst ( .DIN1(_33331), .DIN2(_26529), .Q(_33330) );
  or2s1 _33194_inst ( .DIN1(_33332), .DIN2(_33333), .Q(_33331) );
  nnd2s1 _33195_inst ( .DIN1(_33333), .DIN2(_33332), .Q(_33329) );
  nnd2s1 _33196_inst ( .DIN1(_33334), .DIN2(_33335), .Q(
        _____________________________75________) );
  nor2s1 _33197_inst ( .DIN1(_33336), .DIN2(_33337), .Q(_33334) );
  nor2s1 _33198_inst ( .DIN1(_33338), .DIN2(_33339), .Q(_33337) );
  nnd2s1 _33199_inst ( .DIN1(_33340), .DIN2(_33341), .Q(_33339) );
  nnd2s1 _33200_inst ( .DIN1(_33285), .DIN2(_33342), .Q(_33341) );
  xor2s1 _33201_inst ( .DIN1(_33332), .DIN2(_33343), .Q(_33342) );
  xor2s1 _33202_inst ( .DIN1(_26529), .DIN2(_33344), .Q(_33343) );
  xnr2s1 _33203_inst ( .DIN1(_33345), .DIN2(_30163), .Q(_33332) );
  nnd2s1 _33204_inst ( .DIN1(_33346), .DIN2(_33347), .Q(_33345) );
  nnd2s1 _33205_inst ( .DIN1(_33348), .DIN2(_26287), .Q(_33347) );
  nnd2s1 _33206_inst ( .DIN1(_26801), .DIN2(_33350), .Q(_33348) );
  or2s1 _33207_inst ( .DIN1(_33350), .DIN2(_26801), .Q(_33346) );
  nnd2s1 _33208_inst ( .DIN1(_33351), .DIN2(_33281), .Q(_33340) );
  xor2s1 _33209_inst ( .DIN1(_26520), .DIN2(_33321), .Q(_33351) );
  hi1s1 _33210_inst ( .DIN(_33352), .Q(_33321) );
  nor2s1 _33211_inst ( .DIN1(_53072), .DIN2(_30175), .Q(_33336) );
  nnd2s1 _33212_inst ( .DIN1(_33353), .DIN2(_33354), .Q(
        _____________________________74________) );
  nnd2s1 _33213_inst ( .DIN1(_33355), .DIN2(_33356), .Q(_33354) );
  nnd2s1 _33214_inst ( .DIN1(_53313), .DIN2(_33357), .Q(_33355) );
  nnd2s1 _33215_inst ( .DIN1(_33358), .DIN2(_33359), .Q(_33353) );
  nor2s1 _33216_inst ( .DIN1(_33360), .DIN2(_33361), .Q(_33358) );
  nor2s1 _33217_inst ( .DIN1(_33362), .DIN2(_33363), .Q(_33360) );
  nor2s1 _33218_inst ( .DIN1(_33364), .DIN2(_33365), .Q(_33363) );
  xor2s1 _33219_inst ( .DIN1(_33349), .DIN2(_33366), .Q(_33364) );
  xor2s1 _33220_inst ( .DIN1(_26287), .DIN2(_33350), .Q(_33366) );
  nnd2s1 _33221_inst ( .DIN1(_33367), .DIN2(_33368), .Q(_33350) );
  nnd2s1 _33222_inst ( .DIN1(_33369), .DIN2(_26350), .Q(_33368) );
  xnr2s1 _33223_inst ( .DIN1(_32615), .DIN2(_33370), .Q(_33369) );
  nnd2s1 _33224_inst ( .DIN1(_33371), .DIN2(_33372), .Q(
        _____________________________73________) );
  nor2s1 _33225_inst ( .DIN1(_33298), .DIN2(_33373), .Q(_33372) );
  nor2s1 _33226_inst ( .DIN1(_28100), .DIN2(_33374), .Q(_33373) );
  nnd2s1 _33227_inst ( .DIN1(_33375), .DIN2(_33352), .Q(_33374) );
  nnd2s1 _33228_inst ( .DIN1(_53328), .DIN2(_26550), .Q(_33352) );
  nnd2s1 _33229_inst ( .DIN1(_33376), .DIN2(_33377), .Q(_33375) );
  or2s1 _33230_inst ( .DIN1(_33300), .DIN2(_53333), .Q(_33377) );
  nnd2s1 _33231_inst ( .DIN1(_33378), .DIN2(_33365), .Q(_33300) );
  nnd2s1 _33232_inst ( .DIN1(_33362), .DIN2(_33378), .Q(_33376) );
  nor2s1 _33233_inst ( .DIN1(_26605), .DIN2(_33285), .Q(_33362) );
  hi1s1 _33234_inst ( .DIN(_33379), .Q(_33298) );
  nor2s1 _33235_inst ( .DIN1(_33380), .DIN2(_33381), .Q(_33371) );
  nor2s1 _33236_inst ( .DIN1(_33305), .DIN2(_33382), .Q(_33381) );
  nor2s1 _33237_inst ( .DIN1(_33383), .DIN2(_33384), .Q(_33382) );
  nor2s1 _33238_inst ( .DIN1(_53320), .DIN2(_53327), .Q(_33383) );
  nor2s1 _33239_inst ( .DIN1(_33309), .DIN2(_33385), .Q(_33380) );
  xor2s1 _33240_inst ( .DIN1(_26350), .DIN2(_33386), .Q(_33385) );
  nnd2s1 _33241_inst ( .DIN1(_33370), .DIN2(_33367), .Q(_33386) );
  nnd2s1 _33242_inst ( .DIN1(_33387), .DIN2(_33388), .Q(_33367) );
  nor2s1 _33243_inst ( .DIN1(_33389), .DIN2(_33390), .Q(_33387) );
  nor2s1 _33244_inst ( .DIN1(_53383), .DIN2(_33391), .Q(_33389) );
  nnd2s1 _33245_inst ( .DIN1(_33392), .DIN2(_33393), .Q(_33370) );
  nor2s1 _33246_inst ( .DIN1(_33394), .DIN2(_33391), .Q(_33392) );
  nor2s1 _33247_inst ( .DIN1(_33395), .DIN2(_33396), .Q(_33391) );
  hi1s1 _33248_inst ( .DIN(_33397), .Q(_33395) );
  nor2s1 _33249_inst ( .DIN1(_33390), .DIN2(_26237), .Q(_33394) );
  nor2s1 _33250_inst ( .DIN1(_33398), .DIN2(_33397), .Q(_33390) );
  nnd2s1 _33251_inst ( .DIN1(_33378), .DIN2(_33285), .Q(_33309) );
  nor2s1 _33252_inst ( .DIN1(_33399), .DIN2(_33361), .Q(_33378) );
  nor2s1 _33253_inst ( .DIN1(_33281), .DIN2(_33285), .Q(_33361) );
  nnd2s1 _33254_inst ( .DIN1(_33400), .DIN2(_33401), .Q(
        _____________________________72________) );
  nnd2s1 _33255_inst ( .DIN1(_33402), .DIN2(_33403), .Q(_33401) );
  nor2s1 _33256_inst ( .DIN1(_33404), .DIN2(_27774), .Q(_33402) );
  xor2s1 _33257_inst ( .DIN1(_26375), .DIN2(_53271), .Q(_33404) );
  nnd2s1 _33258_inst ( .DIN1(_33405), .DIN2(_28470), .Q(_33400) );
  nor2s1 _33259_inst ( .DIN1(_33406), .DIN2(_33407), .Q(_33405) );
  nor2s1 _33260_inst ( .DIN1(_33408), .DIN2(_33409), .Q(_33407) );
  nnd2s1 _33261_inst ( .DIN1(______[20]), .DIN2(_33410), .Q(_33409) );
  xor2s1 _33262_inst ( .DIN1(_26490), .DIN2(_33411), .Q(_33408) );
  nor2s1 _33263_inst ( .DIN1(_33412), .DIN2(_33413), .Q(_33406) );
  xor2s1 _33264_inst ( .DIN1(_33398), .DIN2(_33414), .Q(_33412) );
  xor2s1 _33265_inst ( .DIN1(_26237), .DIN2(_33397), .Q(_33414) );
  nnd2s1 _33266_inst ( .DIN1(_33415), .DIN2(_33416), .Q(_33397) );
  nnd2s1 _33267_inst ( .DIN1(_53161), .DIN2(_33417), .Q(_33416) );
  or2s1 _33268_inst ( .DIN1(_33418), .DIN2(_33419), .Q(_33417) );
  nnd2s1 _33269_inst ( .DIN1(_33419), .DIN2(_33418), .Q(_33415) );
  nnd2s1 _33270_inst ( .DIN1(_33420), .DIN2(_33421), .Q(
        _____________________________71________) );
  nnd2s1 _33271_inst ( .DIN1(_33422), .DIN2(_33423), .Q(_33421) );
  xor2s1 _33272_inst ( .DIN1(_53313), .DIN2(_53333), .Q(_33423) );
  nnd2s1 _33273_inst ( .DIN1(_33424), .DIN2(_33359), .Q(_33420) );
  nor2s1 _33274_inst ( .DIN1(_33425), .DIN2(_33426), .Q(_33424) );
  nor2s1 _33275_inst ( .DIN1(_33427), .DIN2(_33428), .Q(_33426) );
  nnd2s1 _33276_inst ( .DIN1(______[0]), .DIN2(_33410), .Q(_33428) );
  xor2s1 _33277_inst ( .DIN1(_26474), .DIN2(_33411), .Q(_33427) );
  nnd2s1 _33278_inst ( .DIN1(_53259), .DIN2(_53337), .Q(_33411) );
  nor2s1 _33279_inst ( .DIN1(_33429), .DIN2(_33413), .Q(_33425) );
  xor2s1 _33280_inst ( .DIN1(_33419), .DIN2(_33430), .Q(_33429) );
  xor2s1 _33281_inst ( .DIN1(_26384), .DIN2(_33418), .Q(_33430) );
  nnd2s1 _33282_inst ( .DIN1(_33431), .DIN2(_33432), .Q(_33418) );
  nnd2s1 _33283_inst ( .DIN1(_53072), .DIN2(_33433), .Q(_33432) );
  or2s1 _33284_inst ( .DIN1(_33434), .DIN2(_26831), .Q(_33433) );
  nnd2s1 _33285_inst ( .DIN1(_26831), .DIN2(_33434), .Q(_33431) );
  nnd2s1 _33286_inst ( .DIN1(_33436), .DIN2(_26993), .Q(
        _____________________________70________) );
  nor2s1 _33287_inst ( .DIN1(_33437), .DIN2(_33438), .Q(_33436) );
  nor2s1 _33288_inst ( .DIN1(_26996), .DIN2(_33439), .Q(_33438) );
  nnd2s1 _33289_inst ( .DIN1(_33440), .DIN2(_33441), .Q(_33439) );
  nnd2s1 _33290_inst ( .DIN1(_33442), .DIN2(_33443), .Q(_33440) );
  xnr2s1 _33291_inst ( .DIN1(_26831), .DIN2(_33444), .Q(_33443) );
  xnr2s1 _33292_inst ( .DIN1(_53072), .DIN2(_33434), .Q(_33444) );
  nnd2s1 _33293_inst ( .DIN1(_33445), .DIN2(_33446), .Q(_33434) );
  nnd2s1 _33294_inst ( .DIN1(_33447), .DIN2(_26232), .Q(_33446) );
  or2s1 _33295_inst ( .DIN1(_33448), .DIN2(_33449), .Q(_33447) );
  nnd2s1 _33296_inst ( .DIN1(_33449), .DIN2(_33448), .Q(_33445) );
  nor2s1 _33297_inst ( .DIN1(_27007), .DIN2(_33450), .Q(_33437) );
  nor2s1 _33298_inst ( .DIN1(_26853), .DIN2(_33451), .Q(_33450) );
  xor2s1 _33299_inst ( .DIN1(_53258), .DIN2(_53260), .Q(_33451) );
  nnd2s1 _33300_inst ( .DIN1(_33452), .DIN2(_33379), .Q(
        _____________________________6________) );
  nor2s1 _33301_inst ( .DIN1(_33453), .DIN2(_33454), .Q(_33452) );
  nor2s1 _33302_inst ( .DIN1(_33305), .DIN2(_33455), .Q(_33454) );
  xor2s1 _33303_inst ( .DIN1(_53035), .DIN2(_53103), .Q(_33455) );
  nor2s1 _33304_inst ( .DIN1(_33456), .DIN2(_33399), .Q(_33453) );
  nor2s1 _33305_inst ( .DIN1(_33457), .DIN2(_33458), .Q(_33456) );
  nor2s1 _33306_inst ( .DIN1(_33459), .DIN2(_33460), .Q(_33458) );
  xor2s1 _33307_inst ( .DIN1(_33461), .DIN2(_33462), .Q(_33459) );
  xnr2s1 _33308_inst ( .DIN1(_53012), .DIN2(_33463), .Q(_33462) );
  nor2s1 _33309_inst ( .DIN1(_33464), .DIN2(_33465), .Q(_33457) );
  nnd2s1 _33310_inst ( .DIN1(______[16]), .DIN2(_33466), .Q(_33465) );
  xor2s1 _33311_inst ( .DIN1(_53315), .DIN2(_33467), .Q(_33466) );
  nnd2s1 _33312_inst ( .DIN1(_33468), .DIN2(_33469), .Q(
        _____________________________69________) );
  nnd2s1 _33313_inst ( .DIN1(_29390), .DIN2(_33470), .Q(_33469) );
  xor2s1 _33314_inst ( .DIN1(_53267), .DIN2(_53268), .Q(_33470) );
  nnd2s1 _33315_inst ( .DIN1(_28250), .DIN2(_33471), .Q(_33468) );
  nnd2s1 _33316_inst ( .DIN1(_33472), .DIN2(_33473), .Q(_33471) );
  nnd2s1 _33317_inst ( .DIN1(_33442), .DIN2(_33474), .Q(_33473) );
  xor2s1 _33318_inst ( .DIN1(_33449), .DIN2(_33475), .Q(_33474) );
  xor2s1 _33319_inst ( .DIN1(_26232), .DIN2(_33448), .Q(_33475) );
  nnd2s1 _33320_inst ( .DIN1(_33476), .DIN2(_33477), .Q(_33448) );
  nnd2s1 _33321_inst ( .DIN1(_53287), .DIN2(_33478), .Q(_33477) );
  or2s1 _33322_inst ( .DIN1(_33479), .DIN2(_26833), .Q(_33478) );
  xor2s1 _33323_inst ( .DIN1(_31947), .DIN2(_33481), .Q(_33476) );
  nnd2s1 _33324_inst ( .DIN1(_26833), .DIN2(_33479), .Q(_33481) );
  nor2s1 _33325_inst ( .DIN1(_33482), .DIN2(_33483), .Q(_33472) );
  nor2s1 _33326_inst ( .DIN1(_26737), .DIN2(_33484), .Q(_33483) );
  or2s1 _33327_inst ( .DIN1(_33485), .DIN2(_53337), .Q(_33484) );
  nor2s1 _33328_inst ( .DIN1(_53259), .DIN2(_33441), .Q(_33482) );
  nnd2s1 _33329_inst ( .DIN1(_53337), .DIN2(_33410), .Q(_33441) );
  nnd2s1 _33330_inst ( .DIN1(_33486), .DIN2(_33487), .Q(
        _____________________________68________) );
  nnd2s1 _33331_inst ( .DIN1(_33488), .DIN2(_29555), .Q(_33487) );
  nnd2s1 _33332_inst ( .DIN1(_29556), .DIN2(_26424), .Q(_33488) );
  nor2s1 _33333_inst ( .DIN1(_33489), .DIN2(_27291), .Q(_29556) );
  nnd2s1 _33334_inst ( .DIN1(_33490), .DIN2(_29560), .Q(_33486) );
  nor2s1 _33335_inst ( .DIN1(_33491), .DIN2(_33492), .Q(_33490) );
  nor2s1 _33336_inst ( .DIN1(_33485), .DIN2(_33493), .Q(_33492) );
  xor2s1 _33337_inst ( .DIN1(_33494), .DIN2(_33495), .Q(_33493) );
  nnd2s1 _33338_inst ( .DIN1(_33496), .DIN2(_33497), .Q(_33494) );
  nnd2s1 _33339_inst ( .DIN1(_53014), .DIN2(_26220), .Q(_33497) );
  nor2s1 _33340_inst ( .DIN1(_33498), .DIN2(_33413), .Q(_33491) );
  xor2s1 _33341_inst ( .DIN1(_26833), .DIN2(_33499), .Q(_33498) );
  xor2s1 _33342_inst ( .DIN1(_26658), .DIN2(_33479), .Q(_33499) );
  nnd2s1 _33343_inst ( .DIN1(_33500), .DIN2(_33501), .Q(_33479) );
  nnd2s1 _33344_inst ( .DIN1(_53047), .DIN2(_33502), .Q(_33501) );
  or2s1 _33345_inst ( .DIN1(_33503), .DIN2(_33504), .Q(_33502) );
  nnd2s1 _33346_inst ( .DIN1(_33504), .DIN2(_33503), .Q(_33500) );
  nnd2s1 _33347_inst ( .DIN1(_33505), .DIN2(_33506), .Q(
        _____________________________67________) );
  nnd2s1 _33348_inst ( .DIN1(_27684), .DIN2(_33507), .Q(_33506) );
  nnd2s1 _33349_inst ( .DIN1(_33508), .DIN2(_33509), .Q(_33507) );
  nnd2s1 _33350_inst ( .DIN1(_33442), .DIN2(_33510), .Q(_33509) );
  xnr2s1 _33351_inst ( .DIN1(_33504), .DIN2(_33511), .Q(_33510) );
  xnr2s1 _33352_inst ( .DIN1(_53047), .DIN2(_33503), .Q(_33511) );
  nnd2s1 _33353_inst ( .DIN1(_33512), .DIN2(_33513), .Q(_33503) );
  nnd2s1 _33354_inst ( .DIN1(_33514), .DIN2(_33515), .Q(_33513) );
  nor2s1 _33355_inst ( .DIN1(_53013), .DIN2(_33516), .Q(_33514) );
  nor2s1 _33356_inst ( .DIN1(_52841), .DIN2(_33517), .Q(_33516) );
  nnd2s1 _33357_inst ( .DIN1(_52841), .DIN2(_33517), .Q(_33512) );
  hi1s1 _33358_inst ( .DIN(_33413), .Q(_33442) );
  nnd2s1 _33359_inst ( .DIN1(_33485), .DIN2(_33518), .Q(_33413) );
  hi1s1 _33360_inst ( .DIN(_33410), .Q(_33485) );
  nnd2s1 _33361_inst ( .DIN1(_53347), .DIN2(_33410), .Q(_33508) );
  nnd2s1 _33362_inst ( .DIN1(_33519), .DIN2(_33520), .Q(_33410) );
  nnd2s1 _33363_inst ( .DIN1(_33521), .DIN2(_27679), .Q(_33505) );
  nor2s1 _33364_inst ( .DIN1(_33522), .DIN2(_26607), .Q(_33521) );
  nnd2s1 _33365_inst ( .DIN1(_33523), .DIN2(_30601), .Q(
        _____________________________66________) );
  nor2s1 _33366_inst ( .DIN1(_33524), .DIN2(_33525), .Q(_33523) );
  nor2s1 _33367_inst ( .DIN1(_27392), .DIN2(_33526), .Q(_33525) );
  nnd2s1 _33368_inst ( .DIN1(_33527), .DIN2(_33528), .Q(_33526) );
  nor2s1 _33369_inst ( .DIN1(_33529), .DIN2(_33530), .Q(_33527) );
  nor2s1 _33370_inst ( .DIN1(_33531), .DIN2(_33532), .Q(_33530) );
  xor2s1 _33371_inst ( .DIN1(_33533), .DIN2(_33534), .Q(_33532) );
  xor2s1 _33372_inst ( .DIN1(_33535), .DIN2(_52841), .Q(_33533) );
  nnd2s1 _33373_inst ( .DIN1(_33515), .DIN2(_26554), .Q(_33535) );
  nor2s1 _33374_inst ( .DIN1(_33536), .DIN2(_33537), .Q(_33529) );
  nor2s1 _33375_inst ( .DIN1(_26220), .DIN2(_28100), .Q(_33537) );
  nor2s1 _33376_inst ( .DIN1(_27397), .DIN2(_33538), .Q(_33524) );
  xnr2s1 _33377_inst ( .DIN1(_52917), .DIN2(_30628), .Q(_33538) );
  nor2s1 _33378_inst ( .DIN1(_26493), .DIN2(_53441), .Q(_30628) );
  nnd2s1 _33379_inst ( .DIN1(_33539), .DIN2(_33540), .Q(
        _____________________________65________) );
  nnd2s1 _33380_inst ( .DIN1(_33541), .DIN2(_27749), .Q(_33540) );
  nnd2s1 _33381_inst ( .DIN1(_33542), .DIN2(______[0]), .Q(_33541) );
  nor2s1 _33382_inst ( .DIN1(_28296), .DIN2(_33543), .Q(_33542) );
  nor2s1 _33383_inst ( .DIN1(_53016), .DIN2(_53017), .Q(_33543) );
  nor2s1 _33384_inst ( .DIN1(_26473), .DIN2(_26251), .Q(_28296) );
  nor2s1 _33385_inst ( .DIN1(_33544), .DIN2(_33545), .Q(_33539) );
  nor2s1 _33386_inst ( .DIN1(_33546), .DIN2(_33547), .Q(_33545) );
  nor2s1 _33387_inst ( .DIN1(_33548), .DIN2(_27241), .Q(_33547) );
  nor2s1 _33388_inst ( .DIN1(_33549), .DIN2(_27749), .Q(_33548) );
  nor2s1 _33389_inst ( .DIN1(_33550), .DIN2(_33551), .Q(_33549) );
  nnd2s1 _33390_inst ( .DIN1(_33552), .DIN2(_33553), .Q(_33551) );
  nnd2s1 _33391_inst ( .DIN1(_33496), .DIN2(_26513), .Q(_33553) );
  nnd2s1 _33392_inst ( .DIN1(_53345), .DIN2(_26441), .Q(_33496) );
  nnd2s1 _33393_inst ( .DIN1(_33495), .DIN2(_26441), .Q(_33552) );
  nor2s1 _33394_inst ( .DIN1(_26513), .DIN2(_26220), .Q(_33495) );
  nor2s1 _33395_inst ( .DIN1(_33554), .DIN2(_33531), .Q(_33546) );
  xor2s1 _33396_inst ( .DIN1(_33515), .DIN2(_53013), .Q(_33554) );
  nnd2s1 _33397_inst ( .DIN1(_33555), .DIN2(_28811), .Q(
        _____________________________64________) );
  nor2s1 _33398_inst ( .DIN1(_33556), .DIN2(_33557), .Q(_33555) );
  nor2s1 _33399_inst ( .DIN1(_28814), .DIN2(_33558), .Q(_33557) );
  nnd2s1 _33400_inst ( .DIN1(_33559), .DIN2(_33560), .Q(_33558) );
  nnd2s1 _33401_inst ( .DIN1(_33561), .DIN2(_53354), .Q(_33560) );
  nor2s1 _33402_inst ( .DIN1(_33562), .DIN2(_33563), .Q(_33559) );
  nor2s1 _33403_inst ( .DIN1(_53208), .DIN2(_33564), .Q(_33563) );
  nor2s1 _33404_inst ( .DIN1(_33561), .DIN2(_33565), .Q(_33564) );
  nnd2s1 _33405_inst ( .DIN1(_33566), .DIN2(_33567), .Q(_33565) );
  nnd2s1 _33406_inst ( .DIN1(_32907), .DIN2(_33568), .Q(_33567) );
  nnd2s1 _33407_inst ( .DIN1(_33569), .DIN2(_32904), .Q(_33566) );
  and2s1 _33408_inst ( .DIN1(_33570), .DIN2(_26849), .Q(_33561) );
  nor2s1 _33409_inst ( .DIN1(_33571), .DIN2(_27241), .Q(_33570) );
  nor2s1 _33410_inst ( .DIN1(_33572), .DIN2(_26600), .Q(_33562) );
  nor2s1 _33411_inst ( .DIN1(_33573), .DIN2(_33574), .Q(_33572) );
  nnd2s1 _33412_inst ( .DIN1(_33575), .DIN2(_33576), .Q(_33574) );
  nnd2s1 _33413_inst ( .DIN1(_32904), .DIN2(_33568), .Q(_33576) );
  hi1s1 _33414_inst ( .DIN(_33577), .Q(_32904) );
  nnd2s1 _33415_inst ( .DIN1(_33569), .DIN2(_32907), .Q(_33575) );
  hi1s1 _33416_inst ( .DIN(_33578), .Q(_32907) );
  hi1s1 _33417_inst ( .DIN(_33568), .Q(_33569) );
  nnd2s1 _33418_inst ( .DIN1(_33579), .DIN2(_33580), .Q(_33568) );
  nnd2s1 _33419_inst ( .DIN1(_33581), .DIN2(_26663), .Q(_33580) );
  or2s1 _33420_inst ( .DIN1(_33582), .DIN2(_26850), .Q(_33581) );
  nnd2s1 _33421_inst ( .DIN1(_33582), .DIN2(_26850), .Q(_33579) );
  nor2s1 _33422_inst ( .DIN1(_33583), .DIN2(_33584), .Q(_33573) );
  nnd2s1 _33423_inst ( .DIN1(______[0]), .DIN2(_32920), .Q(_33584) );
  nnd2s1 _33424_inst ( .DIN1(_26850), .DIN2(_26451), .Q(_33583) );
  nor2s1 _33425_inst ( .DIN1(_53224), .DIN2(_28356), .Q(_33556) );
  nnd2s1 _33426_inst ( .DIN1(_33585), .DIN2(_33586), .Q(
        _____________________________63________) );
  nnd2s1 _33427_inst ( .DIN1(_33587), .DIN2(_33588), .Q(_33586) );
  xor2s1 _33428_inst ( .DIN1(_26432), .DIN2(_53430), .Q(_33588) );
  nor2s1 _33429_inst ( .DIN1(_27448), .DIN2(_33589), .Q(_33587) );
  nnd2s1 _33430_inst ( .DIN1(_33590), .DIN2(_27895), .Q(_33585) );
  nor2s1 _33431_inst ( .DIN1(_33591), .DIN2(_33592), .Q(_33590) );
  nor2s1 _33432_inst ( .DIN1(_53049), .DIN2(_33593), .Q(_33592) );
  nor2s1 _33433_inst ( .DIN1(_33594), .DIN2(_33595), .Q(_33591) );
  xor2s1 _33434_inst ( .DIN1(_33582), .DIN2(_33596), .Q(_33594) );
  xor2s1 _33435_inst ( .DIN1(_53018), .DIN2(_53384), .Q(_33596) );
  nnd2s1 _33436_inst ( .DIN1(_33597), .DIN2(_33598), .Q(_33582) );
  nnd2s1 _33437_inst ( .DIN1(_33599), .DIN2(_26639), .Q(_33598) );
  nnd2s1 _33438_inst ( .DIN1(_32914), .DIN2(_33600), .Q(_33599) );
  or2s1 _33439_inst ( .DIN1(_33600), .DIN2(_32914), .Q(_33597) );
  nnd2s1 _33440_inst ( .DIN1(_33601), .DIN2(_33602), .Q(
        _____________________________62________) );
  nnd2s1 _33441_inst ( .DIN1(_33603), .DIN2(_27875), .Q(_33602) );
  and2s1 _33442_inst ( .DIN1(_33604), .DIN2(_27929), .Q(_27875) );
  nnd2s1 _33443_inst ( .DIN1(_33605), .DIN2(_33606), .Q(_33604) );
  nor2s1 _33444_inst ( .DIN1(_27937), .DIN2(_27936), .Q(_33605) );
  nor2s1 _33445_inst ( .DIN1(_33607), .DIN2(_27393), .Q(_33603) );
  xnr2s1 _33446_inst ( .DIN1(_53074), .DIN2(_53019), .Q(_33607) );
  nnd2s1 _33447_inst ( .DIN1(_33608), .DIN2(_27868), .Q(_33601) );
  hi1s1 _33448_inst ( .DIN(_27929), .Q(_27868) );
  nnd2s1 _33449_inst ( .DIN1(_33609), .DIN2(_33610), .Q(_27929) );
  nor2s1 _33450_inst ( .DIN1(_33611), .DIN2(_33612), .Q(_33610) );
  nnd2s1 _33451_inst ( .DIN1(_33613), .DIN2(_33614), .Q(_33612) );
  nor2s1 _33452_inst ( .DIN1(_27934), .DIN2(_33615), .Q(_33609) );
  or2s1 _33453_inst ( .DIN1(_33616), .DIN2(_33617), .Q(_33615) );
  nor2s1 _33454_inst ( .DIN1(_33618), .DIN2(_33619), .Q(_33608) );
  nor2s1 _33455_inst ( .DIN1(_33620), .DIN2(_33621), .Q(_33619) );
  or2s1 _33456_inst ( .DIN1(_27614), .DIN2(_33593), .Q(_33621) );
  xor2s1 _33457_inst ( .DIN1(_26339), .DIN2(_33622), .Q(_33620) );
  nor2s1 _33458_inst ( .DIN1(_33623), .DIN2(_33595), .Q(_33618) );
  xor2s1 _33459_inst ( .DIN1(_33600), .DIN2(_33624), .Q(_33623) );
  xor2s1 _33460_inst ( .DIN1(_26639), .DIN2(_32914), .Q(_33624) );
  nnd2s1 _33461_inst ( .DIN1(_33625), .DIN2(_33626), .Q(_33600) );
  nnd2s1 _33462_inst ( .DIN1(_33627), .DIN2(_26253), .Q(_33626) );
  or2s1 _33463_inst ( .DIN1(_33628), .DIN2(_32935), .Q(_33627) );
  xor2s1 _33464_inst ( .DIN1(_29599), .DIN2(_33629), .Q(_33625) );
  nnd2s1 _33465_inst ( .DIN1(_32935), .DIN2(_33628), .Q(_33629) );
  nnd2s1 _33466_inst ( .DIN1(_33630), .DIN2(_31127), .Q(
        _____________________________61________) );
  nnd2s1 _33467_inst ( .DIN1(_28733), .DIN2(_33489), .Q(_31127) );
  nor2s1 _33468_inst ( .DIN1(_33631), .DIN2(_33632), .Q(_33630) );
  nor2s1 _33469_inst ( .DIN1(_28733), .DIN2(_33633), .Q(_33632) );
  nnd2s1 _33470_inst ( .DIN1(_33634), .DIN2(_33635), .Q(_33633) );
  nnd2s1 _33471_inst ( .DIN1(_33636), .DIN2(_33637), .Q(_33635) );
  xor2s1 _33472_inst ( .DIN1(_32935), .DIN2(_33638), .Q(_33636) );
  xor2s1 _33473_inst ( .DIN1(_26253), .DIN2(_33628), .Q(_33638) );
  nnd2s1 _33474_inst ( .DIN1(_33639), .DIN2(_33640), .Q(_33628) );
  nnd2s1 _33475_inst ( .DIN1(_53022), .DIN2(_33641), .Q(_33640) );
  xor2s1 _33476_inst ( .DIN1(_31925), .DIN2(_33642), .Q(_33641) );
  nnd2s1 _33477_inst ( .DIN1(_33643), .DIN2(______[0]), .Q(_33634) );
  nor2s1 _33478_inst ( .DIN1(_33644), .DIN2(_33645), .Q(_33643) );
  nor2s1 _33479_inst ( .DIN1(_33646), .DIN2(_33647), .Q(_33645) );
  nor2s1 _33480_inst ( .DIN1(_33593), .DIN2(_26346), .Q(_33646) );
  nor2s1 _33481_inst ( .DIN1(_33648), .DIN2(_33649), .Q(_33644) );
  hi1s1 _33482_inst ( .DIN(_33647), .Q(_33649) );
  xor2s1 _33483_inst ( .DIN1(_26376), .DIN2(_33650), .Q(_33647) );
  nor2s1 _33484_inst ( .DIN1(_53020), .DIN2(_28738), .Q(_33631) );
  nnd2s1 _33485_inst ( .DIN1(_27325), .DIN2(_33651), .Q(
        _____________________________60________) );
  nnd2s1 _33486_inst ( .DIN1(_33652), .DIN2(_33653), .Q(_33651) );
  nnd2s1 _33487_inst ( .DIN1(_33654), .DIN2(_53021), .Q(_33653) );
  nor2s1 _33488_inst ( .DIN1(_33593), .DIN2(_26773), .Q(_33654) );
  nnd2s1 _33489_inst ( .DIN1(_33637), .DIN2(_33655), .Q(_33652) );
  xnr2s1 _33490_inst ( .DIN1(_53022), .DIN2(_33656), .Q(_33655) );
  nnd2s1 _33491_inst ( .DIN1(_33639), .DIN2(_33642), .Q(_33656) );
  nnd2s1 _33492_inst ( .DIN1(_33657), .DIN2(_32973), .Q(_33642) );
  nor2s1 _33493_inst ( .DIN1(_33658), .DIN2(_33659), .Q(_33657) );
  nor2s1 _33494_inst ( .DIN1(_53066), .DIN2(_33660), .Q(_33658) );
  nnd2s1 _33495_inst ( .DIN1(_33661), .DIN2(_32951), .Q(_33639) );
  nor2s1 _33496_inst ( .DIN1(_33662), .DIN2(_33660), .Q(_33661) );
  nor2s1 _33497_inst ( .DIN1(_32979), .DIN2(_33663), .Q(_33660) );
  nor2s1 _33498_inst ( .DIN1(_33659), .DIN2(_26563), .Q(_33662) );
  nor2s1 _33499_inst ( .DIN1(_33664), .DIN2(_32994), .Q(_33659) );
  hi1s1 _33500_inst ( .DIN(_33663), .Q(_33664) );
  nnd2s1 _33501_inst ( .DIN1(_33665), .DIN2(_33666), .Q(
        _____________________________5________) );
  nnd2s1 _33502_inst ( .DIN1(_33667), .DIN2(_33039), .Q(_33666) );
  nor2s1 _33503_inst ( .DIN1(_27039), .DIN2(_26695), .Q(_33667) );
  nnd2s1 _33504_inst ( .DIN1(_33668), .DIN2(_32837), .Q(_33665) );
  nor2s1 _33505_inst ( .DIN1(_33669), .DIN2(_33670), .Q(_33668) );
  nor2s1 _33506_inst ( .DIN1(_33671), .DIN2(_33460), .Q(_33670) );
  xor2s1 _33507_inst ( .DIN1(_33672), .DIN2(_33673), .Q(_33671) );
  xnr2s1 _33508_inst ( .DIN1(_33674), .DIN2(_33675), .Q(_33673) );
  xor2s1 _33509_inst ( .DIN1(_53023), .DIN2(_31925), .Q(_33672) );
  nor2s1 _33510_inst ( .DIN1(_33676), .DIN2(_33677), .Q(_33669) );
  nnd2s1 _33511_inst ( .DIN1(_33678), .DIN2(______[30]), .Q(_33677) );
  xor2s1 _33512_inst ( .DIN1(_53041), .DIN2(_33467), .Q(_33676) );
  nnd2s1 _33513_inst ( .DIN1(_33679), .DIN2(_33680), .Q(
        _____________________________59________) );
  nnd2s1 _33514_inst ( .DIN1(_33681), .DIN2(_33149), .Q(_33680) );
  nnd2s1 _33515_inst ( .DIN1(_33682), .DIN2(_53222), .Q(_33681) );
  nor2s1 _33516_inst ( .DIN1(_33683), .DIN2(_27291), .Q(_33682) );
  nnd2s1 _33517_inst ( .DIN1(_33684), .DIN2(_33132), .Q(_33679) );
  nor2s1 _33518_inst ( .DIN1(_33648), .DIN2(_33685), .Q(_33684) );
  nor2s1 _33519_inst ( .DIN1(_33595), .DIN2(_33686), .Q(_33685) );
  nnd2s1 _33520_inst ( .DIN1(_33687), .DIN2(_33688), .Q(_33686) );
  nnd2s1 _33521_inst ( .DIN1(_33689), .DIN2(_26563), .Q(_33688) );
  xor2s1 _33522_inst ( .DIN1(_33663), .DIN2(_32979), .Q(_33689) );
  nnd2s1 _33523_inst ( .DIN1(_33690), .DIN2(_53066), .Q(_33687) );
  xor2s1 _33524_inst ( .DIN1(_33663), .DIN2(_32994), .Q(_33690) );
  nnd2s1 _33525_inst ( .DIN1(_33691), .DIN2(_33692), .Q(_33663) );
  nnd2s1 _33526_inst ( .DIN1(_53330), .DIN2(_33693), .Q(_33692) );
  or2s1 _33527_inst ( .DIN1(_33694), .DIN2(_33000), .Q(_33693) );
  nnd2s1 _33528_inst ( .DIN1(_33000), .DIN2(_33694), .Q(_33691) );
  nor2s1 _33529_inst ( .DIN1(_33593), .DIN2(_53024), .Q(_33648) );
  nnd2s1 _33530_inst ( .DIN1(_33695), .DIN2(_29181), .Q(
        _____________________________58________) );
  or2s1 _33531_inst ( .DIN1(_33696), .DIN2(_29206), .Q(_29181) );
  nor2s1 _33532_inst ( .DIN1(_33697), .DIN2(_33698), .Q(_33695) );
  nor2s1 _33533_inst ( .DIN1(_29184), .DIN2(_33699), .Q(_33698) );
  nnd2s1 _33534_inst ( .DIN1(_33700), .DIN2(_33701), .Q(_33699) );
  nnd2s1 _33535_inst ( .DIN1(_33702), .DIN2(_33637), .Q(_33701) );
  hi1s1 _33536_inst ( .DIN(_33595), .Q(_33637) );
  xor2s1 _33537_inst ( .DIN1(_33703), .DIN2(_33000), .Q(_33702) );
  xor2s1 _33538_inst ( .DIN1(_33694), .DIN2(_53330), .Q(_33703) );
  nnd2s1 _33539_inst ( .DIN1(_33704), .DIN2(_33705), .Q(_33694) );
  nnd2s1 _33540_inst ( .DIN1(_33706), .DIN2(_26480), .Q(_33705) );
  or2s1 _33541_inst ( .DIN1(_33707), .DIN2(_26828), .Q(_33706) );
  nnd2s1 _33542_inst ( .DIN1(_33017), .DIN2(_33707), .Q(_33704) );
  nnd2s1 _33543_inst ( .DIN1(_33708), .DIN2(_33709), .Q(_33700) );
  nor2s1 _33544_inst ( .DIN1(_33593), .DIN2(_33710), .Q(_33709) );
  nor2s1 _33545_inst ( .DIN1(_53223), .DIN2(_33711), .Q(_33710) );
  nor2s1 _33546_inst ( .DIN1(_53322), .DIN2(_53024), .Q(_33711) );
  nor2s1 _33547_inst ( .DIN1(_33712), .DIN2(_27393), .Q(_33708) );
  nor2s1 _33548_inst ( .DIN1(_53322), .DIN2(_33650), .Q(_33712) );
  nnd2s1 _33549_inst ( .DIN1(_53223), .DIN2(_26346), .Q(_33650) );
  nor2s1 _33550_inst ( .DIN1(_29206), .DIN2(_33713), .Q(_33697) );
  xor2s1 _33551_inst ( .DIN1(_33714), .DIN2(_26342), .Q(_33713) );
  nnd2s1 _33552_inst ( .DIN1(_33715), .DIN2(_33716), .Q(
        _____________________________57________) );
  nor2s1 _33553_inst ( .DIN1(_33717), .DIN2(_33718), .Q(_33716) );
  nor2s1 _33554_inst ( .DIN1(_29828), .DIN2(_33719), .Q(_33718) );
  nor2s1 _33555_inst ( .DIN1(_33720), .DIN2(_33721), .Q(_33719) );
  nor2s1 _33556_inst ( .DIN1(_33722), .DIN2(_33723), .Q(_33721) );
  xor2s1 _33557_inst ( .DIN1(_33017), .DIN2(_33724), .Q(_33723) );
  xor2s1 _33558_inst ( .DIN1(_26480), .DIN2(_33707), .Q(_33724) );
  nnd2s1 _33559_inst ( .DIN1(_33725), .DIN2(_33726), .Q(_33707) );
  nnd2s1 _33560_inst ( .DIN1(_53026), .DIN2(_33727), .Q(_33726) );
  or2s1 _33561_inst ( .DIN1(_33728), .DIN2(_33035), .Q(_33727) );
  nnd2s1 _33562_inst ( .DIN1(_33035), .DIN2(_33728), .Q(_33725) );
  nor2s1 _33563_inst ( .DIN1(_33729), .DIN2(_33730), .Q(_33720) );
  nor2s1 _33564_inst ( .DIN1(_27365), .DIN2(_33731), .Q(_33730) );
  nnd2s1 _33565_inst ( .DIN1(_33732), .DIN2(_33733), .Q(_33731) );
  xor2s1 _33566_inst ( .DIN1(_33734), .DIN2(_33735), .Q(_33732) );
  xor2s1 _33567_inst ( .DIN1(_53203), .DIN2(_53243), .Q(_33735) );
  nnd2s1 _33568_inst ( .DIN1(_53028), .DIN2(_53149), .Q(_33734) );
  nor2s1 _33569_inst ( .DIN1(_29849), .DIN2(_33736), .Q(_33717) );
  nnd2s1 _33570_inst ( .DIN1(_53025), .DIN2(_33737), .Q(_33736) );
  nor2s1 _33571_inst ( .DIN1(_29853), .DIN2(_33738), .Q(_33715) );
  nor2s1 _33572_inst ( .DIN1(_53025), .DIN2(_29855), .Q(_33738) );
  nnd2s1 _33573_inst ( .DIN1(_29852), .DIN2(_29828), .Q(_29855) );
  hi1s1 _33574_inst ( .DIN(_33737), .Q(_29852) );
  nnd2s1 _33575_inst ( .DIN1(_53147), .DIN2(_53149), .Q(_33737) );
  hi1s1 _33576_inst ( .DIN(_33094), .Q(_29853) );
  nnd2s1 _33577_inst ( .DIN1(_33739), .DIN2(_33740), .Q(
        _____________________________56________) );
  nnd2s1 _33578_inst ( .DIN1(_33741), .DIN2(_30853), .Q(_33740) );
  nnd2s1 _33579_inst ( .DIN1(_33742), .DIN2(______[16]), .Q(_33741) );
  nor2s1 _33580_inst ( .DIN1(_33743), .DIN2(_33744), .Q(_33742) );
  xor2s1 _33581_inst ( .DIN1(_53240), .DIN2(_26394), .Q(_33744) );
  nnd2s1 _33582_inst ( .DIN1(_33745), .DIN2(_30856), .Q(_33739) );
  nnd2s1 _33583_inst ( .DIN1(_33746), .DIN2(_33747), .Q(_33745) );
  nnd2s1 _33584_inst ( .DIN1(_33748), .DIN2(_33722), .Q(_33747) );
  nor2s1 _33585_inst ( .DIN1(_26485), .DIN2(_33749), .Q(_33748) );
  nnd2s1 _33586_inst ( .DIN1(______[6]), .DIN2(_33733), .Q(_33749) );
  nnd2s1 _33587_inst ( .DIN1(_33750), .DIN2(_33729), .Q(_33746) );
  xor2s1 _33588_inst ( .DIN1(_33751), .DIN2(_33752), .Q(_33750) );
  xnr2s1 _33589_inst ( .DIN1(_53026), .DIN2(_33728), .Q(_33752) );
  nnd2s1 _33590_inst ( .DIN1(_33753), .DIN2(_33754), .Q(_33728) );
  nnd2s1 _33591_inst ( .DIN1(_53112), .DIN2(_33755), .Q(_33754) );
  or2s1 _33592_inst ( .DIN1(_33756), .DIN2(_26800), .Q(_33755) );
  nnd2s1 _33593_inst ( .DIN1(_33065), .DIN2(_33756), .Q(_33753) );
  hi1s1 _33594_inst ( .DIN(_33035), .Q(_33751) );
  nnd2s1 _33595_inst ( .DIN1(_33757), .DIN2(_28010), .Q(
        _____________________________55________) );
  nor2s1 _33596_inst ( .DIN1(_33758), .DIN2(_33759), .Q(_33757) );
  nor2s1 _33597_inst ( .DIN1(_33760), .DIN2(_33722), .Q(_33759) );
  xor2s1 _33598_inst ( .DIN1(_33082), .DIN2(_33761), .Q(_33760) );
  xnr2s1 _33599_inst ( .DIN1(_53112), .DIN2(_33756), .Q(_33761) );
  nnd2s1 _33600_inst ( .DIN1(_33762), .DIN2(_33763), .Q(_33756) );
  nnd2s1 _33601_inst ( .DIN1(_33764), .DIN2(_26348), .Q(_33763) );
  or2s1 _33602_inst ( .DIN1(_33765), .DIN2(_33088), .Q(_33764) );
  nnd2s1 _33603_inst ( .DIN1(_33088), .DIN2(_33765), .Q(_33762) );
  hi1s1 _33604_inst ( .DIN(_33065), .Q(_33082) );
  nor2s1 _33605_inst ( .DIN1(_33729), .DIN2(_33766), .Q(_33758) );
  nor2s1 _33606_inst ( .DIN1(_26366), .DIN2(_33767), .Q(_33766) );
  nnd2s1 _33607_inst ( .DIN1(______[16]), .DIN2(_33733), .Q(_33767) );
  nnd2s1 _33608_inst ( .DIN1(_33768), .DIN2(_33769), .Q(
        _____________________________54________) );
  nnd2s1 _33609_inst ( .DIN1(_33770), .DIN2(_27717), .Q(_33769) );
  nor2s1 _33610_inst ( .DIN1(_33771), .DIN2(_27611), .Q(_27717) );
  nor2s1 _33611_inst ( .DIN1(_33772), .DIN2(_27774), .Q(_33770) );
  xor2s1 _33612_inst ( .DIN1(_33773), .DIN2(_33774), .Q(_33772) );
  xor2s1 _33613_inst ( .DIN1(_53027), .DIN2(_53200), .Q(_33774) );
  nnd2s1 _33614_inst ( .DIN1(_53111), .DIN2(_53200), .Q(_33773) );
  nnd2s1 _33615_inst ( .DIN1(_33775), .DIN2(_27611), .Q(_33768) );
  nor2s1 _33616_inst ( .DIN1(_33776), .DIN2(_33777), .Q(_33775) );
  nor2s1 _33617_inst ( .DIN1(_33722), .DIN2(_33778), .Q(_33777) );
  xor2s1 _33618_inst ( .DIN1(_33103), .DIN2(_33779), .Q(_33778) );
  xor2s1 _33619_inst ( .DIN1(_26348), .DIN2(_33765), .Q(_33779) );
  nnd2s1 _33620_inst ( .DIN1(_33780), .DIN2(_33781), .Q(_33765) );
  nnd2s1 _33621_inst ( .DIN1(_53399), .DIN2(_33782), .Q(_33781) );
  or2s1 _33622_inst ( .DIN1(_33783), .DIN2(_26797), .Q(_33782) );
  nnd2s1 _33623_inst ( .DIN1(_33108), .DIN2(_33783), .Q(_33780) );
  nor2s1 _33624_inst ( .DIN1(_33729), .DIN2(_33784), .Q(_33776) );
  nnd2s1 _33625_inst ( .DIN1(_33785), .DIN2(______[28]), .Q(_33784) );
  nor2s1 _33626_inst ( .DIN1(_33786), .DIN2(_33787), .Q(_33785) );
  xor2s1 _33627_inst ( .DIN1(_53028), .DIN2(_26366), .Q(_33787) );
  nnd2s1 _33628_inst ( .DIN1(_33788), .DIN2(_27560), .Q(
        _____________________________53________) );
  nor2s1 _33629_inst ( .DIN1(_33789), .DIN2(_33790), .Q(_33788) );
  nor2s1 _33630_inst ( .DIN1(_27563), .DIN2(_33791), .Q(_33790) );
  nor2s1 _33631_inst ( .DIN1(_33792), .DIN2(_33793), .Q(_33791) );
  nor2s1 _33632_inst ( .DIN1(_33794), .DIN2(_33722), .Q(_33793) );
  xor2s1 _33633_inst ( .DIN1(_33123), .DIN2(_33795), .Q(_33794) );
  xor2s1 _33634_inst ( .DIN1(_26362), .DIN2(_33783), .Q(_33795) );
  nnd2s1 _33635_inst ( .DIN1(_33796), .DIN2(_33797), .Q(_33783) );
  nnd2s1 _33636_inst ( .DIN1(_33798), .DIN2(_26244), .Q(_33797) );
  or2s1 _33637_inst ( .DIN1(_33799), .DIN2(_33129), .Q(_33798) );
  nnd2s1 _33638_inst ( .DIN1(_33129), .DIN2(_33799), .Q(_33796) );
  nor2s1 _33639_inst ( .DIN1(_33729), .DIN2(_33800), .Q(_33792) );
  nor2s1 _33640_inst ( .DIN1(_33786), .DIN2(_33801), .Q(_33800) );
  xor2s1 _33641_inst ( .DIN1(_26380), .DIN2(_33802), .Q(_33801) );
  nnd2s1 _33642_inst ( .DIN1(_53427), .DIN2(_26352), .Q(_33802) );
  nor2s1 _33643_inst ( .DIN1(_27571), .DIN2(_33803), .Q(_33789) );
  nor2s1 _33644_inst ( .DIN1(_33804), .DIN2(_28684), .Q(_33803) );
  xor2s1 _33645_inst ( .DIN1(_33805), .DIN2(_53071), .Q(_33804) );
  nnd2s1 _33646_inst ( .DIN1(_53029), .DIN2(_53106), .Q(_33805) );
  nnd2s1 _33647_inst ( .DIN1(_33806), .DIN2(_33807), .Q(
        _____________________________52________) );
  nnd2s1 _33648_inst ( .DIN1(_33808), .DIN2(_33809), .Q(_33807) );
  nnd2s1 _33649_inst ( .DIN1(_33810), .DIN2(_33811), .Q(_33809) );
  nnd2s1 _33650_inst ( .DIN1(_33786), .DIN2(_33722), .Q(_33811) );
  xor2s1 _33651_inst ( .DIN1(_27329), .DIN2(_33812), .Q(_33810) );
  nnd2s1 _33652_inst ( .DIN1(_33813), .DIN2(_33814), .Q(_33812) );
  nnd2s1 _33653_inst ( .DIN1(_33815), .DIN2(_33722), .Q(_33814) );
  hi1s1 _33654_inst ( .DIN(_33729), .Q(_33722) );
  nor2s1 _33655_inst ( .DIN1(_33816), .DIN2(_27448), .Q(_33815) );
  xnr2s1 _33656_inst ( .DIN1(_53029), .DIN2(_53427), .Q(_33816) );
  nnd2s1 _33657_inst ( .DIN1(_33817), .DIN2(_33729), .Q(_33813) );
  nor2s1 _33658_inst ( .DIN1(_33818), .DIN2(_33276), .Q(_33729) );
  nnd2s1 _33659_inst ( .DIN1(_33819), .DIN2(_33820), .Q(_33276) );
  nor2s1 _33660_inst ( .DIN1(_33821), .DIN2(_33822), .Q(_33820) );
  nor2s1 _33661_inst ( .DIN1(_33823), .DIN2(_33824), .Q(_33819) );
  nnd2s1 _33662_inst ( .DIN1(_33139), .DIN2(_33825), .Q(_33818) );
  xor2s1 _33663_inst ( .DIN1(_33129), .DIN2(_33826), .Q(_33817) );
  xor2s1 _33664_inst ( .DIN1(_26244), .DIN2(_33799), .Q(_33826) );
  nnd2s1 _33665_inst ( .DIN1(_33827), .DIN2(_33828), .Q(_33799) );
  nnd2s1 _33666_inst ( .DIN1(_33829), .DIN2(_26404), .Q(_33828) );
  or2s1 _33667_inst ( .DIN1(_33830), .DIN2(_26832), .Q(_33829) );
  nnd2s1 _33668_inst ( .DIN1(_26832), .DIN2(_33830), .Q(_33827) );
  nnd2s1 _33669_inst ( .DIN1(_33831), .DIN2(_53042), .Q(_33806) );
  nnd2s1 _33670_inst ( .DIN1(_33832), .DIN2(_33833), .Q(
        _____________________________51________) );
  nnd2s1 _33671_inst ( .DIN1(_33834), .DIN2(_29082), .Q(_33833) );
  xor2s1 _33672_inst ( .DIN1(_33835), .DIN2(_53417), .Q(_33834) );
  nnd2s1 _33673_inst ( .DIN1(_29083), .DIN2(_33836), .Q(_33832) );
  nnd2s1 _33674_inst ( .DIN1(_33837), .DIN2(_33838), .Q(_33836) );
  nnd2s1 _33675_inst ( .DIN1(_33839), .DIN2(_33840), .Q(_33838) );
  hi1s1 _33676_inst ( .DIN(_33841), .Q(_33840) );
  xor2s1 _33677_inst ( .DIN1(_33147), .DIN2(_33842), .Q(_33839) );
  xor2s1 _33678_inst ( .DIN1(_26404), .DIN2(_33830), .Q(_33842) );
  nnd2s1 _33679_inst ( .DIN1(_33843), .DIN2(_33844), .Q(_33830) );
  nnd2s1 _33680_inst ( .DIN1(_53227), .DIN2(_33845), .Q(_33844) );
  or2s1 _33681_inst ( .DIN1(_33846), .DIN2(_33178), .Q(_33845) );
  nnd2s1 _33682_inst ( .DIN1(_33178), .DIN2(_33846), .Q(_33843) );
  nnd2s1 _33683_inst ( .DIN1(_33847), .DIN2(_26352), .Q(_33837) );
  nnd2s1 _33684_inst ( .DIN1(_33848), .DIN2(_33379), .Q(
        _____________________________50________) );
  nor2s1 _33685_inst ( .DIN1(_33849), .DIN2(_33850), .Q(_33848) );
  nor2s1 _33686_inst ( .DIN1(_33305), .DIN2(_33851), .Q(_33850) );
  nor2s1 _33687_inst ( .DIN1(_28646), .DIN2(_33852), .Q(_33851) );
  xor2s1 _33688_inst ( .DIN1(_53334), .DIN2(_33384), .Q(_33852) );
  nor2s1 _33689_inst ( .DIN1(_26520), .DIN2(_26267), .Q(_33384) );
  nor2s1 _33690_inst ( .DIN1(_33853), .DIN2(_33399), .Q(_33849) );
  nor2s1 _33691_inst ( .DIN1(_33854), .DIN2(_33855), .Q(_33853) );
  nor2s1 _33692_inst ( .DIN1(_33856), .DIN2(_33857), .Q(_33855) );
  xor2s1 _33693_inst ( .DIN1(_53031), .DIN2(_53427), .Q(_33857) );
  nor2s1 _33694_inst ( .DIN1(_33841), .DIN2(_33858), .Q(_33854) );
  xor2s1 _33695_inst ( .DIN1(_33178), .DIN2(_33859), .Q(_33858) );
  xor2s1 _33696_inst ( .DIN1(_26371), .DIN2(_33846), .Q(_33859) );
  nnd2s1 _33697_inst ( .DIN1(_33860), .DIN2(_33861), .Q(_33846) );
  nnd2s1 _33698_inst ( .DIN1(_33862), .DIN2(_26379), .Q(_33861) );
  or2s1 _33699_inst ( .DIN1(_33863), .DIN2(_33196), .Q(_33862) );
  nnd2s1 _33700_inst ( .DIN1(_33196), .DIN2(_33863), .Q(_33860) );
  nor2s1 _33701_inst ( .DIN1(_31037), .DIN2(_33864), .Q(
        _____________________________4________) );
  xor2s1 _33702_inst ( .DIN1(_33865), .DIN2(_33866), .Q(_33864) );
  nnd2s1 _33703_inst ( .DIN1(_33867), .DIN2(_33868), .Q(_33866) );
  nnd2s1 _33704_inst ( .DIN1(_33869), .DIN2(_33678), .Q(_33868) );
  nor2s1 _33705_inst ( .DIN1(_53042), .DIN2(_27365), .Q(_33869) );
  nnd2s1 _33706_inst ( .DIN1(_33870), .DIN2(_33871), .Q(_33867) );
  xor2s1 _33707_inst ( .DIN1(_33872), .DIN2(_33873), .Q(_33870) );
  xor2s1 _33708_inst ( .DIN1(_26479), .DIN2(_33874), .Q(_33873) );
  nnd2s1 _33709_inst ( .DIN1(_33875), .DIN2(_28794), .Q(
        _____________________________49________) );
  nor2s1 _33710_inst ( .DIN1(_33876), .DIN2(_33877), .Q(_33875) );
  nor2s1 _33711_inst ( .DIN1(_33878), .DIN2(_28801), .Q(_33877) );
  nor2s1 _33712_inst ( .DIN1(_33879), .DIN2(_33880), .Q(_33878) );
  nor2s1 _33713_inst ( .DIN1(_33881), .DIN2(_33841), .Q(_33880) );
  xor2s1 _33714_inst ( .DIN1(_33882), .DIN2(_33883), .Q(_33881) );
  xor2s1 _33715_inst ( .DIN1(_26379), .DIN2(_33863), .Q(_33883) );
  nnd2s1 _33716_inst ( .DIN1(_33884), .DIN2(_33885), .Q(_33863) );
  nnd2s1 _33717_inst ( .DIN1(_53228), .DIN2(_33886), .Q(_33885) );
  or2s1 _33718_inst ( .DIN1(_33887), .DIN2(_33213), .Q(_33886) );
  nnd2s1 _33719_inst ( .DIN1(_33213), .DIN2(_33887), .Q(_33884) );
  nor2s1 _33720_inst ( .DIN1(_27448), .DIN2(_33888), .Q(_33879) );
  nnd2s1 _33721_inst ( .DIN1(_33889), .DIN2(_33847), .Q(_33888) );
  xnr2s1 _33722_inst ( .DIN1(_53113), .DIN2(_33890), .Q(_33889) );
  nor2s1 _33723_inst ( .DIN1(_28797), .DIN2(_33891), .Q(_33876) );
  nor2s1 _33724_inst ( .DIN1(_33892), .DIN2(_28799), .Q(_33891) );
  nor2s1 _33725_inst ( .DIN1(_26525), .DIN2(_26259), .Q(_28799) );
  nor2s1 _33726_inst ( .DIN1(_53030), .DIN2(_53039), .Q(_33892) );
  nnd2s1 _33727_inst ( .DIN1(_33893), .DIN2(_33894), .Q(
        _____________________________48________) );
  nor2s1 _33728_inst ( .DIN1(_33895), .DIN2(_33896), .Q(_33893) );
  nor2s1 _33729_inst ( .DIN1(_33897), .DIN2(_33898), .Q(_33896) );
  nor2s1 _33730_inst ( .DIN1(_33899), .DIN2(_33900), .Q(_33897) );
  nor2s1 _33731_inst ( .DIN1(_33901), .DIN2(_33841), .Q(_33900) );
  xor2s1 _33732_inst ( .DIN1(_33213), .DIN2(_33902), .Q(_33901) );
  xnr2s1 _33733_inst ( .DIN1(_53228), .DIN2(_33887), .Q(_33902) );
  nnd2s1 _33734_inst ( .DIN1(_33903), .DIN2(_33904), .Q(_33887) );
  nnd2s1 _33735_inst ( .DIN1(_53231), .DIN2(_33905), .Q(_33904) );
  or2s1 _33736_inst ( .DIN1(_33906), .DIN2(_33907), .Q(_33905) );
  nnd2s1 _33737_inst ( .DIN1(_33907), .DIN2(_33906), .Q(_33903) );
  nor2s1 _33738_inst ( .DIN1(_27066), .DIN2(_33908), .Q(_33899) );
  nnd2s1 _33739_inst ( .DIN1(_33909), .DIN2(_33847), .Q(_33908) );
  xnr2s1 _33740_inst ( .DIN1(_53010), .DIN2(_33890), .Q(_33909) );
  nor2s1 _33741_inst ( .DIN1(_33808), .DIN2(_33910), .Q(_33895) );
  nor2s1 _33742_inst ( .DIN1(_33911), .DIN2(_28100), .Q(_33910) );
  xor2s1 _33743_inst ( .DIN1(_26352), .DIN2(_53042), .Q(_33911) );
  nnd2s1 _33744_inst ( .DIN1(_33912), .DIN2(_27183), .Q(
        _____________________________47________) );
  nor2s1 _33745_inst ( .DIN1(_33913), .DIN2(_33914), .Q(_33912) );
  nor2s1 _33746_inst ( .DIN1(_33856), .DIN2(_26675), .Q(_33914) );
  hi1s1 _33747_inst ( .DIN(_33847), .Q(_33856) );
  nor2s1 _33748_inst ( .DIN1(_33915), .DIN2(_33841), .Q(_33913) );
  xor2s1 _33749_inst ( .DIN1(_26775), .DIN2(_33916), .Q(_33915) );
  xnr2s1 _33750_inst ( .DIN1(_53231), .DIN2(_33906), .Q(_33916) );
  nnd2s1 _33751_inst ( .DIN1(_33917), .DIN2(_33918), .Q(_33906) );
  nnd2s1 _33752_inst ( .DIN1(_53034), .DIN2(_33919), .Q(_33918) );
  or2s1 _33753_inst ( .DIN1(_33920), .DIN2(_26834), .Q(_33919) );
  nnd2s1 _33754_inst ( .DIN1(_26834), .DIN2(_33920), .Q(_33917) );
  nnd2s1 _33755_inst ( .DIN1(_33921), .DIN2(_33922), .Q(
        _____________________________46________) );
  nnd2s1 _33756_inst ( .DIN1(_33923), .DIN2(_33053), .Q(_33922) );
  nnd2s1 _33757_inst ( .DIN1(_29039), .DIN2(_53112), .Q(_33923) );
  nnd2s1 _33758_inst ( .DIN1(_33924), .DIN2(_33069), .Q(_33921) );
  nor2s1 _33759_inst ( .DIN1(_33925), .DIN2(_33926), .Q(_33924) );
  nor2s1 _33760_inst ( .DIN1(_33927), .DIN2(_33841), .Q(_33926) );
  nnd2s1 _33761_inst ( .DIN1(_33928), .DIN2(_33929), .Q(_33841) );
  nor2s1 _33762_inst ( .DIN1(_33930), .DIN2(_33823), .Q(_33929) );
  hi1s1 _33763_inst ( .DIN(_33931), .Q(_33823) );
  nor2s1 _33764_inst ( .DIN1(_33932), .DIN2(_33595), .Q(_33928) );
  nnd2s1 _33765_inst ( .DIN1(_33593), .DIN2(_33933), .Q(_33595) );
  nor2s1 _33766_inst ( .DIN1(_33847), .DIN2(_33934), .Q(_33593) );
  xor2s1 _33767_inst ( .DIN1(_26834), .DIN2(_33935), .Q(_33927) );
  xnr2s1 _33768_inst ( .DIN1(_53034), .DIN2(_33920), .Q(_33935) );
  nnd2s1 _33769_inst ( .DIN1(_33936), .DIN2(_33937), .Q(_33920) );
  nnd2s1 _33770_inst ( .DIN1(_33938), .DIN2(_26521), .Q(_33937) );
  or2s1 _33771_inst ( .DIN1(_33939), .DIN2(_33271), .Q(_33938) );
  nnd2s1 _33772_inst ( .DIN1(_33271), .DIN2(_33939), .Q(_33936) );
  nor2s1 _33773_inst ( .DIN1(_33940), .DIN2(_33941), .Q(_33925) );
  nnd2s1 _33774_inst ( .DIN1(_26860), .DIN2(_33942), .Q(_33941) );
  nnd2s1 _33775_inst ( .DIN1(_26675), .DIN2(_26307), .Q(_33942) );
  nnd2s1 _33776_inst ( .DIN1(_33847), .DIN2(_33890), .Q(_33940) );
  nnd2s1 _33777_inst ( .DIN1(_53033), .DIN2(_53032), .Q(_33890) );
  nnd2s1 _33778_inst ( .DIN1(_33943), .DIN2(_33786), .Q(_33847) );
  hi1s1 _33779_inst ( .DIN(_33733), .Q(_33786) );
  nnd2s1 _33780_inst ( .DIN1(_33944), .DIN2(_33825), .Q(_33733) );
  nor2s1 _33781_inst ( .DIN1(_33945), .DIN2(_33824), .Q(_33944) );
  nor2s1 _33782_inst ( .DIN1(_33946), .DIN2(_33275), .Q(_33943) );
  nnd2s1 _33783_inst ( .DIN1(_33947), .DIN2(_33948), .Q(
        _____________________________45________) );
  nnd2s1 _33784_inst ( .DIN1(_33949), .DIN2(_33053), .Q(_33948) );
  nnd2s1 _33785_inst ( .DIN1(_33950), .DIN2(_33951), .Q(_33949) );
  nor2s1 _33786_inst ( .DIN1(_33952), .DIN2(_33953), .Q(_33950) );
  nor2s1 _33787_inst ( .DIN1(_53112), .DIN2(_53113), .Q(_33953) );
  hi1s1 _33788_inst ( .DIN(_27574), .Q(_33952) );
  nnd2s1 _33789_inst ( .DIN1(_33954), .DIN2(_33069), .Q(_33947) );
  nor2s1 _33790_inst ( .DIN1(_33955), .DIN2(_33956), .Q(_33954) );
  nor2s1 _33791_inst ( .DIN1(_33957), .DIN2(_33958), .Q(_33956) );
  xor2s1 _33792_inst ( .DIN1(_53244), .DIN2(_33959), .Q(_33957) );
  nor2s1 _33793_inst ( .DIN1(_33960), .DIN2(_33961), .Q(_33955) );
  xnr2s1 _33794_inst ( .DIN1(_33271), .DIN2(_33962), .Q(_33960) );
  xor2s1 _33795_inst ( .DIN1(_26521), .DIN2(_33939), .Q(_33962) );
  nnd2s1 _33796_inst ( .DIN1(_33963), .DIN2(_33964), .Q(_33939) );
  nnd2s1 _33797_inst ( .DIN1(_33965), .DIN2(_26290), .Q(_33964) );
  nnd2s1 _33798_inst ( .DIN1(_33966), .DIN2(_33310), .Q(_33965) );
  nnd2s1 _33799_inst ( .DIN1(_33291), .DIN2(_33967), .Q(_33963) );
  nnd2s1 _33800_inst ( .DIN1(_33968), .DIN2(_33894), .Q(
        _____________________________44________) );
  nor2s1 _33801_inst ( .DIN1(_33969), .DIN2(_33970), .Q(_33968) );
  nor2s1 _33802_inst ( .DIN1(_33898), .DIN2(_33971), .Q(_33970) );
  nnd2s1 _33803_inst ( .DIN1(_33972), .DIN2(_33973), .Q(_33971) );
  nor2s1 _33804_inst ( .DIN1(_33974), .DIN2(_33975), .Q(_33972) );
  nor2s1 _33805_inst ( .DIN1(_33961), .DIN2(_33976), .Q(_33975) );
  xor2s1 _33806_inst ( .DIN1(_33310), .DIN2(_33977), .Q(_33976) );
  xor2s1 _33807_inst ( .DIN1(_26290), .DIN2(_33966), .Q(_33977) );
  hi1s1 _33808_inst ( .DIN(_33967), .Q(_33966) );
  nnd2s1 _33809_inst ( .DIN1(_33978), .DIN2(_33979), .Q(_33967) );
  nnd2s1 _33810_inst ( .DIN1(_33980), .DIN2(_26650), .Q(_33979) );
  or2s1 _33811_inst ( .DIN1(_33981), .DIN2(_26822), .Q(_33980) );
  nnd2s1 _33812_inst ( .DIN1(_33982), .DIN2(_33981), .Q(_33978) );
  nor2s1 _33813_inst ( .DIN1(_33983), .DIN2(_33984), .Q(_33974) );
  nor2s1 _33814_inst ( .DIN1(_26774), .DIN2(_33985), .Q(_33984) );
  xor2s1 _33815_inst ( .DIN1(_26374), .DIN2(_33959), .Q(_33985) );
  nor2s1 _33816_inst ( .DIN1(_33808), .DIN2(_33986), .Q(_33969) );
  nor2s1 _33817_inst ( .DIN1(_27241), .DIN2(_33987), .Q(_33986) );
  xor2s1 _33818_inst ( .DIN1(_53047), .DIN2(_33988), .Q(_33987) );
  nnd2s1 _33819_inst ( .DIN1(_33989), .DIN2(_33990), .Q(
        _____________________________43________) );
  nnd2s1 _33820_inst ( .DIN1(_33991), .DIN2(_53279), .Q(_33990) );
  nor2s1 _33821_inst ( .DIN1(_33992), .DIN2(_27614), .Q(_33991) );
  nnd2s1 _33822_inst ( .DIN1(_28356), .DIN2(_33993), .Q(_33989) );
  nnd2s1 _33823_inst ( .DIN1(_33994), .DIN2(_33995), .Q(_33993) );
  nnd2s1 _33824_inst ( .DIN1(_33996), .DIN2(_33983), .Q(_33995) );
  xor2s1 _33825_inst ( .DIN1(_33982), .DIN2(_33997), .Q(_33996) );
  xor2s1 _33826_inst ( .DIN1(_26650), .DIN2(_33981), .Q(_33997) );
  nnd2s1 _33827_inst ( .DIN1(_33998), .DIN2(_33999), .Q(_33981) );
  nnd2s1 _33828_inst ( .DIN1(_53036), .DIN2(_34000), .Q(_33999) );
  nnd2s1 _33829_inst ( .DIN1(_34001), .DIN2(_33333), .Q(_34000) );
  nnd2s1 _33830_inst ( .DIN1(_33344), .DIN2(_34002), .Q(_33998) );
  nnd2s1 _33831_inst ( .DIN1(_34003), .DIN2(_26590), .Q(_33994) );
  nnd2s1 _33832_inst ( .DIN1(_34004), .DIN2(_34005), .Q(
        _____________________________42________) );
  nnd2s1 _33833_inst ( .DIN1(_34006), .DIN2(_33053), .Q(_34005) );
  nnd2s1 _33834_inst ( .DIN1(_29039), .DIN2(_34007), .Q(_34006) );
  xor2s1 _33835_inst ( .DIN1(_53197), .DIN2(_53261), .Q(_34007) );
  nnd2s1 _33836_inst ( .DIN1(_34008), .DIN2(_33069), .Q(_34004) );
  nor2s1 _33837_inst ( .DIN1(_34009), .DIN2(_34010), .Q(_34008) );
  nor2s1 _33838_inst ( .DIN1(_34011), .DIN2(_34012), .Q(_34010) );
  nnd2s1 _33839_inst ( .DIN1(_34003), .DIN2(_26864), .Q(_34012) );
  hi1s1 _33840_inst ( .DIN(_33958), .Q(_34003) );
  nnd2s1 _33841_inst ( .DIN1(_33961), .DIN2(_34013), .Q(_33958) );
  nnd2s1 _33842_inst ( .DIN1(_34014), .DIN2(_34015), .Q(_34013) );
  hi1s1 _33843_inst ( .DIN(_34016), .Q(_34015) );
  nor2s1 _33844_inst ( .DIN1(_34017), .DIN2(_33824), .Q(_34014) );
  nnd2s1 _33845_inst ( .DIN1(_34018), .DIN2(_33959), .Q(_34011) );
  nnd2s1 _33846_inst ( .DIN1(_53278), .DIN2(_26590), .Q(_33959) );
  nnd2s1 _33847_inst ( .DIN1(_53037), .DIN2(_26529), .Q(_34018) );
  nor2s1 _33848_inst ( .DIN1(_33961), .DIN2(_34019), .Q(_34009) );
  xor2s1 _33849_inst ( .DIN1(_34020), .DIN2(_34021), .Q(_34019) );
  xor2s1 _33850_inst ( .DIN1(_33344), .DIN2(_34001), .Q(_34021) );
  hi1s1 _33851_inst ( .DIN(_34002), .Q(_34001) );
  nnd2s1 _33852_inst ( .DIN1(_34022), .DIN2(_34023), .Q(_34002) );
  nnd2s1 _33853_inst ( .DIN1(_53209), .DIN2(_34024), .Q(_34023) );
  or2s1 _33854_inst ( .DIN1(_34025), .DIN2(_26801), .Q(_34024) );
  nnd2s1 _33855_inst ( .DIN1(_33349), .DIN2(_34025), .Q(_34022) );
  xor2s1 _33856_inst ( .DIN1(_34026), .DIN2(_53036), .Q(_34020) );
  nnd2s1 _33857_inst ( .DIN1(_34027), .DIN2(_34028), .Q(
        _____________________________41________) );
  nnd2s1 _33858_inst ( .DIN1(_33808), .DIN2(_34029), .Q(_34028) );
  nnd2s1 _33859_inst ( .DIN1(_34030), .DIN2(_33973), .Q(_34029) );
  nor2s1 _33860_inst ( .DIN1(_34031), .DIN2(_34032), .Q(_34030) );
  nor2s1 _33861_inst ( .DIN1(_33961), .DIN2(_34033), .Q(_34032) );
  xor2s1 _33862_inst ( .DIN1(_34034), .DIN2(_34035), .Q(_34033) );
  xnr2s1 _33863_inst ( .DIN1(_53209), .DIN2(_34025), .Q(_34035) );
  nnd2s1 _33864_inst ( .DIN1(_34036), .DIN2(_34037), .Q(_34025) );
  nnd2s1 _33865_inst ( .DIN1(_34038), .DIN2(_26695), .Q(_34037) );
  nnd2s1 _33866_inst ( .DIN1(_34039), .DIN2(_33393), .Q(_34038) );
  nnd2s1 _33867_inst ( .DIN1(_33388), .DIN2(_34040), .Q(_34036) );
  nor2s1 _33868_inst ( .DIN1(_33983), .DIN2(_34041), .Q(_34031) );
  xor2s1 _33869_inst ( .DIN1(_34042), .DIN2(_34043), .Q(_34041) );
  xor2s1 _33870_inst ( .DIN1(_53072), .DIN2(_53383), .Q(_34043) );
  nnd2s1 _33871_inst ( .DIN1(_34044), .DIN2(_33831), .Q(_34027) );
  nor2s1 _33872_inst ( .DIN1(_34045), .DIN2(_28646), .Q(_34044) );
  xor2s1 _33873_inst ( .DIN1(_26232), .DIN2(_53037), .Q(_34045) );
  nnd2s1 _33874_inst ( .DIN1(_34046), .DIN2(_34047), .Q(
        _____________________________40________) );
  nnd2s1 _33875_inst ( .DIN1(_28098), .DIN2(_34048), .Q(_34047) );
  nnd2s1 _33876_inst ( .DIN1(_34049), .DIN2(_34050), .Q(_34048) );
  nor2s1 _33877_inst ( .DIN1(_34051), .DIN2(_34052), .Q(_34050) );
  nor2s1 _33878_inst ( .DIN1(_34053), .DIN2(_33961), .Q(_34052) );
  nor2s1 _33879_inst ( .DIN1(_34054), .DIN2(_31842), .Q(_34053) );
  xor2s1 _33880_inst ( .DIN1(_33393), .DIN2(_34055), .Q(_34054) );
  xor2s1 _33881_inst ( .DIN1(_53038), .DIN2(_34039), .Q(_34055) );
  hi1s1 _33882_inst ( .DIN(_34040), .Q(_34039) );
  nnd2s1 _33883_inst ( .DIN1(_34056), .DIN2(_34057), .Q(_34040) );
  nnd2s1 _33884_inst ( .DIN1(_34058), .DIN2(_26259), .Q(_34057) );
  or2s1 _33885_inst ( .DIN1(_34059), .DIN2(_26802), .Q(_34058) );
  nnd2s1 _33886_inst ( .DIN1(_26802), .DIN2(_34059), .Q(_34056) );
  nor2s1 _33887_inst ( .DIN1(_33983), .DIN2(_34060), .Q(_34051) );
  nnd2s1 _33888_inst ( .DIN1(_34061), .DIN2(_34062), .Q(_34060) );
  nor2s1 _33889_inst ( .DIN1(_34063), .DIN2(_34064), .Q(_34049) );
  nor2s1 _33890_inst ( .DIN1(_34061), .DIN2(_34062), .Q(_34064) );
  nnd2s1 _33891_inst ( .DIN1(______[22]), .DIN2(_26350), .Q(_34062) );
  hi1s1 _33892_inst ( .DIN(_31842), .Q(_34061) );
  hi1s1 _33893_inst ( .DIN(_33973), .Q(_34063) );
  nnd2s1 _33894_inst ( .DIN1(_34065), .DIN2(_34066), .Q(_33973) );
  nor2s1 _33895_inst ( .DIN1(_33983), .DIN2(_34017), .Q(_34066) );
  hi1s1 _33896_inst ( .DIN(_33961), .Q(_33983) );
  nnd2s1 _33897_inst ( .DIN1(_34067), .DIN2(_33933), .Q(_33961) );
  nor2s1 _33898_inst ( .DIN1(_33930), .DIN2(_33824), .Q(_34067) );
  nor2s1 _33899_inst ( .DIN1(_33824), .DIN2(_34016), .Q(_34065) );
  nnd2s1 _33900_inst ( .DIN1(_34068), .DIN2(_28095), .Q(_34046) );
  nor2s1 _33901_inst ( .DIN1(_28646), .DIN2(_34069), .Q(_34068) );
  nnd2s1 _33902_inst ( .DIN1(_28857), .DIN2(_26211), .Q(_34069) );
  nnd2s1 _33903_inst ( .DIN1(_34070), .DIN2(_34071), .Q(
        _____________________________3________) );
  nor2s1 _33904_inst ( .DIN1(_34072), .DIN2(_34073), .Q(_34071) );
  nor2s1 _33905_inst ( .DIN1(_28533), .DIN2(_34074), .Q(_34073) );
  nnd2s1 _33906_inst ( .DIN1(_34075), .DIN2(_33460), .Q(_34074) );
  nnd2s1 _33907_inst ( .DIN1(_34076), .DIN2(_34077), .Q(_34075) );
  nor2s1 _33908_inst ( .DIN1(_27761), .DIN2(_33467), .Q(_34077) );
  and2s1 _33909_inst ( .DIN1(_53043), .DIN2(_26446), .Q(_33467) );
  nor2s1 _33910_inst ( .DIN1(_34078), .DIN2(_27774), .Q(_34076) );
  nor2s1 _33911_inst ( .DIN1(_53043), .DIN2(_26446), .Q(_34078) );
  nor2s1 _33912_inst ( .DIN1(_28542), .DIN2(_34079), .Q(_34072) );
  xor2s1 _33913_inst ( .DIN1(_52877), .DIN2(_53325), .Q(_34079) );
  nor2s1 _33914_inst ( .DIN1(_34080), .DIN2(_34081), .Q(_34070) );
  nor2s1 _33915_inst ( .DIN1(_34082), .DIN2(_34083), .Q(_34081) );
  xor2s1 _33916_inst ( .DIN1(_34084), .DIN2(_34085), .Q(_34083) );
  xor2s1 _33917_inst ( .DIN1(_26399), .DIN2(_34086), .Q(_34085) );
  hi1s1 _33918_inst ( .DIN(_28530), .Q(_34080) );
  nnd2s1 _33919_inst ( .DIN1(_34087), .DIN2(_34088), .Q(
        _____________________________39________) );
  nnd2s1 _33920_inst ( .DIN1(_34089), .DIN2(______[4]), .Q(_34088) );
  nor2s1 _33921_inst ( .DIN1(_34090), .DIN2(_34091), .Q(_34089) );
  xor2s1 _33922_inst ( .DIN1(_26235), .DIN2(_53162), .Q(_34091) );
  nnd2s1 _33923_inst ( .DIN1(_28792), .DIN2(_34092), .Q(_34087) );
  nnd2s1 _33924_inst ( .DIN1(_34093), .DIN2(_34094), .Q(_34092) );
  nnd2s1 _33925_inst ( .DIN1(_34095), .DIN2(_34096), .Q(_34094) );
  xor2s1 _33926_inst ( .DIN1(_33398), .DIN2(_34097), .Q(_34095) );
  xor2s1 _33927_inst ( .DIN1(_26259), .DIN2(_34059), .Q(_34097) );
  nnd2s1 _33928_inst ( .DIN1(_34098), .DIN2(_34099), .Q(_34059) );
  nnd2s1 _33929_inst ( .DIN1(_34100), .DIN2(_26673), .Q(_34099) );
  nnd2s1 _33930_inst ( .DIN1(_34101), .DIN2(_34102), .Q(_34100) );
  nnd2s1 _33931_inst ( .DIN1(_33419), .DIN2(_34103), .Q(_34098) );
  or2s1 _33932_inst ( .DIN1(_34104), .DIN2(_26237), .Q(_34093) );
  nnd2s1 _33933_inst ( .DIN1(_34105), .DIN2(_33335), .Q(
        _____________________________38________) );
  nor2s1 _33934_inst ( .DIN1(_34106), .DIN2(_34107), .Q(_34105) );
  nor2s1 _33935_inst ( .DIN1(_33338), .DIN2(_34108), .Q(_34107) );
  nor2s1 _33936_inst ( .DIN1(_34109), .DIN2(_34110), .Q(_34108) );
  nor2s1 _33937_inst ( .DIN1(_34111), .DIN2(_34112), .Q(_34110) );
  xor2s1 _33938_inst ( .DIN1(_33419), .DIN2(_34113), .Q(_34112) );
  xor2s1 _33939_inst ( .DIN1(_53041), .DIN2(_34101), .Q(_34113) );
  hi1s1 _33940_inst ( .DIN(_34103), .Q(_34101) );
  nnd2s1 _33941_inst ( .DIN1(_34114), .DIN2(_34115), .Q(_34103) );
  nnd2s1 _33942_inst ( .DIN1(_34116), .DIN2(_26446), .Q(_34115) );
  or2s1 _33943_inst ( .DIN1(_34117), .DIN2(_26831), .Q(_34116) );
  nnd2s1 _33944_inst ( .DIN1(_26831), .DIN2(_34117), .Q(_34114) );
  nor2s1 _33945_inst ( .DIN1(_34096), .DIN2(_34118), .Q(_34109) );
  nor2s1 _33946_inst ( .DIN1(_34119), .DIN2(_34120), .Q(_34118) );
  nnd2s1 _33947_inst ( .DIN1(______[16]), .DIN2(_34121), .Q(_34120) );
  nnd2s1 _33948_inst ( .DIN1(_34042), .DIN2(_53072), .Q(_34121) );
  nor2s1 _33949_inst ( .DIN1(_26237), .DIN2(_26384), .Q(_34042) );
  nnd2s1 _33950_inst ( .DIN1(_34122), .DIN2(_34016), .Q(_34119) );
  nnd2s1 _33951_inst ( .DIN1(_34123), .DIN2(_26384), .Q(_34122) );
  nnd2s1 _33952_inst ( .DIN1(_53383), .DIN2(_53072), .Q(_34123) );
  nor2s1 _33953_inst ( .DIN1(_30175), .DIN2(_34124), .Q(_34106) );
  xor2s1 _33954_inst ( .DIN1(_53040), .DIN2(_53328), .Q(_34124) );
  nnd2s1 _33955_inst ( .DIN1(_34125), .DIN2(_33894), .Q(
        _____________________________37________) );
  nnd2s1 _33956_inst ( .DIN1(_34126), .DIN2(_33898), .Q(_33894) );
  nor2s1 _33957_inst ( .DIN1(_34127), .DIN2(_34128), .Q(_34125) );
  nor2s1 _33958_inst ( .DIN1(_34129), .DIN2(_33898), .Q(_34128) );
  nor2s1 _33959_inst ( .DIN1(_34130), .DIN2(_34131), .Q(_34129) );
  nor2s1 _33960_inst ( .DIN1(_34111), .DIN2(_34132), .Q(_34131) );
  xnr2s1 _33961_inst ( .DIN1(_26831), .DIN2(_34133), .Q(_34132) );
  xor2s1 _33962_inst ( .DIN1(_26446), .DIN2(_34117), .Q(_34133) );
  nnd2s1 _33963_inst ( .DIN1(_34134), .DIN2(_34135), .Q(_34117) );
  nnd2s1 _33964_inst ( .DIN1(_53043), .DIN2(_34136), .Q(_34135) );
  nnd2s1 _33965_inst ( .DIN1(_34137), .DIN2(_34138), .Q(_34136) );
  nnd2s1 _33966_inst ( .DIN1(_34139), .DIN2(_33449), .Q(_34134) );
  hi1s1 _33967_inst ( .DIN(_34137), .Q(_34139) );
  nor2s1 _33968_inst ( .DIN1(_34104), .DIN2(_34140), .Q(_34130) );
  nnd2s1 _33969_inst ( .DIN1(______[22]), .DIN2(_34141), .Q(_34140) );
  xor2s1 _33970_inst ( .DIN1(_52841), .DIN2(_53047), .Q(_34141) );
  nor2s1 _33971_inst ( .DIN1(_33808), .DIN2(_34142), .Q(_34127) );
  nor2s1 _33972_inst ( .DIN1(_27393), .DIN2(_26350), .Q(_34142) );
  nnd2s1 _33973_inst ( .DIN1(_34143), .DIN2(_34144), .Q(
        _____________________________36________) );
  nnd2s1 _33974_inst ( .DIN1(_34145), .DIN2(_30856), .Q(_34144) );
  nor2s1 _33975_inst ( .DIN1(_34146), .DIN2(_34147), .Q(_34145) );
  nor2s1 _33976_inst ( .DIN1(_34111), .DIN2(_34148), .Q(_34147) );
  xor2s1 _33977_inst ( .DIN1(_34137), .DIN2(_34149), .Q(_34148) );
  xor2s1 _33978_inst ( .DIN1(_53043), .DIN2(_33449), .Q(_34149) );
  xnr2s1 _33979_inst ( .DIN1(_34150), .DIN2(_34151), .Q(_34137) );
  nnd2s1 _33980_inst ( .DIN1(_34152), .DIN2(_34153), .Q(_34150) );
  nnd2s1 _33981_inst ( .DIN1(_53315), .DIN2(_34154), .Q(_34153) );
  or2s1 _33982_inst ( .DIN1(_34155), .DIN2(_26833), .Q(_34154) );
  nnd2s1 _33983_inst ( .DIN1(_26833), .DIN2(_34155), .Q(_34152) );
  nor2s1 _33984_inst ( .DIN1(_34096), .DIN2(_34156), .Q(_34146) );
  nnd2s1 _33985_inst ( .DIN1(_34157), .DIN2(_34016), .Q(_34156) );
  xor2s1 _33986_inst ( .DIN1(_34158), .DIN2(_53048), .Q(_34157) );
  nnd2s1 _33987_inst ( .DIN1(_53287), .DIN2(_53047), .Q(_34158) );
  nnd2s1 _33988_inst ( .DIN1(_34159), .DIN2(_31056), .Q(_34143) );
  and2s1 _33989_inst ( .DIN1(_34160), .DIN2(______[14]), .Q(_31056) );
  xor2s1 _33990_inst ( .DIN1(_26366), .DIN2(_34161), .Q(_34159) );
  nor2s1 _33991_inst ( .DIN1(_53287), .DIN2(_53285), .Q(_34161) );
  nnd2s1 _33992_inst ( .DIN1(_34162), .DIN2(_34163), .Q(
        _____________________________35________) );
  nnd2s1 _33993_inst ( .DIN1(_34164), .DIN2(_33808), .Q(_34163) );
  nor2s1 _33994_inst ( .DIN1(_34165), .DIN2(_34166), .Q(_34164) );
  nor2s1 _33995_inst ( .DIN1(_34167), .DIN2(_34111), .Q(_34166) );
  xor2s1 _33996_inst ( .DIN1(_26833), .DIN2(_34168), .Q(_34167) );
  xor2s1 _33997_inst ( .DIN1(_26602), .DIN2(_34155), .Q(_34168) );
  nnd2s1 _33998_inst ( .DIN1(_34169), .DIN2(_34170), .Q(_34155) );
  nnd2s1 _33999_inst ( .DIN1(_34171), .DIN2(_34172), .Q(_34170) );
  nor2s1 _34000_inst ( .DIN1(_53049), .DIN2(_34173), .Q(_34171) );
  nor2s1 _34001_inst ( .DIN1(_53080), .DIN2(_33504), .Q(_34173) );
  nnd2s1 _34002_inst ( .DIN1(_33504), .DIN2(_53080), .Q(_34169) );
  nor2s1 _34003_inst ( .DIN1(_34104), .DIN2(_34174), .Q(_34165) );
  nnd2s1 _34004_inst ( .DIN1(_53287), .DIN2(______[26]), .Q(_34174) );
  nnd2s1 _34005_inst ( .DIN1(_34175), .DIN2(_33831), .Q(_34162) );
  nor2s1 _34006_inst ( .DIN1(_33808), .DIN2(_34126), .Q(_33831) );
  nor2s1 _34007_inst ( .DIN1(_33988), .DIN2(_34176), .Q(_34175) );
  nor2s1 _34008_inst ( .DIN1(_53044), .DIN2(_53048), .Q(_34176) );
  nor2s1 _34009_inst ( .DIN1(_26232), .DIN2(_26350), .Q(_33988) );
  nnd2s1 _34010_inst ( .DIN1(_34177), .DIN2(_34178), .Q(
        _____________________________34________) );
  nnd2s1 _34011_inst ( .DIN1(_34179), .DIN2(______[2]), .Q(_34178) );
  nor2s1 _34012_inst ( .DIN1(_32183), .DIN2(_34180), .Q(_34179) );
  xor2s1 _34013_inst ( .DIN1(_53046), .DIN2(_26429), .Q(_34180) );
  nnd2s1 _34014_inst ( .DIN1(_28056), .DIN2(_34181), .Q(_34177) );
  nnd2s1 _34015_inst ( .DIN1(_34182), .DIN2(_34183), .Q(_34181) );
  nnd2s1 _34016_inst ( .DIN1(_34184), .DIN2(_34185), .Q(_34183) );
  xor2s1 _34017_inst ( .DIN1(_26232), .DIN2(_53047), .Q(_34185) );
  nor2s1 _34018_inst ( .DIN1(_26774), .DIN2(_34104), .Q(_34184) );
  nnd2s1 _34019_inst ( .DIN1(_34111), .DIN2(_34016), .Q(_34104) );
  nnd2s1 _34020_inst ( .DIN1(_34186), .DIN2(_34096), .Q(_34182) );
  hi1s1 _34021_inst ( .DIN(_34111), .Q(_34096) );
  nnd2s1 _34022_inst ( .DIN1(_34187), .DIN2(_34188), .Q(_34111) );
  nor2s1 _34023_inst ( .DIN1(_33275), .DIN2(_34189), .Q(_34188) );
  nnd2s1 _34024_inst ( .DIN1(_34190), .DIN2(_34191), .Q(_34189) );
  nor2s1 _34025_inst ( .DIN1(_33100), .DIN2(_34192), .Q(_34187) );
  nnd2s1 _34026_inst ( .DIN1(_33825), .DIN2(_33931), .Q(_34192) );
  nnd2s1 _34027_inst ( .DIN1(_33933), .DIN2(_34193), .Q(_33100) );
  nor2s1 _34028_inst ( .DIN1(_34017), .DIN2(_33821), .Q(_33933) );
  xnr2s1 _34029_inst ( .DIN1(_34194), .DIN2(_33504), .Q(_34186) );
  xor2s1 _34030_inst ( .DIN1(_34195), .DIN2(_53080), .Q(_34194) );
  nnd2s1 _34031_inst ( .DIN1(_33517), .DIN2(_26719), .Q(_34195) );
  nnd2s1 _34032_inst ( .DIN1(_34196), .DIN2(_34197), .Q(
        _____________________________33________) );
  nnd2s1 _34033_inst ( .DIN1(_28010), .DIN2(_34198), .Q(_34197) );
  nnd2s1 _34034_inst ( .DIN1(_34199), .DIN2(_34200), .Q(_34198) );
  nnd2s1 _34035_inst ( .DIN1(_32929), .DIN2(_34201), .Q(_34200) );
  xor2s1 _34036_inst ( .DIN1(_53049), .DIN2(_33534), .Q(_34201) );
  nor2s1 _34037_inst ( .DIN1(_34202), .DIN2(_33236), .Q(_32929) );
  nnd2s1 _34038_inst ( .DIN1(_34203), .DIN2(_33274), .Q(_33236) );
  nor2s1 _34039_inst ( .DIN1(_33934), .DIN2(_33946), .Q(_33274) );
  nor2s1 _34040_inst ( .DIN1(_33932), .DIN2(_34016), .Q(_34203) );
  nnd2s1 _34041_inst ( .DIN1(_34204), .DIN2(_34190), .Q(_34016) );
  nnd2s1 _34042_inst ( .DIN1(_34205), .DIN2(_34193), .Q(_34202) );
  nor2s1 _34043_inst ( .DIN1(_34206), .DIN2(_34207), .Q(_34199) );
  nor2s1 _34044_inst ( .DIN1(_34208), .DIN2(_32943), .Q(_34207) );
  nnd2s1 _34045_inst ( .DIN1(_53280), .DIN2(_32936), .Q(_32943) );
  hi1s1 _34046_inst ( .DIN(_34209), .Q(_34208) );
  nor2s1 _34047_inst ( .DIN1(_34209), .DIN2(_34210), .Q(_34206) );
  nnd2s1 _34048_inst ( .DIN1(_32936), .DIN2(_26367), .Q(_34210) );
  nnd2s1 _34049_inst ( .DIN1(_34211), .DIN2(_34193), .Q(_32936) );
  xor2s1 _34050_inst ( .DIN1(_32968), .DIN2(_53283), .Q(_34209) );
  nor2s1 _34051_inst ( .DIN1(_26367), .DIN2(_53462), .Q(_32968) );
  nnd2s1 _34052_inst ( .DIN1(_34212), .DIN2(_34213), .Q(_34196) );
  nnd2s1 _34053_inst ( .DIN1(_34214), .DIN2(_34215), .Q(_34213) );
  xor2s1 _34054_inst ( .DIN1(_26347), .DIN2(_34216), .Q(_34212) );
  nor2s1 _34055_inst ( .DIN1(_53188), .DIN2(_26258), .Q(_34216) );
  nnd2s1 _34056_inst ( .DIN1(_34217), .DIN2(_34218), .Q(
        _____________________________32________) );
  nnd2s1 _34057_inst ( .DIN1(_28010), .DIN2(_34219), .Q(_34218) );
  nnd2s1 _34058_inst ( .DIN1(_34220), .DIN2(_34221), .Q(_34219) );
  nnd2s1 _34059_inst ( .DIN1(_34222), .DIN2(_34223), .Q(_34221) );
  nnd2s1 _34060_inst ( .DIN1(_34224), .DIN2(_32920), .Q(_34222) );
  xor2s1 _34061_inst ( .DIN1(_26487), .DIN2(_53354), .Q(_34224) );
  nor2s1 _34062_inst ( .DIN1(_34225), .DIN2(_34226), .Q(_34220) );
  nor2s1 _34063_inst ( .DIN1(_34227), .DIN2(_26669), .Q(_34226) );
  nor2s1 _34064_inst ( .DIN1(_34228), .DIN2(_34229), .Q(_34227) );
  nor2s1 _34065_inst ( .DIN1(_33577), .DIN2(_34230), .Q(_34229) );
  nor2s1 _34066_inst ( .DIN1(_34231), .DIN2(_33578), .Q(_34228) );
  nor2s1 _34067_inst ( .DIN1(_53051), .DIN2(_34232), .Q(_34225) );
  nor2s1 _34068_inst ( .DIN1(_34233), .DIN2(_34234), .Q(_34232) );
  xor2s1 _34069_inst ( .DIN1(_34235), .DIN2(_34236), .Q(_34234) );
  nor2s1 _34070_inst ( .DIN1(_33578), .DIN2(_34230), .Q(_34236) );
  nor2s1 _34071_inst ( .DIN1(_34231), .DIN2(_33577), .Q(_34233) );
  hi1s1 _34072_inst ( .DIN(_34230), .Q(_34231) );
  nnd2s1 _34073_inst ( .DIN1(_34237), .DIN2(_34238), .Q(_34230) );
  nnd2s1 _34074_inst ( .DIN1(_34239), .DIN2(_26690), .Q(_34238) );
  nnd2s1 _34075_inst ( .DIN1(_53384), .DIN2(_34240), .Q(_34239) );
  or2s1 _34076_inst ( .DIN1(_34240), .DIN2(_26849), .Q(_34237) );
  nnd2s1 _34077_inst ( .DIN1(_34241), .DIN2(_28178), .Q(_34217) );
  xor2s1 _34078_inst ( .DIN1(_53158), .DIN2(_26240), .Q(_34241) );
  nnd2s1 _34079_inst ( .DIN1(_34242), .DIN2(_28569), .Q(
        _____________________________31________) );
  nor2s1 _34080_inst ( .DIN1(_34243), .DIN2(_34244), .Q(_34242) );
  nor2s1 _34081_inst ( .DIN1(_28575), .DIN2(_34245), .Q(_34244) );
  nnd2s1 _34082_inst ( .DIN1(_34246), .DIN2(_34247), .Q(_34245) );
  nnd2s1 _34083_inst ( .DIN1(_34248), .DIN2(_27567), .Q(_34247) );
  xor2s1 _34084_inst ( .DIN1(_34240), .DIN2(_34249), .Q(_34248) );
  xor2s1 _34085_inst ( .DIN1(_53132), .DIN2(_53384), .Q(_34249) );
  nnd2s1 _34086_inst ( .DIN1(_34250), .DIN2(_34251), .Q(_34240) );
  nnd2s1 _34087_inst ( .DIN1(_34252), .DIN2(_26530), .Q(_34251) );
  nnd2s1 _34088_inst ( .DIN1(_26850), .DIN2(_34253), .Q(_34252) );
  or2s1 _34089_inst ( .DIN1(_34253), .DIN2(_26850), .Q(_34250) );
  nnd2s1 _34090_inst ( .DIN1(_34254), .DIN2(______[10]), .Q(_34246) );
  nor2s1 _34091_inst ( .DIN1(_34255), .DIN2(_27596), .Q(_34254) );
  xnr2s1 _34092_inst ( .DIN1(_53319), .DIN2(_53053), .Q(_34255) );
  nor2s1 _34093_inst ( .DIN1(_28572), .DIN2(_34256), .Q(_34243) );
  nor2s1 _34094_inst ( .DIN1(_27365), .DIN2(_26276), .Q(_34256) );
  nnd2s1 _34095_inst ( .DIN1(_34257), .DIN2(_34258), .Q(
        _____________________________30________) );
  nnd2s1 _34096_inst ( .DIN1(_34259), .DIN2(______[24]), .Q(_34258) );
  nor2s1 _34097_inst ( .DIN1(_28182), .DIN2(_34260), .Q(_34259) );
  xor2s1 _34098_inst ( .DIN1(_26477), .DIN2(_53225), .Q(_34260) );
  nnd2s1 _34099_inst ( .DIN1(_28144), .DIN2(_34261), .Q(_34257) );
  nnd2s1 _34100_inst ( .DIN1(_34262), .DIN2(_34263), .Q(_34261) );
  nnd2s1 _34101_inst ( .DIN1(_34264), .DIN2(_34265), .Q(_34263) );
  xor2s1 _34102_inst ( .DIN1(_34253), .DIN2(_34266), .Q(_34264) );
  xor2s1 _34103_inst ( .DIN1(_53052), .DIN2(_53384), .Q(_34266) );
  nnd2s1 _34104_inst ( .DIN1(_34267), .DIN2(_34268), .Q(_34253) );
  nnd2s1 _34105_inst ( .DIN1(_34269), .DIN2(_26636), .Q(_34268) );
  nnd2s1 _34106_inst ( .DIN1(_53384), .DIN2(_34270), .Q(_34269) );
  or2s1 _34107_inst ( .DIN1(_34270), .DIN2(_26849), .Q(_34267) );
  nnd2s1 _34108_inst ( .DIN1(_34271), .DIN2(_34272), .Q(_34262) );
  xor2s1 _34109_inst ( .DIN1(_34273), .DIN2(_34274), .Q(_34271) );
  nnd2s1 _34110_inst ( .DIN1(_53022), .DIN2(_26253), .Q(_34274) );
  nnd2s1 _34111_inst ( .DIN1(_34275), .DIN2(_34276), .Q(_34273) );
  nnd2s1 _34112_inst ( .DIN1(_53066), .DIN2(_53102), .Q(_34276) );
  hi1s1 _34113_inst ( .DIN(_28405), .Q(_28144) );
  nnd2s1 _34114_inst ( .DIN1(_34277), .DIN2(_34278), .Q(
        _____________________________2________) );
  nnd2s1 _34115_inst ( .DIN1(_34279), .DIN2(_53023), .Q(_34278) );
  nor2s1 _34116_inst ( .DIN1(_27551), .DIN2(_27393), .Q(_34279) );
  nnd2s1 _34117_inst ( .DIN1(_27164), .DIN2(_34280), .Q(_34277) );
  nnd2s1 _34118_inst ( .DIN1(_34281), .DIN2(_34282), .Q(_34280) );
  nnd2s1 _34119_inst ( .DIN1(_33871), .DIN2(_34283), .Q(_34282) );
  xor2s1 _34120_inst ( .DIN1(_34284), .DIN2(_34285), .Q(_34283) );
  xnr2s1 _34121_inst ( .DIN1(_34286), .DIN2(_34287), .Q(_34285) );
  nnd2s1 _34122_inst ( .DIN1(_53319), .DIN2(_34288), .Q(_34286) );
  xnr2s1 _34123_inst ( .DIN1(_29492), .DIN2(_53053), .Q(_34284) );
  nor2s1 _34124_inst ( .DIN1(_26241), .DIN2(_34289), .Q(_29492) );
  nnd2s1 _34125_inst ( .DIN1(_34290), .DIN2(_34291), .Q(_34281) );
  nor2s1 _34126_inst ( .DIN1(_34292), .DIN2(_34293), .Q(_34291) );
  nor2s1 _34127_inst ( .DIN1(_26339), .DIN2(_33622), .Q(_34293) );
  nnd2s1 _34128_inst ( .DIN1(_53054), .DIN2(_26719), .Q(_33622) );
  nor2s1 _34129_inst ( .DIN1(_53054), .DIN2(_34294), .Q(_34292) );
  nor2s1 _34130_inst ( .DIN1(_53049), .DIN2(_26339), .Q(_34294) );
  nor2s1 _34131_inst ( .DIN1(_27039), .DIN2(_33464), .Q(_34290) );
  nnd2s1 _34132_inst ( .DIN1(_34295), .DIN2(_34296), .Q(
        _____________________________29________) );
  nnd2s1 _34133_inst ( .DIN1(_34297), .DIN2(_34298), .Q(_34296) );
  nnd2s1 _34134_inst ( .DIN1(_34299), .DIN2(_53318), .Q(_34297) );
  nor2s1 _34135_inst ( .DIN1(_34300), .DIN2(_27066), .Q(_34299) );
  nnd2s1 _34136_inst ( .DIN1(_34301), .DIN2(_34302), .Q(_34295) );
  nnd2s1 _34137_inst ( .DIN1(_34303), .DIN2(_34304), .Q(_34302) );
  nnd2s1 _34138_inst ( .DIN1(_34305), .DIN2(_53139), .Q(_34304) );
  nor2s1 _34139_inst ( .DIN1(_34306), .DIN2(_27651), .Q(_34305) );
  nnd2s1 _34140_inst ( .DIN1(_34307), .DIN2(_34265), .Q(_34303) );
  xor2s1 _34141_inst ( .DIN1(_34270), .DIN2(_34308), .Q(_34307) );
  xor2s1 _34142_inst ( .DIN1(_53141), .DIN2(_53384), .Q(_34308) );
  nnd2s1 _34143_inst ( .DIN1(_34309), .DIN2(_34310), .Q(_34270) );
  nnd2s1 _34144_inst ( .DIN1(_34311), .DIN2(_26484), .Q(_34310) );
  or2s1 _34145_inst ( .DIN1(_34312), .DIN2(_34313), .Q(_34311) );
  nnd2s1 _34146_inst ( .DIN1(_34313), .DIN2(_34312), .Q(_34309) );
  nnd2s1 _34147_inst ( .DIN1(_34314), .DIN2(_34315), .Q(
        _____________________________28________) );
  nnd2s1 _34148_inst ( .DIN1(_27116), .DIN2(_34316), .Q(_34315) );
  nnd2s1 _34149_inst ( .DIN1(_34317), .DIN2(_34318), .Q(_34316) );
  nnd2s1 _34150_inst ( .DIN1(_34319), .DIN2(_34265), .Q(_34318) );
  xor2s1 _34151_inst ( .DIN1(_34313), .DIN2(_34320), .Q(_34319) );
  xor2s1 _34152_inst ( .DIN1(_26484), .DIN2(_34312), .Q(_34320) );
  nnd2s1 _34153_inst ( .DIN1(_34321), .DIN2(_34322), .Q(_34313) );
  nnd2s1 _34154_inst ( .DIN1(_53067), .DIN2(_34323), .Q(_34322) );
  or2s1 _34155_inst ( .DIN1(_34324), .DIN2(_34325), .Q(_34323) );
  nnd2s1 _34156_inst ( .DIN1(_34325), .DIN2(_34324), .Q(_34321) );
  nnd2s1 _34157_inst ( .DIN1(_34272), .DIN2(_26253), .Q(_34317) );
  nnd2s1 _34158_inst ( .DIN1(_34326), .DIN2(_27122), .Q(_34314) );
  nor2s1 _34159_inst ( .DIN1(_27123), .DIN2(_26270), .Q(_34326) );
  nnd2s1 _34160_inst ( .DIN1(_34327), .DIN2(_27256), .Q(
        _____________________________288________) );
  nor2s1 _34161_inst ( .DIN1(_34328), .DIN2(_34329), .Q(_34327) );
  nor2s1 _34162_inst ( .DIN1(_27122), .DIN2(_34330), .Q(_34329) );
  nnd2s1 _34163_inst ( .DIN1(_34331), .DIN2(_34332), .Q(_34330) );
  nnd2s1 _34164_inst ( .DIN1(_34333), .DIN2(_34334), .Q(_34332) );
  xnr2s1 _34165_inst ( .DIN1(_28320), .DIN2(_53378), .Q(_34334) );
  nor2s1 _34166_inst ( .DIN1(_28321), .DIN2(_27066), .Q(_34333) );
  nor2s1 _34167_inst ( .DIN1(_34335), .DIN2(_34336), .Q(_34331) );
  nor2s1 _34168_inst ( .DIN1(_26276), .DIN2(_34337), .Q(_34336) );
  xor2s1 _34169_inst ( .DIN1(_34338), .DIN2(_34339), .Q(_34337) );
  nnd2s1 _34170_inst ( .DIN1(_34340), .DIN2(_34341), .Q(_34339) );
  nnd2s1 _34171_inst ( .DIN1(_34342), .DIN2(_34343), .Q(_34341) );
  nnd2s1 _34172_inst ( .DIN1(_34344), .DIN2(_34345), .Q(_34340) );
  nor2s1 _34173_inst ( .DIN1(_53138), .DIN2(_34346), .Q(_34335) );
  nor2s1 _34174_inst ( .DIN1(_34347), .DIN2(_34348), .Q(_34346) );
  nor2s1 _34175_inst ( .DIN1(_34345), .DIN2(_34344), .Q(_34348) );
  nor2s1 _34176_inst ( .DIN1(_34342), .DIN2(_34343), .Q(_34347) );
  hi1s1 _34177_inst ( .DIN(_34344), .Q(_34342) );
  nnd2s1 _34178_inst ( .DIN1(_34349), .DIN2(_34350), .Q(_34344) );
  nnd2s1 _34179_inst ( .DIN1(_34351), .DIN2(_26514), .Q(_34350) );
  nnd2s1 _34180_inst ( .DIN1(_53384), .DIN2(_34352), .Q(_34351) );
  or2s1 _34181_inst ( .DIN1(_34352), .DIN2(_26849), .Q(_34349) );
  nor2s1 _34182_inst ( .DIN1(_27116), .DIN2(_34353), .Q(_34328) );
  nor2s1 _34183_inst ( .DIN1(_27039), .DIN2(_34354), .Q(_34353) );
  xor2s1 _34184_inst ( .DIN1(_53057), .DIN2(_53210), .Q(_34354) );
  nnd2s1 _34185_inst ( .DIN1(_34355), .DIN2(_34356), .Q(
        _____________________________287________) );
  nnd2s1 _34186_inst ( .DIN1(_29139), .DIN2(_34357), .Q(_34356) );
  nnd2s1 _34187_inst ( .DIN1(_34358), .DIN2(_34359), .Q(_34357) );
  xnr2s1 _34188_inst ( .DIN1(_34360), .DIN2(_34352), .Q(_34358) );
  nnd2s1 _34189_inst ( .DIN1(_34361), .DIN2(_34362), .Q(_34352) );
  nnd2s1 _34190_inst ( .DIN1(_34363), .DIN2(_26746), .Q(_34362) );
  or2s1 _34191_inst ( .DIN1(_34364), .DIN2(_26849), .Q(_34363) );
  nnd2s1 _34192_inst ( .DIN1(_53384), .DIN2(_34364), .Q(_34361) );
  xor2s1 _34193_inst ( .DIN1(_26514), .DIN2(_53384), .Q(_34360) );
  nnd2s1 _34194_inst ( .DIN1(_29137), .DIN2(_53061), .Q(_34355) );
  hi1s1 _34195_inst ( .DIN(_34365), .Q(_29137) );
  nnd2s1 _34196_inst ( .DIN1(_34366), .DIN2(_28148), .Q(
        _____________________________286________) );
  nor2s1 _34197_inst ( .DIN1(_34367), .DIN2(_34368), .Q(_34366) );
  nor2s1 _34198_inst ( .DIN1(_34369), .DIN2(_28151), .Q(_34368) );
  nor2s1 _34199_inst ( .DIN1(_34370), .DIN2(_34371), .Q(_34369) );
  xor2s1 _34200_inst ( .DIN1(_34364), .DIN2(_34372), .Q(_34371) );
  xor2s1 _34201_inst ( .DIN1(_53171), .DIN2(_53384), .Q(_34372) );
  nnd2s1 _34202_inst ( .DIN1(_34373), .DIN2(_34374), .Q(_34364) );
  nnd2s1 _34203_inst ( .DIN1(_34375), .DIN2(_26552), .Q(_34374) );
  or2s1 _34204_inst ( .DIN1(_34376), .DIN2(_26849), .Q(_34375) );
  nnd2s1 _34205_inst ( .DIN1(_53384), .DIN2(_34376), .Q(_34373) );
  nor2s1 _34206_inst ( .DIN1(_53059), .DIN2(_28153), .Q(_34367) );
  nnd2s1 _34207_inst ( .DIN1(_34377), .DIN2(_34378), .Q(
        _____________________________285________) );
  nor2s1 _34208_inst ( .DIN1(_34379), .DIN2(_34380), .Q(_34378) );
  nor2s1 _34209_inst ( .DIN1(_28151), .DIN2(_34381), .Q(_34380) );
  xor2s1 _34210_inst ( .DIN1(_34382), .DIN2(_30912), .Q(_34381) );
  nnd2s1 _34211_inst ( .DIN1(_34383), .DIN2(_34359), .Q(_34382) );
  xnr2s1 _34212_inst ( .DIN1(_34376), .DIN2(_34384), .Q(_34383) );
  xor2s1 _34213_inst ( .DIN1(_53100), .DIN2(_53384), .Q(_34384) );
  nnd2s1 _34214_inst ( .DIN1(_34385), .DIN2(_34386), .Q(_34376) );
  nnd2s1 _34215_inst ( .DIN1(_34387), .DIN2(_26683), .Q(_34386) );
  or2s1 _34216_inst ( .DIN1(_34388), .DIN2(_26849), .Q(_34387) );
  nnd2s1 _34217_inst ( .DIN1(_26849), .DIN2(_34388), .Q(_34385) );
  nor2s1 _34218_inst ( .DIN1(_28153), .DIN2(_34389), .Q(_34379) );
  nor2s1 _34219_inst ( .DIN1(_34390), .DIN2(_27241), .Q(_34389) );
  nor2s1 _34220_inst ( .DIN1(_29131), .DIN2(_26630), .Q(_34390) );
  hi1s1 _34221_inst ( .DIN(_28151), .Q(_28153) );
  nor2s1 _34222_inst ( .DIN1(_29132), .DIN2(_34391), .Q(_34377) );
  nor2s1 _34223_inst ( .DIN1(_53058), .DIN2(_29134), .Q(_34391) );
  nnd2s1 _34224_inst ( .DIN1(_29131), .DIN2(_28151), .Q(_29134) );
  and2s1 _34225_inst ( .DIN1(_53059), .DIN2(_53060), .Q(_29131) );
  hi1s1 _34226_inst ( .DIN(_28148), .Q(_29132) );
  nnd2s1 _34227_inst ( .DIN1(_28159), .DIN2(_28151), .Q(_28148) );
  nnd2s1 _34228_inst ( .DIN1(_34392), .DIN2(_34393), .Q(_28151) );
  nor2s1 _34229_inst ( .DIN1(_34394), .DIN2(_34395), .Q(_34393) );
  nnd2s1 _34230_inst ( .DIN1(_34396), .DIN2(_33613), .Q(_34395) );
  nor2s1 _34231_inst ( .DIN1(_34397), .DIN2(_34398), .Q(_34392) );
  nor2s1 _34232_inst ( .DIN1(_27936), .DIN2(_34399), .Q(_28159) );
  nnd2s1 _34233_inst ( .DIN1(_34400), .DIN2(_34401), .Q(
        _____________________________284________) );
  nnd2s1 _34234_inst ( .DIN1(_34402), .DIN2(_34403), .Q(_34401) );
  xor2s1 _34235_inst ( .DIN1(_53062), .DIN2(_26612), .Q(_34403) );
  nor2s1 _34236_inst ( .DIN1(_27082), .DIN2(_34365), .Q(_34402) );
  nnd2s1 _34237_inst ( .DIN1(_28672), .DIN2(_28670), .Q(_34365) );
  nnd2s1 _34238_inst ( .DIN1(_29139), .DIN2(_34404), .Q(_34400) );
  nnd2s1 _34239_inst ( .DIN1(_34405), .DIN2(_34359), .Q(_34404) );
  xnr2s1 _34240_inst ( .DIN1(_34388), .DIN2(_34406), .Q(_34405) );
  xor2s1 _34241_inst ( .DIN1(_53230), .DIN2(_53384), .Q(_34406) );
  nnd2s1 _34242_inst ( .DIN1(_34407), .DIN2(_34408), .Q(_34388) );
  nnd2s1 _34243_inst ( .DIN1(_34409), .DIN2(_26482), .Q(_34408) );
  or2s1 _34244_inst ( .DIN1(_34410), .DIN2(_26849), .Q(_34409) );
  nnd2s1 _34245_inst ( .DIN1(_26849), .DIN2(_34410), .Q(_34407) );
  hi1s1 _34246_inst ( .DIN(_28670), .Q(_29139) );
  nnd2s1 _34247_inst ( .DIN1(_34411), .DIN2(_28887), .Q(_28670) );
  and2s1 _34248_inst ( .DIN1(_34412), .DIN2(_34413), .Q(_28887) );
  nor2s1 _34249_inst ( .DIN1(_34414), .DIN2(_34415), .Q(_34412) );
  nor2s1 _34250_inst ( .DIN1(_30026), .DIN2(_31084), .Q(_34411) );
  nnd2s1 _34251_inst ( .DIN1(_34416), .DIN2(_34417), .Q(_31084) );
  nor2s1 _34252_inst ( .DIN1(_29940), .DIN2(_30027), .Q(_34417) );
  nor2s1 _34253_inst ( .DIN1(_30772), .DIN2(_31077), .Q(_34416) );
  hi1s1 _34254_inst ( .DIN(_30434), .Q(_31077) );
  nnd2s1 _34255_inst ( .DIN1(_34418), .DIN2(_34419), .Q(
        _____________________________283________) );
  nnd2s1 _34256_inst ( .DIN1(_34420), .DIN2(_34421), .Q(_34419) );
  nnd2s1 _34257_inst ( .DIN1(_34422), .DIN2(_34423), .Q(_34421) );
  xor2s1 _34258_inst ( .DIN1(_34424), .DIN2(_53065), .Q(_34422) );
  hi1s1 _34259_inst ( .DIN(_34425), .Q(_34420) );
  nor2s1 _34260_inst ( .DIN1(_34426), .DIN2(_34427), .Q(_34418) );
  nor2s1 _34261_inst ( .DIN1(_34428), .DIN2(_34429), .Q(_34427) );
  xnr2s1 _34262_inst ( .DIN1(_34410), .DIN2(_34430), .Q(_34429) );
  xor2s1 _34263_inst ( .DIN1(_53172), .DIN2(_53384), .Q(_34430) );
  nnd2s1 _34264_inst ( .DIN1(_34431), .DIN2(_34432), .Q(_34410) );
  nnd2s1 _34265_inst ( .DIN1(_53101), .DIN2(_34433), .Q(_34432) );
  or2s1 _34266_inst ( .DIN1(_34434), .DIN2(_26849), .Q(_34433) );
  nnd2s1 _34267_inst ( .DIN1(_26849), .DIN2(_34434), .Q(_34431) );
  nor2s1 _34268_inst ( .DIN1(_27774), .DIN2(_34435), .Q(_34426) );
  nnd2s1 _34269_inst ( .DIN1(_53064), .DIN2(_27498), .Q(_34435) );
  nor2s1 _34270_inst ( .DIN1(_34436), .DIN2(_28998), .Q(
        _____________________________282________) );
  nor2s1 _34271_inst ( .DIN1(_34437), .DIN2(_34438), .Q(_34436) );
  nor2s1 _34272_inst ( .DIN1(_27082), .DIN2(_34439), .Q(_34438) );
  nnd2s1 _34273_inst ( .DIN1(_34440), .DIN2(_34441), .Q(_34439) );
  nnd2s1 _34274_inst ( .DIN1(_34442), .DIN2(_26540), .Q(_34441) );
  nnd2s1 _34275_inst ( .DIN1(_53515), .DIN2(_34443), .Q(_34440) );
  or2s1 _34276_inst ( .DIN1(_34424), .DIN2(_34444), .Q(_34443) );
  nor2s1 _34277_inst ( .DIN1(_34445), .DIN2(_34446), .Q(_34437) );
  xor2s1 _34278_inst ( .DIN1(_34434), .DIN2(_34447), .Q(_34446) );
  xor2s1 _34279_inst ( .DIN1(_53101), .DIN2(_26850), .Q(_34447) );
  nnd2s1 _34280_inst ( .DIN1(_34448), .DIN2(_34449), .Q(_34434) );
  nnd2s1 _34281_inst ( .DIN1(_53363), .DIN2(_34450), .Q(_34449) );
  or2s1 _34282_inst ( .DIN1(_26410), .DIN2(_34451), .Q(_34450) );
  nnd2s1 _34283_inst ( .DIN1(_34451), .DIN2(_26410), .Q(_34448) );
  nnd2s1 _34284_inst ( .DIN1(_34452), .DIN2(_34453), .Q(
        _____________________________281________) );
  nor2s1 _34285_inst ( .DIN1(_34454), .DIN2(_34455), .Q(_34452) );
  nor2s1 _34286_inst ( .DIN1(_34456), .DIN2(_34457), .Q(_34455) );
  nor2s1 _34287_inst ( .DIN1(_34458), .DIN2(_34459), .Q(_34457) );
  nor2s1 _34288_inst ( .DIN1(_34445), .DIN2(_34460), .Q(_34459) );
  xnr2s1 _34289_inst ( .DIN1(_34461), .DIN2(_34451), .Q(_34460) );
  nnd2s1 _34290_inst ( .DIN1(_34462), .DIN2(_34463), .Q(_34451) );
  nnd2s1 _34291_inst ( .DIN1(_34464), .DIN2(_26738), .Q(_34463) );
  or2s1 _34292_inst ( .DIN1(_34465), .DIN2(_53364), .Q(_34464) );
  nnd2s1 _34293_inst ( .DIN1(_53364), .DIN2(_34465), .Q(_34462) );
  xor2s1 _34294_inst ( .DIN1(_26410), .DIN2(_53363), .Q(_34461) );
  nor2s1 _34295_inst ( .DIN1(_34466), .DIN2(_34467), .Q(_34458) );
  nnd2s1 _34296_inst ( .DIN1(_53063), .DIN2(_34423), .Q(_34467) );
  nor2s1 _34297_inst ( .DIN1(_30949), .DIN2(_34468), .Q(_34454) );
  xor2s1 _34298_inst ( .DIN1(_34469), .DIN2(_53081), .Q(_34468) );
  nnd2s1 _34299_inst ( .DIN1(_34470), .DIN2(_34471), .Q(
        _____________________________280________) );
  nnd2s1 _34300_inst ( .DIN1(_34472), .DIN2(_34473), .Q(_34471) );
  hi1s1 _34301_inst ( .DIN(_34428), .Q(_34473) );
  nnd2s1 _34302_inst ( .DIN1(_34466), .DIN2(_27421), .Q(_34428) );
  xor2s1 _34303_inst ( .DIN1(_34465), .DIN2(_34474), .Q(_34472) );
  xor2s1 _34304_inst ( .DIN1(_53109), .DIN2(_53364), .Q(_34474) );
  nnd2s1 _34305_inst ( .DIN1(_34475), .DIN2(_34476), .Q(_34465) );
  nnd2s1 _34306_inst ( .DIN1(_53104), .DIN2(_34477), .Q(_34476) );
  nnd2s1 _34307_inst ( .DIN1(_53362), .DIN2(_34478), .Q(_34477) );
  or2s1 _34308_inst ( .DIN1(_34478), .DIN2(_53362), .Q(_34475) );
  nor2s1 _34309_inst ( .DIN1(_34479), .DIN2(_34480), .Q(_34470) );
  nor2s1 _34310_inst ( .DIN1(_34481), .DIN2(_34482), .Q(_34480) );
  xor2s1 _34311_inst ( .DIN1(_34483), .DIN2(_53515), .Q(_34482) );
  nnd2s1 _34312_inst ( .DIN1(_53065), .DIN2(_53064), .Q(_34483) );
  hi1s1 _34313_inst ( .DIN(_27498), .Q(_34481) );
  nnd2s1 _34314_inst ( .DIN1(_34484), .DIN2(_34485), .Q(_27498) );
  nor2s1 _34315_inst ( .DIN1(_34486), .DIN2(_34425), .Q(_34479) );
  nnd2s1 _34316_inst ( .DIN1(_27421), .DIN2(_34445), .Q(_34425) );
  hi1s1 _34317_inst ( .DIN(_34466), .Q(_34445) );
  hi1s1 _34318_inst ( .DIN(_27408), .Q(_27421) );
  nnd2s1 _34319_inst ( .DIN1(_34487), .DIN2(_34488), .Q(_27408) );
  nor2s1 _34320_inst ( .DIN1(_34489), .DIN2(_34490), .Q(_34487) );
  nor2s1 _34321_inst ( .DIN1(_34491), .DIN2(_34442), .Q(_34486) );
  nnd2s1 _34322_inst ( .DIN1(_34423), .DIN2(_34424), .Q(_34442) );
  nnd2s1 _34323_inst ( .DIN1(_53063), .DIN2(_53068), .Q(_34424) );
  nor2s1 _34324_inst ( .DIN1(_53063), .DIN2(_53068), .Q(_34491) );
  nnd2s1 _34325_inst ( .DIN1(_28769), .DIN2(_34492), .Q(
        _____________________________27________) );
  nnd2s1 _34326_inst ( .DIN1(_34493), .DIN2(_34494), .Q(_34492) );
  nnd2s1 _34327_inst ( .DIN1(_34265), .DIN2(_34495), .Q(_34494) );
  xnr2s1 _34328_inst ( .DIN1(_34325), .DIN2(_34496), .Q(_34495) );
  xor2s1 _34329_inst ( .DIN1(_26593), .DIN2(_34324), .Q(_34496) );
  nnd2s1 _34330_inst ( .DIN1(_34497), .DIN2(_34498), .Q(_34324) );
  nnd2s1 _34331_inst ( .DIN1(_34499), .DIN2(_26451), .Q(_34498) );
  or2s1 _34332_inst ( .DIN1(_34500), .DIN2(_34501), .Q(_34499) );
  xor2s1 _34333_inst ( .DIN1(_31282), .DIN2(_34502), .Q(_34497) );
  nnd2s1 _34334_inst ( .DIN1(_34501), .DIN2(_34500), .Q(_34502) );
  nnd2s1 _34335_inst ( .DIN1(_34503), .DIN2(_34272), .Q(_34493) );
  xnr2s1 _34336_inst ( .DIN1(_53022), .DIN2(_34275), .Q(_34503) );
  nnd2s1 _34337_inst ( .DIN1(_26563), .DIN2(_26253), .Q(_34275) );
  hi1s1 _34338_inst ( .DIN(_28998), .Q(_28769) );
  nnd2s1 _34339_inst ( .DIN1(_34504), .DIN2(_30774), .Q(
        _____________________________279________) );
  nor2s1 _34340_inst ( .DIN1(_34505), .DIN2(_34506), .Q(_34504) );
  nor2s1 _34341_inst ( .DIN1(_30777), .DIN2(_34507), .Q(_34506) );
  nnd2s1 _34342_inst ( .DIN1(_34508), .DIN2(_34509), .Q(_34507) );
  nnd2s1 _34343_inst ( .DIN1(_34510), .DIN2(_34466), .Q(_34509) );
  xnr2s1 _34344_inst ( .DIN1(_34511), .DIN2(_34478), .Q(_34510) );
  nnd2s1 _34345_inst ( .DIN1(_34512), .DIN2(_34513), .Q(_34478) );
  nnd2s1 _34346_inst ( .DIN1(_53105), .DIN2(_34514), .Q(_34513) );
  nnd2s1 _34347_inst ( .DIN1(_34515), .DIN2(_34516), .Q(_34514) );
  nnd2s1 _34348_inst ( .DIN1(_34517), .DIN2(_53361), .Q(_34512) );
  xor2s1 _34349_inst ( .DIN1(_26547), .DIN2(_53362), .Q(_34511) );
  nnd2s1 _34350_inst ( .DIN1(_34518), .DIN2(_34423), .Q(_34508) );
  xnr2s1 _34351_inst ( .DIN1(_34519), .DIN2(_34520), .Q(_34518) );
  nnd2s1 _34352_inst ( .DIN1(_34521), .DIN2(_34522), .Q(_34519) );
  nnd2s1 _34353_inst ( .DIN1(_53179), .DIN2(_26432), .Q(_34522) );
  nor2s1 _34354_inst ( .DIN1(_53079), .DIN2(_27227), .Q(_34505) );
  nnd2s1 _34355_inst ( .DIN1(_34523), .DIN2(_31861), .Q(
        _____________________________278________) );
  nor2s1 _34356_inst ( .DIN1(_34524), .DIN2(_34525), .Q(_34523) );
  nor2s1 _34357_inst ( .DIN1(_31864), .DIN2(_34526), .Q(_34525) );
  nnd2s1 _34358_inst ( .DIN1(_34527), .DIN2(_34528), .Q(_34526) );
  nnd2s1 _34359_inst ( .DIN1(_53083), .DIN2(_34423), .Q(_34528) );
  nnd2s1 _34360_inst ( .DIN1(_34529), .DIN2(_34466), .Q(_34527) );
  nor2s1 _34361_inst ( .DIN1(_34530), .DIN2(_34531), .Q(_34466) );
  nor2s1 _34362_inst ( .DIN1(_34532), .DIN2(_34533), .Q(_34529) );
  nor2s1 _34363_inst ( .DIN1(_26735), .DIN2(_34534), .Q(_34533) );
  xor2s1 _34364_inst ( .DIN1(_34515), .DIN2(_34516), .Q(_34534) );
  nor2s1 _34365_inst ( .DIN1(_53105), .DIN2(_26762), .Q(_34532) );
  hi1s1 _34366_inst ( .DIN(_34516), .Q(_34517) );
  nnd2s1 _34367_inst ( .DIN1(_34535), .DIN2(_34536), .Q(_34516) );
  nnd2s1 _34368_inst ( .DIN1(_34537), .DIN2(_26748), .Q(_34536) );
  or2s1 _34369_inst ( .DIN1(_34538), .DIN2(_53365), .Q(_34537) );
  nnd2s1 _34370_inst ( .DIN1(_53365), .DIN2(_34538), .Q(_34535) );
  nor2s1 _34371_inst ( .DIN1(_31907), .DIN2(_34539), .Q(_34524) );
  xor2s1 _34372_inst ( .DIN1(_53342), .DIN2(_26344), .Q(_34539) );
  nnd2s1 _34373_inst ( .DIN1(_34540), .DIN2(_34541), .Q(
        _____________________________277________) );
  nnd2s1 _34374_inst ( .DIN1(_34542), .DIN2(_34456), .Q(_34541) );
  nor2s1 _34375_inst ( .DIN1(_27365), .DIN2(_34543), .Q(_34542) );
  nnd2s1 _34376_inst ( .DIN1(_34544), .DIN2(_31083), .Q(_34543) );
  xor2s1 _34377_inst ( .DIN1(_34469), .DIN2(_53068), .Q(_34544) );
  nnd2s1 _34378_inst ( .DIN1(_53077), .DIN2(_53078), .Q(_34469) );
  nnd2s1 _34379_inst ( .DIN1(_34545), .DIN2(_30949), .Q(_34540) );
  nnd2s1 _34380_inst ( .DIN1(_34546), .DIN2(_34547), .Q(_34545) );
  nnd2s1 _34381_inst ( .DIN1(_34548), .DIN2(_34549), .Q(_34547) );
  nnd2s1 _34382_inst ( .DIN1(_34550), .DIN2(______[28]), .Q(_34548) );
  nor2s1 _34383_inst ( .DIN1(_53179), .DIN2(_34551), .Q(_34550) );
  nnd2s1 _34384_inst ( .DIN1(_34552), .DIN2(_34553), .Q(_34546) );
  xor2s1 _34385_inst ( .DIN1(_34538), .DIN2(_34554), .Q(_34553) );
  xor2s1 _34386_inst ( .DIN1(_53108), .DIN2(_53365), .Q(_34554) );
  nnd2s1 _34387_inst ( .DIN1(_34555), .DIN2(_34556), .Q(_34538) );
  nnd2s1 _34388_inst ( .DIN1(_53071), .DIN2(_34557), .Q(_34556) );
  or2s1 _34389_inst ( .DIN1(_34558), .DIN2(_26781), .Q(_34557) );
  nnd2s1 _34390_inst ( .DIN1(_26781), .DIN2(_34558), .Q(_34555) );
  nnd2s1 _34391_inst ( .DIN1(_34559), .DIN2(_34560), .Q(
        _____________________________276________) );
  nnd2s1 _34392_inst ( .DIN1(_34561), .DIN2(_34562), .Q(_34560) );
  xor2s1 _34393_inst ( .DIN1(_26339), .DIN2(_53430), .Q(_34562) );
  nor2s1 _34394_inst ( .DIN1(_33589), .DIN2(_28100), .Q(_34561) );
  nnd2s1 _34395_inst ( .DIN1(_34563), .DIN2(_27895), .Q(_34559) );
  nor2s1 _34396_inst ( .DIN1(_34564), .DIN2(_34565), .Q(_34563) );
  nor2s1 _34397_inst ( .DIN1(_34549), .DIN2(_34566), .Q(_34565) );
  xor2s1 _34398_inst ( .DIN1(_34558), .DIN2(_34567), .Q(_34566) );
  xor2s1 _34399_inst ( .DIN1(_53071), .DIN2(_53368), .Q(_34567) );
  nnd2s1 _34400_inst ( .DIN1(_34568), .DIN2(_34569), .Q(_34558) );
  nnd2s1 _34401_inst ( .DIN1(_34570), .DIN2(_26713), .Q(_34569) );
  or2s1 _34402_inst ( .DIN1(_34571), .DIN2(_53367), .Q(_34570) );
  nnd2s1 _34403_inst ( .DIN1(_53367), .DIN2(_34571), .Q(_34568) );
  nor2s1 _34404_inst ( .DIN1(_34552), .DIN2(_34572), .Q(_34564) );
  nor2s1 _34405_inst ( .DIN1(_34573), .DIN2(_34574), .Q(_34572) );
  nnd2s1 _34406_inst ( .DIN1(______[28]), .DIN2(_34575), .Q(_34574) );
  nnd2s1 _34407_inst ( .DIN1(_53077), .DIN2(_34521), .Q(_34575) );
  or2s1 _34408_inst ( .DIN1(_26432), .DIN2(_53179), .Q(_34521) );
  nnd2s1 _34409_inst ( .DIN1(_34576), .DIN2(_34577), .Q(_34573) );
  nnd2s1 _34410_inst ( .DIN1(_34520), .DIN2(_53070), .Q(_34576) );
  nor2s1 _34411_inst ( .DIN1(_53077), .DIN2(_53179), .Q(_34520) );
  nnd2s1 _34412_inst ( .DIN1(_34578), .DIN2(_28941), .Q(
        _____________________________275________) );
  or2s1 _34413_inst ( .DIN1(_31001), .DIN2(_28944), .Q(_28941) );
  nnd2s1 _34414_inst ( .DIN1(_34579), .DIN2(_34580), .Q(_31001) );
  nor2s1 _34415_inst ( .DIN1(_33617), .DIN2(_34394), .Q(_34579) );
  nor2s1 _34416_inst ( .DIN1(_34581), .DIN2(_34582), .Q(_34578) );
  nor2s1 _34417_inst ( .DIN1(_28949), .DIN2(_34583), .Q(_34582) );
  nor2s1 _34418_inst ( .DIN1(_34584), .DIN2(_34585), .Q(_34583) );
  nor2s1 _34419_inst ( .DIN1(_34586), .DIN2(_34549), .Q(_34585) );
  xnr2s1 _34420_inst ( .DIN1(_34571), .DIN2(_34587), .Q(_34586) );
  xor2s1 _34421_inst ( .DIN1(_53110), .DIN2(_53367), .Q(_34587) );
  nnd2s1 _34422_inst ( .DIN1(_34588), .DIN2(_34589), .Q(_34571) );
  nnd2s1 _34423_inst ( .DIN1(_53309), .DIN2(_34590), .Q(_34589) );
  or2s1 _34424_inst ( .DIN1(_34591), .DIN2(_53355), .Q(_34590) );
  nnd2s1 _34425_inst ( .DIN1(_53355), .DIN2(_34591), .Q(_34588) );
  nor2s1 _34426_inst ( .DIN1(_34552), .DIN2(_34592), .Q(_34584) );
  nor2s1 _34427_inst ( .DIN1(_34593), .DIN2(_34594), .Q(_34592) );
  nnd2s1 _34428_inst ( .DIN1(_34595), .DIN2(_34577), .Q(_34594) );
  nnd2s1 _34429_inst ( .DIN1(_53078), .DIN2(_26556), .Q(_34595) );
  nnd2s1 _34430_inst ( .DIN1(_34596), .DIN2(_34597), .Q(_34593) );
  nnd2s1 _34431_inst ( .DIN1(_34598), .DIN2(_53073), .Q(_34597) );
  nnd2s1 _34432_inst ( .DIN1(_53078), .DIN2(_26708), .Q(_34596) );
  nor2s1 _34433_inst ( .DIN1(_28944), .DIN2(_34599), .Q(_34581) );
  nor2s1 _34434_inst ( .DIN1(_27393), .DIN2(_26586), .Q(_34599) );
  hi1s1 _34435_inst ( .DIN(_28949), .Q(_28944) );
  nnd2s1 _34436_inst ( .DIN1(_34600), .DIN2(_34601), .Q(_28949) );
  nor2s1 _34437_inst ( .DIN1(_34602), .DIN2(_34397), .Q(_34600) );
  nnd2s1 _34438_inst ( .DIN1(_34603), .DIN2(_34604), .Q(
        _____________________________274________) );
  nnd2s1 _34439_inst ( .DIN1(_31809), .DIN2(_34605), .Q(_34604) );
  xor2s1 _34440_inst ( .DIN1(_53072), .DIN2(_53328), .Q(_34605) );
  nnd2s1 _34441_inst ( .DIN1(_34606), .DIN2(_30175), .Q(_34603) );
  nor2s1 _34442_inst ( .DIN1(_34607), .DIN2(_34608), .Q(_34606) );
  nor2s1 _34443_inst ( .DIN1(_34552), .DIN2(_34609), .Q(_34608) );
  nnd2s1 _34444_inst ( .DIN1(_53082), .DIN2(_34577), .Q(_34609) );
  nor2s1 _34445_inst ( .DIN1(_34610), .DIN2(_34549), .Q(_34607) );
  xor2s1 _34446_inst ( .DIN1(_34591), .DIN2(_34611), .Q(_34610) );
  xor2s1 _34447_inst ( .DIN1(_26449), .DIN2(_53309), .Q(_34611) );
  nnd2s1 _34448_inst ( .DIN1(_34612), .DIN2(_34613), .Q(_34591) );
  nnd2s1 _34449_inst ( .DIN1(_53131), .DIN2(_34614), .Q(_34613) );
  or2s1 _34450_inst ( .DIN1(_34615), .DIN2(_53314), .Q(_34614) );
  nnd2s1 _34451_inst ( .DIN1(_53314), .DIN2(_34615), .Q(_34612) );
  nor2s1 _34452_inst ( .DIN1(_28084), .DIN2(_34616), .Q(
        _____________________________273________) );
  nnd2s1 _34453_inst ( .DIN1(_34617), .DIN2(_34618), .Q(_34616) );
  nnd2s1 _34454_inst ( .DIN1(_34619), .DIN2(_34549), .Q(_34618) );
  nnd2s1 _34455_inst ( .DIN1(_34620), .DIN2(_52901), .Q(_34619) );
  nor2s1 _34456_inst ( .DIN1(_34551), .DIN2(_28100), .Q(_34620) );
  nnd2s1 _34457_inst ( .DIN1(_34621), .DIN2(_34552), .Q(_34617) );
  xnr2s1 _34458_inst ( .DIN1(_34615), .DIN2(_34622), .Q(_34621) );
  xor2s1 _34459_inst ( .DIN1(_53131), .DIN2(_53314), .Q(_34622) );
  nnd2s1 _34460_inst ( .DIN1(_34623), .DIN2(_34624), .Q(_34615) );
  nnd2s1 _34461_inst ( .DIN1(_53371), .DIN2(_34625), .Q(_34624) );
  or2s1 _34462_inst ( .DIN1(_34626), .DIN2(_53523), .Q(_34625) );
  nnd2s1 _34463_inst ( .DIN1(_53523), .DIN2(_34626), .Q(_34623) );
  nnd2s1 _34464_inst ( .DIN1(_34627), .DIN2(_34453), .Q(
        _____________________________272________) );
  hi1s1 _34465_inst ( .DIN(_34628), .Q(_34453) );
  nor2s1 _34466_inst ( .DIN1(_34629), .DIN2(_34630), .Q(_34627) );
  nor2s1 _34467_inst ( .DIN1(_34456), .DIN2(_34631), .Q(_34630) );
  nor2s1 _34468_inst ( .DIN1(_34632), .DIN2(_34633), .Q(_34631) );
  nor2s1 _34469_inst ( .DIN1(_34552), .DIN2(_34634), .Q(_34633) );
  nnd2s1 _34470_inst ( .DIN1(_34635), .DIN2(______[30]), .Q(_34634) );
  nor2s1 _34471_inst ( .DIN1(_34551), .DIN2(_34636), .Q(_34635) );
  xor2s1 _34472_inst ( .DIN1(_53073), .DIN2(_34598), .Q(_34636) );
  nor2s1 _34473_inst ( .DIN1(_26556), .DIN2(_53078), .Q(_34598) );
  hi1s1 _34474_inst ( .DIN(_34577), .Q(_34551) );
  nnd2s1 _34475_inst ( .DIN1(_34637), .DIN2(_34638), .Q(_34577) );
  hi1s1 _34476_inst ( .DIN(_34549), .Q(_34552) );
  nor2s1 _34477_inst ( .DIN1(_34639), .DIN2(_34549), .Q(_34632) );
  nnd2s1 _34478_inst ( .DIN1(_34640), .DIN2(_34641), .Q(_34549) );
  nor2s1 _34479_inst ( .DIN1(_34642), .DIN2(_34530), .Q(_34640) );
  xor2s1 _34480_inst ( .DIN1(_34626), .DIN2(_34643), .Q(_34639) );
  xor2s1 _34481_inst ( .DIN1(_26258), .DIN2(_53371), .Q(_34643) );
  nnd2s1 _34482_inst ( .DIN1(_34644), .DIN2(_34645), .Q(_34626) );
  nnd2s1 _34483_inst ( .DIN1(_34646), .DIN2(_26694), .Q(_34645) );
  or2s1 _34484_inst ( .DIN1(_34647), .DIN2(_53370), .Q(_34646) );
  nnd2s1 _34485_inst ( .DIN1(_53370), .DIN2(_34647), .Q(_34644) );
  nor2s1 _34486_inst ( .DIN1(_53077), .DIN2(_30949), .Q(_34629) );
  nnd2s1 _34487_inst ( .DIN1(_34648), .DIN2(_34649), .Q(
        _____________________________271________) );
  nnd2s1 _34488_inst ( .DIN1(_34650), .DIN2(_26863), .Q(_34649) );
  nor2s1 _34489_inst ( .DIN1(_53054), .DIN2(_32239), .Q(_34650) );
  hi1s1 _34490_inst ( .DIN(_34651), .Q(_32239) );
  nnd2s1 _34491_inst ( .DIN1(_27064), .DIN2(_34652), .Q(_34648) );
  nnd2s1 _34492_inst ( .DIN1(_34653), .DIN2(_34654), .Q(_34652) );
  nnd2s1 _34493_inst ( .DIN1(_34655), .DIN2(_34656), .Q(_34654) );
  xnr2s1 _34494_inst ( .DIN1(_34647), .DIN2(_34657), .Q(_34655) );
  xor2s1 _34495_inst ( .DIN1(_53117), .DIN2(_53370), .Q(_34657) );
  nnd2s1 _34496_inst ( .DIN1(_34658), .DIN2(_34659), .Q(_34647) );
  nnd2s1 _34497_inst ( .DIN1(_53118), .DIN2(_34660), .Q(_34659) );
  or2s1 _34498_inst ( .DIN1(_34661), .DIN2(_53517), .Q(_34660) );
  nnd2s1 _34499_inst ( .DIN1(_53517), .DIN2(_34661), .Q(_34658) );
  nnd2s1 _34500_inst ( .DIN1(_34662), .DIN2(_34663), .Q(_34653) );
  xor2s1 _34501_inst ( .DIN1(_34664), .DIN2(_34665), .Q(_34663) );
  nor2s1 _34502_inst ( .DIN1(_53074), .DIN2(_26516), .Q(_34665) );
  xor2s1 _34503_inst ( .DIN1(_26631), .DIN2(_53075), .Q(_34664) );
  nor2s1 _34504_inst ( .DIN1(_27039), .DIN2(_34666), .Q(_34662) );
  hi1s1 _34505_inst ( .DIN(_27053), .Q(_27064) );
  nnd2s1 _34506_inst ( .DIN1(_34667), .DIN2(_34668), .Q(_27053) );
  nor2s1 _34507_inst ( .DIN1(_34669), .DIN2(_34670), .Q(_34668) );
  nnd2s1 _34508_inst ( .DIN1(_34671), .DIN2(_34672), .Q(_34670) );
  nor2s1 _34509_inst ( .DIN1(_34673), .DIN2(_34651), .Q(_34667) );
  nnd2s1 _34510_inst ( .DIN1(_34674), .DIN2(_34675), .Q(_34651) );
  nor2s1 _34511_inst ( .DIN1(_34676), .DIN2(_34677), .Q(_34675) );
  nor2s1 _34512_inst ( .DIN1(_34678), .DIN2(_34394), .Q(_34674) );
  nor2s1 _34513_inst ( .DIN1(_34679), .DIN2(_27235), .Q(
        _____________________________270________) );
  nor2s1 _34514_inst ( .DIN1(_34680), .DIN2(_34681), .Q(_34679) );
  nor2s1 _34515_inst ( .DIN1(_34682), .DIN2(_34683), .Q(_34681) );
  xor2s1 _34516_inst ( .DIN1(_34661), .DIN2(_34684), .Q(_34683) );
  xor2s1 _34517_inst ( .DIN1(_26452), .DIN2(_53517), .Q(_34684) );
  nnd2s1 _34518_inst ( .DIN1(_34685), .DIN2(_34686), .Q(_34661) );
  nnd2s1 _34519_inst ( .DIN1(_34687), .DIN2(_26574), .Q(_34686) );
  nnd2s1 _34520_inst ( .DIN1(_53375), .DIN2(_34688), .Q(_34687) );
  or2s1 _34521_inst ( .DIN1(_34688), .DIN2(_53375), .Q(_34685) );
  nor2s1 _34522_inst ( .DIN1(_34666), .DIN2(_34689), .Q(_34680) );
  or2s1 _34523_inst ( .DIN1(_27082), .DIN2(_53074), .Q(_34689) );
  nnd2s1 _34524_inst ( .DIN1(_28010), .DIN2(_34690), .Q(
        _____________________________26________) );
  nnd2s1 _34525_inst ( .DIN1(_34691), .DIN2(_34692), .Q(_34690) );
  nnd2s1 _34526_inst ( .DIN1(_34693), .DIN2(_34694), .Q(_34692) );
  xor2s1 _34527_inst ( .DIN1(_34695), .DIN2(_34696), .Q(_34694) );
  xor2s1 _34528_inst ( .DIN1(_53112), .DIN2(_53114), .Q(_34696) );
  nnd2s1 _34529_inst ( .DIN1(_53330), .DIN2(_53026), .Q(_34695) );
  nor2s1 _34530_inst ( .DIN1(_34306), .DIN2(_26773), .Q(_34693) );
  nnd2s1 _34531_inst ( .DIN1(_34265), .DIN2(_34697), .Q(_34691) );
  xor2s1 _34532_inst ( .DIN1(_34501), .DIN2(_34698), .Q(_34697) );
  xor2s1 _34533_inst ( .DIN1(_26451), .DIN2(_34500), .Q(_34698) );
  nnd2s1 _34534_inst ( .DIN1(_34699), .DIN2(_34700), .Q(_34500) );
  nnd2s1 _34535_inst ( .DIN1(_34701), .DIN2(_26644), .Q(_34700) );
  or2s1 _34536_inst ( .DIN1(_34702), .DIN2(_34703), .Q(_34701) );
  nnd2s1 _34537_inst ( .DIN1(_34703), .DIN2(_34702), .Q(_34699) );
  nnd2s1 _34538_inst ( .DIN1(_34704), .DIN2(_34705), .Q(
        _____________________________269________) );
  nnd2s1 _34539_inst ( .DIN1(_34706), .DIN2(_34707), .Q(_34705) );
  or2s1 _34540_inst ( .DIN1(_26720), .DIN2(_27123), .Q(_34706) );
  nnd2s1 _34541_inst ( .DIN1(_34708), .DIN2(_29096), .Q(_34704) );
  nnd2s1 _34542_inst ( .DIN1(_34709), .DIN2(_34710), .Q(_34708) );
  nnd2s1 _34543_inst ( .DIN1(_34682), .DIN2(_34711), .Q(_34710) );
  nnd2s1 _34544_inst ( .DIN1(_53076), .DIN2(_34712), .Q(_34711) );
  nnd2s1 _34545_inst ( .DIN1(_34713), .DIN2(_34656), .Q(_34709) );
  xor2s1 _34546_inst ( .DIN1(_34688), .DIN2(_34714), .Q(_34713) );
  xor2s1 _34547_inst ( .DIN1(_53129), .DIN2(_53375), .Q(_34714) );
  nnd2s1 _34548_inst ( .DIN1(_34715), .DIN2(_34716), .Q(_34688) );
  nnd2s1 _34549_inst ( .DIN1(_34717), .DIN2(_26373), .Q(_34716) );
  nnd2s1 _34550_inst ( .DIN1(_53373), .DIN2(_34718), .Q(_34717) );
  or2s1 _34551_inst ( .DIN1(_34718), .DIN2(_53373), .Q(_34715) );
  nnd2s1 _34552_inst ( .DIN1(_34719), .DIN2(_34720), .Q(
        _____________________________268________) );
  nnd2s1 _34553_inst ( .DIN1(_27233), .DIN2(_34721), .Q(_34720) );
  xnr2s1 _34554_inst ( .DIN1(_53190), .DIN2(_34722), .Q(_34721) );
  nnd2s1 _34555_inst ( .DIN1(_53075), .DIN2(_53237), .Q(_34722) );
  nnd2s1 _34556_inst ( .DIN1(_34723), .DIN2(_27227), .Q(_34719) );
  nor2s1 _34557_inst ( .DIN1(_34724), .DIN2(_34725), .Q(_34723) );
  nor2s1 _34558_inst ( .DIN1(_34682), .DIN2(_34726), .Q(_34725) );
  xor2s1 _34559_inst ( .DIN1(_34718), .DIN2(_34727), .Q(_34726) );
  xor2s1 _34560_inst ( .DIN1(_26373), .DIN2(_53373), .Q(_34727) );
  nnd2s1 _34561_inst ( .DIN1(_34728), .DIN2(_34729), .Q(_34718) );
  nnd2s1 _34562_inst ( .DIN1(_53120), .DIN2(_34730), .Q(_34729) );
  nnd2s1 _34563_inst ( .DIN1(_34731), .DIN2(_26322), .Q(_34730) );
  or2s1 _34564_inst ( .DIN1(_34731), .DIN2(_26322), .Q(_34728) );
  nor2s1 _34565_inst ( .DIN1(_34666), .DIN2(_34732), .Q(_34724) );
  nnd2s1 _34566_inst ( .DIN1(______[30]), .DIN2(_34733), .Q(_34732) );
  xor2s1 _34567_inst ( .DIN1(_53076), .DIN2(_53121), .Q(_34733) );
  nnd2s1 _34568_inst ( .DIN1(_34734), .DIN2(_34735), .Q(
        _____________________________267________) );
  nnd2s1 _34569_inst ( .DIN1(_34736), .DIN2(_34456), .Q(_34735) );
  hi1s1 _34570_inst ( .DIN(_30949), .Q(_34456) );
  nor2s1 _34571_inst ( .DIN1(_26987), .DIN2(_34737), .Q(_34736) );
  nnd2s1 _34572_inst ( .DIN1(_34738), .DIN2(_31083), .Q(_34737) );
  xor2s1 _34573_inst ( .DIN1(_53077), .DIN2(_53078), .Q(_34738) );
  nnd2s1 _34574_inst ( .DIN1(_34739), .DIN2(_30949), .Q(_34734) );
  nnd2s1 _34575_inst ( .DIN1(_34740), .DIN2(_34741), .Q(_34739) );
  nnd2s1 _34576_inst ( .DIN1(_34682), .DIN2(_34742), .Q(_34741) );
  nnd2s1 _34577_inst ( .DIN1(_34743), .DIN2(_34712), .Q(_34742) );
  xor2s1 _34578_inst ( .DIN1(_34744), .DIN2(_53079), .Q(_34743) );
  nnd2s1 _34579_inst ( .DIN1(_34745), .DIN2(_34656), .Q(_34740) );
  xor2s1 _34580_inst ( .DIN1(_34731), .DIN2(_34746), .Q(_34745) );
  xor2s1 _34581_inst ( .DIN1(_53120), .DIN2(_53374), .Q(_34746) );
  xnr2s1 _34582_inst ( .DIN1(_34747), .DIN2(_30787), .Q(_34731) );
  nnd2s1 _34583_inst ( .DIN1(_34748), .DIN2(_34749), .Q(_34747) );
  nnd2s1 _34584_inst ( .DIN1(_34750), .DIN2(_26336), .Q(_34749) );
  or2s1 _34585_inst ( .DIN1(_34751), .DIN2(_26453), .Q(_34750) );
  nnd2s1 _34586_inst ( .DIN1(_34751), .DIN2(_26453), .Q(_34748) );
  nnd2s1 _34587_inst ( .DIN1(_34752), .DIN2(_34753), .Q(
        _____________________________266________) );
  nnd2s1 _34588_inst ( .DIN1(_34754), .DIN2(______[26]), .Q(_34753) );
  and2s1 _34589_inst ( .DIN1(_27177), .DIN2(_53080), .Q(_34754) );
  nnd2s1 _34590_inst ( .DIN1(_27164), .DIN2(_34755), .Q(_34752) );
  nnd2s1 _34591_inst ( .DIN1(_34756), .DIN2(_34757), .Q(_34755) );
  nnd2s1 _34592_inst ( .DIN1(_34758), .DIN2(_34759), .Q(_34757) );
  xor2s1 _34593_inst ( .DIN1(_53081), .DIN2(_53085), .Q(_34759) );
  hi1s1 _34594_inst ( .DIN(_34666), .Q(_34758) );
  nnd2s1 _34595_inst ( .DIN1(_34682), .DIN2(_34712), .Q(_34666) );
  nnd2s1 _34596_inst ( .DIN1(_34760), .DIN2(_34656), .Q(_34756) );
  hi1s1 _34597_inst ( .DIN(_34682), .Q(_34656) );
  xor2s1 _34598_inst ( .DIN1(_34761), .DIN2(_2064), .Q(_34682) );
  nnd2s1 _34599_inst ( .DIN1(_27842), .DIN2(_34762), .Q(_34761) );
  and2s1 _34600_inst ( .DIN1(_34763), .DIN2(_34764), .Q(_27842) );
  nor2s1 _34601_inst ( .DIN1(_34765), .DIN2(_34766), .Q(_34763) );
  xnr2s1 _34602_inst ( .DIN1(_34751), .DIN2(_34767), .Q(_34760) );
  xor2s1 _34603_inst ( .DIN1(_53372), .DIN2(_53430), .Q(_34767) );
  nnd2s1 _34604_inst ( .DIN1(_34768), .DIN2(_34769), .Q(_34751) );
  nnd2s1 _34605_inst ( .DIN1(_34770), .DIN2(_26754), .Q(_34769) );
  or2s1 _34606_inst ( .DIN1(_34771), .DIN2(_26319), .Q(_34770) );
  nnd2s1 _34607_inst ( .DIN1(_34771), .DIN2(_26319), .Q(_34768) );
  nnd2s1 _34608_inst ( .DIN1(_34772), .DIN2(_30112), .Q(
        _____________________________265________) );
  nor2s1 _34609_inst ( .DIN1(_34773), .DIN2(_34774), .Q(_34772) );
  nor2s1 _34610_inst ( .DIN1(_34775), .DIN2(_28032), .Q(_34774) );
  nor2s1 _34611_inst ( .DIN1(_34776), .DIN2(_34777), .Q(_34775) );
  nnd2s1 _34612_inst ( .DIN1(_34778), .DIN2(_34779), .Q(_34777) );
  nnd2s1 _34613_inst ( .DIN1(_34780), .DIN2(_26313), .Q(_34779) );
  nnd2s1 _34614_inst ( .DIN1(_34781), .DIN2(_34782), .Q(_34778) );
  xor2s1 _34615_inst ( .DIN1(_34771), .DIN2(_34783), .Q(_34781) );
  xor2s1 _34616_inst ( .DIN1(_53124), .DIN2(_53338), .Q(_34783) );
  nnd2s1 _34617_inst ( .DIN1(_34784), .DIN2(_34785), .Q(_34771) );
  nnd2s1 _34618_inst ( .DIN1(_34786), .DIN2(_26230), .Q(_34785) );
  nnd2s1 _34619_inst ( .DIN1(_34787), .DIN2(_34788), .Q(_34786) );
  or2s1 _34620_inst ( .DIN1(_34788), .DIN2(_34787), .Q(_34784) );
  hi1s1 _34621_inst ( .DIN(_34789), .Q(_34776) );
  nor2s1 _34622_inst ( .DIN1(_53436), .DIN2(_28037), .Q(_34773) );
  nnd2s1 _34623_inst ( .DIN1(_34790), .DIN2(_34791), .Q(
        _____________________________264________) );
  nnd2s1 _34624_inst ( .DIN1(_27227), .DIN2(_34792), .Q(_34791) );
  nnd2s1 _34625_inst ( .DIN1(_34793), .DIN2(_34789), .Q(_34792) );
  nor2s1 _34626_inst ( .DIN1(_34794), .DIN2(_34795), .Q(_34793) );
  nor2s1 _34627_inst ( .DIN1(_34780), .DIN2(_34796), .Q(_34795) );
  xor2s1 _34628_inst ( .DIN1(_34788), .DIN2(_34797), .Q(_34796) );
  xor2s1 _34629_inst ( .DIN1(_26230), .DIN2(_53376), .Q(_34797) );
  nnd2s1 _34630_inst ( .DIN1(_34798), .DIN2(_34799), .Q(_34788) );
  nnd2s1 _34631_inst ( .DIN1(_53119), .DIN2(_34800), .Q(_34799) );
  nnd2s1 _34632_inst ( .DIN1(_26318), .DIN2(_34801), .Q(_34800) );
  or2s1 _34633_inst ( .DIN1(_34801), .DIN2(_26318), .Q(_34798) );
  nor2s1 _34634_inst ( .DIN1(_34782), .DIN2(_34802), .Q(_34794) );
  nor2s1 _34635_inst ( .DIN1(_27082), .DIN2(_34803), .Q(_34802) );
  nnd2s1 _34636_inst ( .DIN1(_34804), .DIN2(_34744), .Q(_34803) );
  nnd2s1 _34637_inst ( .DIN1(_53085), .DIN2(_53084), .Q(_34744) );
  nnd2s1 _34638_inst ( .DIN1(_26751), .DIN2(_26313), .Q(_34804) );
  nnd2s1 _34639_inst ( .DIN1(_27233), .DIN2(_34805), .Q(_34790) );
  xor2s1 _34640_inst ( .DIN1(_34806), .DIN2(_34807), .Q(_34805) );
  nnd2s1 _34641_inst ( .DIN1(_53082), .DIN2(_53083), .Q(_34807) );
  nnd2s1 _34642_inst ( .DIN1(_31136), .DIN2(_34808), .Q(_34806) );
  nnd2s1 _34643_inst ( .DIN1(_52947), .DIN2(_26586), .Q(_34808) );
  or2s1 _34644_inst ( .DIN1(_26586), .DIN2(_52947), .Q(_31136) );
  nor2s1 _34645_inst ( .DIN1(_27227), .DIN2(_34809), .Q(_27233) );
  nnd2s1 _34646_inst ( .DIN1(_34810), .DIN2(_34811), .Q(
        _____________________________263________) );
  nnd2s1 _34647_inst ( .DIN1(_27298), .DIN2(_34812), .Q(_34811) );
  nnd2s1 _34648_inst ( .DIN1(_34813), .DIN2(_34814), .Q(_34812) );
  nnd2s1 _34649_inst ( .DIN1(_34782), .DIN2(_34815), .Q(_34814) );
  xor2s1 _34650_inst ( .DIN1(_34801), .DIN2(_34816), .Q(_34815) );
  xor2s1 _34651_inst ( .DIN1(_53119), .DIN2(_26318), .Q(_34816) );
  nnd2s1 _34652_inst ( .DIN1(_34817), .DIN2(_34818), .Q(_34801) );
  nnd2s1 _34653_inst ( .DIN1(_34819), .DIN2(_26332), .Q(_34818) );
  nnd2s1 _34654_inst ( .DIN1(_26579), .DIN2(_34820), .Q(_34819) );
  or2s1 _34655_inst ( .DIN1(_26579), .DIN2(_34820), .Q(_34817) );
  nnd2s1 _34656_inst ( .DIN1(_34821), .DIN2(_34822), .Q(_34813) );
  xor2s1 _34657_inst ( .DIN1(_34823), .DIN2(_34824), .Q(_34821) );
  xor2s1 _34658_inst ( .DIN1(_26239), .DIN2(_53091), .Q(_34823) );
  hi1s1 _34659_inst ( .DIN(_27284), .Q(_27298) );
  nnd2s1 _34660_inst ( .DIN1(_34825), .DIN2(_34826), .Q(_27284) );
  and2s1 _34661_inst ( .DIN1(_34827), .DIN2(_34828), .Q(_34825) );
  nnd2s1 _34662_inst ( .DIN1(_34829), .DIN2(_27903), .Q(_34810) );
  nor2s1 _34663_inst ( .DIN1(_34830), .DIN2(_34831), .Q(_34829) );
  nor2s1 _34664_inst ( .DIN1(_34832), .DIN2(_34833), .Q(_34831) );
  nor2s1 _34665_inst ( .DIN1(_53513), .DIN2(_27448), .Q(_34833) );
  hi1s1 _34666_inst ( .DIN(_34834), .Q(_34832) );
  nor2s1 _34667_inst ( .DIN1(_27900), .DIN2(_34834), .Q(_34830) );
  nnd2s1 _34668_inst ( .DIN1(_26660), .DIN2(_26306), .Q(_34834) );
  nor2s1 _34669_inst ( .DIN1(_27448), .DIN2(_26454), .Q(_27900) );
  nnd2s1 _34670_inst ( .DIN1(_34835), .DIN2(_34836), .Q(
        _____________________________262________) );
  nor2s1 _34671_inst ( .DIN1(_34628), .DIN2(_34837), .Q(_34836) );
  nor2s1 _34672_inst ( .DIN1(_34838), .DIN2(_34839), .Q(_34837) );
  nnd2s1 _34673_inst ( .DIN1(_53086), .DIN2(_34780), .Q(_34839) );
  nor2s1 _34674_inst ( .DIN1(_34840), .DIN2(_34841), .Q(_34835) );
  nor2s1 _34675_inst ( .DIN1(_30949), .DIN2(_34842), .Q(_34841) );
  xor2s1 _34676_inst ( .DIN1(_53087), .DIN2(_53090), .Q(_34842) );
  nor2s1 _34677_inst ( .DIN1(_34843), .DIN2(_34844), .Q(_34840) );
  xor2s1 _34678_inst ( .DIN1(_34820), .DIN2(_34845), .Q(_34843) );
  xor2s1 _34679_inst ( .DIN1(_53379), .DIN2(_53431), .Q(_34845) );
  nnd2s1 _34680_inst ( .DIN1(_34846), .DIN2(_34847), .Q(_34820) );
  nnd2s1 _34681_inst ( .DIN1(_53307), .DIN2(_34848), .Q(_34847) );
  nnd2s1 _34682_inst ( .DIN1(_27558), .DIN2(_34849), .Q(_34848) );
  or2s1 _34683_inst ( .DIN1(_34849), .DIN2(_27558), .Q(_34846) );
  nnd2s1 _34684_inst ( .DIN1(_34850), .DIN2(_34851), .Q(
        _____________________________261________) );
  nor2s1 _34685_inst ( .DIN1(_34628), .DIN2(_34852), .Q(_34851) );
  nor2s1 _34686_inst ( .DIN1(_34838), .DIN2(_34853), .Q(_34852) );
  nnd2s1 _34687_inst ( .DIN1(_34780), .DIN2(_26256), .Q(_34853) );
  nor2s1 _34688_inst ( .DIN1(_31083), .DIN2(_30949), .Q(_34628) );
  nnd2s1 _34689_inst ( .DIN1(_34854), .DIN2(_34855), .Q(_31083) );
  nor2s1 _34690_inst ( .DIN1(_30026), .DIN2(_30029), .Q(_34854) );
  nor2s1 _34691_inst ( .DIN1(_34856), .DIN2(_34857), .Q(_34850) );
  nor2s1 _34692_inst ( .DIN1(_30949), .DIN2(_34858), .Q(_34857) );
  nor2s1 _34693_inst ( .DIN1(_34824), .DIN2(_34859), .Q(_34858) );
  nnd2s1 _34694_inst ( .DIN1(_34860), .DIN2(_34861), .Q(_34859) );
  nnd2s1 _34695_inst ( .DIN1(_26256), .DIN2(_26677), .Q(_34861) );
  nnd2s1 _34696_inst ( .DIN1(_34862), .DIN2(_53087), .Q(_34860) );
  nor2s1 _34697_inst ( .DIN1(_26355), .DIN2(_26256), .Q(_34862) );
  hi1s1 _34698_inst ( .DIN(_34863), .Q(_34824) );
  nor2s1 _34699_inst ( .DIN1(_34864), .DIN2(_34844), .Q(_34856) );
  or2s1 _34700_inst ( .DIN1(_34838), .DIN2(_34780), .Q(_34844) );
  nnd2s1 _34701_inst ( .DIN1(_30949), .DIN2(_34789), .Q(_34838) );
  nnd2s1 _34702_inst ( .DIN1(_34865), .DIN2(_34866), .Q(_34789) );
  nor2s1 _34703_inst ( .DIN1(_34782), .DIN2(_27843), .Q(_34865) );
  nor2s1 _34704_inst ( .DIN1(_34867), .DIN2(_28672), .Q(_30949) );
  nnd2s1 _34705_inst ( .DIN1(_34868), .DIN2(_34869), .Q(_28672) );
  nor2s1 _34706_inst ( .DIN1(_30029), .DIN2(_30027), .Q(_34868) );
  nnd2s1 _34707_inst ( .DIN1(_32091), .DIN2(_34870), .Q(_34867) );
  xor2s1 _34708_inst ( .DIN1(_34849), .DIN2(_34871), .Q(_34864) );
  xor2s1 _34709_inst ( .DIN1(_53307), .DIN2(_53346), .Q(_34871) );
  nnd2s1 _34710_inst ( .DIN1(_34872), .DIN2(_34873), .Q(_34849) );
  nnd2s1 _34711_inst ( .DIN1(_34874), .DIN2(_26424), .Q(_34873) );
  nnd2s1 _34712_inst ( .DIN1(_53381), .DIN2(_34875), .Q(_34874) );
  or2s1 _34713_inst ( .DIN1(_34875), .DIN2(_53381), .Q(_34872) );
  nnd2s1 _34714_inst ( .DIN1(_34876), .DIN2(_29686), .Q(
        _____________________________260________) );
  nor2s1 _34715_inst ( .DIN1(_34877), .DIN2(_34878), .Q(_34876) );
  nor2s1 _34716_inst ( .DIN1(_29689), .DIN2(_34879), .Q(_34878) );
  nnd2s1 _34717_inst ( .DIN1(_34880), .DIN2(_34881), .Q(_34879) );
  nnd2s1 _34718_inst ( .DIN1(_34882), .DIN2(_34822), .Q(_34881) );
  and2s1 _34719_inst ( .DIN1(_34780), .DIN2(_34883), .Q(_34822) );
  nnd2s1 _34720_inst ( .DIN1(_34866), .DIN2(_34884), .Q(_34883) );
  nor2s1 _34721_inst ( .DIN1(_34885), .DIN2(_34886), .Q(_34882) );
  nor2s1 _34722_inst ( .DIN1(_26239), .DIN2(_34863), .Q(_34886) );
  nnd2s1 _34723_inst ( .DIN1(_26256), .DIN2(_26355), .Q(_34863) );
  nor2s1 _34724_inst ( .DIN1(_34887), .DIN2(_26355), .Q(_34885) );
  nor2s1 _34725_inst ( .DIN1(_53091), .DIN2(_26239), .Q(_34887) );
  nnd2s1 _34726_inst ( .DIN1(_34888), .DIN2(_34782), .Q(_34880) );
  hi1s1 _34727_inst ( .DIN(_34780), .Q(_34782) );
  nnd2s1 _34728_inst ( .DIN1(_34889), .DIN2(_34444), .Q(_34780) );
  hi1s1 _34729_inst ( .DIN(_34423), .Q(_34444) );
  nnd2s1 _34730_inst ( .DIN1(_34884), .DIN2(_34890), .Q(_34423) );
  hi1s1 _34731_inst ( .DIN(_27843), .Q(_34884) );
  nor2s1 _34732_inst ( .DIN1(_34891), .DIN2(_27708), .Q(_34889) );
  nnd2s1 _34733_inst ( .DIN1(_34892), .DIN2(_34893), .Q(_27708) );
  nor2s1 _34734_inst ( .DIN1(_34894), .DIN2(_34765), .Q(_34892) );
  xnr2s1 _34735_inst ( .DIN1(_34895), .DIN2(_34875), .Q(_34888) );
  nnd2s1 _34736_inst ( .DIN1(_34896), .DIN2(_34897), .Q(_34875) );
  nnd2s1 _34737_inst ( .DIN1(_53116), .DIN2(_34898), .Q(_34897) );
  or2s1 _34738_inst ( .DIN1(_34899), .DIN2(_53380), .Q(_34898) );
  nnd2s1 _34739_inst ( .DIN1(_53380), .DIN2(_34899), .Q(_34896) );
  xor2s1 _34740_inst ( .DIN1(_26424), .DIN2(_53381), .Q(_34895) );
  and2s1 _34741_inst ( .DIN1(_29689), .DIN2(_53412), .Q(_34877) );
  nnd2s1 _34742_inst ( .DIN1(_34900), .DIN2(_34901), .Q(
        _____________________________25________) );
  nnd2s1 _34743_inst ( .DIN1(_34902), .DIN2(_27246), .Q(_34901) );
  nor2s1 _34744_inst ( .DIN1(_33158), .DIN2(_27247), .Q(_27246) );
  xnr2s1 _34745_inst ( .DIN1(_53302), .DIN2(_33159), .Q(_34902) );
  nor2s1 _34746_inst ( .DIN1(_53089), .DIN2(_53306), .Q(_33159) );
  nnd2s1 _34747_inst ( .DIN1(_27247), .DIN2(_34903), .Q(_34900) );
  nnd2s1 _34748_inst ( .DIN1(_34904), .DIN2(_34905), .Q(_34903) );
  nnd2s1 _34749_inst ( .DIN1(_34265), .DIN2(_34906), .Q(_34905) );
  xor2s1 _34750_inst ( .DIN1(_34703), .DIN2(_34907), .Q(_34906) );
  xor2s1 _34751_inst ( .DIN1(_26644), .DIN2(_34702), .Q(_34907) );
  nnd2s1 _34752_inst ( .DIN1(_34908), .DIN2(_34909), .Q(_34702) );
  nnd2s1 _34753_inst ( .DIN1(_34910), .DIN2(_26657), .Q(_34909) );
  or2s1 _34754_inst ( .DIN1(_34911), .DIN2(_34912), .Q(_34910) );
  nnd2s1 _34755_inst ( .DIN1(_34912), .DIN2(_34911), .Q(_34908) );
  and2s1 _34756_inst ( .DIN1(_34306), .DIN2(_34913), .Q(_34265) );
  nnd2s1 _34757_inst ( .DIN1(_53330), .DIN2(_34272), .Q(_34904) );
  nnd2s1 _34758_inst ( .DIN1(_34914), .DIN2(_34915), .Q(
        _____________________________259________) );
  nor2s1 _34759_inst ( .DIN1(_34916), .DIN2(_34917), .Q(_34915) );
  nor2s1 _34760_inst ( .DIN1(_34918), .DIN2(_34919), .Q(_34917) );
  nor2s1 _34761_inst ( .DIN1(_34920), .DIN2(_34921), .Q(_34918) );
  nnd2s1 _34762_inst ( .DIN1(______[16]), .DIN2(_34922), .Q(_34921) );
  nnd2s1 _34763_inst ( .DIN1(_53090), .DIN2(_26221), .Q(_34922) );
  nnd2s1 _34764_inst ( .DIN1(_34923), .DIN2(_34924), .Q(_34920) );
  nnd2s1 _34765_inst ( .DIN1(_34925), .DIN2(_26406), .Q(_34924) );
  nnd2s1 _34766_inst ( .DIN1(_53351), .DIN2(_26221), .Q(_34923) );
  nor2s1 _34767_inst ( .DIN1(_34926), .DIN2(_34927), .Q(_34916) );
  xor2s1 _34768_inst ( .DIN1(_34899), .DIN2(_34928), .Q(_34926) );
  xor2s1 _34769_inst ( .DIN1(_53116), .DIN2(_53380), .Q(_34928) );
  nnd2s1 _34770_inst ( .DIN1(_34929), .DIN2(_34930), .Q(_34899) );
  nnd2s1 _34771_inst ( .DIN1(_53133), .DIN2(_34931), .Q(_34930) );
  nnd2s1 _34772_inst ( .DIN1(_26320), .DIN2(_34932), .Q(_34931) );
  or2s1 _34773_inst ( .DIN1(_34932), .DIN2(_26320), .Q(_34929) );
  nor2s1 _34774_inst ( .DIN1(_34933), .DIN2(_34934), .Q(_34914) );
  nor2s1 _34775_inst ( .DIN1(_28137), .DIN2(_34935), .Q(_34934) );
  nor2s1 _34776_inst ( .DIN1(_27881), .DIN2(_26355), .Q(_34933) );
  nnd2s1 _34777_inst ( .DIN1(_34936), .DIN2(_34937), .Q(
        _____________________________258________) );
  nnd2s1 _34778_inst ( .DIN1(_34938), .DIN2(_34935), .Q(_34937) );
  nnd2s1 _34779_inst ( .DIN1(_34939), .DIN2(_34940), .Q(_34938) );
  nnd2s1 _34780_inst ( .DIN1(_34941), .DIN2(_34942), .Q(_34940) );
  hi1s1 _34781_inst ( .DIN(_34919), .Q(_34942) );
  nnd2s1 _34782_inst ( .DIN1(_27882), .DIN2(_34943), .Q(_34919) );
  nor2s1 _34783_inst ( .DIN1(_53087), .DIN2(_27066), .Q(_34941) );
  nnd2s1 _34784_inst ( .DIN1(_34944), .DIN2(_34945), .Q(_34939) );
  xor2s1 _34785_inst ( .DIN1(_34932), .DIN2(_34946), .Q(_34945) );
  xor2s1 _34786_inst ( .DIN1(_26450), .DIN2(_53350), .Q(_34946) );
  nnd2s1 _34787_inst ( .DIN1(_53092), .DIN2(_53352), .Q(_34932) );
  hi1s1 _34788_inst ( .DIN(_34927), .Q(_34944) );
  nnd2s1 _34789_inst ( .DIN1(_34947), .DIN2(_27882), .Q(_34927) );
  nnd2s1 _34790_inst ( .DIN1(_34948), .DIN2(_28137), .Q(_34936) );
  nnd2s1 _34791_inst ( .DIN1(_34949), .DIN2(_28139), .Q(_34948) );
  xor2s1 _34792_inst ( .DIN1(_53087), .DIN2(_53091), .Q(_34949) );
  nnd2s1 _34793_inst ( .DIN1(_34950), .DIN2(_29686), .Q(
        _____________________________257________) );
  nor2s1 _34794_inst ( .DIN1(_34951), .DIN2(_34952), .Q(_34950) );
  nor2s1 _34795_inst ( .DIN1(_29689), .DIN2(_34953), .Q(_34952) );
  nnd2s1 _34796_inst ( .DIN1(_34954), .DIN2(_34955), .Q(_34953) );
  nnd2s1 _34797_inst ( .DIN1(_34947), .DIN2(_34956), .Q(_34955) );
  xor2s1 _34798_inst ( .DIN1(_53092), .DIN2(_53352), .Q(_34956) );
  nnd2s1 _34799_inst ( .DIN1(_26701), .DIN2(_34957), .Q(_34954) );
  nnd2s1 _34800_inst ( .DIN1(_34958), .DIN2(_34959), .Q(_34957) );
  nor2s1 _34801_inst ( .DIN1(_34960), .DIN2(_34766), .Q(_34958) );
  nor2s1 _34802_inst ( .DIN1(_27154), .DIN2(_34961), .Q(_34951) );
  xor2s1 _34803_inst ( .DIN1(_26442), .DIN2(_53093), .Q(_34961) );
  nnd2s1 _34804_inst ( .DIN1(_34962), .DIN2(_34963), .Q(
        _____________________________256________) );
  nnd2s1 _34805_inst ( .DIN1(_28572), .DIN2(_34964), .Q(_34963) );
  nnd2s1 _34806_inst ( .DIN1(_34965), .DIN2(_34966), .Q(_34964) );
  nnd2s1 _34807_inst ( .DIN1(_34967), .DIN2(_53137), .Q(_34966) );
  nor2s1 _34808_inst ( .DIN1(_28321), .DIN2(_28684), .Q(_34967) );
  nor2s1 _34809_inst ( .DIN1(_34968), .DIN2(_34969), .Q(_34965) );
  nor2s1 _34810_inst ( .DIN1(_26596), .DIN2(_34970), .Q(_34969) );
  nor2s1 _34811_inst ( .DIN1(_34971), .DIN2(_34972), .Q(_34970) );
  nor2s1 _34812_inst ( .DIN1(_34345), .DIN2(_34973), .Q(_34972) );
  nor2s1 _34813_inst ( .DIN1(_34974), .DIN2(_34343), .Q(_34971) );
  nor2s1 _34814_inst ( .DIN1(_53096), .DIN2(_34975), .Q(_34968) );
  nor2s1 _34815_inst ( .DIN1(_34976), .DIN2(_34977), .Q(_34975) );
  nor2s1 _34816_inst ( .DIN1(_34343), .DIN2(_34973), .Q(_34977) );
  nor2s1 _34817_inst ( .DIN1(_34974), .DIN2(_34345), .Q(_34976) );
  hi1s1 _34818_inst ( .DIN(_34973), .Q(_34974) );
  nnd2s1 _34819_inst ( .DIN1(_34978), .DIN2(_34979), .Q(_34973) );
  nnd2s1 _34820_inst ( .DIN1(_34980), .DIN2(_26629), .Q(_34979) );
  nnd2s1 _34821_inst ( .DIN1(_26849), .DIN2(_34981), .Q(_34980) );
  hi1s1 _34822_inst ( .DIN(_34982), .Q(_34981) );
  nnd2s1 _34823_inst ( .DIN1(_34982), .DIN2(_26850), .Q(_34978) );
  nnd2s1 _34824_inst ( .DIN1(_34983), .DIN2(_28575), .Q(_34962) );
  nor2s1 _34825_inst ( .DIN1(_26405), .DIN2(_34984), .Q(_34983) );
  nnd2s1 _34826_inst ( .DIN1(______[24]), .DIN2(_34985), .Q(_34984) );
  nnd2s1 _34827_inst ( .DIN1(_34986), .DIN2(_28782), .Q(
        _____________________________255________) );
  nor2s1 _34828_inst ( .DIN1(_34987), .DIN2(_34988), .Q(_34986) );
  nor2s1 _34829_inst ( .DIN1(_28786), .DIN2(_34989), .Q(_34988) );
  nnd2s1 _34830_inst ( .DIN1(_34990), .DIN2(_34991), .Q(_34989) );
  nnd2s1 _34831_inst ( .DIN1(_34992), .DIN2(_34993), .Q(_34991) );
  nor2s1 _34832_inst ( .DIN1(_34994), .DIN2(_34995), .Q(_34993) );
  nor2s1 _34833_inst ( .DIN1(_34996), .DIN2(_27448), .Q(_34992) );
  xor2s1 _34834_inst ( .DIN1(_34997), .DIN2(_34998), .Q(_34996) );
  xor2s1 _34835_inst ( .DIN1(_53171), .DIN2(_53230), .Q(_34998) );
  nnd2s1 _34836_inst ( .DIN1(_53097), .DIN2(_26552), .Q(_34997) );
  xor2s1 _34837_inst ( .DIN1(_30349), .DIN2(_34999), .Q(_34990) );
  nnd2s1 _34838_inst ( .DIN1(_34994), .DIN2(_35000), .Q(_34999) );
  xor2s1 _34839_inst ( .DIN1(_34982), .DIN2(_35001), .Q(_35000) );
  xor2s1 _34840_inst ( .DIN1(_26629), .DIN2(_53384), .Q(_35001) );
  xor2s1 _34841_inst ( .DIN1(_35002), .DIN2(_28088), .Q(_34982) );
  nnd2s1 _34842_inst ( .DIN1(_35003), .DIN2(_35004), .Q(_35002) );
  nnd2s1 _34843_inst ( .DIN1(_53225), .DIN2(_35005), .Q(_35004) );
  nnd2s1 _34844_inst ( .DIN1(_26850), .DIN2(_35006), .Q(_35005) );
  or2s1 _34845_inst ( .DIN1(_35006), .DIN2(_26850), .Q(_35003) );
  nor2s1 _34846_inst ( .DIN1(_28792), .DIN2(_35007), .Q(_34987) );
  xnr2s1 _34847_inst ( .DIN1(_53225), .DIN2(_35008), .Q(_35007) );
  nnd2s1 _34848_inst ( .DIN1(_53097), .DIN2(_53504), .Q(_35008) );
  nnd2s1 _34849_inst ( .DIN1(_35009), .DIN2(_35010), .Q(
        _____________________________254________) );
  nnd2s1 _34850_inst ( .DIN1(_35011), .DIN2(_35012), .Q(_35010) );
  xor2s1 _34851_inst ( .DIN1(_35013), .DIN2(_53170), .Q(_35011) );
  nnd2s1 _34852_inst ( .DIN1(_35014), .DIN2(_35015), .Q(_35009) );
  nor2s1 _34853_inst ( .DIN1(_35016), .DIN2(_35017), .Q(_35014) );
  nor2s1 _34854_inst ( .DIN1(_35018), .DIN2(_35019), .Q(_35017) );
  xor2s1 _34855_inst ( .DIN1(_35006), .DIN2(_35020), .Q(_35019) );
  xor2s1 _34856_inst ( .DIN1(_53225), .DIN2(_53384), .Q(_35020) );
  nnd2s1 _34857_inst ( .DIN1(_35021), .DIN2(_35022), .Q(_35006) );
  nnd2s1 _34858_inst ( .DIN1(_53155), .DIN2(_35023), .Q(_35022) );
  nnd2s1 _34859_inst ( .DIN1(_26849), .DIN2(_35024), .Q(_35023) );
  or2s1 _34860_inst ( .DIN1(_35024), .DIN2(_26849), .Q(_35021) );
  nor2s1 _34861_inst ( .DIN1(_34994), .DIN2(_35025), .Q(_35016) );
  nnd2s1 _34862_inst ( .DIN1(_35026), .DIN2(_53097), .Q(_35025) );
  nor2s1 _34863_inst ( .DIN1(_34995), .DIN2(_28684), .Q(_35026) );
  nnd2s1 _34864_inst ( .DIN1(_35027), .DIN2(_35028), .Q(
        _____________________________253________) );
  nnd2s1 _34865_inst ( .DIN1(_35029), .DIN2(_35030), .Q(_35028) );
  xor2s1 _34866_inst ( .DIN1(_52881), .DIN2(_53180), .Q(_35030) );
  nnd2s1 _34867_inst ( .DIN1(_35031), .DIN2(_29206), .Q(_35027) );
  nor2s1 _34868_inst ( .DIN1(_35032), .DIN2(_35033), .Q(_35031) );
  nor2s1 _34869_inst ( .DIN1(_35018), .DIN2(_35034), .Q(_35033) );
  xor2s1 _34870_inst ( .DIN1(_35035), .DIN2(_35024), .Q(_35034) );
  xnr2s1 _34871_inst ( .DIN1(_35036), .DIN2(_35037), .Q(_35024) );
  nnd2s1 _34872_inst ( .DIN1(_35038), .DIN2(_35039), .Q(_35036) );
  nnd2s1 _34873_inst ( .DIN1(_35040), .DIN2(_26616), .Q(_35039) );
  or2s1 _34874_inst ( .DIN1(_35041), .DIN2(_34312), .Q(_35040) );
  nnd2s1 _34875_inst ( .DIN1(_35041), .DIN2(_34312), .Q(_35038) );
  xor2s1 _34876_inst ( .DIN1(_26455), .DIN2(_53384), .Q(_35035) );
  nor2s1 _34877_inst ( .DIN1(_34994), .DIN2(_35042), .Q(_35032) );
  nor2s1 _34878_inst ( .DIN1(_53171), .DIN2(_34995), .Q(_35042) );
  nnd2s1 _34879_inst ( .DIN1(_35043), .DIN2(_35044), .Q(
        _____________________________252________) );
  nor2s1 _34880_inst ( .DIN1(_35045), .DIN2(_35046), .Q(_35044) );
  nor2s1 _34881_inst ( .DIN1(_28016), .DIN2(_35047), .Q(_35046) );
  nor2s1 _34882_inst ( .DIN1(_35048), .DIN2(_35049), .Q(_35047) );
  nor2s1 _34883_inst ( .DIN1(_35018), .DIN2(_35050), .Q(_35049) );
  xnr2s1 _34884_inst ( .DIN1(_35051), .DIN2(_35041), .Q(_35050) );
  nnd2s1 _34885_inst ( .DIN1(_35052), .DIN2(_35053), .Q(_35041) );
  nnd2s1 _34886_inst ( .DIN1(_35054), .DIN2(_26422), .Q(_35053) );
  or2s1 _34887_inst ( .DIN1(_35055), .DIN2(_34325), .Q(_35054) );
  nnd2s1 _34888_inst ( .DIN1(_34325), .DIN2(_35055), .Q(_35052) );
  xor2s1 _34889_inst ( .DIN1(_34312), .DIN2(_53098), .Q(_35051) );
  nnd2s1 _34890_inst ( .DIN1(_35056), .DIN2(_35057), .Q(_34312) );
  nnd2s1 _34891_inst ( .DIN1(_35058), .DIN2(_35059), .Q(_35057) );
  nor2s1 _34892_inst ( .DIN1(_34994), .DIN2(_35060), .Q(_35048) );
  nor2s1 _34893_inst ( .DIN1(_34995), .DIN2(_35061), .Q(_35060) );
  xor2s1 _34894_inst ( .DIN1(_26552), .DIN2(_53171), .Q(_35061) );
  nor2s1 _34895_inst ( .DIN1(_28024), .DIN2(_35062), .Q(_35045) );
  nnd2s1 _34896_inst ( .DIN1(_53099), .DIN2(_35063), .Q(_35062) );
  nor2s1 _34897_inst ( .DIN1(_35064), .DIN2(_35065), .Q(_35043) );
  nor2s1 _34898_inst ( .DIN1(_53099), .DIN2(_28027), .Q(_35065) );
  nnd2s1 _34899_inst ( .DIN1(_35066), .DIN2(_35067), .Q(
        _____________________________251________) );
  nnd2s1 _34900_inst ( .DIN1(_35068), .DIN2(_35069), .Q(_35067) );
  nnd2s1 _34901_inst ( .DIN1(_35070), .DIN2(_53171), .Q(_35068) );
  nor2s1 _34902_inst ( .DIN1(_35071), .DIN2(_27066), .Q(_35070) );
  nor2s1 _34903_inst ( .DIN1(_35072), .DIN2(_35073), .Q(_35066) );
  nor2s1 _34904_inst ( .DIN1(_35074), .DIN2(_35075), .Q(_35073) );
  xnr2s1 _34905_inst ( .DIN1(_34325), .DIN2(_35076), .Q(_35075) );
  xor2s1 _34906_inst ( .DIN1(_26422), .DIN2(_35055), .Q(_35076) );
  nnd2s1 _34907_inst ( .DIN1(_35077), .DIN2(_35078), .Q(_35055) );
  nnd2s1 _34908_inst ( .DIN1(_53428), .DIN2(_35079), .Q(_35078) );
  or2s1 _34909_inst ( .DIN1(_35080), .DIN2(_34501), .Q(_35079) );
  nnd2s1 _34910_inst ( .DIN1(_34501), .DIN2(_35080), .Q(_35077) );
  hi1s1 _34911_inst ( .DIN(_35081), .Q(_34501) );
  xnr2s1 _34912_inst ( .DIN1(_35058), .DIN2(_35082), .Q(_34325) );
  nnd2s1 _34913_inst ( .DIN1(_35083), .DIN2(_35084), .Q(_35058) );
  nnd2s1 _34914_inst ( .DIN1(_53364), .DIN2(_35085), .Q(_35084) );
  or2s1 _34915_inst ( .DIN1(_35086), .DIN2(_35087), .Q(_35085) );
  nnd2s1 _34916_inst ( .DIN1(_35087), .DIN2(_35086), .Q(_35083) );
  nor2s1 _34917_inst ( .DIN1(_35088), .DIN2(_35089), .Q(_35072) );
  nnd2s1 _34918_inst ( .DIN1(_35090), .DIN2(_35091), .Q(_35089) );
  xor2s1 _34919_inst ( .DIN1(_53109), .DIN2(_53415), .Q(_35090) );
  nnd2s1 _34920_inst ( .DIN1(_35092), .DIN2(_35093), .Q(
        _____________________________250________) );
  nnd2s1 _34921_inst ( .DIN1(_35094), .DIN2(_35095), .Q(_35093) );
  nnd2s1 _34922_inst ( .DIN1(_35096), .DIN2(_35097), .Q(_35095) );
  xor2s1 _34923_inst ( .DIN1(_26482), .DIN2(_35098), .Q(_35097) );
  and2s1 _34924_inst ( .DIN1(_26410), .DIN2(_53101), .Q(_35098) );
  nor2s1 _34925_inst ( .DIN1(_34995), .DIN2(_27651), .Q(_35096) );
  hi1s1 _34926_inst ( .DIN(_35091), .Q(_34995) );
  nnd2s1 _34927_inst ( .DIN1(_35099), .DIN2(_35100), .Q(_35091) );
  nor2s1 _34928_inst ( .DIN1(_35101), .DIN2(_35102), .Q(_35100) );
  nnd2s1 _34929_inst ( .DIN1(_35103), .DIN2(_35104), .Q(_35102) );
  hi1s1 _34930_inst ( .DIN(_35088), .Q(_35094) );
  nnd2s1 _34931_inst ( .DIN1(_35105), .DIN2(_35018), .Q(_35088) );
  nor2s1 _34932_inst ( .DIN1(_35106), .DIN2(_35107), .Q(_35092) );
  nor2s1 _34933_inst ( .DIN1(_35108), .DIN2(_35109), .Q(_35107) );
  xor2s1 _34934_inst ( .DIN1(_26482), .DIN2(_53171), .Q(_35108) );
  nor2s1 _34935_inst ( .DIN1(_35110), .DIN2(_35074), .Q(_35106) );
  nnd2s1 _34936_inst ( .DIN1(_35105), .DIN2(_34994), .Q(_35074) );
  hi1s1 _34937_inst ( .DIN(_35018), .Q(_34994) );
  nnd2s1 _34938_inst ( .DIN1(_35111), .DIN2(_35112), .Q(_35018) );
  nor2s1 _34939_inst ( .DIN1(_35113), .DIN2(_35114), .Q(_35112) );
  nor2s1 _34940_inst ( .DIN1(_35115), .DIN2(_35116), .Q(_35111) );
  xor2s1 _34941_inst ( .DIN1(_35081), .DIN2(_35117), .Q(_35110) );
  xor2s1 _34942_inst ( .DIN1(_26500), .DIN2(_35080), .Q(_35117) );
  nnd2s1 _34943_inst ( .DIN1(_35118), .DIN2(_35119), .Q(_35080) );
  nnd2s1 _34944_inst ( .DIN1(_35120), .DIN2(_26263), .Q(_35119) );
  nnd2s1 _34945_inst ( .DIN1(_35121), .DIN2(_35122), .Q(_35120) );
  xor2s1 _34946_inst ( .DIN1(_35037), .DIN2(_35123), .Q(_35118) );
  nor2s1 _34947_inst ( .DIN1(_35121), .DIN2(_35122), .Q(_35123) );
  xor2s1 _34948_inst ( .DIN1(_35087), .DIN2(_35124), .Q(_35081) );
  xor2s1 _34949_inst ( .DIN1(_27620), .DIN2(_35086), .Q(_35124) );
  nnd2s1 _34950_inst ( .DIN1(_35125), .DIN2(_35126), .Q(_35086) );
  nnd2s1 _34951_inst ( .DIN1(_35127), .DIN2(_26338), .Q(_35126) );
  nnd2s1 _34952_inst ( .DIN1(_35128), .DIN2(_35129), .Q(_35127) );
  xor2s1 _34953_inst ( .DIN1(_31752), .DIN2(_35130), .Q(_35125) );
  nor2s1 _34954_inst ( .DIN1(_35128), .DIN2(_35129), .Q(_35130) );
  nnd2s1 _34955_inst ( .DIN1(_35131), .DIN2(_35132), .Q(
        _____________________________24________) );
  nor2s1 _34956_inst ( .DIN1(_35133), .DIN2(_35134), .Q(_35132) );
  nor2s1 _34957_inst ( .DIN1(_35135), .DIN2(_35136), .Q(_35134) );
  xor2s1 _34958_inst ( .DIN1(_34912), .DIN2(_35137), .Q(_35135) );
  xor2s1 _34959_inst ( .DIN1(_26657), .DIN2(_34911), .Q(_35137) );
  nnd2s1 _34960_inst ( .DIN1(_35138), .DIN2(_35139), .Q(_34911) );
  nnd2s1 _34961_inst ( .DIN1(_35140), .DIN2(_26717), .Q(_35139) );
  or2s1 _34962_inst ( .DIN1(_35141), .DIN2(_35142), .Q(_35140) );
  nnd2s1 _34963_inst ( .DIN1(_35142), .DIN2(_35141), .Q(_35138) );
  nor2s1 _34964_inst ( .DIN1(_35143), .DIN2(_35144), .Q(_35131) );
  nor2s1 _34965_inst ( .DIN1(_34300), .DIN2(_35145), .Q(_35144) );
  xor2s1 _34966_inst ( .DIN1(_26399), .DIN2(_53102), .Q(_35145) );
  nor2s1 _34967_inst ( .DIN1(_35146), .DIN2(_35147), .Q(_35143) );
  nor2s1 _34968_inst ( .DIN1(_53114), .DIN2(_27365), .Q(_35146) );
  nnd2s1 _34969_inst ( .DIN1(_35148), .DIN2(_35149), .Q(
        _____________________________249________) );
  nnd2s1 _34970_inst ( .DIN1(_35150), .DIN2(_35069), .Q(_35149) );
  nnd2s1 _34971_inst ( .DIN1(_35151), .DIN2(______[4]), .Q(_35150) );
  nor2s1 _34972_inst ( .DIN1(_35071), .DIN2(_35152), .Q(_35151) );
  xor2s1 _34973_inst ( .DIN1(_35153), .DIN2(_35154), .Q(_35152) );
  xor2s1 _34974_inst ( .DIN1(_53109), .DIN2(_53110), .Q(_35154) );
  nnd2s1 _34975_inst ( .DIN1(_53108), .DIN2(_53109), .Q(_35153) );
  nor2s1 _34976_inst ( .DIN1(_35155), .DIN2(_35156), .Q(_35148) );
  nor2s1 _34977_inst ( .DIN1(_35157), .DIN2(_35158), .Q(_35156) );
  xor2s1 _34978_inst ( .DIN1(_34703), .DIN2(_35159), .Q(_35158) );
  xor2s1 _34979_inst ( .DIN1(_26263), .DIN2(_35122), .Q(_35159) );
  nnd2s1 _34980_inst ( .DIN1(_35160), .DIN2(_35161), .Q(_35122) );
  nnd2s1 _34981_inst ( .DIN1(_53398), .DIN2(_35162), .Q(_35161) );
  nnd2s1 _34982_inst ( .DIN1(_34912), .DIN2(_35163), .Q(_35162) );
  or2s1 _34983_inst ( .DIN1(_35163), .DIN2(_34912), .Q(_35160) );
  hi1s1 _34984_inst ( .DIN(_35121), .Q(_34703) );
  xor2s1 _34985_inst ( .DIN1(_35129), .DIN2(_35164), .Q(_35121) );
  xor2s1 _34986_inst ( .DIN1(_53362), .DIN2(_35128), .Q(_35164) );
  and2s1 _34987_inst ( .DIN1(_35165), .DIN2(_35166), .Q(_35128) );
  nnd2s1 _34988_inst ( .DIN1(_35167), .DIN2(_34515), .Q(_35166) );
  or2s1 _34989_inst ( .DIN1(_35168), .DIN2(_35169), .Q(_35167) );
  nnd2s1 _34990_inst ( .DIN1(_35169), .DIN2(_35168), .Q(_35165) );
  nor2s1 _34991_inst ( .DIN1(_35170), .DIN2(_35171), .Q(_35155) );
  nnd2s1 _34992_inst ( .DIN1(_35172), .DIN2(_53101), .Q(_35171) );
  nnd2s1 _34993_inst ( .DIN1(______[18]), .DIN2(_35116), .Q(_35170) );
  nnd2s1 _34994_inst ( .DIN1(_35173), .DIN2(_35174), .Q(
        _____________________________248________) );
  nnd2s1 _34995_inst ( .DIN1(_35172), .DIN2(_35175), .Q(_35174) );
  nnd2s1 _34996_inst ( .DIN1(_35176), .DIN2(_35116), .Q(_35175) );
  xor2s1 _34997_inst ( .DIN1(_53172), .DIN2(_53415), .Q(_35176) );
  hi1s1 _34998_inst ( .DIN(_35177), .Q(_35172) );
  nor2s1 _34999_inst ( .DIN1(_35178), .DIN2(_35179), .Q(_35173) );
  nor2s1 _35000_inst ( .DIN1(_35180), .DIN2(_35157), .Q(_35179) );
  xor2s1 _35001_inst ( .DIN1(_34912), .DIN2(_35181), .Q(_35180) );
  xor2s1 _35002_inst ( .DIN1(_26543), .DIN2(_35163), .Q(_35181) );
  nnd2s1 _35003_inst ( .DIN1(_35182), .DIN2(_35183), .Q(_35163) );
  nnd2s1 _35004_inst ( .DIN1(_53145), .DIN2(_35184), .Q(_35183) );
  or2s1 _35005_inst ( .DIN1(_35185), .DIN2(_35142), .Q(_35184) );
  nnd2s1 _35006_inst ( .DIN1(_35142), .DIN2(_35185), .Q(_35182) );
  xor2s1 _35007_inst ( .DIN1(_35169), .DIN2(_26763), .Q(_34912) );
  nnd2s1 _35008_inst ( .DIN1(_35186), .DIN2(_35187), .Q(_35168) );
  nnd2s1 _35009_inst ( .DIN1(_53365), .DIN2(_35188), .Q(_35187) );
  or2s1 _35010_inst ( .DIN1(_35189), .DIN2(_35190), .Q(_35188) );
  nnd2s1 _35011_inst ( .DIN1(_35190), .DIN2(_35189), .Q(_35186) );
  nor2s1 _35012_inst ( .DIN1(_35109), .DIN2(_35191), .Q(_35178) );
  nnd2s1 _35013_inst ( .DIN1(_53415), .DIN2(______[28]), .Q(_35191) );
  nnd2s1 _35014_inst ( .DIN1(_35192), .DIN2(_27983), .Q(
        _____________________________247________) );
  nor2s1 _35015_inst ( .DIN1(_35193), .DIN2(_35194), .Q(_35192) );
  nor2s1 _35016_inst ( .DIN1(_27500), .DIN2(_35195), .Q(_35194) );
  nor2s1 _35017_inst ( .DIN1(_35196), .DIN2(_35197), .Q(_35195) );
  nor2s1 _35018_inst ( .DIN1(_35198), .DIN2(_35199), .Q(_35197) );
  xnr2s1 _35019_inst ( .DIN1(_35142), .DIN2(_35200), .Q(_35199) );
  xor2s1 _35020_inst ( .DIN1(_26236), .DIN2(_35185), .Q(_35200) );
  nnd2s1 _35021_inst ( .DIN1(_35201), .DIN2(_35202), .Q(_35185) );
  nnd2s1 _35022_inst ( .DIN1(_53146), .DIN2(_35203), .Q(_35202) );
  or2s1 _35023_inst ( .DIN1(_35204), .DIN2(_35205), .Q(_35203) );
  nnd2s1 _35024_inst ( .DIN1(_35205), .DIN2(_35204), .Q(_35201) );
  nor2s1 _35025_inst ( .DIN1(_35206), .DIN2(_35207), .Q(_35196) );
  nor2s1 _35026_inst ( .DIN1(_35208), .DIN2(_35209), .Q(_35207) );
  xor2s1 _35027_inst ( .DIN1(_53071), .DIN2(_53108), .Q(_35209) );
  nor2s1 _35028_inst ( .DIN1(_27994), .DIN2(_26265), .Q(_35193) );
  nor2s1 _35029_inst ( .DIN1(_35210), .DIN2(_31037), .Q(
        _____________________________246________) );
  nor2s1 _35030_inst ( .DIN1(_35211), .DIN2(_35212), .Q(_35210) );
  nnd2s1 _35031_inst ( .DIN1(_35213), .DIN2(_35214), .Q(_35212) );
  or2s1 _35032_inst ( .DIN1(_35215), .DIN2(_53105), .Q(_35213) );
  nnd2s1 _35033_inst ( .DIN1(_35216), .DIN2(_35217), .Q(_35211) );
  nnd2s1 _35034_inst ( .DIN1(_35218), .DIN2(_35198), .Q(_35217) );
  nnd2s1 _35035_inst ( .DIN1(______[28]), .DIN2(_35219), .Q(_35218) );
  nnd2s1 _35036_inst ( .DIN1(_53105), .DIN2(_26547), .Q(_35219) );
  nnd2s1 _35037_inst ( .DIN1(_35220), .DIN2(_35206), .Q(_35216) );
  xor2s1 _35038_inst ( .DIN1(_35205), .DIN2(_35221), .Q(_35220) );
  xor2s1 _35039_inst ( .DIN1(_26517), .DIN2(_35204), .Q(_35221) );
  nnd2s1 _35040_inst ( .DIN1(_35222), .DIN2(_35223), .Q(_35204) );
  nnd2s1 _35041_inst ( .DIN1(_35224), .DIN2(_26460), .Q(_35223) );
  or2s1 _35042_inst ( .DIN1(_35225), .DIN2(_35226), .Q(_35224) );
  xor2s1 _35043_inst ( .DIN1(_29544), .DIN2(_35227), .Q(_35222) );
  nnd2s1 _35044_inst ( .DIN1(_35226), .DIN2(_35225), .Q(_35227) );
  nnd2s1 _35045_inst ( .DIN1(_35228), .DIN2(_35229), .Q(
        _____________________________245________) );
  nnd2s1 _35046_inst ( .DIN1(_35230), .DIN2(_53109), .Q(_35229) );
  nor2s1 _35047_inst ( .DIN1(_35231), .DIN2(_35232), .Q(_35228) );
  nor2s1 _35048_inst ( .DIN1(_35233), .DIN2(_35157), .Q(_35232) );
  nnd2s1 _35049_inst ( .DIN1(_35206), .DIN2(_35105), .Q(_35157) );
  xor2s1 _35050_inst ( .DIN1(_35226), .DIN2(_35234), .Q(_35233) );
  xor2s1 _35051_inst ( .DIN1(_26460), .DIN2(_35225), .Q(_35234) );
  nnd2s1 _35052_inst ( .DIN1(_35235), .DIN2(_35236), .Q(_35225) );
  nnd2s1 _35053_inst ( .DIN1(_53147), .DIN2(_35237), .Q(_35236) );
  or2s1 _35054_inst ( .DIN1(_35238), .DIN2(_35239), .Q(_35237) );
  xor2s1 _35055_inst ( .DIN1(_33328), .DIN2(_35240), .Q(_35235) );
  nnd2s1 _35056_inst ( .DIN1(_35239), .DIN2(_35238), .Q(_35240) );
  nor2s1 _35057_inst ( .DIN1(_35241), .DIN2(_35177), .Q(_35231) );
  nnd2s1 _35058_inst ( .DIN1(_35105), .DIN2(_35198), .Q(_35177) );
  nor2s1 _35059_inst ( .DIN1(_35208), .DIN2(_53105), .Q(_35241) );
  hi1s1 _35060_inst ( .DIN(_35116), .Q(_35208) );
  nnd2s1 _35061_inst ( .DIN1(_35242), .DIN2(_27560), .Q(
        _____________________________244________) );
  nnd2s1 _35062_inst ( .DIN1(_28744), .DIN2(_27563), .Q(_27560) );
  nor2s1 _35063_inst ( .DIN1(_35243), .DIN2(_35244), .Q(_35242) );
  nor2s1 _35064_inst ( .DIN1(_27571), .DIN2(_35245), .Q(_35244) );
  xor2s1 _35065_inst ( .DIN1(_53106), .DIN2(_53107), .Q(_35245) );
  nor2s1 _35066_inst ( .DIN1(_35246), .DIN2(_27563), .Q(_35243) );
  nor2s1 _35067_inst ( .DIN1(_35247), .DIN2(_35248), .Q(_35246) );
  nnd2s1 _35068_inst ( .DIN1(_35215), .DIN2(_35214), .Q(_35248) );
  nnd2s1 _35069_inst ( .DIN1(_35249), .DIN2(_35198), .Q(_35214) );
  nnd2s1 _35070_inst ( .DIN1(_35116), .DIN2(_35250), .Q(_35249) );
  nnd2s1 _35071_inst ( .DIN1(_53108), .DIN2(_26547), .Q(_35250) );
  nnd2s1 _35072_inst ( .DIN1(_35251), .DIN2(_35252), .Q(_35116) );
  nor2s1 _35073_inst ( .DIN1(_35253), .DIN2(_35254), .Q(_35252) );
  nor2s1 _35074_inst ( .DIN1(_35255), .DIN2(_35256), .Q(_35251) );
  nnd2s1 _35075_inst ( .DIN1(_35257), .DIN2(_53104), .Q(_35215) );
  nor2s1 _35076_inst ( .DIN1(_53108), .DIN2(_35206), .Q(_35257) );
  hi1s1 _35077_inst ( .DIN(_35198), .Q(_35206) );
  nor2s1 _35078_inst ( .DIN1(_35198), .DIN2(_35258), .Q(_35247) );
  xor2s1 _35079_inst ( .DIN1(_35259), .DIN2(_35260), .Q(_35258) );
  xnr2s1 _35080_inst ( .DIN1(_53147), .DIN2(_35238), .Q(_35260) );
  nnd2s1 _35081_inst ( .DIN1(_35261), .DIN2(_35262), .Q(_35238) );
  nnd2s1 _35082_inst ( .DIN1(_35263), .DIN2(_26648), .Q(_35262) );
  or2s1 _35083_inst ( .DIN1(_35264), .DIN2(_35265), .Q(_35263) );
  nnd2s1 _35084_inst ( .DIN1(_35265), .DIN2(_35264), .Q(_35261) );
  hi1s1 _35085_inst ( .DIN(_35239), .Q(_35259) );
  nnd2s1 _35086_inst ( .DIN1(_35266), .DIN2(_35267), .Q(_35198) );
  nor2s1 _35087_inst ( .DIN1(_35255), .DIN2(_35268), .Q(_35267) );
  nnd2s1 _35088_inst ( .DIN1(_35269), .DIN2(_35270), .Q(_35268) );
  hi1s1 _35089_inst ( .DIN(_35271), .Q(_35255) );
  nor2s1 _35090_inst ( .DIN1(_35272), .DIN2(_35273), .Q(_35266) );
  nnd2s1 _35091_inst ( .DIN1(_35274), .DIN2(_35275), .Q(
        _____________________________243________) );
  nnd2s1 _35092_inst ( .DIN1(_35276), .DIN2(_35230), .Q(_35275) );
  hi1s1 _35093_inst ( .DIN(_35109), .Q(_35230) );
  nnd2s1 _35094_inst ( .DIN1(_35277), .DIN2(_35069), .Q(_35109) );
  nor2s1 _35095_inst ( .DIN1(_35278), .DIN2(_28684), .Q(_35276) );
  xor2s1 _35096_inst ( .DIN1(_35279), .DIN2(_53108), .Q(_35278) );
  nnd2s1 _35097_inst ( .DIN1(_53110), .DIN2(_53109), .Q(_35279) );
  nnd2s1 _35098_inst ( .DIN1(_35105), .DIN2(_35280), .Q(_35274) );
  nnd2s1 _35099_inst ( .DIN1(_35281), .DIN2(_35282), .Q(_35280) );
  nor2s1 _35100_inst ( .DIN1(_35283), .DIN2(_35284), .Q(_35281) );
  nor2s1 _35101_inst ( .DIN1(_35285), .DIN2(_35286), .Q(_35284) );
  xor2s1 _35102_inst ( .DIN1(_35265), .DIN2(_35287), .Q(_35286) );
  xor2s1 _35103_inst ( .DIN1(_26648), .DIN2(_35264), .Q(_35287) );
  nnd2s1 _35104_inst ( .DIN1(_35288), .DIN2(_35289), .Q(_35264) );
  nnd2s1 _35105_inst ( .DIN1(_35290), .DIN2(_53148), .Q(_35289) );
  xor2s1 _35106_inst ( .DIN1(_35291), .DIN2(_35292), .Q(_35290) );
  nnd2s1 _35107_inst ( .DIN1(_35293), .DIN2(_35294), .Q(_35288) );
  nor2s1 _35108_inst ( .DIN1(_35295), .DIN2(_35296), .Q(_35283) );
  xnr2s1 _35109_inst ( .DIN1(_35297), .DIN2(_35298), .Q(_35296) );
  xor2s1 _35110_inst ( .DIN1(_53355), .DIN2(_53523), .Q(_35298) );
  hi1s1 _35111_inst ( .DIN(_35069), .Q(_35105) );
  nnd2s1 _35112_inst ( .DIN1(_35299), .DIN2(_35300), .Q(_35069) );
  nor2s1 _35113_inst ( .DIN1(_35301), .DIN2(_35302), .Q(_35299) );
  nnd2s1 _35114_inst ( .DIN1(_35303), .DIN2(_27644), .Q(
        _____________________________242________) );
  nor2s1 _35115_inst ( .DIN1(_35304), .DIN2(_35305), .Q(_35303) );
  nor2s1 _35116_inst ( .DIN1(_27648), .DIN2(_35306), .Q(_35305) );
  nnd2s1 _35117_inst ( .DIN1(_35307), .DIN2(_35308), .Q(_35306) );
  nnd2s1 _35118_inst ( .DIN1(_35309), .DIN2(_26713), .Q(_35308) );
  nnd2s1 _35119_inst ( .DIN1(_35310), .DIN2(_35295), .Q(_35307) );
  nor2s1 _35120_inst ( .DIN1(_35311), .DIN2(_35312), .Q(_35310) );
  nor2s1 _35121_inst ( .DIN1(_26609), .DIN2(_35313), .Q(_35312) );
  xor2s1 _35122_inst ( .DIN1(_35294), .DIN2(_35314), .Q(_35313) );
  nor2s1 _35123_inst ( .DIN1(_53148), .DIN2(_35315), .Q(_35311) );
  nor2s1 _35124_inst ( .DIN1(_35316), .DIN2(_35292), .Q(_35315) );
  nor2s1 _35125_inst ( .DIN1(_35294), .DIN2(_35293), .Q(_35292) );
  and2s1 _35126_inst ( .DIN1(_35294), .DIN2(_35293), .Q(_35316) );
  nnd2s1 _35127_inst ( .DIN1(_35317), .DIN2(_35318), .Q(_35294) );
  nnd2s1 _35128_inst ( .DIN1(_35319), .DIN2(_26661), .Q(_35318) );
  nnd2s1 _35129_inst ( .DIN1(_35320), .DIN2(_35321), .Q(_35319) );
  hi1s1 _35130_inst ( .DIN(_35322), .Q(_35321) );
  nnd2s1 _35131_inst ( .DIN1(_35322), .DIN2(_35323), .Q(_35317) );
  nor2s1 _35132_inst ( .DIN1(_27655), .DIN2(_35324), .Q(_35304) );
  xor2s1 _35133_inst ( .DIN1(_53277), .DIN2(_53356), .Q(_35324) );
  nnd2s1 _35134_inst ( .DIN1(_35325), .DIN2(_27676), .Q(
        _____________________________241________) );
  nnd2s1 _35135_inst ( .DIN1(_33522), .DIN2(_27679), .Q(_27676) );
  nor2s1 _35136_inst ( .DIN1(_35326), .DIN2(_35327), .Q(_35325) );
  nor2s1 _35137_inst ( .DIN1(_27679), .DIN2(_35328), .Q(_35327) );
  nnd2s1 _35138_inst ( .DIN1(_35329), .DIN2(_35330), .Q(_35328) );
  nnd2s1 _35139_inst ( .DIN1(_35309), .DIN2(_53355), .Q(_35330) );
  hi1s1 _35140_inst ( .DIN(_35331), .Q(_35309) );
  nnd2s1 _35141_inst ( .DIN1(_35332), .DIN2(_35295), .Q(_35329) );
  xor2s1 _35142_inst ( .DIN1(_35322), .DIN2(_35333), .Q(_35332) );
  xor2s1 _35143_inst ( .DIN1(_53111), .DIN2(_35320), .Q(_35333) );
  hi1s1 _35144_inst ( .DIN(_35323), .Q(_35320) );
  nnd2s1 _35145_inst ( .DIN1(_35334), .DIN2(_35335), .Q(_35323) );
  nnd2s1 _35146_inst ( .DIN1(_35336), .DIN2(_26495), .Q(_35335) );
  or2s1 _35147_inst ( .DIN1(_35337), .DIN2(_35338), .Q(_35336) );
  nnd2s1 _35148_inst ( .DIN1(_35338), .DIN2(_35337), .Q(_35334) );
  nor2s1 _35149_inst ( .DIN1(_27684), .DIN2(_35339), .Q(_35326) );
  nor2s1 _35150_inst ( .DIN1(_26988), .DIN2(_26690), .Q(_35339) );
  nnd2s1 _35151_inst ( .DIN1(_35340), .DIN2(_27998), .Q(
        _____________________________240________) );
  hi1s1 _35152_inst ( .DIN(_33544), .Q(_27998) );
  nor2s1 _35153_inst ( .DIN1(_35341), .DIN2(_35342), .Q(_33544) );
  nor2s1 _35154_inst ( .DIN1(_35343), .DIN2(_35344), .Q(_35340) );
  nor2s1 _35155_inst ( .DIN1(_27749), .DIN2(_35345), .Q(_35344) );
  nnd2s1 _35156_inst ( .DIN1(_35346), .DIN2(_35347), .Q(_35345) );
  nnd2s1 _35157_inst ( .DIN1(_35348), .DIN2(_35295), .Q(_35347) );
  xor2s1 _35158_inst ( .DIN1(_35338), .DIN2(_35349), .Q(_35348) );
  xor2s1 _35159_inst ( .DIN1(_26495), .DIN2(_35337), .Q(_35349) );
  nnd2s1 _35160_inst ( .DIN1(_35350), .DIN2(_35351), .Q(_35337) );
  nnd2s1 _35161_inst ( .DIN1(_53152), .DIN2(_35352), .Q(_35351) );
  nnd2s1 _35162_inst ( .DIN1(_35353), .DIN2(_35354), .Q(_35352) );
  hi1s1 _35163_inst ( .DIN(_35355), .Q(_35354) );
  nnd2s1 _35164_inst ( .DIN1(_35355), .DIN2(_35356), .Q(_35350) );
  nnd2s1 _35165_inst ( .DIN1(_35357), .DIN2(_35358), .Q(_35346) );
  nor2s1 _35166_inst ( .DIN1(_35359), .DIN2(_35360), .Q(_35358) );
  nor2s1 _35167_inst ( .DIN1(_26258), .DIN2(_35297), .Q(_35360) );
  nnd2s1 _35168_inst ( .DIN1(_53355), .DIN2(_53131), .Q(_35297) );
  nor2s1 _35169_inst ( .DIN1(_53131), .DIN2(_35361), .Q(_35359) );
  nor2s1 _35170_inst ( .DIN1(_26258), .DIN2(_26449), .Q(_35361) );
  nor2s1 _35171_inst ( .DIN1(_26987), .DIN2(_35331), .Q(_35357) );
  nor2s1 _35172_inst ( .DIN1(_28010), .DIN2(_35362), .Q(_35343) );
  nor2s1 _35173_inst ( .DIN1(_53188), .DIN2(_27365), .Q(_35362) );
  nnd2s1 _35174_inst ( .DIN1(_35363), .DIN2(_35364), .Q(
        _____________________________23________) );
  nnd2s1 _35175_inst ( .DIN1(_35365), .DIN2(_35366), .Q(_35364) );
  xor2s1 _35176_inst ( .DIN1(_27574), .DIN2(_53317), .Q(_35366) );
  nnd2s1 _35177_inst ( .DIN1(_53112), .DIN2(_53113), .Q(_27574) );
  nor2s1 _35178_inst ( .DIN1(_28744), .DIN2(_27651), .Q(_35365) );
  nnd2s1 _35179_inst ( .DIN1(_35367), .DIN2(_27571), .Q(_35363) );
  hi1s1 _35180_inst ( .DIN(_27563), .Q(_27571) );
  nnd2s1 _35181_inst ( .DIN1(_33158), .DIN2(_35368), .Q(_27563) );
  hi1s1 _35182_inst ( .DIN(_31027), .Q(_33158) );
  nnd2s1 _35183_inst ( .DIN1(_28744), .DIN2(_35369), .Q(_31027) );
  nor2s1 _35184_inst ( .DIN1(_30854), .DIN2(_35370), .Q(_28744) );
  nor2s1 _35185_inst ( .DIN1(_35371), .DIN2(_35372), .Q(_35367) );
  nor2s1 _35186_inst ( .DIN1(_35373), .DIN2(_35374), .Q(_35372) );
  xnr2s1 _35187_inst ( .DIN1(_35142), .DIN2(_35375), .Q(_35374) );
  xor2s1 _35188_inst ( .DIN1(_35141), .DIN2(_53115), .Q(_35375) );
  nnd2s1 _35189_inst ( .DIN1(_35376), .DIN2(_35377), .Q(_35141) );
  nnd2s1 _35190_inst ( .DIN1(_35378), .DIN2(_26535), .Q(_35377) );
  or2s1 _35191_inst ( .DIN1(_35379), .DIN2(_35205), .Q(_35378) );
  nnd2s1 _35192_inst ( .DIN1(_35205), .DIN2(_35379), .Q(_35376) );
  xnr2s1 _35193_inst ( .DIN1(_35190), .DIN2(_35380), .Q(_35142) );
  xor2s1 _35194_inst ( .DIN1(_53365), .DIN2(_35381), .Q(_35380) );
  nnd2s1 _35195_inst ( .DIN1(_35382), .DIN2(_35383), .Q(_35190) );
  nnd2s1 _35196_inst ( .DIN1(_26781), .DIN2(_35384), .Q(_35383) );
  or2s1 _35197_inst ( .DIN1(_35385), .DIN2(_35386), .Q(_35384) );
  nnd2s1 _35198_inst ( .DIN1(_35386), .DIN2(_35385), .Q(_35382) );
  nor2s1 _35199_inst ( .DIN1(_35387), .DIN2(_35388), .Q(_35371) );
  nor2s1 _35200_inst ( .DIN1(_35389), .DIN2(_35390), .Q(_35388) );
  nnd2s1 _35201_inst ( .DIN1(______[28]), .DIN2(_35391), .Q(_35390) );
  nnd2s1 _35202_inst ( .DIN1(_34306), .DIN2(_27596), .Q(_35391) );
  xor2s1 _35203_inst ( .DIN1(_53026), .DIN2(_53114), .Q(_35389) );
  nnd2s1 _35204_inst ( .DIN1(_35392), .DIN2(_35393), .Q(
        _____________________________239________) );
  nnd2s1 _35205_inst ( .DIN1(_35394), .DIN2(_35395), .Q(_35393) );
  nnd2s1 _35206_inst ( .DIN1(_35396), .DIN2(_35282), .Q(_35395) );
  nnd2s1 _35207_inst ( .DIN1(_35397), .DIN2(_35398), .Q(_35282) );
  nor2s1 _35208_inst ( .DIN1(_35295), .DIN2(_28598), .Q(_35397) );
  nor2s1 _35209_inst ( .DIN1(_35399), .DIN2(_35400), .Q(_35396) );
  nor2s1 _35210_inst ( .DIN1(_35285), .DIN2(_35401), .Q(_35400) );
  xor2s1 _35211_inst ( .DIN1(_35355), .DIN2(_35402), .Q(_35401) );
  xor2s1 _35212_inst ( .DIN1(_53152), .DIN2(_35356), .Q(_35402) );
  xor2s1 _35213_inst ( .DIN1(_35403), .DIN2(_29231), .Q(_35355) );
  nnd2s1 _35214_inst ( .DIN1(_35404), .DIN2(_35405), .Q(_35403) );
  nnd2s1 _35215_inst ( .DIN1(_35406), .DIN2(_26684), .Q(_35405) );
  nnd2s1 _35216_inst ( .DIN1(_35407), .DIN2(_35408), .Q(_35406) );
  or2s1 _35217_inst ( .DIN1(_35408), .DIN2(_35407), .Q(_35404) );
  nor2s1 _35218_inst ( .DIN1(_35295), .DIN2(_35409), .Q(_35399) );
  nor2s1 _35219_inst ( .DIN1(_35410), .DIN2(_27448), .Q(_35409) );
  xor2s1 _35220_inst ( .DIN1(_26373), .DIN2(_35411), .Q(_35410) );
  nor2s1 _35221_inst ( .DIN1(_53129), .DIN2(_26452), .Q(_35411) );
  hi1s1 _35222_inst ( .DIN(_35285), .Q(_35295) );
  nor2s1 _35223_inst ( .DIN1(_35412), .DIN2(_35413), .Q(_35392) );
  and2s1 _35224_inst ( .DIN1(_35414), .DIN2(_35415), .Q(_35413) );
  nor2s1 _35225_inst ( .DIN1(_35414), .DIN2(_35416), .Q(_35412) );
  nnd2s1 _35226_inst ( .DIN1(_28350), .DIN2(_26574), .Q(_35416) );
  xnr2s1 _35227_inst ( .DIN1(_35417), .DIN2(_53116), .Q(_35414) );
  nnd2s1 _35228_inst ( .DIN1(_53130), .DIN2(_53117), .Q(_35417) );
  nor2s1 _35229_inst ( .DIN1(_35418), .DIN2(_27500), .Q(
        _____________________________238________) );
  nor2s1 _35230_inst ( .DIN1(_35419), .DIN2(_35420), .Q(_35418) );
  nor2s1 _35231_inst ( .DIN1(_35285), .DIN2(_35421), .Q(_35420) );
  xor2s1 _35232_inst ( .DIN1(_35407), .DIN2(_35422), .Q(_35421) );
  xor2s1 _35233_inst ( .DIN1(_26684), .DIN2(_35408), .Q(_35422) );
  nnd2s1 _35234_inst ( .DIN1(_35423), .DIN2(_35424), .Q(_35408) );
  nnd2s1 _35235_inst ( .DIN1(_35425), .DIN2(_26627), .Q(_35424) );
  or2s1 _35236_inst ( .DIN1(_35426), .DIN2(_35427), .Q(_35425) );
  nnd2s1 _35237_inst ( .DIN1(_35427), .DIN2(_35426), .Q(_35423) );
  nor2s1 _35238_inst ( .DIN1(_35331), .DIN2(_35428), .Q(_35419) );
  nnd2s1 _35239_inst ( .DIN1(______[2]), .DIN2(_35429), .Q(_35428) );
  xor2s1 _35240_inst ( .DIN1(_53117), .DIN2(_53129), .Q(_35429) );
  nnd2s1 _35241_inst ( .DIN1(_35285), .DIN2(_35430), .Q(_35331) );
  nnd2s1 _35242_inst ( .DIN1(_35398), .DIN2(_28442), .Q(_35430) );
  nnd2s1 _35243_inst ( .DIN1(_35431), .DIN2(_35432), .Q(_35285) );
  nor2s1 _35244_inst ( .DIN1(_35433), .DIN2(_28603), .Q(_35431) );
  nnd2s1 _35245_inst ( .DIN1(_35434), .DIN2(_35435), .Q(
        _____________________________237________) );
  nnd2s1 _35246_inst ( .DIN1(_35436), .DIN2(_35437), .Q(_35435) );
  xor2s1 _35247_inst ( .DIN1(_35427), .DIN2(_35438), .Q(_35436) );
  xor2s1 _35248_inst ( .DIN1(_26627), .DIN2(_35426), .Q(_35438) );
  nnd2s1 _35249_inst ( .DIN1(_35439), .DIN2(_35440), .Q(_35426) );
  nnd2s1 _35250_inst ( .DIN1(_53157), .DIN2(_35441), .Q(_35440) );
  or2s1 _35251_inst ( .DIN1(_35442), .DIN2(_35443), .Q(_35441) );
  nnd2s1 _35252_inst ( .DIN1(_35443), .DIN2(_35442), .Q(_35439) );
  nor2s1 _35253_inst ( .DIN1(_35444), .DIN2(_35445), .Q(_35434) );
  nor2s1 _35254_inst ( .DIN1(_28629), .DIN2(_35446), .Q(_35445) );
  nnd2s1 _35255_inst ( .DIN1(_53118), .DIN2(_35447), .Q(_35446) );
  nor2s1 _35256_inst ( .DIN1(_35394), .DIN2(_35448), .Q(_35444) );
  nor2s1 _35257_inst ( .DIN1(_26694), .DIN2(_35449), .Q(_35448) );
  nnd2s1 _35258_inst ( .DIN1(______[10]), .DIN2(_28350), .Q(_35449) );
  nnd2s1 _35259_inst ( .DIN1(_35450), .DIN2(_35451), .Q(
        _____________________________236________) );
  nnd2s1 _35260_inst ( .DIN1(_35437), .DIN2(_35452), .Q(_35451) );
  xor2s1 _35261_inst ( .DIN1(_35453), .DIN2(_35454), .Q(_35452) );
  xnr2s1 _35262_inst ( .DIN1(_53157), .DIN2(_35442), .Q(_35454) );
  nnd2s1 _35263_inst ( .DIN1(_35455), .DIN2(_35456), .Q(_35442) );
  nnd2s1 _35264_inst ( .DIN1(_35457), .DIN2(_26469), .Q(_35456) );
  or2s1 _35265_inst ( .DIN1(_35458), .DIN2(_35459), .Q(_35457) );
  nnd2s1 _35266_inst ( .DIN1(_35459), .DIN2(_35458), .Q(_35455) );
  hi1s1 _35267_inst ( .DIN(_35443), .Q(_35453) );
  nor2s1 _35268_inst ( .DIN1(_35460), .DIN2(_28629), .Q(_35437) );
  nor2s1 _35269_inst ( .DIN1(_35415), .DIN2(_35461), .Q(_35450) );
  nor2s1 _35270_inst ( .DIN1(_35462), .DIN2(_35463), .Q(_35461) );
  nnd2s1 _35271_inst ( .DIN1(_35464), .DIN2(_35394), .Q(_35463) );
  xor2s1 _35272_inst ( .DIN1(_26452), .DIN2(_53129), .Q(_35464) );
  nnd2s1 _35273_inst ( .DIN1(______[22]), .DIN2(_35447), .Q(_35462) );
  nor2s1 _35274_inst ( .DIN1(_26574), .DIN2(_35465), .Q(_35415) );
  nnd2s1 _35275_inst ( .DIN1(_35466), .DIN2(_35467), .Q(
        _____________________________235________) );
  nnd2s1 _35276_inst ( .DIN1(_35468), .DIN2(_34707), .Q(_35467) );
  nnd2s1 _35277_inst ( .DIN1(_35469), .DIN2(______[30]), .Q(_35468) );
  nor2s1 _35278_inst ( .DIN1(_27123), .DIN2(_35470), .Q(_35469) );
  xor2s1 _35279_inst ( .DIN1(_35471), .DIN2(_53119), .Q(_35470) );
  nnd2s1 _35280_inst ( .DIN1(_53120), .DIN2(_53121), .Q(_35471) );
  nnd2s1 _35281_inst ( .DIN1(_35472), .DIN2(_29096), .Q(_35466) );
  nor2s1 _35282_inst ( .DIN1(_35473), .DIN2(_35474), .Q(_35472) );
  nor2s1 _35283_inst ( .DIN1(_35475), .DIN2(_35476), .Q(_35474) );
  nnd2s1 _35284_inst ( .DIN1(_35477), .DIN2(_35447), .Q(_35476) );
  nnd2s1 _35285_inst ( .DIN1(_35478), .DIN2(_26230), .Q(_35477) );
  nnd2s1 _35286_inst ( .DIN1(_53430), .DIN2(_35479), .Q(_35478) );
  and2s1 _35287_inst ( .DIN1(_35479), .DIN2(_35480), .Q(_35475) );
  nor2s1 _35288_inst ( .DIN1(_35481), .DIN2(_35460), .Q(_35473) );
  xor2s1 _35289_inst ( .DIN1(_35482), .DIN2(_35483), .Q(_35481) );
  xor2s1 _35290_inst ( .DIN1(_26469), .DIN2(_35458), .Q(_35483) );
  nnd2s1 _35291_inst ( .DIN1(_35484), .DIN2(_35485), .Q(_35458) );
  nnd2s1 _35292_inst ( .DIN1(_53164), .DIN2(_35486), .Q(_35485) );
  or2s1 _35293_inst ( .DIN1(_35487), .DIN2(_35488), .Q(_35486) );
  xor2s1 _35294_inst ( .DIN1(_34235), .DIN2(_35489), .Q(_35484) );
  nnd2s1 _35295_inst ( .DIN1(_35488), .DIN2(_35487), .Q(_35489) );
  nnd2s1 _35296_inst ( .DIN1(_35490), .DIN2(_35491), .Q(
        _____________________________234________) );
  nnd2s1 _35297_inst ( .DIN1(_35492), .DIN2(_27895), .Q(_35491) );
  nor2s1 _35298_inst ( .DIN1(_35493), .DIN2(_35494), .Q(_35492) );
  nor2s1 _35299_inst ( .DIN1(_35460), .DIN2(_35495), .Q(_35494) );
  xor2s1 _35300_inst ( .DIN1(_35488), .DIN2(_35496), .Q(_35495) );
  xor2s1 _35301_inst ( .DIN1(_26390), .DIN2(_35487), .Q(_35496) );
  nnd2s1 _35302_inst ( .DIN1(_35497), .DIN2(_35498), .Q(_35487) );
  nnd2s1 _35303_inst ( .DIN1(_53154), .DIN2(_35499), .Q(_35498) );
  or2s1 _35304_inst ( .DIN1(_35500), .DIN2(_32840), .Q(_35499) );
  nnd2s1 _35305_inst ( .DIN1(_32840), .DIN2(_35500), .Q(_35497) );
  nor2s1 _35306_inst ( .DIN1(_35398), .DIN2(_26720), .Q(_35493) );
  nnd2s1 _35307_inst ( .DIN1(_27894), .DIN2(_53453), .Q(_35490) );
  hi1s1 _35308_inst ( .DIN(_33589), .Q(_27894) );
  nnd2s1 _35309_inst ( .DIN1(_35501), .DIN2(_35502), .Q(_33589) );
  nnd2s1 _35310_inst ( .DIN1(_35503), .DIN2(_35504), .Q(
        _____________________________233________) );
  nnd2s1 _35311_inst ( .DIN1(_35505), .DIN2(_35506), .Q(_35504) );
  xor2s1 _35312_inst ( .DIN1(_53122), .DIN2(_26365), .Q(_35506) );
  nor2s1 _35313_inst ( .DIN1(_27551), .DIN2(_27614), .Q(_35505) );
  hi1s1 _35314_inst ( .DIN(_27177), .Q(_27551) );
  nnd2s1 _35315_inst ( .DIN1(_35507), .DIN2(_34214), .Q(_27177) );
  nnd2s1 _35316_inst ( .DIN1(_35508), .DIN2(_27164), .Q(_35503) );
  hi1s1 _35317_inst ( .DIN(_27546), .Q(_27164) );
  nnd2s1 _35318_inst ( .DIN1(_35509), .DIN2(_28253), .Q(_27546) );
  nor2s1 _35319_inst ( .DIN1(_35510), .DIN2(_35511), .Q(_35509) );
  nor2s1 _35320_inst ( .DIN1(_35512), .DIN2(_35513), .Q(_35508) );
  nor2s1 _35321_inst ( .DIN1(_35460), .DIN2(_35514), .Q(_35513) );
  xor2s1 _35322_inst ( .DIN1(_32840), .DIN2(_35515), .Q(_35514) );
  xor2s1 _35323_inst ( .DIN1(_26463), .DIN2(_35500), .Q(_35515) );
  nnd2s1 _35324_inst ( .DIN1(_35516), .DIN2(_35517), .Q(_35500) );
  nnd2s1 _35325_inst ( .DIN1(_35518), .DIN2(_26252), .Q(_35517) );
  or2s1 _35326_inst ( .DIN1(_35519), .DIN2(_35520), .Q(_35518) );
  nnd2s1 _35327_inst ( .DIN1(_35520), .DIN2(_35519), .Q(_35516) );
  nor2s1 _35328_inst ( .DIN1(_26453), .DIN2(_35521), .Q(_35512) );
  nnd2s1 _35329_inst ( .DIN1(______[20]), .DIN2(_35447), .Q(_35521) );
  nnd2s1 _35330_inst ( .DIN1(_35522), .DIN2(_28445), .Q(
        _____________________________232________) );
  nor2s1 _35331_inst ( .DIN1(_35523), .DIN2(_35524), .Q(_35522) );
  nor2s1 _35332_inst ( .DIN1(_27845), .DIN2(_35525), .Q(_35524) );
  nnd2s1 _35333_inst ( .DIN1(_35526), .DIN2(_35527), .Q(_35525) );
  nnd2s1 _35334_inst ( .DIN1(_35528), .DIN2(_35529), .Q(_35527) );
  hi1s1 _35335_inst ( .DIN(_35460), .Q(_35529) );
  nnd2s1 _35336_inst ( .DIN1(_35530), .DIN2(_35531), .Q(_35460) );
  nor2s1 _35337_inst ( .DIN1(_35433), .DIN2(_35532), .Q(_35531) );
  nnd2s1 _35338_inst ( .DIN1(_35533), .DIN2(_35534), .Q(_35532) );
  nor2s1 _35339_inst ( .DIN1(_28597), .DIN2(_28233), .Q(_35530) );
  nnd2s1 _35340_inst ( .DIN1(_35535), .DIN2(_28321), .Q(_28233) );
  nor2s1 _35341_inst ( .DIN1(_28599), .DIN2(_28603), .Q(_35535) );
  xor2s1 _35342_inst ( .DIN1(_35520), .DIN2(_35536), .Q(_35528) );
  xor2s1 _35343_inst ( .DIN1(_26252), .DIN2(_35519), .Q(_35536) );
  nnd2s1 _35344_inst ( .DIN1(_35537), .DIN2(_35538), .Q(_35519) );
  nnd2s1 _35345_inst ( .DIN1(_35539), .DIN2(_26501), .Q(_35538) );
  or2s1 _35346_inst ( .DIN1(_35540), .DIN2(_33253), .Q(_35539) );
  nnd2s1 _35347_inst ( .DIN1(_33253), .DIN2(_35540), .Q(_35537) );
  nnd2s1 _35348_inst ( .DIN1(_35541), .DIN2(_35542), .Q(_35526) );
  or2s1 _35349_inst ( .DIN1(_35479), .DIN2(_26230), .Q(_35542) );
  nnd2s1 _35350_inst ( .DIN1(_53124), .DIN2(_53430), .Q(_35479) );
  nor2s1 _35351_inst ( .DIN1(_35398), .DIN2(_35543), .Q(_35541) );
  nor2s1 _35352_inst ( .DIN1(_53124), .DIN2(_35480), .Q(_35543) );
  nor2s1 _35353_inst ( .DIN1(_26453), .DIN2(_26230), .Q(_35480) );
  nor2s1 _35354_inst ( .DIN1(_27836), .DIN2(_35544), .Q(_35523) );
  xor2s1 _35355_inst ( .DIN1(_35545), .DIN2(_35546), .Q(_35544) );
  xor2s1 _35356_inst ( .DIN1(_53125), .DIN2(_53316), .Q(_35546) );
  nor2s1 _35357_inst ( .DIN1(_26607), .DIN2(_26220), .Q(_35545) );
  nnd2s1 _35358_inst ( .DIN1(_35547), .DIN2(_35548), .Q(
        _____________________________231________) );
  nnd2s1 _35359_inst ( .DIN1(_29096), .DIN2(_35549), .Q(_35548) );
  nnd2s1 _35360_inst ( .DIN1(_35550), .DIN2(_35551), .Q(_35549) );
  nnd2s1 _35361_inst ( .DIN1(_35552), .DIN2(_35553), .Q(_35551) );
  xor2s1 _35362_inst ( .DIN1(_35554), .DIN2(_35555), .Q(_35553) );
  xnr2s1 _35363_inst ( .DIN1(_35540), .DIN2(_33253), .Q(_35555) );
  nnd2s1 _35364_inst ( .DIN1(_35556), .DIN2(_35557), .Q(_35540) );
  nnd2s1 _35365_inst ( .DIN1(_35558), .DIN2(_26625), .Q(_35557) );
  nnd2s1 _35366_inst ( .DIN1(_35559), .DIN2(_35560), .Q(_35558) );
  hi1s1 _35367_inst ( .DIN(_33461), .Q(_35560) );
  nnd2s1 _35368_inst ( .DIN1(_33461), .DIN2(_35561), .Q(_35556) );
  xor2s1 _35369_inst ( .DIN1(_26501), .DIN2(_31459), .Q(_35554) );
  nnd2s1 _35370_inst ( .DIN1(_35562), .DIN2(_35563), .Q(_35550) );
  nor2s1 _35371_inst ( .DIN1(_35564), .DIN2(_35565), .Q(_35563) );
  nor2s1 _35372_inst ( .DIN1(_53088), .DIN2(_35566), .Q(_35565) );
  nor2s1 _35373_inst ( .DIN1(_53431), .DIN2(_53307), .Q(_35566) );
  nor2s1 _35374_inst ( .DIN1(_35567), .DIN2(_26773), .Q(_35562) );
  and2s1 _35375_inst ( .DIN1(_26427), .DIN2(_35568), .Q(_35567) );
  nnd2s1 _35376_inst ( .DIN1(_29094), .DIN2(_35569), .Q(_35547) );
  xor2s1 _35377_inst ( .DIN1(_53121), .DIN2(_53126), .Q(_35569) );
  nnd2s1 _35378_inst ( .DIN1(_35570), .DIN2(_27970), .Q(
        _____________________________230________) );
  nor2s1 _35379_inst ( .DIN1(_35571), .DIN2(_35572), .Q(_35570) );
  nor2s1 _35380_inst ( .DIN1(_27973), .DIN2(_35573), .Q(_35572) );
  nnd2s1 _35381_inst ( .DIN1(_35574), .DIN2(_35575), .Q(_35573) );
  nor2s1 _35382_inst ( .DIN1(_35576), .DIN2(_35577), .Q(_35574) );
  nor2s1 _35383_inst ( .DIN1(_35578), .DIN2(_35579), .Q(_35577) );
  xor2s1 _35384_inst ( .DIN1(_35580), .DIN2(_35581), .Q(_35579) );
  xor2s1 _35385_inst ( .DIN1(_33461), .DIN2(_35559), .Q(_35581) );
  hi1s1 _35386_inst ( .DIN(_35561), .Q(_35559) );
  nnd2s1 _35387_inst ( .DIN1(_35582), .DIN2(_35583), .Q(_35561) );
  nnd2s1 _35388_inst ( .DIN1(_35584), .DIN2(_26483), .Q(_35583) );
  or2s1 _35389_inst ( .DIN1(_35585), .DIN2(_33675), .Q(_35584) );
  nnd2s1 _35390_inst ( .DIN1(_33675), .DIN2(_35585), .Q(_35582) );
  xor2s1 _35391_inst ( .DIN1(_31222), .DIN2(_53168), .Q(_35580) );
  nor2s1 _35392_inst ( .DIN1(_53119), .DIN2(_35552), .Q(_35576) );
  nor2s1 _35393_inst ( .DIN1(_27915), .DIN2(_35586), .Q(_35571) );
  xnr2s1 _35394_inst ( .DIN1(_53506), .DIN2(_35587), .Q(_35586) );
  nor2s1 _35395_inst ( .DIN1(_53455), .DIN2(_26579), .Q(_35587) );
  nnd2s1 _35396_inst ( .DIN1(_35588), .DIN2(_35589), .Q(
        _____________________________22________) );
  nor2s1 _35397_inst ( .DIN1(_35133), .DIN2(_35590), .Q(_35589) );
  nor2s1 _35398_inst ( .DIN1(_35136), .DIN2(_35591), .Q(_35590) );
  xor2s1 _35399_inst ( .DIN1(_35205), .DIN2(_35592), .Q(_35591) );
  xor2s1 _35400_inst ( .DIN1(_26535), .DIN2(_35379), .Q(_35592) );
  nnd2s1 _35401_inst ( .DIN1(_35593), .DIN2(_35594), .Q(_35379) );
  nnd2s1 _35402_inst ( .DIN1(_53142), .DIN2(_35595), .Q(_35594) );
  or2s1 _35403_inst ( .DIN1(_35596), .DIN2(_35226), .Q(_35595) );
  nnd2s1 _35404_inst ( .DIN1(_35226), .DIN2(_35596), .Q(_35593) );
  xnr2s1 _35405_inst ( .DIN1(_35597), .DIN2(_35598), .Q(_35205) );
  xor2s1 _35406_inst ( .DIN1(_35385), .DIN2(_53368), .Q(_35597) );
  nnd2s1 _35407_inst ( .DIN1(_35599), .DIN2(_35600), .Q(_35385) );
  nnd2s1 _35408_inst ( .DIN1(_53367), .DIN2(_35601), .Q(_35600) );
  or2s1 _35409_inst ( .DIN1(_35602), .DIN2(_35603), .Q(_35601) );
  nnd2s1 _35410_inst ( .DIN1(_35603), .DIN2(_35602), .Q(_35599) );
  nor2s1 _35411_inst ( .DIN1(_35604), .DIN2(_35605), .Q(_35588) );
  nor2s1 _35412_inst ( .DIN1(_35606), .DIN2(_35147), .Q(_35605) );
  nor2s1 _35413_inst ( .DIN1(_27082), .DIN2(_35607), .Q(_35606) );
  nnd2s1 _35414_inst ( .DIN1(_35608), .DIN2(_35609), .Q(_35607) );
  nnd2s1 _35415_inst ( .DIN1(_26244), .DIN2(_26404), .Q(_35608) );
  nor2s1 _35416_inst ( .DIN1(_34300), .DIN2(_35610), .Q(_35604) );
  xnr2s1 _35417_inst ( .DIN1(_35611), .DIN2(_35609), .Q(_35610) );
  nnd2s1 _35418_inst ( .DIN1(_53194), .DIN2(_53196), .Q(_35609) );
  nnd2s1 _35419_inst ( .DIN1(_35612), .DIN2(_35613), .Q(_35611) );
  nnd2s1 _35420_inst ( .DIN1(_26244), .DIN2(_26379), .Q(_35613) );
  hi1s1 _35421_inst ( .DIN(_35614), .Q(_34300) );
  nnd2s1 _35422_inst ( .DIN1(_35615), .DIN2(_27126), .Q(
        _____________________________229________) );
  nnd2s1 _35423_inst ( .DIN1(_35616), .DIN2(_34826), .Q(_27126) );
  nor2s1 _35424_inst ( .DIN1(_27129), .DIN2(_35617), .Q(_35616) );
  nor2s1 _35425_inst ( .DIN1(_35618), .DIN2(_35619), .Q(_35615) );
  nor2s1 _35426_inst ( .DIN1(_27132), .DIN2(_35620), .Q(_35619) );
  nnd2s1 _35427_inst ( .DIN1(_35621), .DIN2(_35575), .Q(_35620) );
  xor2s1 _35428_inst ( .DIN1(_31307), .DIN2(_35622), .Q(_35621) );
  nnd2s1 _35429_inst ( .DIN1(_35623), .DIN2(_35624), .Q(_35622) );
  nnd2s1 _35430_inst ( .DIN1(_35625), .DIN2(_35578), .Q(_35624) );
  nor2s1 _35431_inst ( .DIN1(_53431), .DIN2(_27448), .Q(_35625) );
  nnd2s1 _35432_inst ( .DIN1(_35626), .DIN2(_35552), .Q(_35623) );
  xor2s1 _35433_inst ( .DIN1(_33675), .DIN2(_35627), .Q(_35626) );
  xor2s1 _35434_inst ( .DIN1(_26483), .DIN2(_35585), .Q(_35627) );
  nnd2s1 _35435_inst ( .DIN1(_35628), .DIN2(_35629), .Q(_35585) );
  nnd2s1 _35436_inst ( .DIN1(_53391), .DIN2(_35630), .Q(_35629) );
  or2s1 _35437_inst ( .DIN1(_35631), .DIN2(_33872), .Q(_35630) );
  nnd2s1 _35438_inst ( .DIN1(_33872), .DIN2(_35631), .Q(_35628) );
  nor2s1 _35439_inst ( .DIN1(_27129), .DIN2(_35632), .Q(_35618) );
  nor2s1 _35440_inst ( .DIN1(_28100), .DIN2(_35633), .Q(_35632) );
  xor2s1 _35441_inst ( .DIN1(_53248), .DIN2(_29787), .Q(_35633) );
  hi1s1 _35442_inst ( .DIN(_27132), .Q(_27129) );
  nnd2s1 _35443_inst ( .DIN1(_35634), .DIN2(_30228), .Q(
        _____________________________228________) );
  nor2s1 _35444_inst ( .DIN1(_35635), .DIN2(_35636), .Q(_35634) );
  nor2s1 _35445_inst ( .DIN1(_29555), .DIN2(_35637), .Q(_35636) );
  nnd2s1 _35446_inst ( .DIN1(_35638), .DIN2(_35575), .Q(_35637) );
  nor2s1 _35447_inst ( .DIN1(_35639), .DIN2(_35640), .Q(_35638) );
  nor2s1 _35448_inst ( .DIN1(_35578), .DIN2(_35641), .Q(_35640) );
  xnr2s1 _35449_inst ( .DIN1(_33872), .DIN2(_35642), .Q(_35641) );
  xor2s1 _35450_inst ( .DIN1(_26386), .DIN2(_35631), .Q(_35642) );
  nnd2s1 _35451_inst ( .DIN1(_35643), .DIN2(_35644), .Q(_35631) );
  nnd2s1 _35452_inst ( .DIN1(_53356), .DIN2(_35645), .Q(_35644) );
  or2s1 _35453_inst ( .DIN1(_35646), .DIN2(_34084), .Q(_35645) );
  nnd2s1 _35454_inst ( .DIN1(_34084), .DIN2(_35646), .Q(_35643) );
  nor2s1 _35455_inst ( .DIN1(_35552), .DIN2(_35647), .Q(_35639) );
  nor2s1 _35456_inst ( .DIN1(_35648), .DIN2(_26773), .Q(_35647) );
  xor2s1 _35457_inst ( .DIN1(_26427), .DIN2(_35568), .Q(_35648) );
  nor2s1 _35458_inst ( .DIN1(_26424), .DIN2(_53431), .Q(_35568) );
  nor2s1 _35459_inst ( .DIN1(_29560), .DIN2(_35649), .Q(_35635) );
  nor2s1 _35460_inst ( .DIN1(_35650), .DIN2(_26987), .Q(_35649) );
  xor2s1 _35461_inst ( .DIN1(_35651), .DIN2(_35652), .Q(_35650) );
  nor2s1 _35462_inst ( .DIN1(_26519), .DIN2(_26292), .Q(_35652) );
  nnd2s1 _35463_inst ( .DIN1(_29558), .DIN2(_35653), .Q(_35651) );
  nnd2s1 _35464_inst ( .DIN1(_53128), .DIN2(_26519), .Q(_35653) );
  nnd2s1 _35465_inst ( .DIN1(_53347), .DIN2(_26561), .Q(_29558) );
  nnd2s1 _35466_inst ( .DIN1(_35654), .DIN2(_35655), .Q(
        _____________________________227________) );
  nnd2s1 _35467_inst ( .DIN1(_35656), .DIN2(______[4]), .Q(_35655) );
  nor2s1 _35468_inst ( .DIN1(_35465), .DIN2(_35657), .Q(_35656) );
  xor2s1 _35469_inst ( .DIN1(_26373), .DIN2(_53129), .Q(_35657) );
  nnd2s1 _35470_inst ( .DIN1(_35394), .DIN2(_35658), .Q(_35654) );
  xor2s1 _35471_inst ( .DIN1(_29994), .DIN2(_35659), .Q(_35658) );
  nnd2s1 _35472_inst ( .DIN1(_35660), .DIN2(_35575), .Q(_35659) );
  nnd2s1 _35473_inst ( .DIN1(_35564), .DIN2(_35578), .Q(_35575) );
  hi1s1 _35474_inst ( .DIN(_35661), .Q(_35564) );
  nor2s1 _35475_inst ( .DIN1(_35662), .DIN2(_35663), .Q(_35660) );
  nor2s1 _35476_inst ( .DIN1(_35578), .DIN2(_35664), .Q(_35663) );
  xor2s1 _35477_inst ( .DIN1(_35665), .DIN2(_35666), .Q(_35664) );
  xnr2s1 _35478_inst ( .DIN1(_53356), .DIN2(_35646), .Q(_35666) );
  nnd2s1 _35479_inst ( .DIN1(_35667), .DIN2(_35668), .Q(_35646) );
  xor2s1 _35480_inst ( .DIN1(_33328), .DIN2(_35669), .Q(_35667) );
  nnd2s1 _35481_inst ( .DIN1(_35670), .DIN2(_35671), .Q(_35669) );
  nor2s1 _35482_inst ( .DIN1(_35552), .DIN2(_35672), .Q(_35662) );
  xor2s1 _35483_inst ( .DIN1(_35673), .DIN2(_35674), .Q(_35672) );
  xor2s1 _35484_inst ( .DIN1(_53133), .DIN2(_53135), .Q(_35674) );
  nnd2s1 _35485_inst ( .DIN1(_53116), .DIN2(_53092), .Q(_35673) );
  nnd2s1 _35486_inst ( .DIN1(_35675), .DIN2(_35676), .Q(
        _____________________________226________) );
  nnd2s1 _35487_inst ( .DIN1(_27684), .DIN2(_35677), .Q(_35676) );
  nnd2s1 _35488_inst ( .DIN1(_35678), .DIN2(_35679), .Q(_35677) );
  nnd2s1 _35489_inst ( .DIN1(_35552), .DIN2(_35680), .Q(_35679) );
  xnr2s1 _35490_inst ( .DIN1(_35670), .DIN2(_35681), .Q(_35680) );
  nnd2s1 _35491_inst ( .DIN1(_35671), .DIN2(_35668), .Q(_35681) );
  nnd2s1 _35492_inst ( .DIN1(_53170), .DIN2(_34287), .Q(_35668) );
  or2s1 _35493_inst ( .DIN1(_34287), .DIN2(_53170), .Q(_35671) );
  hi1s1 _35494_inst ( .DIN(_35578), .Q(_35552) );
  nnd2s1 _35495_inst ( .DIN1(_35682), .DIN2(_28441), .Q(_35578) );
  hi1s1 _35496_inst ( .DIN(_28528), .Q(_28441) );
  nnd2s1 _35497_inst ( .DIN1(_35683), .DIN2(_35684), .Q(_28528) );
  nor2s1 _35498_inst ( .DIN1(_35433), .DIN2(_28597), .Q(_35683) );
  nor2s1 _35499_inst ( .DIN1(_28596), .DIN2(_35685), .Q(_35682) );
  nnd2s1 _35500_inst ( .DIN1(_53116), .DIN2(_35661), .Q(_35678) );
  nnd2s1 _35501_inst ( .DIN1(_35398), .DIN2(_35686), .Q(_35661) );
  hi1s1 _35502_inst ( .DIN(_35447), .Q(_35398) );
  nnd2s1 _35503_inst ( .DIN1(_35687), .DIN2(_35688), .Q(_35447) );
  nor2s1 _35504_inst ( .DIN1(_28599), .DIN2(_35433), .Q(_35687) );
  hi1s1 _35505_inst ( .DIN(_27679), .Q(_27684) );
  nnd2s1 _35506_inst ( .DIN1(_35689), .DIN2(_27679), .Q(_35675) );
  nnd2s1 _35507_inst ( .DIN1(_35690), .DIN2(_35691), .Q(_27679) );
  nor2s1 _35508_inst ( .DIN1(_35692), .DIN2(_35693), .Q(_35691) );
  nnd2s1 _35509_inst ( .DIN1(_35694), .DIN2(_35695), .Q(_35693) );
  nnd2s1 _35510_inst ( .DIN1(_35696), .DIN2(_33614), .Q(_35692) );
  nor2s1 _35511_inst ( .DIN1(_35697), .DIN2(_35698), .Q(_35690) );
  or2s1 _35512_inst ( .DIN1(_35699), .DIN2(_35700), .Q(_35698) );
  nor2s1 _35513_inst ( .DIN1(_27774), .DIN2(_35701), .Q(_35689) );
  nnd2s1 _35514_inst ( .DIN1(_35702), .DIN2(_35703), .Q(_35701) );
  hi1s1 _35515_inst ( .DIN(_33522), .Q(_35703) );
  nor2s1 _35516_inst ( .DIN1(_35704), .DIN2(_35697), .Q(_33522) );
  nnd2s1 _35517_inst ( .DIN1(_35705), .DIN2(_33606), .Q(_35697) );
  hi1s1 _35518_inst ( .DIN(_27934), .Q(_33606) );
  nor2s1 _35519_inst ( .DIN1(_35706), .DIN2(_33617), .Q(_35705) );
  nnd2s1 _35520_inst ( .DIN1(_35707), .DIN2(_35708), .Q(_35704) );
  xor2s1 _35521_inst ( .DIN1(_53131), .DIN2(_53132), .Q(_35702) );
  nnd2s1 _35522_inst ( .DIN1(_35709), .DIN2(_35710), .Q(
        _____________________________225________) );
  nnd2s1 _35523_inst ( .DIN1(_35711), .DIN2(_28289), .Q(_35710) );
  nnd2s1 _35524_inst ( .DIN1(_28442), .DIN2(_28292), .Q(_28289) );
  nnd2s1 _35525_inst ( .DIN1(_35712), .DIN2(_35713), .Q(_35711) );
  nnd2s1 _35526_inst ( .DIN1(_35714), .DIN2(_35715), .Q(_35713) );
  nor2s1 _35527_inst ( .DIN1(_35670), .DIN2(_35716), .Q(_35715) );
  nor2s1 _35528_inst ( .DIN1(_52835), .DIN2(_34288), .Q(_35716) );
  and2s1 _35529_inst ( .DIN1(_52835), .DIN2(_34288), .Q(_35670) );
  nor2s1 _35530_inst ( .DIN1(_28292), .DIN2(_28629), .Q(_35714) );
  nnd2s1 _35531_inst ( .DIN1(_28625), .DIN2(______[26]), .Q(_35712) );
  and2s1 _35532_inst ( .DIN1(_35717), .DIN2(_35394), .Q(_28625) );
  hi1s1 _35533_inst ( .DIN(_28629), .Q(_35394) );
  nor2s1 _35534_inst ( .DIN1(_28293), .DIN2(_26450), .Q(_35717) );
  hi1s1 _35535_inst ( .DIN(_28292), .Q(_28293) );
  nnd2s1 _35536_inst ( .DIN1(_35718), .DIN2(_35432), .Q(_28292) );
  nor2s1 _35537_inst ( .DIN1(_28595), .DIN2(_28597), .Q(_35718) );
  nnd2s1 _35538_inst ( .DIN1(_35719), .DIN2(_28629), .Q(_35709) );
  nnd2s1 _35539_inst ( .DIN1(_28589), .DIN2(_35720), .Q(_28629) );
  hi1s1 _35540_inst ( .DIN(_28347), .Q(_28589) );
  nnd2s1 _35541_inst ( .DIN1(_35071), .DIN2(_35721), .Q(_28347) );
  hi1s1 _35542_inst ( .DIN(_35277), .Q(_35071) );
  nnd2s1 _35543_inst ( .DIN1(_35722), .DIN2(_35723), .Q(_35277) );
  nor2s1 _35544_inst ( .DIN1(_35301), .DIN2(_35724), .Q(_35722) );
  nnd2s1 _35545_inst ( .DIN1(_35725), .DIN2(_35726), .Q(_35719) );
  xor2s1 _35546_inst ( .DIN1(_28351), .DIN2(_53134), .Q(_35726) );
  nnd2s1 _35547_inst ( .DIN1(_53135), .DIN2(_53511), .Q(_28351) );
  nor2s1 _35548_inst ( .DIN1(_35465), .DIN2(_27365), .Q(_35725) );
  nnd2s1 _35549_inst ( .DIN1(_35727), .DIN2(_35728), .Q(
        _____________________________224________) );
  nnd2s1 _35550_inst ( .DIN1(_35729), .DIN2(_52942), .Q(_35728) );
  nor2s1 _35551_inst ( .DIN1(_27774), .DIN2(_30068), .Q(_35729) );
  nnd2s1 _35552_inst ( .DIN1(_28329), .DIN2(_35730), .Q(_30068) );
  nnd2s1 _35553_inst ( .DIN1(_28338), .DIN2(_35731), .Q(_35727) );
  nnd2s1 _35554_inst ( .DIN1(_35732), .DIN2(_35733), .Q(_35731) );
  nnd2s1 _35555_inst ( .DIN1(_35734), .DIN2(_35735), .Q(_35733) );
  nnd2s1 _35556_inst ( .DIN1(_35736), .DIN2(_35737), .Q(_35734) );
  nnd2s1 _35557_inst ( .DIN1(_26276), .DIN2(_26712), .Q(_35737) );
  nor2s1 _35558_inst ( .DIN1(_28321), .DIN2(_28320), .Q(_35736) );
  nor2s1 _35559_inst ( .DIN1(_26276), .DIN2(_26712), .Q(_28320) );
  nor2s1 _35560_inst ( .DIN1(_35738), .DIN2(_35739), .Q(_35732) );
  nor2s1 _35561_inst ( .DIN1(_26524), .DIN2(_35740), .Q(_35739) );
  nor2s1 _35562_inst ( .DIN1(_35741), .DIN2(_35742), .Q(_35740) );
  nor2s1 _35563_inst ( .DIN1(_34345), .DIN2(_35743), .Q(_35742) );
  nor2s1 _35564_inst ( .DIN1(_35744), .DIN2(_34343), .Q(_35741) );
  nor2s1 _35565_inst ( .DIN1(_53136), .DIN2(_35745), .Q(_35738) );
  nor2s1 _35566_inst ( .DIN1(_35746), .DIN2(_35747), .Q(_35745) );
  nor2s1 _35567_inst ( .DIN1(_34343), .DIN2(_35743), .Q(_35747) );
  nnd2s1 _35568_inst ( .DIN1(_28317), .DIN2(_26849), .Q(_34343) );
  nor2s1 _35569_inst ( .DIN1(_35744), .DIN2(_34345), .Q(_35746) );
  nnd2s1 _35570_inst ( .DIN1(_28317), .DIN2(_26850), .Q(_34345) );
  hi1s1 _35571_inst ( .DIN(_35743), .Q(_35744) );
  nnd2s1 _35572_inst ( .DIN1(_35748), .DIN2(_35749), .Q(_35743) );
  nnd2s1 _35573_inst ( .DIN1(_35750), .DIN2(_26632), .Q(_35749) );
  or2s1 _35574_inst ( .DIN1(_35751), .DIN2(_26850), .Q(_35750) );
  nnd2s1 _35575_inst ( .DIN1(_35751), .DIN2(_26850), .Q(_35748) );
  nnd2s1 _35576_inst ( .DIN1(_35752), .DIN2(_28569), .Q(
        _____________________________223________) );
  or2s1 _35577_inst ( .DIN1(_34985), .DIN2(_28572), .Q(_28569) );
  nnd2s1 _35578_inst ( .DIN1(_35753), .DIN2(_35754), .Q(_34985) );
  nor2s1 _35579_inst ( .DIN1(_35755), .DIN2(_35756), .Q(_35754) );
  nnd2s1 _35580_inst ( .DIN1(_35757), .DIN2(_35758), .Q(_35756) );
  nor2s1 _35581_inst ( .DIN1(_35700), .DIN2(_33616), .Q(_35753) );
  nor2s1 _35582_inst ( .DIN1(_35759), .DIN2(_35760), .Q(_35752) );
  nor2s1 _35583_inst ( .DIN1(_28575), .DIN2(_35761), .Q(_35760) );
  nor2s1 _35584_inst ( .DIN1(_35762), .DIN2(_35763), .Q(_35761) );
  nor2s1 _35585_inst ( .DIN1(_35764), .DIN2(_35765), .Q(_35763) );
  xor2s1 _35586_inst ( .DIN1(_35751), .DIN2(_35766), .Q(_35765) );
  xor2s1 _35587_inst ( .DIN1(_26632), .DIN2(_53384), .Q(_35766) );
  nnd2s1 _35588_inst ( .DIN1(_35767), .DIN2(_35768), .Q(_35751) );
  nnd2s1 _35589_inst ( .DIN1(_35769), .DIN2(_26681), .Q(_35768) );
  nnd2s1 _35590_inst ( .DIN1(_32914), .DIN2(_35770), .Q(_35769) );
  or2s1 _35591_inst ( .DIN1(_35770), .DIN2(_32914), .Q(_35767) );
  nor2s1 _35592_inst ( .DIN1(_35771), .DIN2(_35772), .Q(_35762) );
  nor2s1 _35593_inst ( .DIN1(_27614), .DIN2(_35773), .Q(_35772) );
  nnd2s1 _35594_inst ( .DIN1(_35774), .DIN2(_35775), .Q(_35773) );
  xor2s1 _35595_inst ( .DIN1(_53222), .DIN2(_35776), .Q(_35774) );
  nor2s1 _35596_inst ( .DIN1(_53275), .DIN2(_28572), .Q(_35759) );
  hi1s1 _35597_inst ( .DIN(_28575), .Q(_28572) );
  nnd2s1 _35598_inst ( .DIN1(_35777), .DIN2(_35778), .Q(_28575) );
  nor2s1 _35599_inst ( .DIN1(_35779), .DIN2(_35780), .Q(_35778) );
  nnd2s1 _35600_inst ( .DIN1(_35757), .DIN2(_35781), .Q(_35780) );
  nnd2s1 _35601_inst ( .DIN1(_33614), .DIN2(_35758), .Q(_35779) );
  nor2s1 _35602_inst ( .DIN1(_35782), .DIN2(_35783), .Q(_35777) );
  nnd2s1 _35603_inst ( .DIN1(_34601), .DIN2(_35784), .Q(_35783) );
  nnd2s1 _35604_inst ( .DIN1(_35785), .DIN2(_33613), .Q(_35782) );
  nnd2s1 _35605_inst ( .DIN1(_35786), .DIN2(_28782), .Q(
        _____________________________222________) );
  nnd2s1 _35606_inst ( .DIN1(_34090), .DIN2(_28786), .Q(_28782) );
  nor2s1 _35607_inst ( .DIN1(_35787), .DIN2(_35788), .Q(_35786) );
  nor2s1 _35608_inst ( .DIN1(_28792), .DIN2(_35789), .Q(_35788) );
  xor2s1 _35609_inst ( .DIN1(_53139), .DIN2(_53504), .Q(_35789) );
  nor2s1 _35610_inst ( .DIN1(_35790), .DIN2(_28786), .Q(_35787) );
  nor2s1 _35611_inst ( .DIN1(_35791), .DIN2(_35792), .Q(_35790) );
  nnd2s1 _35612_inst ( .DIN1(_35793), .DIN2(_35794), .Q(_35792) );
  nnd2s1 _35613_inst ( .DIN1(_35795), .DIN2(_35796), .Q(_35794) );
  nnd2s1 _35614_inst ( .DIN1(_53224), .DIN2(______[28]), .Q(_35795) );
  nnd2s1 _35615_inst ( .DIN1(_35797), .DIN2(_35798), .Q(_35793) );
  xor2s1 _35616_inst ( .DIN1(_35770), .DIN2(_35799), .Q(_35798) );
  xor2s1 _35617_inst ( .DIN1(_26681), .DIN2(_32914), .Q(_35799) );
  nnd2s1 _35618_inst ( .DIN1(_35800), .DIN2(_35801), .Q(_35770) );
  nnd2s1 _35619_inst ( .DIN1(_53185), .DIN2(_35802), .Q(_35801) );
  or2s1 _35620_inst ( .DIN1(_35803), .DIN2(_32935), .Q(_35802) );
  nnd2s1 _35621_inst ( .DIN1(_32935), .DIN2(_35803), .Q(_35800) );
  nnd2s1 _35622_inst ( .DIN1(_35804), .DIN2(_27660), .Q(
        _____________________________221________) );
  nor2s1 _35623_inst ( .DIN1(_35805), .DIN2(_35806), .Q(_35804) );
  nor2s1 _35624_inst ( .DIN1(_27663), .DIN2(_35807), .Q(_35806) );
  nnd2s1 _35625_inst ( .DIN1(_35808), .DIN2(_35809), .Q(_35807) );
  nor2s1 _35626_inst ( .DIN1(_35810), .DIN2(_35811), .Q(_35808) );
  nor2s1 _35627_inst ( .DIN1(_35796), .DIN2(_35812), .Q(_35811) );
  xor2s1 _35628_inst ( .DIN1(_35813), .DIN2(_35814), .Q(_35812) );
  xor2s1 _35629_inst ( .DIN1(_35803), .DIN2(_32935), .Q(_35814) );
  nnd2s1 _35630_inst ( .DIN1(_35815), .DIN2(_35816), .Q(_35803) );
  nnd2s1 _35631_inst ( .DIN1(_53186), .DIN2(_35817), .Q(_35816) );
  or2s1 _35632_inst ( .DIN1(_35818), .DIN2(_32951), .Q(_35817) );
  nnd2s1 _35633_inst ( .DIN1(_32951), .DIN2(_35818), .Q(_35815) );
  xor2s1 _35634_inst ( .DIN1(_29518), .DIN2(_53185), .Q(_35813) );
  nor2s1 _35635_inst ( .DIN1(_35797), .DIN2(_35819), .Q(_35810) );
  xor2s1 _35636_inst ( .DIN1(_35820), .DIN2(_35821), .Q(_35819) );
  nnd2s1 _35637_inst ( .DIN1(_35822), .DIN2(______[22]), .Q(_35820) );
  nor2s1 _35638_inst ( .DIN1(_35776), .DIN2(_35823), .Q(_35822) );
  nor2s1 _35639_inst ( .DIN1(_53224), .DIN2(_53225), .Q(_35823) );
  hi1s1 _35640_inst ( .DIN(_35824), .Q(_35776) );
  nor2s1 _35641_inst ( .DIN1(_27672), .DIN2(_35825), .Q(_35805) );
  nor2s1 _35642_inst ( .DIN1(_26988), .DIN2(_35826), .Q(_35825) );
  xor2s1 _35643_inst ( .DIN1(_26636), .DIN2(_27815), .Q(_35826) );
  nnd2s1 _35644_inst ( .DIN1(_53155), .DIN2(_53157), .Q(_27815) );
  nnd2s1 _35645_inst ( .DIN1(_35827), .DIN2(_35828), .Q(
        _____________________________220________) );
  nnd2s1 _35646_inst ( .DIN1(_35829), .DIN2(_35830), .Q(_35828) );
  nnd2s1 _35647_inst ( .DIN1(_35831), .DIN2(_35809), .Q(_35830) );
  nor2s1 _35648_inst ( .DIN1(_35832), .DIN2(_35833), .Q(_35831) );
  nor2s1 _35649_inst ( .DIN1(_35834), .DIN2(_35796), .Q(_35833) );
  xor2s1 _35650_inst ( .DIN1(_32973), .DIN2(_35835), .Q(_35834) );
  xnr2s1 _35651_inst ( .DIN1(_53186), .DIN2(_35818), .Q(_35835) );
  nnd2s1 _35652_inst ( .DIN1(_35836), .DIN2(_35837), .Q(_35818) );
  nnd2s1 _35653_inst ( .DIN1(_53180), .DIN2(_35838), .Q(_35837) );
  or2s1 _35654_inst ( .DIN1(_35839), .DIN2(_32979), .Q(_35838) );
  xnr2s1 _35655_inst ( .DIN1(_32615), .DIN2(_35840), .Q(_35836) );
  nnd2s1 _35656_inst ( .DIN1(_32979), .DIN2(_35839), .Q(_35840) );
  nor2s1 _35657_inst ( .DIN1(_35797), .DIN2(_35841), .Q(_35832) );
  nor2s1 _35658_inst ( .DIN1(_27291), .DIN2(_35842), .Q(_35841) );
  xor2s1 _35659_inst ( .DIN1(_53219), .DIN2(_53428), .Q(_35842) );
  nnd2s1 _35660_inst ( .DIN1(_35843), .DIN2(_53218), .Q(_35827) );
  nnd2s1 _35661_inst ( .DIN1(_35844), .DIN2(_35341), .Q(
        _____________________________21________) );
  nor2s1 _35662_inst ( .DIN1(_35845), .DIN2(_35846), .Q(_35844) );
  nor2s1 _35663_inst ( .DIN1(_27749), .DIN2(_35847), .Q(_35846) );
  nor2s1 _35664_inst ( .DIN1(_35848), .DIN2(_35849), .Q(_35847) );
  nor2s1 _35665_inst ( .DIN1(_35373), .DIN2(_35850), .Q(_35849) );
  xor2s1 _35666_inst ( .DIN1(_35226), .DIN2(_35851), .Q(_35850) );
  xor2s1 _35667_inst ( .DIN1(_26397), .DIN2(_35596), .Q(_35851) );
  nnd2s1 _35668_inst ( .DIN1(_35852), .DIN2(_35853), .Q(_35596) );
  nnd2s1 _35669_inst ( .DIN1(_35854), .DIN2(_26638), .Q(_35853) );
  or2s1 _35670_inst ( .DIN1(_35855), .DIN2(_35239), .Q(_35854) );
  nnd2s1 _35671_inst ( .DIN1(_35239), .DIN2(_35855), .Q(_35852) );
  xnr2s1 _35672_inst ( .DIN1(_35856), .DIN2(_35603), .Q(_35226) );
  xor2s1 _35673_inst ( .DIN1(_26209), .DIN2(_35602), .Q(_35856) );
  nnd2s1 _35674_inst ( .DIN1(_35857), .DIN2(_35858), .Q(_35602) );
  nnd2s1 _35675_inst ( .DIN1(_53309), .DIN2(_35859), .Q(_35858) );
  or2s1 _35676_inst ( .DIN1(_35860), .DIN2(_35861), .Q(_35859) );
  nnd2s1 _35677_inst ( .DIN1(_35861), .DIN2(_35860), .Q(_35857) );
  nor2s1 _35678_inst ( .DIN1(_35387), .DIN2(_35862), .Q(_35848) );
  nnd2s1 _35679_inst ( .DIN1(_35863), .DIN2(_35864), .Q(_35862) );
  xor2s1 _35680_inst ( .DIN1(_26348), .DIN2(_35865), .Q(_35863) );
  nor2s1 _35681_inst ( .DIN1(_53196), .DIN2(_26362), .Q(_35865) );
  nor2s1 _35682_inst ( .DIN1(_28010), .DIN2(_35866), .Q(_35845) );
  nor2s1 _35683_inst ( .DIN1(_26772), .DIN2(_35867), .Q(_35866) );
  xor2s1 _35684_inst ( .DIN1(_53208), .DIN2(_35868), .Q(_35867) );
  nor2s1 _35685_inst ( .DIN1(_53405), .DIN2(_53399), .Q(_35868) );
  nnd2s1 _35686_inst ( .DIN1(_35869), .DIN2(_35870), .Q(
        _____________________________219________) );
  nnd2s1 _35687_inst ( .DIN1(_35871), .DIN2(_35872), .Q(_35870) );
  xor2s1 _35688_inst ( .DIN1(_26528), .DIN2(_53152), .Q(_35872) );
  nor2s1 _35689_inst ( .DIN1(_35873), .DIN2(_27082), .Q(_35871) );
  nnd2s1 _35690_inst ( .DIN1(_35874), .DIN2(_27512), .Q(_35869) );
  nor2s1 _35691_inst ( .DIN1(_35875), .DIN2(_35876), .Q(_35874) );
  nor2s1 _35692_inst ( .DIN1(_35796), .DIN2(_35877), .Q(_35876) );
  xor2s1 _35693_inst ( .DIN1(_32994), .DIN2(_35878), .Q(_35877) );
  xnr2s1 _35694_inst ( .DIN1(_53180), .DIN2(_35839), .Q(_35878) );
  nnd2s1 _35695_inst ( .DIN1(_35879), .DIN2(_35880), .Q(_35839) );
  nnd2s1 _35696_inst ( .DIN1(_35881), .DIN2(_26347), .Q(_35880) );
  or2s1 _35697_inst ( .DIN1(_35882), .DIN2(_33000), .Q(_35881) );
  nnd2s1 _35698_inst ( .DIN1(_33000), .DIN2(_35882), .Q(_35879) );
  nor2s1 _35699_inst ( .DIN1(_35797), .DIN2(_35883), .Q(_35875) );
  nor2s1 _35700_inst ( .DIN1(_35884), .DIN2(_35885), .Q(_35883) );
  xor2s1 _35701_inst ( .DIN1(_26616), .DIN2(_35886), .Q(_35885) );
  nnd2s1 _35702_inst ( .DIN1(_53428), .DIN2(_26422), .Q(_35886) );
  nor2s1 _35703_inst ( .DIN1(_35887), .DIN2(_35888), .Q(_35884) );
  nnd2s1 _35704_inst ( .DIN1(_35889), .DIN2(_35890), .Q(
        _____________________________218________) );
  nnd2s1 _35705_inst ( .DIN1(_29083), .DIN2(_35891), .Q(_35890) );
  nnd2s1 _35706_inst ( .DIN1(_35892), .DIN2(_35809), .Q(_35891) );
  hi1s1 _35707_inst ( .DIN(_35791), .Q(_35809) );
  nor2s1 _35708_inst ( .DIN1(_35893), .DIN2(_35894), .Q(_35892) );
  nor2s1 _35709_inst ( .DIN1(_35895), .DIN2(_35796), .Q(_35894) );
  xor2s1 _35710_inst ( .DIN1(_33000), .DIN2(_35896), .Q(_35895) );
  xor2s1 _35711_inst ( .DIN1(_26347), .DIN2(_35882), .Q(_35896) );
  nnd2s1 _35712_inst ( .DIN1(_35897), .DIN2(_35898), .Q(_35882) );
  nnd2s1 _35713_inst ( .DIN1(_53342), .DIN2(_35899), .Q(_35898) );
  or2s1 _35714_inst ( .DIN1(_35900), .DIN2(_26828), .Q(_35899) );
  nnd2s1 _35715_inst ( .DIN1(_33017), .DIN2(_35900), .Q(_35897) );
  nor2s1 _35716_inst ( .DIN1(_35797), .DIN2(_26422), .Q(_35893) );
  nnd2s1 _35717_inst ( .DIN1(_35901), .DIN2(_35902), .Q(_35889) );
  nnd2s1 _35718_inst ( .DIN1(_35903), .DIN2(_53427), .Q(_35901) );
  nor2s1 _35719_inst ( .DIN1(_30866), .DIN2(_28646), .Q(_35903) );
  nnd2s1 _35720_inst ( .DIN1(_35904), .DIN2(_35905), .Q(
        _____________________________217________) );
  nor2s1 _35721_inst ( .DIN1(_35906), .DIN2(_35907), .Q(_35905) );
  nor2s1 _35722_inst ( .DIN1(_35908), .DIN2(_35909), .Q(_35907) );
  nor2s1 _35723_inst ( .DIN1(_35910), .DIN2(_35911), .Q(_35909) );
  nor2s1 _35724_inst ( .DIN1(_35796), .DIN2(_35912), .Q(_35911) );
  xor2s1 _35725_inst ( .DIN1(_33017), .DIN2(_35913), .Q(_35912) );
  xnr2s1 _35726_inst ( .DIN1(_53342), .DIN2(_35900), .Q(_35913) );
  nnd2s1 _35727_inst ( .DIN1(_35914), .DIN2(_35915), .Q(_35900) );
  nnd2s1 _35728_inst ( .DIN1(_35916), .DIN2(_26643), .Q(_35915) );
  or2s1 _35729_inst ( .DIN1(_35917), .DIN2(_33035), .Q(_35916) );
  nnd2s1 _35730_inst ( .DIN1(_33035), .DIN2(_35917), .Q(_35914) );
  nor2s1 _35731_inst ( .DIN1(_35797), .DIN2(_35918), .Q(_35910) );
  nnd2s1 _35732_inst ( .DIN1(_35919), .DIN2(_53098), .Q(_35918) );
  nor2s1 _35733_inst ( .DIN1(_35791), .DIN2(_26500), .Q(_35919) );
  nor2s1 _35734_inst ( .DIN1(______[22]), .DIN2(_35920), .Q(_35906) );
  nor2s1 _35735_inst ( .DIN1(_35921), .DIN2(_35922), .Q(_35904) );
  nor2s1 _35736_inst ( .DIN1(_53098), .DIN2(_35923), .Q(_35922) );
  nor2s1 _35737_inst ( .DIN1(_35924), .DIN2(_35908), .Q(_35923) );
  nor2s1 _35738_inst ( .DIN1(_35791), .DIN2(_35925), .Q(_35924) );
  nnd2s1 _35739_inst ( .DIN1(_35796), .DIN2(_26500), .Q(_35925) );
  nor2s1 _35740_inst ( .DIN1(_35926), .DIN2(_35888), .Q(_35791) );
  or2s1 _35741_inst ( .DIN1(_35797), .DIN2(_35887), .Q(_35926) );
  hi1s1 _35742_inst ( .DIN(_35796), .Q(_35797) );
  nnd2s1 _35743_inst ( .DIN1(_35927), .DIN2(_35928), .Q(_35796) );
  nor2s1 _35744_inst ( .DIN1(_35929), .DIN2(_35254), .Q(_35928) );
  nnd2s1 _35745_inst ( .DIN1(_35930), .DIN2(_35103), .Q(_35254) );
  nor2s1 _35746_inst ( .DIN1(_35931), .DIN2(_35932), .Q(_35927) );
  or2s1 _35747_inst ( .DIN1(_35933), .DIN2(_35887), .Q(_35932) );
  hi1s1 _35748_inst ( .DIN(_35934), .Q(_35921) );
  nnd2s1 _35749_inst ( .DIN1(_35935), .DIN2(_35936), .Q(
        _____________________________216________) );
  nnd2s1 _35750_inst ( .DIN1(_35937), .DIN2(_35938), .Q(_35936) );
  xor2s1 _35751_inst ( .DIN1(_26515), .DIN2(_35939), .Q(_35937) );
  nnd2s1 _35752_inst ( .DIN1(_35940), .DIN2(_35941), .Q(_35935) );
  nnd2s1 _35753_inst ( .DIN1(_35942), .DIN2(_35943), .Q(_35941) );
  nnd2s1 _35754_inst ( .DIN1(_35944), .DIN2(_26460), .Q(_35943) );
  nor2s1 _35755_inst ( .DIN1(_35945), .DIN2(_35946), .Q(_35942) );
  nor2s1 _35756_inst ( .DIN1(_35947), .DIN2(_35948), .Q(_35946) );
  xor2s1 _35757_inst ( .DIN1(_33035), .DIN2(_35949), .Q(_35948) );
  xor2s1 _35758_inst ( .DIN1(_26643), .DIN2(_35917), .Q(_35949) );
  nnd2s1 _35759_inst ( .DIN1(_35950), .DIN2(_35951), .Q(_35917) );
  nnd2s1 _35760_inst ( .DIN1(_53191), .DIN2(_35952), .Q(_35951) );
  or2s1 _35761_inst ( .DIN1(_35953), .DIN2(_26800), .Q(_35952) );
  nnd2s1 _35762_inst ( .DIN1(_33065), .DIN2(_35953), .Q(_35950) );
  nor2s1 _35763_inst ( .DIN1(_35954), .DIN2(_35955), .Q(_35945) );
  nor2s1 _35764_inst ( .DIN1(_27393), .DIN2(_35956), .Q(_35955) );
  nnd2s1 _35765_inst ( .DIN1(_35957), .DIN2(_35958), .Q(_35956) );
  or2s1 _35766_inst ( .DIN1(_26460), .DIN2(_35959), .Q(_35957) );
  nnd2s1 _35767_inst ( .DIN1(_35960), .DIN2(_26993), .Q(
        _____________________________215________) );
  nnd2s1 _35768_inst ( .DIN1(_35961), .DIN2(_26996), .Q(_26993) );
  nor2s1 _35769_inst ( .DIN1(_35962), .DIN2(_35963), .Q(_35960) );
  nor2s1 _35770_inst ( .DIN1(_35964), .DIN2(_26996), .Q(_35963) );
  nor2s1 _35771_inst ( .DIN1(_35965), .DIN2(_35966), .Q(_35964) );
  nor2s1 _35772_inst ( .DIN1(_35967), .DIN2(_35947), .Q(_35966) );
  xor2s1 _35773_inst ( .DIN1(_33065), .DIN2(_35968), .Q(_35967) );
  xor2s1 _35774_inst ( .DIN1(_26458), .DIN2(_35953), .Q(_35968) );
  nnd2s1 _35775_inst ( .DIN1(_35969), .DIN2(_35970), .Q(_35953) );
  nnd2s1 _35776_inst ( .DIN1(_53232), .DIN2(_35971), .Q(_35970) );
  nnd2s1 _35777_inst ( .DIN1(_33103), .DIN2(_35972), .Q(_35971) );
  xor2s1 _35778_inst ( .DIN1(_35821), .DIN2(_35973), .Q(_35969) );
  nor2s1 _35779_inst ( .DIN1(_33103), .DIN2(_35972), .Q(_35973) );
  nor2s1 _35780_inst ( .DIN1(_35974), .DIN2(_35975), .Q(_35965) );
  nnd2s1 _35781_inst ( .DIN1(_35976), .DIN2(_35977), .Q(_35974) );
  nnd2s1 _35782_inst ( .DIN1(_35944), .DIN2(_26543), .Q(_35977) );
  nnd2s1 _35783_inst ( .DIN1(_35978), .DIN2(_35979), .Q(_35976) );
  nnd2s1 _35784_inst ( .DIN1(_35947), .DIN2(_26543), .Q(_35978) );
  nor2s1 _35785_inst ( .DIN1(_27007), .DIN2(_35980), .Q(_35962) );
  nor2s1 _35786_inst ( .DIN1(_35981), .DIN2(_27291), .Q(_35980) );
  xor2s1 _35787_inst ( .DIN1(_26640), .DIN2(_53259), .Q(_35981) );
  nor2s1 _35788_inst ( .DIN1(_28998), .DIN2(_35982), .Q(
        _____________________________214________) );
  nnd2s1 _35789_inst ( .DIN1(_35983), .DIN2(_35984), .Q(_35982) );
  nnd2s1 _35790_inst ( .DIN1(_35985), .DIN2(_35947), .Q(_35984) );
  nor2s1 _35791_inst ( .DIN1(_26236), .DIN2(_35975), .Q(_35985) );
  nnd2s1 _35792_inst ( .DIN1(______[10]), .DIN2(_35958), .Q(_35975) );
  nnd2s1 _35793_inst ( .DIN1(_35986), .DIN2(_35954), .Q(_35983) );
  xor2s1 _35794_inst ( .DIN1(_33088), .DIN2(_35987), .Q(_35986) );
  xnr2s1 _35795_inst ( .DIN1(_53232), .DIN2(_35972), .Q(_35987) );
  nnd2s1 _35796_inst ( .DIN1(_35988), .DIN2(_35989), .Q(_35972) );
  nnd2s1 _35797_inst ( .DIN1(_35990), .DIN2(_26489), .Q(_35989) );
  nnd2s1 _35798_inst ( .DIN1(_33108), .DIN2(_35991), .Q(_35990) );
  or2s1 _35799_inst ( .DIN1(_35991), .DIN2(_26797), .Q(_35988) );
  nnd2s1 _35800_inst ( .DIN1(_35992), .DIN2(_35993), .Q(_28998) );
  and2s1 _35801_inst ( .DIN1(_34215), .DIN2(_35994), .Q(_35992) );
  nnd2s1 _35802_inst ( .DIN1(_35995), .DIN2(_28326), .Q(
        _____________________________213________) );
  hi1s1 _35803_inst ( .DIN(_30400), .Q(_28326) );
  nor2s1 _35804_inst ( .DIN1(_35730), .DIN2(_28338), .Q(_30400) );
  nnd2s1 _35805_inst ( .DIN1(_35996), .DIN2(_34090), .Q(_35730) );
  nor2s1 _35806_inst ( .DIN1(_35997), .DIN2(_35998), .Q(_35996) );
  nor2s1 _35807_inst ( .DIN1(_35999), .DIN2(_36000), .Q(_35995) );
  nor2s1 _35808_inst ( .DIN1(_28329), .DIN2(_36001), .Q(_36000) );
  nnd2s1 _35809_inst ( .DIN1(_36002), .DIN2(_36003), .Q(_36001) );
  nor2s1 _35810_inst ( .DIN1(_36004), .DIN2(_36005), .Q(_36003) );
  nor2s1 _35811_inst ( .DIN1(_35954), .DIN2(_35958), .Q(_36005) );
  hi1s1 _35812_inst ( .DIN(_36006), .Q(_35958) );
  nor2s1 _35813_inst ( .DIN1(_35947), .DIN2(_36007), .Q(_36004) );
  xor2s1 _35814_inst ( .DIN1(_33123), .DIN2(_36008), .Q(_36007) );
  xor2s1 _35815_inst ( .DIN1(_26489), .DIN2(_35991), .Q(_36008) );
  nnd2s1 _35816_inst ( .DIN1(_36009), .DIN2(_36010), .Q(_35991) );
  nnd2s1 _35817_inst ( .DIN1(_53150), .DIN2(_36011), .Q(_36010) );
  or2s1 _35818_inst ( .DIN1(_36012), .DIN2(_33129), .Q(_36011) );
  nnd2s1 _35819_inst ( .DIN1(_33129), .DIN2(_36012), .Q(_36009) );
  hi1s1 _35820_inst ( .DIN(_33108), .Q(_33123) );
  nor2s1 _35821_inst ( .DIN1(_35944), .DIN2(_36013), .Q(_36002) );
  nor2s1 _35822_inst ( .DIN1(_35954), .DIN2(_36014), .Q(_36013) );
  nnd2s1 _35823_inst ( .DIN1(_26517), .DIN2(_26236), .Q(_36014) );
  hi1s1 _35824_inst ( .DIN(_35979), .Q(_35944) );
  nnd2s1 _35825_inst ( .DIN1(_35959), .DIN2(_35947), .Q(_35979) );
  nor2s1 _35826_inst ( .DIN1(_26236), .DIN2(_26517), .Q(_35959) );
  nor2s1 _35827_inst ( .DIN1(_28338), .DIN2(_36015), .Q(_35999) );
  nor2s1 _35828_inst ( .DIN1(_36016), .DIN2(_27066), .Q(_36015) );
  xor2s1 _35829_inst ( .DIN1(_26486), .DIN2(_53096), .Q(_36016) );
  hi1s1 _35830_inst ( .DIN(_28329), .Q(_28338) );
  nnd2s1 _35831_inst ( .DIN1(_36017), .DIN2(_36018), .Q(_28329) );
  nor2s1 _35832_inst ( .DIN1(_36019), .DIN2(_36020), .Q(_36018) );
  nnd2s1 _35833_inst ( .DIN1(_36021), .DIN2(_36022), .Q(_36020) );
  nor2s1 _35834_inst ( .DIN1(_36023), .DIN2(_36024), .Q(_36017) );
  nnd2s1 _35835_inst ( .DIN1(_36025), .DIN2(_33094), .Q(
        _____________________________212________) );
  nnd2s1 _35836_inst ( .DIN1(_28381), .DIN2(_29828), .Q(_33094) );
  nor2s1 _35837_inst ( .DIN1(_36026), .DIN2(_36027), .Q(_36025) );
  nor2s1 _35838_inst ( .DIN1(_29828), .DIN2(_36028), .Q(_36027) );
  nor2s1 _35839_inst ( .DIN1(_36029), .DIN2(_36030), .Q(_36028) );
  nor2s1 _35840_inst ( .DIN1(_35947), .DIN2(_36031), .Q(_36030) );
  xor2s1 _35841_inst ( .DIN1(_33141), .DIN2(_36032), .Q(_36031) );
  xor2s1 _35842_inst ( .DIN1(_26261), .DIN2(_36012), .Q(_36032) );
  nnd2s1 _35843_inst ( .DIN1(_36033), .DIN2(_36034), .Q(_36012) );
  nnd2s1 _35844_inst ( .DIN1(_36035), .DIN2(_26741), .Q(_36034) );
  or2s1 _35845_inst ( .DIN1(_36036), .DIN2(_26832), .Q(_36035) );
  nnd2s1 _35846_inst ( .DIN1(_33147), .DIN2(_36036), .Q(_36033) );
  nor2s1 _35847_inst ( .DIN1(_35954), .DIN2(_36037), .Q(_36029) );
  nor2s1 _35848_inst ( .DIN1(_36038), .DIN2(_36039), .Q(_36037) );
  xor2s1 _35849_inst ( .DIN1(_30081), .DIN2(_36006), .Q(_36039) );
  xor2s1 _35850_inst ( .DIN1(_36040), .DIN2(_36041), .Q(_36038) );
  xor2s1 _35851_inst ( .DIN1(_53111), .DIN2(_53217), .Q(_36041) );
  nnd2s1 _35852_inst ( .DIN1(_53148), .DIN2(_53147), .Q(_36040) );
  nor2s1 _35853_inst ( .DIN1(_29849), .DIN2(_36042), .Q(_36026) );
  nor2s1 _35854_inst ( .DIN1(_27365), .DIN2(_26485), .Q(_36042) );
  nnd2s1 _35855_inst ( .DIN1(_36043), .DIN2(_35934), .Q(
        _____________________________211________) );
  nor2s1 _35856_inst ( .DIN1(_36044), .DIN2(_36045), .Q(_36043) );
  nor2s1 _35857_inst ( .DIN1(_35908), .DIN2(_36046), .Q(_36045) );
  nor2s1 _35858_inst ( .DIN1(_36047), .DIN2(_36048), .Q(_36046) );
  nor2s1 _35859_inst ( .DIN1(_35947), .DIN2(_36049), .Q(_36048) );
  xor2s1 _35860_inst ( .DIN1(_36050), .DIN2(_36036), .Q(_36049) );
  xor2s1 _35861_inst ( .DIN1(_36051), .DIN2(_34151), .Q(_36036) );
  nnd2s1 _35862_inst ( .DIN1(_36052), .DIN2(_36053), .Q(_36051) );
  nnd2s1 _35863_inst ( .DIN1(_36054), .DIN2(_26381), .Q(_36053) );
  nnd2s1 _35864_inst ( .DIN1(_33190), .DIN2(_36055), .Q(_36054) );
  or2s1 _35865_inst ( .DIN1(_36055), .DIN2(_33190), .Q(_36052) );
  xor2s1 _35866_inst ( .DIN1(_33147), .DIN2(_53201), .Q(_36050) );
  nor2s1 _35867_inst ( .DIN1(_35954), .DIN2(_36056), .Q(_36047) );
  nnd2s1 _35868_inst ( .DIN1(_36057), .DIN2(_53147), .Q(_36056) );
  nor2s1 _35869_inst ( .DIN1(_36006), .DIN2(_26771), .Q(_36057) );
  nor2s1 _35870_inst ( .DIN1(_36058), .DIN2(_36059), .Q(_36006) );
  or2s1 _35871_inst ( .DIN1(_35272), .DIN2(_36060), .Q(_36058) );
  hi1s1 _35872_inst ( .DIN(_35947), .Q(_35954) );
  nnd2s1 _35873_inst ( .DIN1(_36061), .DIN2(_36062), .Q(_35947) );
  nor2s1 _35874_inst ( .DIN1(_36063), .DIN2(_36064), .Q(_36062) );
  nnd2s1 _35875_inst ( .DIN1(_36065), .DIN2(_36066), .Q(_36064) );
  nor2s1 _35876_inst ( .DIN1(_35273), .DIN2(_36067), .Q(_36061) );
  nor2s1 _35877_inst ( .DIN1(_35920), .DIN2(_36068), .Q(_36044) );
  nor2s1 _35878_inst ( .DIN1(_36069), .DIN2(_27291), .Q(_36068) );
  xor2s1 _35879_inst ( .DIN1(_26263), .DIN2(_53098), .Q(_36069) );
  nnd2s1 _35880_inst ( .DIN1(_36070), .DIN2(_36071), .Q(
        _____________________________210________) );
  nnd2s1 _35881_inst ( .DIN1(_36072), .DIN2(_36073), .Q(_36071) );
  nnd2s1 _35882_inst ( .DIN1(_36074), .DIN2(______[2]), .Q(_36073) );
  nor2s1 _35883_inst ( .DIN1(_53217), .DIN2(_36075), .Q(_36074) );
  nor2s1 _35884_inst ( .DIN1(_36076), .DIN2(_36077), .Q(_36070) );
  nor2s1 _35885_inst ( .DIN1(_36078), .DIN2(_36079), .Q(_36077) );
  xor2s1 _35886_inst ( .DIN1(_36055), .DIN2(_36080), .Q(_36079) );
  xor2s1 _35887_inst ( .DIN1(_26381), .DIN2(_33190), .Q(_36080) );
  xnr2s1 _35888_inst ( .DIN1(_35291), .DIN2(_36081), .Q(_36055) );
  nor2s1 _35889_inst ( .DIN1(_36082), .DIN2(_36083), .Q(_36081) );
  and2s1 _35890_inst ( .DIN1(_36084), .DIN2(_33196), .Q(_36083) );
  nor2s1 _35891_inst ( .DIN1(_53202), .DIN2(_36085), .Q(_36082) );
  nor2s1 _35892_inst ( .DIN1(_33196), .DIN2(_36084), .Q(_36085) );
  nor2s1 _35893_inst ( .DIN1(_36086), .DIN2(_36087), .Q(_36076) );
  nnd2s1 _35894_inst ( .DIN1(_36088), .DIN2(______[2]), .Q(_36087) );
  xor2s1 _35895_inst ( .DIN1(_26390), .DIN2(_36089), .Q(_36086) );
  nnd2s1 _35896_inst ( .DIN1(_36090), .DIN2(_36091), .Q(
        _____________________________20________) );
  nnd2s1 _35897_inst ( .DIN1(_36092), .DIN2(_35864), .Q(_36091) );
  nnd2s1 _35898_inst ( .DIN1(_36093), .DIN2(_36094), .Q(_36092) );
  nnd2s1 _35899_inst ( .DIN1(_36095), .DIN2(_36096), .Q(_36094) );
  nor2s1 _35900_inst ( .DIN1(_26988), .DIN2(_26362), .Q(_36095) );
  nnd2s1 _35901_inst ( .DIN1(_36097), .DIN2(_36098), .Q(_36093) );
  hi1s1 _35902_inst ( .DIN(_35136), .Q(_36098) );
  xor2s1 _35903_inst ( .DIN1(_35239), .DIN2(_36099), .Q(_36097) );
  xor2s1 _35904_inst ( .DIN1(_26638), .DIN2(_35855), .Q(_36099) );
  nnd2s1 _35905_inst ( .DIN1(_36100), .DIN2(_36101), .Q(_35855) );
  nnd2s1 _35906_inst ( .DIN1(_36102), .DIN2(_26439), .Q(_36101) );
  nnd2s1 _35907_inst ( .DIN1(_36103), .DIN2(_36104), .Q(_36102) );
  nnd2s1 _35908_inst ( .DIN1(_35265), .DIN2(_36105), .Q(_36100) );
  hi1s1 _35909_inst ( .DIN(_36104), .Q(_35265) );
  xnr2s1 _35910_inst ( .DIN1(_35861), .DIN2(_26761), .Q(_35239) );
  nnd2s1 _35911_inst ( .DIN1(_36106), .DIN2(_36107), .Q(_35860) );
  nnd2s1 _35912_inst ( .DIN1(_53314), .DIN2(_36108), .Q(_36107) );
  nnd2s1 _35913_inst ( .DIN1(_36109), .DIN2(_36110), .Q(_36108) );
  nnd2s1 _35914_inst ( .DIN1(_36111), .DIN2(_36112), .Q(_36106) );
  hi1s1 _35915_inst ( .DIN(_36109), .Q(_36112) );
  nnd2s1 _35916_inst ( .DIN1(_36113), .DIN2(_34298), .Q(_36090) );
  nnd2s1 _35917_inst ( .DIN1(_53166), .DIN2(_35614), .Q(_36113) );
  nnd2s1 _35918_inst ( .DIN1(_36114), .DIN2(_27608), .Q(
        _____________________________209________) );
  nor2s1 _35919_inst ( .DIN1(_36115), .DIN2(_36116), .Q(_36114) );
  nor2s1 _35920_inst ( .DIN1(_27611), .DIN2(_36117), .Q(_36116) );
  nor2s1 _35921_inst ( .DIN1(_27066), .DIN2(_26504), .Q(_36117) );
  nor2s1 _35922_inst ( .DIN1(_36118), .DIN2(_27616), .Q(_36115) );
  nor2s1 _35923_inst ( .DIN1(_36119), .DIN2(_36120), .Q(_36118) );
  nor2s1 _35924_inst ( .DIN1(_36075), .DIN2(_36121), .Q(_36120) );
  xor2s1 _35925_inst ( .DIN1(_53148), .DIN2(_53217), .Q(_36121) );
  hi1s1 _35926_inst ( .DIN(_36122), .Q(_36075) );
  nor2s1 _35927_inst ( .DIN1(_36123), .DIN2(_36124), .Q(_36119) );
  xor2s1 _35928_inst ( .DIN1(_33882), .DIN2(_36125), .Q(_36123) );
  xnr2s1 _35929_inst ( .DIN1(_53202), .DIN2(_36084), .Q(_36125) );
  nnd2s1 _35930_inst ( .DIN1(_36126), .DIN2(_36127), .Q(_36084) );
  nnd2s1 _35931_inst ( .DIN1(_53205), .DIN2(_36128), .Q(_36127) );
  or2s1 _35932_inst ( .DIN1(_36129), .DIN2(_33213), .Q(_36128) );
  nnd2s1 _35933_inst ( .DIN1(_33213), .DIN2(_36129), .Q(_36126) );
  nnd2s1 _35934_inst ( .DIN1(_36130), .DIN2(_36131), .Q(
        _____________________________208________) );
  nor2s1 _35935_inst ( .DIN1(_36132), .DIN2(_36133), .Q(_36131) );
  nor2s1 _35936_inst ( .DIN1(_30360), .DIN2(_36134), .Q(_36133) );
  or2s1 _35937_inst ( .DIN1(_36078), .DIN2(_36135), .Q(_36134) );
  nor2s1 _35938_inst ( .DIN1(_30912), .DIN2(_36136), .Q(_36132) );
  nnd2s1 _35939_inst ( .DIN1(_35920), .DIN2(_36135), .Q(_36136) );
  xnr2s1 _35940_inst ( .DIN1(_33213), .DIN2(_36137), .Q(_36135) );
  xnr2s1 _35941_inst ( .DIN1(_53205), .DIN2(_36129), .Q(_36137) );
  nnd2s1 _35942_inst ( .DIN1(_36138), .DIN2(_36139), .Q(_36129) );
  nnd2s1 _35943_inst ( .DIN1(_53151), .DIN2(_36140), .Q(_36139) );
  or2s1 _35944_inst ( .DIN1(_36141), .DIN2(_33907), .Q(_36140) );
  nnd2s1 _35945_inst ( .DIN1(_33907), .DIN2(_36141), .Q(_36138) );
  nor2s1 _35946_inst ( .DIN1(_36142), .DIN2(_36143), .Q(_36130) );
  nor2s1 _35947_inst ( .DIN1(_36144), .DIN2(_36145), .Q(_36143) );
  nor2s1 _35948_inst ( .DIN1(_36146), .DIN2(_36147), .Q(_36144) );
  nnd2s1 _35949_inst ( .DIN1(_30912), .DIN2(_36122), .Q(_36147) );
  xor2s1 _35950_inst ( .DIN1(_53153), .DIN2(_53160), .Q(_36146) );
  nor2s1 _35951_inst ( .DIN1(_36148), .DIN2(_36149), .Q(_36142) );
  nnd2s1 _35952_inst ( .DIN1(_36088), .DIN2(______[14]), .Q(_36149) );
  xor2s1 _35953_inst ( .DIN1(_26609), .DIN2(_36089), .Q(_36148) );
  nnd2s1 _35954_inst ( .DIN1(_36150), .DIN2(_33229), .Q(
        _____________________________207________) );
  nor2s1 _35955_inst ( .DIN1(_36151), .DIN2(_36152), .Q(_36150) );
  nor2s1 _35956_inst ( .DIN1(_27509), .DIN2(_36153), .Q(_36152) );
  nnd2s1 _35957_inst ( .DIN1(_36154), .DIN2(_36155), .Q(_36153) );
  nnd2s1 _35958_inst ( .DIN1(_36156), .DIN2(_36157), .Q(_36155) );
  xor2s1 _35959_inst ( .DIN1(_33225), .DIN2(_36158), .Q(_36157) );
  xor2s1 _35960_inst ( .DIN1(_26606), .DIN2(_36141), .Q(_36158) );
  nnd2s1 _35961_inst ( .DIN1(_36159), .DIN2(_36160), .Q(_36141) );
  nnd2s1 _35962_inst ( .DIN1(_36161), .DIN2(_26504), .Q(_36160) );
  or2s1 _35963_inst ( .DIN1(_36162), .DIN2(_26834), .Q(_36161) );
  nnd2s1 _35964_inst ( .DIN1(_26834), .DIN2(_36162), .Q(_36159) );
  nnd2s1 _35965_inst ( .DIN1(_36163), .DIN2(_36122), .Q(_36154) );
  xor2s1 _35966_inst ( .DIN1(_36164), .DIN2(_53159), .Q(_36163) );
  nnd2s1 _35967_inst ( .DIN1(_53153), .DIN2(_53152), .Q(_36164) );
  nor2s1 _35968_inst ( .DIN1(_27512), .DIN2(_36165), .Q(_36151) );
  nor2s1 _35969_inst ( .DIN1(_53465), .DIN2(_26773), .Q(_36165) );
  nor2s1 _35970_inst ( .DIN1(_28218), .DIN2(_36166), .Q(
        _____________________________206________) );
  nor2s1 _35971_inst ( .DIN1(_36167), .DIN2(_36168), .Q(_36166) );
  nnd2s1 _35972_inst ( .DIN1(_36169), .DIN2(_36170), .Q(_36168) );
  nnd2s1 _35973_inst ( .DIN1(_36171), .DIN2(_27329), .Q(_36169) );
  nnd2s1 _35974_inst ( .DIN1(_36172), .DIN2(_36173), .Q(_36167) );
  nnd2s1 _35975_inst ( .DIN1(_36174), .DIN2(_36156), .Q(_36173) );
  nor2s1 _35976_inst ( .DIN1(_36171), .DIN2(_27329), .Q(_36174) );
  xor2s1 _35977_inst ( .DIN1(_26834), .DIN2(_36175), .Q(_36171) );
  xor2s1 _35978_inst ( .DIN1(_26504), .DIN2(_36162), .Q(_36175) );
  nnd2s1 _35979_inst ( .DIN1(_36176), .DIN2(_36177), .Q(_36162) );
  nnd2s1 _35980_inst ( .DIN1(_36178), .DIN2(_26372), .Q(_36177) );
  or2s1 _35981_inst ( .DIN1(_36179), .DIN2(_33271), .Q(_36178) );
  nnd2s1 _35982_inst ( .DIN1(_33271), .DIN2(_36179), .Q(_36176) );
  nnd2s1 _35983_inst ( .DIN1(_36180), .DIN2(_36124), .Q(_36172) );
  nnd2s1 _35984_inst ( .DIN1(_53152), .DIN2(_27338), .Q(_36180) );
  nnd2s1 _35985_inst ( .DIN1(_36181), .DIN2(_36182), .Q(
        _____________________________205________) );
  nor2s1 _35986_inst ( .DIN1(_36183), .DIN2(_36184), .Q(_36182) );
  nor2s1 _35987_inst ( .DIN1(_53159), .DIN2(_36185), .Q(_36184) );
  nnd2s1 _35988_inst ( .DIN1(_36072), .DIN2(_53153), .Q(_36185) );
  hi1s1 _35989_inst ( .DIN(_36145), .Q(_36072) );
  nor2s1 _35990_inst ( .DIN1(_36186), .DIN2(_26495), .Q(_36183) );
  nor2s1 _35991_inst ( .DIN1(_36187), .DIN2(_36088), .Q(_36186) );
  nor2s1 _35992_inst ( .DIN1(_35920), .DIN2(_35465), .Q(_36088) );
  nor2s1 _35993_inst ( .DIN1(_53153), .DIN2(_36145), .Q(_36187) );
  nnd2s1 _35994_inst ( .DIN1(_35920), .DIN2(_36124), .Q(_36145) );
  nor2s1 _35995_inst ( .DIN1(_36188), .DIN2(_36189), .Q(_36181) );
  nor2s1 _35996_inst ( .DIN1(_35908), .DIN2(_36170), .Q(_36189) );
  nnd2s1 _35997_inst ( .DIN1(_36190), .DIN2(_36124), .Q(_36170) );
  nnd2s1 _35998_inst ( .DIN1(______[16]), .DIN2(_36122), .Q(_36190) );
  nor2s1 _35999_inst ( .DIN1(_36078), .DIN2(_36191), .Q(_36188) );
  xor2s1 _36000_inst ( .DIN1(_33271), .DIN2(_36192), .Q(_36191) );
  xor2s1 _36001_inst ( .DIN1(_26372), .DIN2(_36179), .Q(_36192) );
  nnd2s1 _36002_inst ( .DIN1(_36193), .DIN2(_36194), .Q(_36179) );
  nnd2s1 _36003_inst ( .DIN1(_53206), .DIN2(_36195), .Q(_36194) );
  or2s1 _36004_inst ( .DIN1(_36196), .DIN2(_33291), .Q(_36195) );
  nnd2s1 _36005_inst ( .DIN1(_33291), .DIN2(_36196), .Q(_36193) );
  nnd2s1 _36006_inst ( .DIN1(_36156), .DIN2(_35920), .Q(_36078) );
  hi1s1 _36007_inst ( .DIN(_36124), .Q(_36156) );
  nnd2s1 _36008_inst ( .DIN1(_36197), .DIN2(_36198), .Q(_36124) );
  nor2s1 _36009_inst ( .DIN1(_36199), .DIN2(_36200), .Q(_36198) );
  nnd2s1 _36010_inst ( .DIN1(_36201), .DIN2(_36202), .Q(_36200) );
  nor2s1 _36011_inst ( .DIN1(_36203), .DIN2(_36122), .Q(_36197) );
  nnd2s1 _36012_inst ( .DIN1(_36204), .DIN2(_36205), .Q(_36122) );
  nor2s1 _36013_inst ( .DIN1(_35253), .DIN2(_36206), .Q(_36205) );
  nnd2s1 _36014_inst ( .DIN1(_36207), .DIN2(_35270), .Q(_36206) );
  nor2s1 _36015_inst ( .DIN1(_36208), .DIN2(_36209), .Q(_36204) );
  nnd2s1 _36016_inst ( .DIN1(_36210), .DIN2(_27660), .Q(
        _____________________________204________) );
  nor2s1 _36017_inst ( .DIN1(_36211), .DIN2(_36212), .Q(_36210) );
  nor2s1 _36018_inst ( .DIN1(_27663), .DIN2(_36213), .Q(_36212) );
  nor2s1 _36019_inst ( .DIN1(_36214), .DIN2(_36215), .Q(_36213) );
  nor2s1 _36020_inst ( .DIN1(_36216), .DIN2(_36217), .Q(_36215) );
  xor2s1 _36021_inst ( .DIN1(_33310), .DIN2(_36218), .Q(_36217) );
  xor2s1 _36022_inst ( .DIN1(_26265), .DIN2(_36196), .Q(_36218) );
  nnd2s1 _36023_inst ( .DIN1(_36219), .DIN2(_36220), .Q(_36196) );
  nnd2s1 _36024_inst ( .DIN1(_53158), .DIN2(_36221), .Q(_36220) );
  or2s1 _36025_inst ( .DIN1(_36222), .DIN2(_26822), .Q(_36221) );
  nnd2s1 _36026_inst ( .DIN1(_33982), .DIN2(_36222), .Q(_36219) );
  nor2s1 _36027_inst ( .DIN1(_36223), .DIN2(_36224), .Q(_36214) );
  nor2s1 _36028_inst ( .DIN1(_28646), .DIN2(_36225), .Q(_36224) );
  xor2s1 _36029_inst ( .DIN1(_34026), .DIN2(_36226), .Q(_36225) );
  nnd2s1 _36030_inst ( .DIN1(_36227), .DIN2(_36228), .Q(_36226) );
  xor2s1 _36031_inst ( .DIN1(_53154), .DIN2(_36229), .Q(_36227) );
  nor2s1 _36032_inst ( .DIN1(_27672), .DIN2(_36230), .Q(_36211) );
  nor2s1 _36033_inst ( .DIN1(_27365), .DIN2(_26455), .Q(_36230) );
  nnd2s1 _36034_inst ( .DIN1(_36231), .DIN2(_35341), .Q(
        _____________________________203________) );
  nnd2s1 _36035_inst ( .DIN1(_27749), .DIN2(_34214), .Q(_35341) );
  nor2s1 _36036_inst ( .DIN1(_36232), .DIN2(_36233), .Q(_36231) );
  nor2s1 _36037_inst ( .DIN1(_27749), .DIN2(_36234), .Q(_36233) );
  nor2s1 _36038_inst ( .DIN1(_36235), .DIN2(_36236), .Q(_36234) );
  nor2s1 _36039_inst ( .DIN1(_36216), .DIN2(_36237), .Q(_36236) );
  xor2s1 _36040_inst ( .DIN1(_33315), .DIN2(_36238), .Q(_36237) );
  xnr2s1 _36041_inst ( .DIN1(_53158), .DIN2(_36222), .Q(_36238) );
  nnd2s1 _36042_inst ( .DIN1(_36239), .DIN2(_36240), .Q(_36222) );
  nnd2s1 _36043_inst ( .DIN1(_53207), .DIN2(_36241), .Q(_36240) );
  or2s1 _36044_inst ( .DIN1(_36242), .DIN2(_33344), .Q(_36241) );
  nnd2s1 _36045_inst ( .DIN1(_33344), .DIN2(_36242), .Q(_36239) );
  hi1s1 _36046_inst ( .DIN(_33982), .Q(_33315) );
  nor2s1 _36047_inst ( .DIN1(_36223), .DIN2(_36243), .Q(_36235) );
  nor2s1 _36048_inst ( .DIN1(_27393), .DIN2(_36244), .Q(_36243) );
  nnd2s1 _36049_inst ( .DIN1(_36245), .DIN2(_36228), .Q(_36244) );
  xor2s1 _36050_inst ( .DIN1(_53157), .DIN2(_36229), .Q(_36245) );
  nor2s1 _36051_inst ( .DIN1(_28010), .DIN2(_36246), .Q(_36232) );
  xor2s1 _36052_inst ( .DIN1(_52847), .DIN2(_53156), .Q(_36246) );
  nnd2s1 _36053_inst ( .DIN1(_36247), .DIN2(_35934), .Q(
        _____________________________202________) );
  nnd2s1 _36054_inst ( .DIN1(_35465), .DIN2(_35908), .Q(_35934) );
  hi1s1 _36055_inst ( .DIN(_28350), .Q(_35465) );
  nnd2s1 _36056_inst ( .DIN1(_35720), .DIN2(_36248), .Q(_28350) );
  nor2s1 _36057_inst ( .DIN1(_36249), .DIN2(_36250), .Q(_36247) );
  nor2s1 _36058_inst ( .DIN1(_35908), .DIN2(_36251), .Q(_36250) );
  nor2s1 _36059_inst ( .DIN1(_36252), .DIN2(_36253), .Q(_36251) );
  nor2s1 _36060_inst ( .DIN1(_36216), .DIN2(_36254), .Q(_36253) );
  xor2s1 _36061_inst ( .DIN1(_26790), .DIN2(_36255), .Q(_36254) );
  xor2s1 _36062_inst ( .DIN1(_26407), .DIN2(_36242), .Q(_36255) );
  nnd2s1 _36063_inst ( .DIN1(_36256), .DIN2(_36257), .Q(_36242) );
  nnd2s1 _36064_inst ( .DIN1(_53210), .DIN2(_36258), .Q(_36257) );
  or2s1 _36065_inst ( .DIN1(_36259), .DIN2(_26801), .Q(_36258) );
  nnd2s1 _36066_inst ( .DIN1(_33349), .DIN2(_36259), .Q(_36256) );
  nor2s1 _36067_inst ( .DIN1(_36223), .DIN2(_36260), .Q(_36252) );
  nnd2s1 _36068_inst ( .DIN1(_36261), .DIN2(______[30]), .Q(_36260) );
  nor2s1 _36069_inst ( .DIN1(_53397), .DIN2(_36262), .Q(_36261) );
  nor2s1 _36070_inst ( .DIN1(_35920), .DIN2(_36263), .Q(_36249) );
  nor2s1 _36071_inst ( .DIN1(_36264), .DIN2(_36265), .Q(_36263) );
  hi1s1 _36072_inst ( .DIN(_36089), .Q(_36265) );
  nnd2s1 _36073_inst ( .DIN1(_53160), .DIN2(_53159), .Q(_36089) );
  nor2s1 _36074_inst ( .DIN1(_53159), .DIN2(_53160), .Q(_36264) );
  hi1s1 _36075_inst ( .DIN(_35908), .Q(_35920) );
  nnd2s1 _36076_inst ( .DIN1(_36266), .DIN2(_35720), .Q(_35908) );
  nnd2s1 _36077_inst ( .DIN1(_36267), .DIN2(_36268), .Q(
        _____________________________201________) );
  nnd2s1 _36078_inst ( .DIN1(_36269), .DIN2(_36024), .Q(_36268) );
  xor2s1 _36079_inst ( .DIN1(_26384), .DIN2(_30168), .Q(_36269) );
  nnd2s1 _36080_inst ( .DIN1(_53162), .DIN2(_53163), .Q(_30168) );
  nnd2s1 _36081_inst ( .DIN1(_36270), .DIN2(_28792), .Q(_36267) );
  nor2s1 _36082_inst ( .DIN1(_36271), .DIN2(_36272), .Q(_36270) );
  nor2s1 _36083_inst ( .DIN1(_36216), .DIN2(_36273), .Q(_36272) );
  xor2s1 _36084_inst ( .DIN1(_33349), .DIN2(_36274), .Q(_36273) );
  xnr2s1 _36085_inst ( .DIN1(_53210), .DIN2(_36259), .Q(_36274) );
  nnd2s1 _36086_inst ( .DIN1(_36275), .DIN2(_36276), .Q(_36259) );
  nnd2s1 _36087_inst ( .DIN1(_36277), .DIN2(_26351), .Q(_36276) );
  or2s1 _36088_inst ( .DIN1(_36278), .DIN2(_33388), .Q(_36277) );
  nnd2s1 _36089_inst ( .DIN1(_33388), .DIN2(_36278), .Q(_36275) );
  nor2s1 _36090_inst ( .DIN1(_36223), .DIN2(_36279), .Q(_36271) );
  nnd2s1 _36091_inst ( .DIN1(_36280), .DIN2(_36281), .Q(_36279) );
  nnd2s1 _36092_inst ( .DIN1(_53397), .DIN2(_26390), .Q(_36281) );
  nor2s1 _36093_inst ( .DIN1(_36229), .DIN2(_36262), .Q(_36280) );
  nor2s1 _36094_inst ( .DIN1(_26390), .DIN2(_53397), .Q(_36229) );
  nnd2s1 _36095_inst ( .DIN1(_36282), .DIN2(_36283), .Q(
        _____________________________200________) );
  nnd2s1 _36096_inst ( .DIN1(_36284), .DIN2(_36285), .Q(_36283) );
  nnd2s1 _36097_inst ( .DIN1(_36286), .DIN2(______[24]), .Q(_36285) );
  nor2s1 _36098_inst ( .DIN1(_36262), .DIN2(_36287), .Q(_36286) );
  hi1s1 _36099_inst ( .DIN(_36288), .Q(_36284) );
  nor2s1 _36100_inst ( .DIN1(_36289), .DIN2(_36290), .Q(_36282) );
  nor2s1 _36101_inst ( .DIN1(_36287), .DIN2(_36291), .Q(_36290) );
  xor2s1 _36102_inst ( .DIN1(_26483), .DIN2(_53168), .Q(_36287) );
  nor2s1 _36103_inst ( .DIN1(_36292), .DIN2(_36293), .Q(_36289) );
  xor2s1 _36104_inst ( .DIN1(_33388), .DIN2(_36294), .Q(_36293) );
  xor2s1 _36105_inst ( .DIN1(_26351), .DIN2(_36278), .Q(_36294) );
  nnd2s1 _36106_inst ( .DIN1(_36295), .DIN2(_36296), .Q(_36278) );
  nnd2s1 _36107_inst ( .DIN1(_36297), .DIN2(_26716), .Q(_36296) );
  or2s1 _36108_inst ( .DIN1(_36298), .DIN2(_26802), .Q(_36297) );
  nnd2s1 _36109_inst ( .DIN1(_26802), .DIN2(_36298), .Q(_36295) );
  nnd2s1 _36110_inst ( .DIN1(_36299), .DIN2(_36300), .Q(
        _____________________________1________) );
  nnd2s1 _36111_inst ( .DIN1(_36301), .DIN2(_36302), .Q(_36300) );
  xor2s1 _36112_inst ( .DIN1(_53315), .DIN2(_53325), .Q(_36301) );
  nor2s1 _36113_inst ( .DIN1(_36303), .DIN2(_36304), .Q(_36299) );
  nor2s1 _36114_inst ( .DIN1(_36305), .DIN2(_34082), .Q(_36304) );
  nnd2s1 _36115_inst ( .DIN1(_33871), .DIN2(_28542), .Q(_34082) );
  xor2s1 _36116_inst ( .DIN1(_53319), .DIN2(_36306), .Q(_36305) );
  nor2s1 _36117_inst ( .DIN1(_33464), .DIN2(_36307), .Q(_36303) );
  nnd2s1 _36118_inst ( .DIN1(_28542), .DIN2(_53080), .Q(_36307) );
  hi1s1 _36119_inst ( .DIN(_33678), .Q(_33464) );
  nor2s1 _36120_inst ( .DIN1(_27761), .DIN2(_33871), .Q(_33678) );
  hi1s1 _36121_inst ( .DIN(_33460), .Q(_33871) );
  nnd2s1 _36122_inst ( .DIN1(_33044), .DIN2(_36308), .Q(_33460) );
  and2s1 _36123_inst ( .DIN1(_36309), .DIN2(_34306), .Q(_27761) );
  nor2s1 _36124_inst ( .DIN1(_36310), .DIN2(_27683), .Q(_36309) );
  nnd2s1 _36125_inst ( .DIN1(_36311), .DIN2(_36312), .Q(
        _____________________________19________) );
  nor2s1 _36126_inst ( .DIN1(_36313), .DIN2(_36314), .Q(_36312) );
  nor2s1 _36127_inst ( .DIN1(_53196), .DIN2(_36315), .Q(_36314) );
  nnd2s1 _36128_inst ( .DIN1(_36096), .DIN2(_26348), .Q(_36315) );
  hi1s1 _36129_inst ( .DIN(_35147), .Q(_36096) );
  nor2s1 _36130_inst ( .DIN1(_36316), .DIN2(_26244), .Q(_36313) );
  nor2s1 _36131_inst ( .DIN1(_36317), .DIN2(_35614), .Q(_36316) );
  nor2s1 _36132_inst ( .DIN1(_26348), .DIN2(_35147), .Q(_36317) );
  nnd2s1 _36133_inst ( .DIN1(_34301), .DIN2(_35373), .Q(_35147) );
  nor2s1 _36134_inst ( .DIN1(_35133), .DIN2(_36318), .Q(_36311) );
  nor2s1 _36135_inst ( .DIN1(_35136), .DIN2(_36319), .Q(_36318) );
  xor2s1 _36136_inst ( .DIN1(_36104), .DIN2(_36320), .Q(_36319) );
  xor2s1 _36137_inst ( .DIN1(_26439), .DIN2(_36103), .Q(_36320) );
  hi1s1 _36138_inst ( .DIN(_36105), .Q(_36103) );
  nnd2s1 _36139_inst ( .DIN1(_36321), .DIN2(_36322), .Q(_36105) );
  nnd2s1 _36140_inst ( .DIN1(_36323), .DIN2(_26499), .Q(_36322) );
  or2s1 _36141_inst ( .DIN1(_36324), .DIN2(_35293), .Q(_36323) );
  nnd2s1 _36142_inst ( .DIN1(_35293), .DIN2(_36324), .Q(_36321) );
  xor2s1 _36143_inst ( .DIN1(_36109), .DIN2(_36325), .Q(_36104) );
  xor2s1 _36144_inst ( .DIN1(_26343), .DIN2(_36110), .Q(_36325) );
  xor2s1 _36145_inst ( .DIN1(_36326), .DIN2(_36327), .Q(_36109) );
  xor2s1 _36146_inst ( .DIN1(_30367), .DIN2(_36328), .Q(_36327) );
  nnd2s1 _36147_inst ( .DIN1(_36329), .DIN2(_36330), .Q(_36326) );
  nnd2s1 _36148_inst ( .DIN1(_36331), .DIN2(_36332), .Q(_36330) );
  nnd2s1 _36149_inst ( .DIN1(_36333), .DIN2(_36334), .Q(_36331) );
  or2s1 _36150_inst ( .DIN1(_36334), .DIN2(_36333), .Q(_36329) );
  nnd2s1 _36151_inst ( .DIN1(_35387), .DIN2(_34301), .Q(_35136) );
  nor2s1 _36152_inst ( .DIN1(_35864), .DIN2(_34298), .Q(_35133) );
  nnd2s1 _36153_inst ( .DIN1(_36335), .DIN2(_34306), .Q(_35864) );
  hi1s1 _36154_inst ( .DIN(_34272), .Q(_34306) );
  nnd2s1 _36155_inst ( .DIN1(_36336), .DIN2(_36337), .Q(_34272) );
  nor2s1 _36156_inst ( .DIN1(_35387), .DIN2(_27683), .Q(_36335) );
  hi1s1 _36157_inst ( .DIN(_35373), .Q(_35387) );
  nnd2s1 _36158_inst ( .DIN1(_27536), .DIN2(_36308), .Q(_35373) );
  hi1s1 _36159_inst ( .DIN(_27503), .Q(_27536) );
  nnd2s1 _36160_inst ( .DIN1(_27567), .DIN2(_36337), .Q(_27503) );
  nnd2s1 _36161_inst ( .DIN1(_36338), .DIN2(_36339), .Q(
        _____________________________199________) );
  nnd2s1 _36162_inst ( .DIN1(_36340), .DIN2(_36341), .Q(_36339) );
  hi1s1 _36163_inst ( .DIN(_36292), .Q(_36341) );
  nnd2s1 _36164_inst ( .DIN1(_36223), .DIN2(_35015), .Q(_36292) );
  hi1s1 _36165_inst ( .DIN(_36216), .Q(_36223) );
  xor2s1 _36166_inst ( .DIN1(_36342), .DIN2(_36343), .Q(_36340) );
  xor2s1 _36167_inst ( .DIN1(_36298), .DIN2(_33398), .Q(_36343) );
  nnd2s1 _36168_inst ( .DIN1(_36344), .DIN2(_36345), .Q(_36298) );
  nnd2s1 _36169_inst ( .DIN1(_53256), .DIN2(_36346), .Q(_36345) );
  or2s1 _36170_inst ( .DIN1(_36347), .DIN2(_33419), .Q(_36346) );
  nnd2s1 _36171_inst ( .DIN1(_33419), .DIN2(_36347), .Q(_36344) );
  xor2s1 _36172_inst ( .DIN1(_34338), .DIN2(_53214), .Q(_36342) );
  nor2s1 _36173_inst ( .DIN1(_36348), .DIN2(_36349), .Q(_36338) );
  nor2s1 _36174_inst ( .DIN1(_36350), .DIN2(_36288), .Q(_36349) );
  nnd2s1 _36175_inst ( .DIN1(_35015), .DIN2(_36216), .Q(_36288) );
  nor2s1 _36176_inst ( .DIN1(_36262), .DIN2(_36351), .Q(_36350) );
  xor2s1 _36177_inst ( .DIN1(_53169), .DIN2(_36352), .Q(_36351) );
  nor2s1 _36178_inst ( .DIN1(_53168), .DIN2(_53167), .Q(_36352) );
  hi1s1 _36179_inst ( .DIN(_36228), .Q(_36262) );
  nor2s1 _36180_inst ( .DIN1(_36291), .DIN2(_36353), .Q(_36348) );
  nnd2s1 _36181_inst ( .DIN1(______[10]), .DIN2(_36354), .Q(_36353) );
  xor2s1 _36182_inst ( .DIN1(_26252), .DIN2(_36355), .Q(_36354) );
  nnd2s1 _36183_inst ( .DIN1(_53168), .DIN2(_53167), .Q(_36355) );
  nnd2s1 _36184_inst ( .DIN1(_36356), .DIN2(_36357), .Q(
        _____________________________198________) );
  or2s1 _36185_inst ( .DIN1(_36358), .DIN2(_36359), .Q(_36357) );
  nor2s1 _36186_inst ( .DIN1(_36360), .DIN2(_36361), .Q(_36356) );
  nor2s1 _36187_inst ( .DIN1(_36362), .DIN2(_26501), .Q(_36361) );
  nor2s1 _36188_inst ( .DIN1(_36363), .DIN2(_36364), .Q(_36362) );
  nor2s1 _36189_inst ( .DIN1(_26774), .DIN2(_36291), .Q(_36363) );
  nor2s1 _36190_inst ( .DIN1(_36365), .DIN2(_36366), .Q(_36360) );
  xor2s1 _36191_inst ( .DIN1(_34102), .DIN2(_36367), .Q(_36366) );
  xor2s1 _36192_inst ( .DIN1(_26272), .DIN2(_36347), .Q(_36367) );
  nnd2s1 _36193_inst ( .DIN1(_36368), .DIN2(_36369), .Q(_36347) );
  nnd2s1 _36194_inst ( .DIN1(_36370), .DIN2(_26533), .Q(_36369) );
  or2s1 _36195_inst ( .DIN1(_36371), .DIN2(_26831), .Q(_36370) );
  nnd2s1 _36196_inst ( .DIN1(_26831), .DIN2(_36371), .Q(_36368) );
  hi1s1 _36197_inst ( .DIN(_33419), .Q(_34102) );
  nnd2s1 _36198_inst ( .DIN1(_36372), .DIN2(_36373), .Q(
        _____________________________197________) );
  nnd2s1 _36199_inst ( .DIN1(_36374), .DIN2(_36375), .Q(_36373) );
  xnr2s1 _36200_inst ( .DIN1(_26831), .DIN2(_36376), .Q(_36375) );
  xor2s1 _36201_inst ( .DIN1(_26533), .DIN2(_36371), .Q(_36376) );
  nnd2s1 _36202_inst ( .DIN1(_36377), .DIN2(_36378), .Q(_36371) );
  nnd2s1 _36203_inst ( .DIN1(_53220), .DIN2(_36379), .Q(_36378) );
  or2s1 _36204_inst ( .DIN1(_36380), .DIN2(_33449), .Q(_36379) );
  nnd2s1 _36205_inst ( .DIN1(_33449), .DIN2(_36380), .Q(_36377) );
  hi1s1 _36206_inst ( .DIN(_34138), .Q(_33449) );
  hi1s1 _36207_inst ( .DIN(_36365), .Q(_36374) );
  nor2s1 _36208_inst ( .DIN1(_36381), .DIN2(_36382), .Q(_36372) );
  nor2s1 _36209_inst ( .DIN1(_36383), .DIN2(_36359), .Q(_36382) );
  and2s1 _36210_inst ( .DIN1(_36358), .DIN2(_36384), .Q(_36383) );
  nor2s1 _36211_inst ( .DIN1(_36291), .DIN2(_36385), .Q(_36381) );
  nnd2s1 _36212_inst ( .DIN1(______[0]), .DIN2(_36384), .Q(_36385) );
  xor2s1 _36213_inst ( .DIN1(_26252), .DIN2(_26625), .Q(_36384) );
  hi1s1 _36214_inst ( .DIN(_35012), .Q(_36291) );
  nor2s1 _36215_inst ( .DIN1(_35015), .DIN2(_36386), .Q(_35012) );
  nnd2s1 _36216_inst ( .DIN1(_36387), .DIN2(_27450), .Q(
        _____________________________196________) );
  nnd2s1 _36217_inst ( .DIN1(_36388), .DIN2(_27453), .Q(_27450) );
  nor2s1 _36218_inst ( .DIN1(_36389), .DIN2(_36390), .Q(_36387) );
  nor2s1 _36219_inst ( .DIN1(_27453), .DIN2(_36391), .Q(_36390) );
  nnd2s1 _36220_inst ( .DIN1(_36392), .DIN2(_36393), .Q(_36391) );
  nnd2s1 _36221_inst ( .DIN1(_36394), .DIN2(_36395), .Q(_36393) );
  xor2s1 _36222_inst ( .DIN1(_34138), .DIN2(_36396), .Q(_36394) );
  xor2s1 _36223_inst ( .DIN1(_26594), .DIN2(_36380), .Q(_36396) );
  nnd2s1 _36224_inst ( .DIN1(_36397), .DIN2(_36398), .Q(_36380) );
  nnd2s1 _36225_inst ( .DIN1(_36399), .DIN2(_26268), .Q(_36398) );
  or2s1 _36226_inst ( .DIN1(_36400), .DIN2(_26833), .Q(_36399) );
  nnd2s1 _36227_inst ( .DIN1(_26833), .DIN2(_36400), .Q(_36397) );
  nnd2s1 _36228_inst ( .DIN1(_36401), .DIN2(_36402), .Q(_36392) );
  xnr2s1 _36229_inst ( .DIN1(_52835), .DIN2(_36403), .Q(_36402) );
  nor2s1 _36230_inst ( .DIN1(_27476), .DIN2(_36404), .Q(_36389) );
  xor2s1 _36231_inst ( .DIN1(_26381), .DIN2(_36405), .Q(_36404) );
  hi1s1 _36232_inst ( .DIN(_27480), .Q(_36405) );
  nnd2s1 _36233_inst ( .DIN1(_36406), .DIN2(_27644), .Q(
        _____________________________195________) );
  or2s1 _36234_inst ( .DIN1(_36407), .DIN2(_27655), .Q(_27644) );
  nor2s1 _36235_inst ( .DIN1(_36408), .DIN2(_36409), .Q(_36406) );
  nor2s1 _36236_inst ( .DIN1(_27648), .DIN2(_36410), .Q(_36409) );
  nnd2s1 _36237_inst ( .DIN1(_36411), .DIN2(_36412), .Q(_36410) );
  nnd2s1 _36238_inst ( .DIN1(_36395), .DIN2(_36413), .Q(_36412) );
  xor2s1 _36239_inst ( .DIN1(_36400), .DIN2(_36414), .Q(_36413) );
  xor2s1 _36240_inst ( .DIN1(_26268), .DIN2(_26833), .Q(_36414) );
  xnr2s1 _36241_inst ( .DIN1(_36415), .DIN2(_32762), .Q(_36400) );
  nnd2s1 _36242_inst ( .DIN1(_36416), .DIN2(_36417), .Q(_36415) );
  nnd2s1 _36243_inst ( .DIN1(_53218), .DIN2(_33504), .Q(_36417) );
  nnd2s1 _36244_inst ( .DIN1(_36418), .DIN2(_53222), .Q(_36416) );
  nor2s1 _36245_inst ( .DIN1(_36419), .DIN2(_33534), .Q(_36418) );
  nor2s1 _36246_inst ( .DIN1(_53218), .DIN2(_33504), .Q(_36419) );
  nnd2s1 _36247_inst ( .DIN1(_36401), .DIN2(_36420), .Q(_36411) );
  xor2s1 _36248_inst ( .DIN1(_26386), .DIN2(_36403), .Q(_36420) );
  nnd2s1 _36249_inst ( .DIN1(_53356), .DIN2(_53170), .Q(_36403) );
  nor2s1 _36250_inst ( .DIN1(_27655), .DIN2(_36421), .Q(_36408) );
  nor2s1 _36251_inst ( .DIN1(_26335), .DIN2(_28100), .Q(_36421) );
  nnd2s1 _36252_inst ( .DIN1(_36422), .DIN2(_36423), .Q(
        _____________________________194________) );
  nnd2s1 _36253_inst ( .DIN1(_36424), .DIN2(_36425), .Q(_36423) );
  nnd2s1 _36254_inst ( .DIN1(_36426), .DIN2(_36427), .Q(_36424) );
  xor2s1 _36255_inst ( .DIN1(_35013), .DIN2(_53101), .Q(_36427) );
  nnd2s1 _36256_inst ( .DIN1(_53172), .DIN2(_53171), .Q(_35013) );
  nor2s1 _36257_inst ( .DIN1(_36386), .DIN2(_27393), .Q(_36426) );
  nor2s1 _36258_inst ( .DIN1(_36428), .DIN2(_36429), .Q(_36422) );
  nor2s1 _36259_inst ( .DIN1(_36365), .DIN2(_36430), .Q(_36429) );
  xnr2s1 _36260_inst ( .DIN1(_33504), .DIN2(_36431), .Q(_36430) );
  xor2s1 _36261_inst ( .DIN1(_26595), .DIN2(_36432), .Q(_36431) );
  nnd2s1 _36262_inst ( .DIN1(_53222), .DIN2(_33517), .Q(_36432) );
  nnd2s1 _36263_inst ( .DIN1(_36395), .DIN2(_35015), .Q(_36365) );
  nor2s1 _36264_inst ( .DIN1(_36433), .DIN2(_36434), .Q(_36428) );
  nnd2s1 _36265_inst ( .DIN1(_36364), .DIN2(_53356), .Q(_36434) );
  hi1s1 _36266_inst ( .DIN(_36359), .Q(_36364) );
  nnd2s1 _36267_inst ( .DIN1(_35015), .DIN2(_36435), .Q(_36359) );
  hi1s1 _36268_inst ( .DIN(_36425), .Q(_35015) );
  nnd2s1 _36269_inst ( .DIN1(_36436), .DIN2(_35300), .Q(_36425) );
  nnd2s1 _36270_inst ( .DIN1(______[20]), .DIN2(_36358), .Q(_36433) );
  nnd2s1 _36271_inst ( .DIN1(_36437), .DIN2(_36438), .Q(
        _____________________________193________) );
  nnd2s1 _36272_inst ( .DIN1(_36439), .DIN2(_30298), .Q(_36438) );
  xor2s1 _36273_inst ( .DIN1(_53173), .DIN2(_26457), .Q(_36439) );
  nnd2s1 _36274_inst ( .DIN1(_27183), .DIN2(_36440), .Q(_36437) );
  nnd2s1 _36275_inst ( .DIN1(_36441), .DIN2(_36442), .Q(_36440) );
  nnd2s1 _36276_inst ( .DIN1(_36401), .DIN2(_36443), .Q(_36442) );
  xor2s1 _36277_inst ( .DIN1(_53170), .DIN2(_53356), .Q(_36443) );
  xor2s1 _36278_inst ( .DIN1(_36444), .DIN2(_36445), .Q(_36401) );
  nnd2s1 _36279_inst ( .DIN1(_36435), .DIN2(_36358), .Q(_36444) );
  nnd2s1 _36280_inst ( .DIN1(_35099), .DIN2(_36446), .Q(_36358) );
  and2s1 _36281_inst ( .DIN1(_36207), .DIN2(_36065), .Q(_36446) );
  nor2s1 _36282_inst ( .DIN1(_35256), .DIN2(_36228), .Q(_35099) );
  nnd2s1 _36283_inst ( .DIN1(_36447), .DIN2(_36395), .Q(_36441) );
  hi1s1 _36284_inst ( .DIN(_36435), .Q(_36395) );
  nnd2s1 _36285_inst ( .DIN1(_36448), .DIN2(_36449), .Q(_36435) );
  nor2s1 _36286_inst ( .DIN1(_36208), .DIN2(_36450), .Q(_36449) );
  nnd2s1 _36287_inst ( .DIN1(_36065), .DIN2(_35270), .Q(_36450) );
  nor2s1 _36288_inst ( .DIN1(_36216), .DIN2(_36451), .Q(_36448) );
  or2s1 _36289_inst ( .DIN1(_35931), .DIN2(_35115), .Q(_36451) );
  nnd2s1 _36290_inst ( .DIN1(_36452), .DIN2(_36453), .Q(_36216) );
  nor2s1 _36291_inst ( .DIN1(_35929), .DIN2(_36454), .Q(_36453) );
  nnd2s1 _36292_inst ( .DIN1(_36455), .DIN2(_36202), .Q(_36454) );
  nor2s1 _36293_inst ( .DIN1(_36456), .DIN2(_35256), .Q(_36452) );
  xor2s1 _36294_inst ( .DIN1(_53222), .DIN2(_34172), .Q(_36447) );
  nnd2s1 _36295_inst ( .DIN1(_36457), .DIN2(_30580), .Q(
        _____________________________192________) );
  nor2s1 _36296_inst ( .DIN1(_36458), .DIN2(_36459), .Q(_36457) );
  nor2s1 _36297_inst ( .DIN1(_27967), .DIN2(_36460), .Q(_36459) );
  nnd2s1 _36298_inst ( .DIN1(_36461), .DIN2(_36462), .Q(_36460) );
  nor2s1 _36299_inst ( .DIN1(_36463), .DIN2(_36464), .Q(_36462) );
  nor2s1 _36300_inst ( .DIN1(_26619), .DIN2(_36465), .Q(_36464) );
  nor2s1 _36301_inst ( .DIN1(_36466), .DIN2(_36467), .Q(_36465) );
  nor2s1 _36302_inst ( .DIN1(_33578), .DIN2(_36468), .Q(_36467) );
  nor2s1 _36303_inst ( .DIN1(_36469), .DIN2(_33577), .Q(_36466) );
  nor2s1 _36304_inst ( .DIN1(_53277), .DIN2(_36470), .Q(_36463) );
  nor2s1 _36305_inst ( .DIN1(_36471), .DIN2(_36472), .Q(_36470) );
  nor2s1 _36306_inst ( .DIN1(_33577), .DIN2(_36468), .Q(_36472) );
  nor2s1 _36307_inst ( .DIN1(_36469), .DIN2(_33578), .Q(_36471) );
  hi1s1 _36308_inst ( .DIN(_36468), .Q(_36469) );
  nnd2s1 _36309_inst ( .DIN1(_36473), .DIN2(_36474), .Q(_36468) );
  nnd2s1 _36310_inst ( .DIN1(_36475), .DIN2(_26518), .Q(_36474) );
  nnd2s1 _36311_inst ( .DIN1(_36476), .DIN2(_32914), .Q(_36475) );
  or2s1 _36312_inst ( .DIN1(_36476), .DIN2(_32914), .Q(_36473) );
  xor2s1 _36313_inst ( .DIN1(_28521), .DIN2(_36477), .Q(_36461) );
  nnd2s1 _36314_inst ( .DIN1(_36478), .DIN2(_32920), .Q(_36477) );
  xor2s1 _36315_inst ( .DIN1(_36479), .DIN2(_36480), .Q(_36478) );
  xor2s1 _36316_inst ( .DIN1(_53276), .DIN2(_53277), .Q(_36480) );
  nor2s1 _36317_inst ( .DIN1(_26300), .DIN2(_26619), .Q(_36479) );
  nor2s1 _36318_inst ( .DIN1(_28755), .DIN2(_36481), .Q(_36458) );
  nor2s1 _36319_inst ( .DIN1(_36482), .DIN2(_36483), .Q(_36481) );
  nor2s1 _36320_inst ( .DIN1(_26524), .DIN2(_30598), .Q(_36483) );
  nnd2s1 _36321_inst ( .DIN1(_53174), .DIN2(_53175), .Q(_30598) );
  nor2s1 _36322_inst ( .DIN1(_53174), .DIN2(_36484), .Q(_36482) );
  nor2s1 _36323_inst ( .DIN1(_26295), .DIN2(_26524), .Q(_36484) );
  nnd2s1 _36324_inst ( .DIN1(_36485), .DIN2(_36486), .Q(
        _____________________________191________) );
  nnd2s1 _36325_inst ( .DIN1(_36487), .DIN2(_36488), .Q(_36486) );
  nor2s1 _36326_inst ( .DIN1(_36489), .DIN2(_28405), .Q(_36487) );
  nnd2s1 _36327_inst ( .DIN1(_36490), .DIN2(_36491), .Q(_28405) );
  nor2s1 _36328_inst ( .DIN1(_36492), .DIN2(_36493), .Q(_36491) );
  nor2s1 _36329_inst ( .DIN1(_35997), .DIN2(_28146), .Q(_36490) );
  xor2s1 _36330_inst ( .DIN1(_36476), .DIN2(_36494), .Q(_36489) );
  xor2s1 _36331_inst ( .DIN1(_26518), .DIN2(_32914), .Q(_36494) );
  nnd2s1 _36332_inst ( .DIN1(_35056), .DIN2(_36495), .Q(_32914) );
  nnd2s1 _36333_inst ( .DIN1(_35059), .DIN2(_36496), .Q(_36495) );
  nnd2s1 _36334_inst ( .DIN1(_36497), .DIN2(_36498), .Q(_36476) );
  nnd2s1 _36335_inst ( .DIN1(_53267), .DIN2(_36499), .Q(_36498) );
  nnd2s1 _36336_inst ( .DIN1(_36500), .DIN2(_32945), .Q(_36499) );
  hi1s1 _36337_inst ( .DIN(_36501), .Q(_36500) );
  nnd2s1 _36338_inst ( .DIN1(_36501), .DIN2(_32935), .Q(_36497) );
  nnd2s1 _36339_inst ( .DIN1(_36502), .DIN2(_28146), .Q(_36485) );
  xor2s1 _36340_inst ( .DIN1(_26604), .DIN2(_28413), .Q(_36502) );
  nnd2s1 _36341_inst ( .DIN1(_53177), .DIN2(_53493), .Q(_28413) );
  nnd2s1 _36342_inst ( .DIN1(_36503), .DIN2(_36504), .Q(
        _____________________________190________) );
  nor2s1 _36343_inst ( .DIN1(_36505), .DIN2(_36506), .Q(_36503) );
  nor2s1 _36344_inst ( .DIN1(_35940), .DIN2(_36507), .Q(_36506) );
  nor2s1 _36345_inst ( .DIN1(_36508), .DIN2(_36509), .Q(_36507) );
  nor2s1 _36346_inst ( .DIN1(_26445), .DIN2(_26224), .Q(_36508) );
  nor2s1 _36347_inst ( .DIN1(_36510), .DIN2(_36511), .Q(_36505) );
  nor2s1 _36348_inst ( .DIN1(_36512), .DIN2(_36513), .Q(_36510) );
  xor2s1 _36349_inst ( .DIN1(_36501), .DIN2(_36514), .Q(_36512) );
  xor2s1 _36350_inst ( .DIN1(_53267), .DIN2(_32945), .Q(_36514) );
  hi1s1 _36351_inst ( .DIN(_32935), .Q(_32945) );
  xnr2s1 _36352_inst ( .DIN1(_36496), .DIN2(_35082), .Q(_32935) );
  nnd2s1 _36353_inst ( .DIN1(_36515), .DIN2(_36516), .Q(_36496) );
  nnd2s1 _36354_inst ( .DIN1(_53364), .DIN2(_36517), .Q(_36516) );
  or2s1 _36355_inst ( .DIN1(_36518), .DIN2(_26849), .Q(_36517) );
  nnd2s1 _36356_inst ( .DIN1(_26849), .DIN2(_36518), .Q(_36515) );
  xor2s1 _36357_inst ( .DIN1(_36519), .DIN2(_31888), .Q(_36501) );
  nnd2s1 _36358_inst ( .DIN1(_36520), .DIN2(_36521), .Q(_36519) );
  nnd2s1 _36359_inst ( .DIN1(_53234), .DIN2(_36522), .Q(_36521) );
  or2s1 _36360_inst ( .DIN1(_36523), .DIN2(_32951), .Q(_36522) );
  nnd2s1 _36361_inst ( .DIN1(_32951), .DIN2(_36523), .Q(_36520) );
  nnd2s1 _36362_inst ( .DIN1(_36524), .DIN2(_31861), .Q(
        _____________________________18________) );
  nor2s1 _36363_inst ( .DIN1(_36525), .DIN2(_36526), .Q(_36524) );
  nor2s1 _36364_inst ( .DIN1(_31864), .DIN2(_36527), .Q(_36526) );
  nnd2s1 _36365_inst ( .DIN1(_36528), .DIN2(_36529), .Q(_36527) );
  nnd2s1 _36366_inst ( .DIN1(_36530), .DIN2(_36531), .Q(_36529) );
  xor2s1 _36367_inst ( .DIN1(_53228), .DIN2(_53231), .Q(_36531) );
  nnd2s1 _36368_inst ( .DIN1(_36532), .DIN2(_36533), .Q(_36528) );
  nor2s1 _36369_inst ( .DIN1(_36534), .DIN2(_36535), .Q(_36532) );
  nor2s1 _36370_inst ( .DIN1(_36536), .DIN2(_26499), .Q(_36535) );
  xor2s1 _36371_inst ( .DIN1(_36324), .DIN2(_35293), .Q(_36536) );
  nor2s1 _36372_inst ( .DIN1(_53178), .DIN2(_36537), .Q(_36534) );
  xor2s1 _36373_inst ( .DIN1(_36324), .DIN2(_35314), .Q(_36537) );
  hi1s1 _36374_inst ( .DIN(_35293), .Q(_35314) );
  xnr2s1 _36375_inst ( .DIN1(_36333), .DIN2(_26814), .Q(_35293) );
  nnd2s1 _36376_inst ( .DIN1(_36539), .DIN2(_36540), .Q(_36334) );
  nnd2s1 _36377_inst ( .DIN1(_53370), .DIN2(_36541), .Q(_36540) );
  or2s1 _36378_inst ( .DIN1(_36542), .DIN2(_36543), .Q(_36541) );
  nnd2s1 _36379_inst ( .DIN1(_36543), .DIN2(_36542), .Q(_36539) );
  nnd2s1 _36380_inst ( .DIN1(_36544), .DIN2(_36545), .Q(_36324) );
  nnd2s1 _36381_inst ( .DIN1(_53193), .DIN2(_36546), .Q(_36545) );
  or2s1 _36382_inst ( .DIN1(_36547), .DIN2(_35322), .Q(_36546) );
  nnd2s1 _36383_inst ( .DIN1(_35322), .DIN2(_36547), .Q(_36544) );
  nor2s1 _36384_inst ( .DIN1(_31907), .DIN2(_36548), .Q(_36525) );
  xor2s1 _36385_inst ( .DIN1(_36549), .DIN2(_36550), .Q(_36548) );
  nor2s1 _36386_inst ( .DIN1(_53348), .DIN2(_26371), .Q(_36550) );
  xnr2s1 _36387_inst ( .DIN1(_53342), .DIN2(_53179), .Q(_36549) );
  nnd2s1 _36388_inst ( .DIN1(_36551), .DIN2(_30601), .Q(
        _____________________________189________) );
  nnd2s1 _36389_inst ( .DIN1(_36552), .DIN2(_27392), .Q(_30601) );
  nor2s1 _36390_inst ( .DIN1(_36553), .DIN2(_36554), .Q(_36551) );
  nor2s1 _36391_inst ( .DIN1(_27392), .DIN2(_36555), .Q(_36554) );
  nnd2s1 _36392_inst ( .DIN1(_36556), .DIN2(_36557), .Q(_36555) );
  nnd2s1 _36393_inst ( .DIN1(_36558), .DIN2(_36559), .Q(_36557) );
  xor2s1 _36394_inst ( .DIN1(_32973), .DIN2(_36560), .Q(_36559) );
  xor2s1 _36395_inst ( .DIN1(_26292), .DIN2(_36523), .Q(_36560) );
  nnd2s1 _36396_inst ( .DIN1(_36561), .DIN2(_36562), .Q(_36523) );
  nnd2s1 _36397_inst ( .DIN1(_53323), .DIN2(_36563), .Q(_36562) );
  or2s1 _36398_inst ( .DIN1(_36564), .DIN2(_32979), .Q(_36563) );
  nnd2s1 _36399_inst ( .DIN1(_32979), .DIN2(_36564), .Q(_36561) );
  hi1s1 _36400_inst ( .DIN(_32994), .Q(_32979) );
  hi1s1 _36401_inst ( .DIN(_32951), .Q(_32973) );
  xnr2s1 _36402_inst ( .DIN1(_36565), .DIN2(_36518), .Q(_32951) );
  nnd2s1 _36403_inst ( .DIN1(_36566), .DIN2(_36567), .Q(_36518) );
  nnd2s1 _36404_inst ( .DIN1(_36568), .DIN2(_26338), .Q(_36567) );
  or2s1 _36405_inst ( .DIN1(_36569), .DIN2(_26849), .Q(_36568) );
  nnd2s1 _36406_inst ( .DIN1(_26849), .DIN2(_36569), .Q(_36566) );
  nnd2s1 _36407_inst ( .DIN1(_36570), .DIN2(_36571), .Q(_36556) );
  nor2s1 _36408_inst ( .DIN1(_36572), .DIN2(_36573), .Q(_36571) );
  and2s1 _36409_inst ( .DIN1(_53180), .DIN2(_53189), .Q(_36573) );
  nor2s1 _36410_inst ( .DIN1(_53180), .DIN2(_36574), .Q(_36572) );
  nor2s1 _36411_inst ( .DIN1(_36575), .DIN2(_36576), .Q(_36570) );
  nor2s1 _36412_inst ( .DIN1(_53186), .DIN2(_26347), .Q(_36575) );
  nor2s1 _36413_inst ( .DIN1(_27397), .DIN2(_36577), .Q(_36553) );
  nor2s1 _36414_inst ( .DIN1(_27066), .DIN2(_36578), .Q(_36577) );
  xnr2s1 _36415_inst ( .DIN1(_53181), .DIN2(_36579), .Q(_36578) );
  nnd2s1 _36416_inst ( .DIN1(_53182), .DIN2(_53183), .Q(_36579) );
  nnd2s1 _36417_inst ( .DIN1(_36580), .DIN2(_28445), .Q(
        _____________________________188________) );
  nnd2s1 _36418_inst ( .DIN1(_27855), .DIN2(_27845), .Q(_28445) );
  hi1s1 _36419_inst ( .DIN(_27849), .Q(_27855) );
  nnd2s1 _36420_inst ( .DIN1(_34601), .DIN2(_35708), .Q(_27849) );
  and2s1 _36421_inst ( .DIN1(_36581), .DIN2(_36582), .Q(_34601) );
  nor2s1 _36422_inst ( .DIN1(_34399), .DIN2(_36583), .Q(_36582) );
  nor2s1 _36423_inst ( .DIN1(_35700), .DIN2(_34398), .Q(_36581) );
  nnd2s1 _36424_inst ( .DIN1(_36584), .DIN2(_36585), .Q(_34398) );
  nor2s1 _36425_inst ( .DIN1(_36586), .DIN2(_36587), .Q(_36584) );
  nor2s1 _36426_inst ( .DIN1(_36588), .DIN2(_36589), .Q(_36580) );
  nor2s1 _36427_inst ( .DIN1(_27845), .DIN2(_36590), .Q(_36589) );
  nnd2s1 _36428_inst ( .DIN1(_36591), .DIN2(_36592), .Q(_36590) );
  nnd2s1 _36429_inst ( .DIN1(_36593), .DIN2(_36594), .Q(_36592) );
  and2s1 _36430_inst ( .DIN1(______[4]), .DIN2(_53185), .Q(_36593) );
  nnd2s1 _36431_inst ( .DIN1(_36595), .DIN2(_36558), .Q(_36591) );
  xor2s1 _36432_inst ( .DIN1(_26779), .DIN2(_36596), .Q(_36595) );
  xor2s1 _36433_inst ( .DIN1(_26260), .DIN2(_36564), .Q(_36596) );
  nnd2s1 _36434_inst ( .DIN1(_36597), .DIN2(_36598), .Q(_36564) );
  nnd2s1 _36435_inst ( .DIN1(_36599), .DIN2(_26476), .Q(_36598) );
  or2s1 _36436_inst ( .DIN1(_36600), .DIN2(_33000), .Q(_36599) );
  nnd2s1 _36437_inst ( .DIN1(_33000), .DIN2(_36600), .Q(_36597) );
  xor2s1 _36438_inst ( .DIN1(_36569), .DIN2(_36601), .Q(_32994) );
  xor2s1 _36439_inst ( .DIN1(_53362), .DIN2(_53384), .Q(_36601) );
  nnd2s1 _36440_inst ( .DIN1(_36602), .DIN2(_36603), .Q(_36569) );
  nnd2s1 _36441_inst ( .DIN1(_26849), .DIN2(_36604), .Q(_36603) );
  nnd2s1 _36442_inst ( .DIN1(_53361), .DIN2(_36605), .Q(_36604) );
  xor2s1 _36443_inst ( .DIN1(_36606), .DIN2(_36607), .Q(_36605) );
  nnd2s1 _36444_inst ( .DIN1(_36607), .DIN2(_34515), .Q(_36602) );
  nor2s1 _36445_inst ( .DIN1(_53184), .DIN2(_27836), .Q(_36588) );
  hi1s1 _36446_inst ( .DIN(_27845), .Q(_27836) );
  nnd2s1 _36447_inst ( .DIN1(_36608), .DIN2(_36609), .Q(_27845) );
  nor2s1 _36448_inst ( .DIN1(_36583), .DIN2(_36610), .Q(_36609) );
  nnd2s1 _36449_inst ( .DIN1(_36611), .DIN2(_35696), .Q(_36610) );
  nor2s1 _36450_inst ( .DIN1(_36612), .DIN2(_36613), .Q(_36608) );
  nnd2s1 _36451_inst ( .DIN1(_36614), .DIN2(_36615), .Q(
        _____________________________187________) );
  nnd2s1 _36452_inst ( .DIN1(_29206), .DIN2(_36616), .Q(_36615) );
  nnd2s1 _36453_inst ( .DIN1(_36617), .DIN2(_36618), .Q(_36616) );
  nnd2s1 _36454_inst ( .DIN1(_36619), .DIN2(_36594), .Q(_36618) );
  and2s1 _36455_inst ( .DIN1(_53186), .DIN2(______[30]), .Q(_36619) );
  nnd2s1 _36456_inst ( .DIN1(_36558), .DIN2(_36620), .Q(_36617) );
  xor2s1 _36457_inst ( .DIN1(_33000), .DIN2(_36621), .Q(_36620) );
  xor2s1 _36458_inst ( .DIN1(_26476), .DIN2(_36600), .Q(_36621) );
  nnd2s1 _36459_inst ( .DIN1(_36622), .DIN2(_36623), .Q(_36600) );
  nnd2s1 _36460_inst ( .DIN1(_53187), .DIN2(_36624), .Q(_36623) );
  or2s1 _36461_inst ( .DIN1(_36625), .DIN2(_26828), .Q(_36624) );
  nnd2s1 _36462_inst ( .DIN1(_33017), .DIN2(_36625), .Q(_36622) );
  xnr2s1 _36463_inst ( .DIN1(_36626), .DIN2(_36627), .Q(_33000) );
  xor2s1 _36464_inst ( .DIN1(_27956), .DIN2(_36607), .Q(_36627) );
  xor2s1 _36465_inst ( .DIN1(_36628), .DIN2(_35291), .Q(_36607) );
  nnd2s1 _36466_inst ( .DIN1(_36629), .DIN2(_36630), .Q(_36628) );
  nnd2s1 _36467_inst ( .DIN1(_36631), .DIN2(_26335), .Q(_36630) );
  nnd2s1 _36468_inst ( .DIN1(_53365), .DIN2(_36632), .Q(_36631) );
  or2s1 _36469_inst ( .DIN1(_36632), .DIN2(_53365), .Q(_36629) );
  xor2s1 _36470_inst ( .DIN1(_34515), .DIN2(_53384), .Q(_36626) );
  nnd2s1 _36471_inst ( .DIN1(_35029), .DIN2(_52859), .Q(_36614) );
  hi1s1 _36472_inst ( .DIN(_36633), .Q(_35029) );
  nnd2s1 _36473_inst ( .DIN1(_36634), .DIN2(_36635), .Q(
        _____________________________186________) );
  nnd2s1 _36474_inst ( .DIN1(_28010), .DIN2(_36636), .Q(_36635) );
  nnd2s1 _36475_inst ( .DIN1(_36637), .DIN2(_36638), .Q(_36636) );
  nnd2s1 _36476_inst ( .DIN1(_36639), .DIN2(_36594), .Q(_36638) );
  nor2s1 _36477_inst ( .DIN1(_36640), .DIN2(_27291), .Q(_36639) );
  xor2s1 _36478_inst ( .DIN1(_36574), .DIN2(_53180), .Q(_36640) );
  nnd2s1 _36479_inst ( .DIN1(_53186), .DIN2(_26347), .Q(_36574) );
  nnd2s1 _36480_inst ( .DIN1(_36558), .DIN2(_36641), .Q(_36637) );
  xor2s1 _36481_inst ( .DIN1(_33029), .DIN2(_36642), .Q(_36641) );
  xnr2s1 _36482_inst ( .DIN1(_53187), .DIN2(_36625), .Q(_36642) );
  nnd2s1 _36483_inst ( .DIN1(_36643), .DIN2(_36644), .Q(_36625) );
  nnd2s1 _36484_inst ( .DIN1(_36645), .DIN2(_26656), .Q(_36644) );
  or2s1 _36485_inst ( .DIN1(_36646), .DIN2(_33035), .Q(_36645) );
  nnd2s1 _36486_inst ( .DIN1(_33035), .DIN2(_36646), .Q(_36643) );
  hi1s1 _36487_inst ( .DIN(_33017), .Q(_33029) );
  xor2s1 _36488_inst ( .DIN1(_36632), .DIN2(_36647), .Q(_33017) );
  xor2s1 _36489_inst ( .DIN1(_53363), .DIN2(_53365), .Q(_36647) );
  nnd2s1 _36490_inst ( .DIN1(_36648), .DIN2(_36649), .Q(_36632) );
  nnd2s1 _36491_inst ( .DIN1(_53364), .DIN2(_36650), .Q(_36649) );
  or2s1 _36492_inst ( .DIN1(_36651), .DIN2(_26781), .Q(_36650) );
  nnd2s1 _36493_inst ( .DIN1(_26781), .DIN2(_36651), .Q(_36648) );
  nnd2s1 _36494_inst ( .DIN1(_36652), .DIN2(_36653), .Q(_36634) );
  xor2s1 _36495_inst ( .DIN1(_26434), .DIN2(_53523), .Q(_36653) );
  nor2s1 _36496_inst ( .DIN1(_36654), .DIN2(_28646), .Q(_36652) );
  nor2s1 _36497_inst ( .DIN1(_35342), .DIN2(_28178), .Q(_36654) );
  nnd2s1 _36498_inst ( .DIN1(_36655), .DIN2(_36656), .Q(
        _____________________________185________) );
  nnd2s1 _36499_inst ( .DIN1(_31907), .DIN2(_36657), .Q(_36656) );
  nnd2s1 _36500_inst ( .DIN1(_36658), .DIN2(_36659), .Q(_36657) );
  nnd2s1 _36501_inst ( .DIN1(_36594), .DIN2(_36660), .Q(_36659) );
  xor2s1 _36502_inst ( .DIN1(_53191), .DIN2(_53232), .Q(_36660) );
  hi1s1 _36503_inst ( .DIN(_36576), .Q(_36594) );
  nnd2s1 _36504_inst ( .DIN1(_36661), .DIN2(_36662), .Q(_36576) );
  nnd2s1 _36505_inst ( .DIN1(_36663), .DIN2(_36558), .Q(_36658) );
  xor2s1 _36506_inst ( .DIN1(_33035), .DIN2(_36664), .Q(_36663) );
  xor2s1 _36507_inst ( .DIN1(_26656), .DIN2(_36646), .Q(_36664) );
  nnd2s1 _36508_inst ( .DIN1(_36665), .DIN2(_36666), .Q(_36646) );
  nnd2s1 _36509_inst ( .DIN1(_53301), .DIN2(_36667), .Q(_36666) );
  or2s1 _36510_inst ( .DIN1(_36668), .DIN2(_26800), .Q(_36667) );
  nnd2s1 _36511_inst ( .DIN1(_33065), .DIN2(_36668), .Q(_36665) );
  xnr2s1 _36512_inst ( .DIN1(_36669), .DIN2(_36651), .Q(_33035) );
  nnd2s1 _36513_inst ( .DIN1(_36670), .DIN2(_36671), .Q(_36651) );
  nnd2s1 _36514_inst ( .DIN1(_36672), .DIN2(_26338), .Q(_36671) );
  or2s1 _36515_inst ( .DIN1(_36673), .DIN2(_53367), .Q(_36672) );
  nnd2s1 _36516_inst ( .DIN1(_53367), .DIN2(_36673), .Q(_36670) );
  xor2s1 _36517_inst ( .DIN1(_27620), .DIN2(_53368), .Q(_36669) );
  nnd2s1 _36518_inst ( .DIN1(_36674), .DIN2(_31864), .Q(_36655) );
  nor2s1 _36519_inst ( .DIN1(_36675), .DIN2(_26371), .Q(_36674) );
  and2s1 _36520_inst ( .DIN1(_33683), .DIN2(_36676), .Q(_36675) );
  nnd2s1 _36521_inst ( .DIN1(_36677), .DIN2(_36678), .Q(
        _____________________________184________) );
  nor2s1 _36522_inst ( .DIN1(_36679), .DIN2(_36680), .Q(_36677) );
  nor2s1 _36523_inst ( .DIN1(_36681), .DIN2(_36682), .Q(_36680) );
  xor2s1 _36524_inst ( .DIN1(_30081), .DIN2(_36683), .Q(_36682) );
  nnd2s1 _36525_inst ( .DIN1(_36684), .DIN2(_36685), .Q(_36683) );
  nnd2s1 _36526_inst ( .DIN1(_36686), .DIN2(_36661), .Q(_36685) );
  nnd2s1 _36527_inst ( .DIN1(_36687), .DIN2(______[4]), .Q(_36686) );
  nor2s1 _36528_inst ( .DIN1(_36688), .DIN2(_36689), .Q(_36687) );
  xnr2s1 _36529_inst ( .DIN1(_53342), .DIN2(_36690), .Q(_36689) );
  nor2s1 _36530_inst ( .DIN1(_53270), .DIN2(_26458), .Q(_36690) );
  nnd2s1 _36531_inst ( .DIN1(_36691), .DIN2(_36558), .Q(_36684) );
  hi1s1 _36532_inst ( .DIN(_36661), .Q(_36558) );
  nnd2s1 _36533_inst ( .DIN1(_36692), .DIN2(_36693), .Q(_36661) );
  nor2s1 _36534_inst ( .DIN1(_36694), .DIN2(_36695), .Q(_36692) );
  xor2s1 _36535_inst ( .DIN1(_33065), .DIN2(_36696), .Q(_36691) );
  xnr2s1 _36536_inst ( .DIN1(_53301), .DIN2(_36668), .Q(_36696) );
  nnd2s1 _36537_inst ( .DIN1(_36697), .DIN2(_36698), .Q(_36668) );
  nnd2s1 _36538_inst ( .DIN1(_53190), .DIN2(_36699), .Q(_36698) );
  or2s1 _36539_inst ( .DIN1(_36700), .DIN2(_33088), .Q(_36699) );
  nnd2s1 _36540_inst ( .DIN1(_33088), .DIN2(_36700), .Q(_36697) );
  xor2s1 _36541_inst ( .DIN1(_36701), .DIN2(_36702), .Q(_33065) );
  xor2s1 _36542_inst ( .DIN1(_53362), .DIN2(_53367), .Q(_36702) );
  xnr2s1 _36543_inst ( .DIN1(_36673), .DIN2(_34151), .Q(_36701) );
  nnd2s1 _36544_inst ( .DIN1(_36703), .DIN2(_36704), .Q(_36673) );
  nnd2s1 _36545_inst ( .DIN1(_53309), .DIN2(_36705), .Q(_36704) );
  or2s1 _36546_inst ( .DIN1(_36706), .DIN2(_34515), .Q(_36705) );
  nnd2s1 _36547_inst ( .DIN1(_36706), .DIN2(_34515), .Q(_36703) );
  nor2s1 _36548_inst ( .DIN1(_33292), .DIN2(_36707), .Q(_36679) );
  nor2s1 _36549_inst ( .DIN1(_27039), .DIN2(_26385), .Q(_36707) );
  nnd2s1 _36550_inst ( .DIN1(_36708), .DIN2(_36709), .Q(
        _____________________________183________) );
  nnd2s1 _36551_inst ( .DIN1(_36710), .DIN2(_36711), .Q(_36709) );
  xor2s1 _36552_inst ( .DIN1(_33088), .DIN2(_36712), .Q(_36711) );
  xnr2s1 _36553_inst ( .DIN1(_53190), .DIN2(_36700), .Q(_36712) );
  nnd2s1 _36554_inst ( .DIN1(_36713), .DIN2(_36714), .Q(_36700) );
  nnd2s1 _36555_inst ( .DIN1(_36715), .DIN2(_26557), .Q(_36714) );
  or2s1 _36556_inst ( .DIN1(_36716), .DIN2(_33108), .Q(_36715) );
  nnd2s1 _36557_inst ( .DIN1(_33108), .DIN2(_36716), .Q(_36713) );
  hi1s1 _36558_inst ( .DIN(_33103), .Q(_33088) );
  xnr2s1 _36559_inst ( .DIN1(_36717), .DIN2(_36706), .Q(_33103) );
  nnd2s1 _36560_inst ( .DIN1(_36718), .DIN2(_36719), .Q(_36706) );
  nnd2s1 _36561_inst ( .DIN1(_53314), .DIN2(_36720), .Q(_36719) );
  or2s1 _36562_inst ( .DIN1(_36721), .DIN2(_53365), .Q(_36720) );
  nnd2s1 _36563_inst ( .DIN1(_53365), .DIN2(_36721), .Q(_36718) );
  xor2s1 _36564_inst ( .DIN1(_26526), .DIN2(_53361), .Q(_36717) );
  hi1s1 _36565_inst ( .DIN(_36722), .Q(_36710) );
  nor2s1 _36566_inst ( .DIN1(_36723), .DIN2(_36724), .Q(_36708) );
  nor2s1 _36567_inst ( .DIN1(_36725), .DIN2(_36726), .Q(_36724) );
  nor2s1 _36568_inst ( .DIN1(_36688), .DIN2(_53270), .Q(_36725) );
  nor2s1 _36569_inst ( .DIN1(_36727), .DIN2(_36728), .Q(_36723) );
  nnd2s1 _36570_inst ( .DIN1(______[18]), .DIN2(_36729), .Q(_36728) );
  xor2s1 _36571_inst ( .DIN1(_53269), .DIN2(_53270), .Q(_36729) );
  nnd2s1 _36572_inst ( .DIN1(_36730), .DIN2(_28026), .Q(
        _____________________________182________) );
  nor2s1 _36573_inst ( .DIN1(_36731), .DIN2(_36732), .Q(_36730) );
  nor2s1 _36574_inst ( .DIN1(_28016), .DIN2(_36733), .Q(_36732) );
  nor2s1 _36575_inst ( .DIN1(_36734), .DIN2(_36735), .Q(_36733) );
  nor2s1 _36576_inst ( .DIN1(_36736), .DIN2(_36737), .Q(_36735) );
  xor2s1 _36577_inst ( .DIN1(_33108), .DIN2(_36738), .Q(_36737) );
  xor2s1 _36578_inst ( .DIN1(_26557), .DIN2(_36716), .Q(_36738) );
  nnd2s1 _36579_inst ( .DIN1(_36739), .DIN2(_36740), .Q(_36716) );
  nnd2s1 _36580_inst ( .DIN1(_53240), .DIN2(_36741), .Q(_36740) );
  or2s1 _36581_inst ( .DIN1(_36742), .DIN2(_33129), .Q(_36741) );
  nnd2s1 _36582_inst ( .DIN1(_33129), .DIN2(_36742), .Q(_36739) );
  hi1s1 _36583_inst ( .DIN(_33141), .Q(_33129) );
  xor2s1 _36584_inst ( .DIN1(_36721), .DIN2(_36743), .Q(_33108) );
  xor2s1 _36585_inst ( .DIN1(_53314), .DIN2(_53365), .Q(_36743) );
  nnd2s1 _36586_inst ( .DIN1(_36744), .DIN2(_36745), .Q(_36721) );
  nnd2s1 _36587_inst ( .DIN1(_26781), .DIN2(_36746), .Q(_36745) );
  or2s1 _36588_inst ( .DIN1(_36747), .DIN2(_53371), .Q(_36746) );
  nnd2s1 _36589_inst ( .DIN1(_53371), .DIN2(_36747), .Q(_36744) );
  nor2s1 _36590_inst ( .DIN1(_36748), .DIN2(_36749), .Q(_36734) );
  nor2s1 _36591_inst ( .DIN1(_36688), .DIN2(_36750), .Q(_36749) );
  xor2s1 _36592_inst ( .DIN1(_53342), .DIN2(_26458), .Q(_36750) );
  nor2s1 _36593_inst ( .DIN1(_53231), .DIN2(_28024), .Q(_36731) );
  nnd2s1 _36594_inst ( .DIN1(_36751), .DIN2(_36752), .Q(
        _____________________________181________) );
  nnd2s1 _36595_inst ( .DIN1(_36753), .DIN2(_36754), .Q(_36752) );
  nnd2s1 _36596_inst ( .DIN1(_36755), .DIN2(_36662), .Q(_36754) );
  xor2s1 _36597_inst ( .DIN1(_36756), .DIN2(_36757), .Q(_36755) );
  nnd2s1 _36598_inst ( .DIN1(_36758), .DIN2(______[0]), .Q(_36756) );
  xor2s1 _36599_inst ( .DIN1(_26381), .DIN2(_36759), .Q(_36758) );
  nor2s1 _36600_inst ( .DIN1(_53201), .DIN2(_26261), .Q(_36759) );
  nor2s1 _36601_inst ( .DIN1(_36760), .DIN2(_36761), .Q(_36751) );
  nor2s1 _36602_inst ( .DIN1(_36762), .DIN2(_36722), .Q(_36761) );
  xor2s1 _36603_inst ( .DIN1(_33141), .DIN2(_36763), .Q(_36762) );
  xnr2s1 _36604_inst ( .DIN1(_53240), .DIN2(_36742), .Q(_36763) );
  nnd2s1 _36605_inst ( .DIN1(_36764), .DIN2(_36765), .Q(_36742) );
  nnd2s1 _36606_inst ( .DIN1(_36766), .DIN2(_26676), .Q(_36765) );
  or2s1 _36607_inst ( .DIN1(_36767), .DIN2(_26832), .Q(_36766) );
  nnd2s1 _36608_inst ( .DIN1(_33147), .DIN2(_36767), .Q(_36764) );
  xor2s1 _36609_inst ( .DIN1(_36768), .DIN2(_36769), .Q(_33141) );
  xor2s1 _36610_inst ( .DIN1(_31947), .DIN2(_36747), .Q(_36769) );
  nnd2s1 _36611_inst ( .DIN1(_36770), .DIN2(_36771), .Q(_36747) );
  nnd2s1 _36612_inst ( .DIN1(_53367), .DIN2(_36772), .Q(_36771) );
  or2s1 _36613_inst ( .DIN1(_36773), .DIN2(_53370), .Q(_36772) );
  nnd2s1 _36614_inst ( .DIN1(_53370), .DIN2(_36773), .Q(_36770) );
  xor2s1 _36615_inst ( .DIN1(_36332), .DIN2(_53368), .Q(_36768) );
  nor2s1 _36616_inst ( .DIN1(_36727), .DIN2(_36774), .Q(_36760) );
  nnd2s1 _36617_inst ( .DIN1(_36775), .DIN2(______[24]), .Q(_36774) );
  xor2s1 _36618_inst ( .DIN1(_36776), .DIN2(_53205), .Q(_36775) );
  nnd2s1 _36619_inst ( .DIN1(_36681), .DIN2(_36777), .Q(_36727) );
  nnd2s1 _36620_inst ( .DIN1(_36778), .DIN2(_30580), .Q(
        _____________________________180________) );
  nnd2s1 _36621_inst ( .DIN1(_30992), .DIN2(_27967), .Q(_30580) );
  nor2s1 _36622_inst ( .DIN1(_36779), .DIN2(_36780), .Q(_36778) );
  nor2s1 _36623_inst ( .DIN1(_27967), .DIN2(_36781), .Q(_36780) );
  nnd2s1 _36624_inst ( .DIN1(_36782), .DIN2(_36783), .Q(_36781) );
  nnd2s1 _36625_inst ( .DIN1(_36784), .DIN2(_36785), .Q(_36783) );
  nor2s1 _36626_inst ( .DIN1(_36748), .DIN2(_36688), .Q(_36785) );
  nor2s1 _36627_inst ( .DIN1(_27774), .DIN2(_36786), .Q(_36784) );
  xor2s1 _36628_inst ( .DIN1(_53198), .DIN2(_53201), .Q(_36786) );
  xor2s1 _36629_inst ( .DIN1(_34338), .DIN2(_36787), .Q(_36782) );
  nnd2s1 _36630_inst ( .DIN1(_36788), .DIN2(_36748), .Q(_36787) );
  xor2s1 _36631_inst ( .DIN1(_33147), .DIN2(_36789), .Q(_36788) );
  xor2s1 _36632_inst ( .DIN1(_26676), .DIN2(_36767), .Q(_36789) );
  nnd2s1 _36633_inst ( .DIN1(_36790), .DIN2(_36791), .Q(_36767) );
  nnd2s1 _36634_inst ( .DIN1(_53197), .DIN2(_36792), .Q(_36791) );
  or2s1 _36635_inst ( .DIN1(_36793), .DIN2(_33178), .Q(_36792) );
  nnd2s1 _36636_inst ( .DIN1(_33178), .DIN2(_36793), .Q(_36790) );
  xor2s1 _36637_inst ( .DIN1(_36773), .DIN2(_36794), .Q(_33147) );
  xor2s1 _36638_inst ( .DIN1(_53367), .DIN2(_53370), .Q(_36794) );
  nnd2s1 _36639_inst ( .DIN1(_36795), .DIN2(_36796), .Q(_36773) );
  nnd2s1 _36640_inst ( .DIN1(_53309), .DIN2(_36797), .Q(_36796) );
  or2s1 _36641_inst ( .DIN1(_36798), .DIN2(_53517), .Q(_36797) );
  nnd2s1 _36642_inst ( .DIN1(_53517), .DIN2(_36798), .Q(_36795) );
  nor2s1 _36643_inst ( .DIN1(_53192), .DIN2(_28755), .Q(_36779) );
  nnd2s1 _36644_inst ( .DIN1(_36799), .DIN2(_36800), .Q(
        _____________________________17________) );
  nnd2s1 _36645_inst ( .DIN1(_34301), .DIN2(_36801), .Q(_36800) );
  nnd2s1 _36646_inst ( .DIN1(_36802), .DIN2(_36803), .Q(_36801) );
  nnd2s1 _36647_inst ( .DIN1(_36804), .DIN2(_36805), .Q(_36803) );
  nnd2s1 _36648_inst ( .DIN1(______[6]), .DIN2(_36806), .Q(_36805) );
  xor2s1 _36649_inst ( .DIN1(_26371), .DIN2(_36807), .Q(_36806) );
  nnd2s1 _36650_inst ( .DIN1(_53228), .DIN2(_26379), .Q(_36807) );
  nor2s1 _36651_inst ( .DIN1(_36808), .DIN2(_36809), .Q(_36802) );
  nor2s1 _36652_inst ( .DIN1(_36810), .DIN2(_36811), .Q(_36809) );
  xor2s1 _36653_inst ( .DIN1(_35322), .DIN2(_36812), .Q(_36811) );
  xor2s1 _36654_inst ( .DIN1(_53193), .DIN2(_36547), .Q(_36812) );
  nnd2s1 _36655_inst ( .DIN1(_36813), .DIN2(_36814), .Q(_36547) );
  nnd2s1 _36656_inst ( .DIN1(_36815), .DIN2(_26534), .Q(_36814) );
  or2s1 _36657_inst ( .DIN1(_36816), .DIN2(_35338), .Q(_36815) );
  nnd2s1 _36658_inst ( .DIN1(_35338), .DIN2(_36816), .Q(_36813) );
  xnr2s1 _36659_inst ( .DIN1(_36543), .DIN2(_36817), .Q(_35322) );
  xor2s1 _36660_inst ( .DIN1(_26778), .DIN2(_36542), .Q(_36817) );
  nnd2s1 _36661_inst ( .DIN1(_36818), .DIN2(_36819), .Q(_36542) );
  nnd2s1 _36662_inst ( .DIN1(_53517), .DIN2(_36820), .Q(_36819) );
  or2s1 _36663_inst ( .DIN1(_36821), .DIN2(_36822), .Q(_36820) );
  nnd2s1 _36664_inst ( .DIN1(_36822), .DIN2(_36821), .Q(_36818) );
  hi1s1 _36665_inst ( .DIN(_34298), .Q(_34301) );
  nnd2s1 _36666_inst ( .DIN1(_36823), .DIN2(_33808), .Q(_34298) );
  hi1s1 _36667_inst ( .DIN(_33898), .Q(_33808) );
  nnd2s1 _36668_inst ( .DIN1(_36824), .DIN2(_36825), .Q(_33898) );
  nor2s1 _36669_inst ( .DIN1(_36826), .DIN2(_36827), .Q(_36825) );
  nor2s1 _36670_inst ( .DIN1(_36828), .DIN2(_33295), .Q(_36824) );
  nor2s1 _36671_inst ( .DIN1(_27821), .DIN2(_36829), .Q(_36823) );
  nnd2s1 _36672_inst ( .DIN1(_36830), .DIN2(_35614), .Q(_36799) );
  nnd2s1 _36673_inst ( .DIN1(_36831), .DIN2(_36832), .Q(_35614) );
  nor2s1 _36674_inst ( .DIN1(_36833), .DIN2(_36828), .Q(_36831) );
  xor2s1 _36675_inst ( .DIN1(_26404), .DIN2(_35612), .Q(_36830) );
  nnd2s1 _36676_inst ( .DIN1(_53195), .DIN2(_53196), .Q(_35612) );
  nnd2s1 _36677_inst ( .DIN1(_36834), .DIN2(_36835), .Q(
        _____________________________179________) );
  nor2s1 _36678_inst ( .DIN1(_36836), .DIN2(_36837), .Q(_36835) );
  nor2s1 _36679_inst ( .DIN1(_36838), .DIN2(_36839), .Q(_36837) );
  nnd2s1 _36680_inst ( .DIN1(_36753), .DIN2(_53150), .Q(_36839) );
  hi1s1 _36681_inst ( .DIN(_36726), .Q(_36753) );
  nnd2s1 _36682_inst ( .DIN1(_33292), .DIN2(_36736), .Q(_36726) );
  nnd2s1 _36683_inst ( .DIN1(______[30]), .DIN2(_36662), .Q(_36838) );
  hi1s1 _36684_inst ( .DIN(_36678), .Q(_36836) );
  nor2s1 _36685_inst ( .DIN1(_36840), .DIN2(_36841), .Q(_36834) );
  nor2s1 _36686_inst ( .DIN1(_33292), .DIN2(_36842), .Q(_36841) );
  nor2s1 _36687_inst ( .DIN1(_28684), .DIN2(_36843), .Q(_36842) );
  xor2s1 _36688_inst ( .DIN1(_26489), .DIN2(_36776), .Q(_36843) );
  nor2s1 _36689_inst ( .DIN1(_36722), .DIN2(_36844), .Q(_36840) );
  xor2s1 _36690_inst ( .DIN1(_33178), .DIN2(_36845), .Q(_36844) );
  xor2s1 _36691_inst ( .DIN1(_26734), .DIN2(_36793), .Q(_36845) );
  nnd2s1 _36692_inst ( .DIN1(_36846), .DIN2(_36847), .Q(_36793) );
  nnd2s1 _36693_inst ( .DIN1(_36848), .DIN2(_26649), .Q(_36847) );
  or2s1 _36694_inst ( .DIN1(_36849), .DIN2(_33196), .Q(_36848) );
  nnd2s1 _36695_inst ( .DIN1(_33196), .DIN2(_36849), .Q(_36846) );
  hi1s1 _36696_inst ( .DIN(_33190), .Q(_33178) );
  xor2s1 _36697_inst ( .DIN1(_36850), .DIN2(_36798), .Q(_33190) );
  xnr2s1 _36698_inst ( .DIN1(_36851), .DIN2(_31802), .Q(_36798) );
  nnd2s1 _36699_inst ( .DIN1(_36852), .DIN2(_36853), .Q(_36851) );
  nnd2s1 _36700_inst ( .DIN1(_53314), .DIN2(_36854), .Q(_36853) );
  or2s1 _36701_inst ( .DIN1(_36855), .DIN2(_27731), .Q(_36854) );
  nnd2s1 _36702_inst ( .DIN1(_36855), .DIN2(_27731), .Q(_36852) );
  xor2s1 _36703_inst ( .DIN1(_26526), .DIN2(_53517), .Q(_36850) );
  nnd2s1 _36704_inst ( .DIN1(_33292), .DIN2(_36748), .Q(_36722) );
  nnd2s1 _36705_inst ( .DIN1(_36856), .DIN2(_36857), .Q(
        _____________________________178________) );
  nnd2s1 _36706_inst ( .DIN1(_36858), .DIN2(_27476), .Q(_36857) );
  nor2s1 _36707_inst ( .DIN1(_36859), .DIN2(_36860), .Q(_36858) );
  nor2s1 _36708_inst ( .DIN1(_36736), .DIN2(_36861), .Q(_36860) );
  xor2s1 _36709_inst ( .DIN1(_33196), .DIN2(_36862), .Q(_36861) );
  xor2s1 _36710_inst ( .DIN1(_26649), .DIN2(_36849), .Q(_36862) );
  nnd2s1 _36711_inst ( .DIN1(_36863), .DIN2(_36864), .Q(_36849) );
  nnd2s1 _36712_inst ( .DIN1(_53251), .DIN2(_36865), .Q(_36864) );
  or2s1 _36713_inst ( .DIN1(_36866), .DIN2(_33213), .Q(_36865) );
  nnd2s1 _36714_inst ( .DIN1(_33213), .DIN2(_36866), .Q(_36863) );
  hi1s1 _36715_inst ( .DIN(_33882), .Q(_33196) );
  xor2s1 _36716_inst ( .DIN1(_36855), .DIN2(_36867), .Q(_33882) );
  xor2s1 _36717_inst ( .DIN1(_53314), .DIN2(_53375), .Q(_36867) );
  nnd2s1 _36718_inst ( .DIN1(_36868), .DIN2(_36869), .Q(_36855) );
  nnd2s1 _36719_inst ( .DIN1(_53371), .DIN2(_36870), .Q(_36869) );
  or2s1 _36720_inst ( .DIN1(_36871), .DIN2(_53373), .Q(_36870) );
  nnd2s1 _36721_inst ( .DIN1(_53373), .DIN2(_36871), .Q(_36868) );
  nor2s1 _36722_inst ( .DIN1(_36748), .DIN2(_36872), .Q(_36859) );
  nor2s1 _36723_inst ( .DIN1(_36873), .DIN2(_36874), .Q(_36872) );
  nnd2s1 _36724_inst ( .DIN1(______[26]), .DIN2(_36662), .Q(_36874) );
  xor2s1 _36725_inst ( .DIN1(_53150), .DIN2(_53201), .Q(_36873) );
  nnd2s1 _36726_inst ( .DIN1(_36875), .DIN2(_36876), .Q(_36856) );
  xor2s1 _36727_inst ( .DIN1(_53199), .DIN2(_27480), .Q(_36876) );
  nnd2s1 _36728_inst ( .DIN1(_53391), .DIN2(_26587), .Q(_27480) );
  and2s1 _36729_inst ( .DIN1(______[4]), .DIN2(_29658), .Q(_36875) );
  nnd2s1 _36730_inst ( .DIN1(_36877), .DIN2(_36678), .Q(
        _____________________________177________) );
  nor2s1 _36731_inst ( .DIN1(_36878), .DIN2(_36879), .Q(_36877) );
  nor2s1 _36732_inst ( .DIN1(_36681), .DIN2(_36880), .Q(_36879) );
  nnd2s1 _36733_inst ( .DIN1(_36881), .DIN2(_36882), .Q(_36880) );
  nor2s1 _36734_inst ( .DIN1(_36883), .DIN2(_36884), .Q(_36881) );
  nor2s1 _36735_inst ( .DIN1(_36885), .DIN2(_36886), .Q(_36884) );
  xor2s1 _36736_inst ( .DIN1(_36887), .DIN2(_36888), .Q(_36886) );
  xor2s1 _36737_inst ( .DIN1(_36866), .DIN2(_33213), .Q(_36888) );
  xnr2s1 _36738_inst ( .DIN1(_36871), .DIN2(_36889), .Q(_33213) );
  nnd2s1 _36739_inst ( .DIN1(_36890), .DIN2(_36891), .Q(_36871) );
  nnd2s1 _36740_inst ( .DIN1(_53370), .DIN2(_36892), .Q(_36891) );
  or2s1 _36741_inst ( .DIN1(_36893), .DIN2(_53374), .Q(_36892) );
  nnd2s1 _36742_inst ( .DIN1(_53374), .DIN2(_36893), .Q(_36890) );
  nnd2s1 _36743_inst ( .DIN1(_36894), .DIN2(_36895), .Q(_36866) );
  nnd2s1 _36744_inst ( .DIN1(_53246), .DIN2(_36896), .Q(_36895) );
  or2s1 _36745_inst ( .DIN1(_36897), .DIN2(_33907), .Q(_36896) );
  nnd2s1 _36746_inst ( .DIN1(_33907), .DIN2(_36897), .Q(_36894) );
  xor2s1 _36747_inst ( .DIN1(_53251), .DIN2(_31925), .Q(_36887) );
  nnd2s1 _36748_inst ( .DIN1(_32762), .DIN2(_36898), .Q(_31925) );
  nor2s1 _36749_inst ( .DIN1(_36899), .DIN2(_36900), .Q(_36883) );
  nor2s1 _36750_inst ( .DIN1(_28100), .DIN2(_36901), .Q(_36900) );
  xor2s1 _36751_inst ( .DIN1(_36902), .DIN2(_36903), .Q(_36901) );
  xor2s1 _36752_inst ( .DIN1(_53200), .DIN2(_53205), .Q(_36903) );
  nor2s1 _36753_inst ( .DIN1(_53202), .DIN2(_26606), .Q(_36902) );
  nor2s1 _36754_inst ( .DIN1(_53201), .DIN2(_33292), .Q(_36878) );
  nnd2s1 _36755_inst ( .DIN1(_36904), .DIN2(_36678), .Q(
        _____________________________176________) );
  nnd2s1 _36756_inst ( .DIN1(_32834), .DIN2(_36681), .Q(_36678) );
  nor2s1 _36757_inst ( .DIN1(_36905), .DIN2(_36906), .Q(_36904) );
  nor2s1 _36758_inst ( .DIN1(_36681), .DIN2(_36907), .Q(_36906) );
  nnd2s1 _36759_inst ( .DIN1(_36908), .DIN2(_36882), .Q(_36907) );
  nor2s1 _36760_inst ( .DIN1(_36909), .DIN2(_36910), .Q(_36908) );
  nor2s1 _36761_inst ( .DIN1(_36885), .DIN2(_36911), .Q(_36910) );
  xor2s1 _36762_inst ( .DIN1(_33225), .DIN2(_36912), .Q(_36911) );
  xor2s1 _36763_inst ( .DIN1(_26549), .DIN2(_36897), .Q(_36912) );
  nnd2s1 _36764_inst ( .DIN1(_36913), .DIN2(_36914), .Q(_36897) );
  nnd2s1 _36765_inst ( .DIN1(_36915), .DIN2(_26342), .Q(_36914) );
  or2s1 _36766_inst ( .DIN1(_36916), .DIN2(_26834), .Q(_36915) );
  nnd2s1 _36767_inst ( .DIN1(_26834), .DIN2(_36916), .Q(_36913) );
  hi1s1 _36768_inst ( .DIN(_33907), .Q(_33225) );
  xor2s1 _36769_inst ( .DIN1(_36893), .DIN2(_36917), .Q(_33907) );
  xor2s1 _36770_inst ( .DIN1(_53370), .DIN2(_53374), .Q(_36917) );
  nnd2s1 _36771_inst ( .DIN1(_36918), .DIN2(_36919), .Q(_36893) );
  nnd2s1 _36772_inst ( .DIN1(_53372), .DIN2(_36920), .Q(_36919) );
  or2s1 _36773_inst ( .DIN1(_36921), .DIN2(_53517), .Q(_36920) );
  nnd2s1 _36774_inst ( .DIN1(_53517), .DIN2(_36921), .Q(_36918) );
  nor2s1 _36775_inst ( .DIN1(_36899), .DIN2(_36922), .Q(_36909) );
  nor2s1 _36776_inst ( .DIN1(_53202), .DIN2(_28646), .Q(_36922) );
  nor2s1 _36777_inst ( .DIN1(_33292), .DIN2(_36923), .Q(_36905) );
  nor2s1 _36778_inst ( .DIN1(_36924), .DIN2(_36925), .Q(_36923) );
  hi1s1 _36779_inst ( .DIN(_36776), .Q(_36925) );
  nnd2s1 _36780_inst ( .DIN1(_53202), .DIN2(_53201), .Q(_36776) );
  nor2s1 _36781_inst ( .DIN1(_53201), .DIN2(_53202), .Q(_36924) );
  hi1s1 _36782_inst ( .DIN(_36681), .Q(_33292) );
  nnd2s1 _36783_inst ( .DIN1(_36926), .DIN2(_36927), .Q(_36681) );
  nnd2s1 _36784_inst ( .DIN1(_36928), .DIN2(_36929), .Q(
        _____________________________175________) );
  nor2s1 _36785_inst ( .DIN1(_36930), .DIN2(_36931), .Q(_36928) );
  nor2s1 _36786_inst ( .DIN1(_36932), .DIN2(_33149), .Q(_36931) );
  xor2s1 _36787_inst ( .DIN1(_36933), .DIN2(_31768), .Q(_36932) );
  nnd2s1 _36788_inst ( .DIN1(_36934), .DIN2(_36935), .Q(_36933) );
  nnd2s1 _36789_inst ( .DIN1(_36936), .DIN2(_36899), .Q(_36935) );
  xor2s1 _36790_inst ( .DIN1(_26834), .DIN2(_36937), .Q(_36936) );
  xor2s1 _36791_inst ( .DIN1(_26342), .DIN2(_36916), .Q(_36937) );
  nnd2s1 _36792_inst ( .DIN1(_36938), .DIN2(_36939), .Q(_36916) );
  nnd2s1 _36793_inst ( .DIN1(_53204), .DIN2(_36940), .Q(_36939) );
  xor2s1 _36794_inst ( .DIN1(_34235), .DIN2(_36941), .Q(_36940) );
  xor2s1 _36795_inst ( .DIN1(_53372), .DIN2(_53517), .Q(_36942) );
  nnd2s1 _36796_inst ( .DIN1(_36943), .DIN2(_36944), .Q(_36921) );
  nnd2s1 _36797_inst ( .DIN1(_53338), .DIN2(_36945), .Q(_36944) );
  or2s1 _36798_inst ( .DIN1(_36946), .DIN2(_27731), .Q(_36945) );
  nnd2s1 _36799_inst ( .DIN1(_36946), .DIN2(_27731), .Q(_36943) );
  nnd2s1 _36800_inst ( .DIN1(_36947), .DIN2(_53205), .Q(_36934) );
  nor2s1 _36801_inst ( .DIN1(_36948), .DIN2(_26987), .Q(_36947) );
  and2s1 _36802_inst ( .DIN1(_36949), .DIN2(_36950), .Q(_36948) );
  nor2s1 _36803_inst ( .DIN1(_33132), .DIN2(_36951), .Q(_36930) );
  nor2s1 _36804_inst ( .DIN1(_27774), .DIN2(_36952), .Q(_36951) );
  nnd2s1 _36805_inst ( .DIN1(_36953), .DIN2(_27608), .Q(
        _____________________________174________) );
  nnd2s1 _36806_inst ( .DIN1(_33771), .DIN2(_27616), .Q(_27608) );
  nor2s1 _36807_inst ( .DIN1(_36954), .DIN2(_36955), .Q(_36953) );
  nor2s1 _36808_inst ( .DIN1(_27616), .DIN2(_36956), .Q(_36955) );
  nnd2s1 _36809_inst ( .DIN1(_36957), .DIN2(_36882), .Q(_36956) );
  nor2s1 _36810_inst ( .DIN1(_36958), .DIN2(_36959), .Q(_36957) );
  nor2s1 _36811_inst ( .DIN1(_36885), .DIN2(_36960), .Q(_36959) );
  xor2s1 _36812_inst ( .DIN1(_26597), .DIN2(_36961), .Q(_36960) );
  nnd2s1 _36813_inst ( .DIN1(_36941), .DIN2(_36938), .Q(_36961) );
  nnd2s1 _36814_inst ( .DIN1(_33271), .DIN2(_36962), .Q(_36938) );
  or2s1 _36815_inst ( .DIN1(_36962), .DIN2(_33271), .Q(_36941) );
  xnr2s1 _36816_inst ( .DIN1(_36946), .DIN2(_36963), .Q(_33271) );
  xor2s1 _36817_inst ( .DIN1(_53338), .DIN2(_53375), .Q(_36963) );
  nnd2s1 _36818_inst ( .DIN1(_36964), .DIN2(_36965), .Q(_36946) );
  nnd2s1 _36819_inst ( .DIN1(_53373), .DIN2(_36966), .Q(_36965) );
  or2s1 _36820_inst ( .DIN1(_36967), .DIN2(_34787), .Q(_36966) );
  nnd2s1 _36821_inst ( .DIN1(_36967), .DIN2(_34787), .Q(_36964) );
  nnd2s1 _36822_inst ( .DIN1(_36968), .DIN2(_36969), .Q(_36962) );
  nnd2s1 _36823_inst ( .DIN1(_36970), .DIN2(_26671), .Q(_36969) );
  or2s1 _36824_inst ( .DIN1(_36971), .DIN2(_33291), .Q(_36970) );
  nnd2s1 _36825_inst ( .DIN1(_33291), .DIN2(_36971), .Q(_36968) );
  nor2s1 _36826_inst ( .DIN1(_36899), .DIN2(_36972), .Q(_36958) );
  xor2s1 _36827_inst ( .DIN1(_53151), .DIN2(_53205), .Q(_36972) );
  nor2s1 _36828_inst ( .DIN1(_27611), .DIN2(_36973), .Q(_36954) );
  nor2s1 _36829_inst ( .DIN1(_27241), .DIN2(_26505), .Q(_36973) );
  hi1s1 _36830_inst ( .DIN(_27616), .Q(_27611) );
  nnd2s1 _36831_inst ( .DIN1(_36974), .DIN2(_36975), .Q(_27616) );
  nor2s1 _36832_inst ( .DIN1(_36976), .DIN2(_36977), .Q(_36975) );
  nor2s1 _36833_inst ( .DIN1(_36492), .DIN2(_35998), .Q(_36974) );
  nnd2s1 _36834_inst ( .DIN1(_36978), .DIN2(_36979), .Q(
        _____________________________173________) );
  nnd2s1 _36835_inst ( .DIN1(_35829), .DIN2(_36980), .Q(_36979) );
  nnd2s1 _36836_inst ( .DIN1(_36981), .DIN2(_36882), .Q(_36980) );
  nor2s1 _36837_inst ( .DIN1(_36982), .DIN2(_36983), .Q(_36981) );
  nor2s1 _36838_inst ( .DIN1(_36885), .DIN2(_36984), .Q(_36983) );
  xor2s1 _36839_inst ( .DIN1(_33291), .DIN2(_36985), .Q(_36984) );
  xor2s1 _36840_inst ( .DIN1(_26671), .DIN2(_36971), .Q(_36985) );
  nnd2s1 _36841_inst ( .DIN1(_36986), .DIN2(_36987), .Q(_36971) );
  nnd2s1 _36842_inst ( .DIN1(_36988), .DIN2(_26523), .Q(_36987) );
  or2s1 _36843_inst ( .DIN1(_36989), .DIN2(_26822), .Q(_36988) );
  nnd2s1 _36844_inst ( .DIN1(_33982), .DIN2(_36989), .Q(_36986) );
  hi1s1 _36845_inst ( .DIN(_33310), .Q(_33291) );
  xor2s1 _36846_inst ( .DIN1(_36967), .DIN2(_36990), .Q(_33310) );
  xor2s1 _36847_inst ( .DIN1(_53373), .DIN2(_53376), .Q(_36990) );
  nnd2s1 _36848_inst ( .DIN1(_36991), .DIN2(_36992), .Q(_36967) );
  nnd2s1 _36849_inst ( .DIN1(_53374), .DIN2(_36993), .Q(_36992) );
  or2s1 _36850_inst ( .DIN1(_36994), .DIN2(_53377), .Q(_36993) );
  nnd2s1 _36851_inst ( .DIN1(_53377), .DIN2(_36994), .Q(_36991) );
  nor2s1 _36852_inst ( .DIN1(_36899), .DIN2(_36995), .Q(_36982) );
  nor2s1 _36853_inst ( .DIN1(_36996), .DIN2(_36997), .Q(_36995) );
  nnd2s1 _36854_inst ( .DIN1(______[12]), .DIN2(_36998), .Q(_36997) );
  nnd2s1 _36855_inst ( .DIN1(_26407), .DIN2(_26265), .Q(_36998) );
  nnd2s1 _36856_inst ( .DIN1(_36999), .DIN2(_37000), .Q(_36996) );
  nnd2s1 _36857_inst ( .DIN1(_37001), .DIN2(_37002), .Q(_37000) );
  or2s1 _36858_inst ( .DIN1(_37002), .DIN2(_53207), .Q(_36999) );
  nnd2s1 _36859_inst ( .DIN1(_35843), .DIN2(_37003), .Q(_36978) );
  xor2s1 _36860_inst ( .DIN1(_53214), .DIN2(_53216), .Q(_37003) );
  hi1s1 _36861_inst ( .DIN(_37004), .Q(_35843) );
  nnd2s1 _36862_inst ( .DIN1(_37005), .DIN2(_27983), .Q(
        _____________________________172________) );
  nnd2s1 _36863_inst ( .DIN1(_27500), .DIN2(_37006), .Q(_27983) );
  nor2s1 _36864_inst ( .DIN1(_37007), .DIN2(_37008), .Q(_37005) );
  nor2s1 _36865_inst ( .DIN1(_27500), .DIN2(_37009), .Q(_37008) );
  nnd2s1 _36866_inst ( .DIN1(_37010), .DIN2(_36882), .Q(_37009) );
  nnd2s1 _36867_inst ( .DIN1(_37011), .DIN2(_36950), .Q(_36882) );
  nor2s1 _36868_inst ( .DIN1(_37012), .DIN2(_36899), .Q(_37011) );
  nor2s1 _36869_inst ( .DIN1(_37013), .DIN2(_37014), .Q(_37010) );
  nor2s1 _36870_inst ( .DIN1(_36885), .DIN2(_37015), .Q(_37014) );
  xor2s1 _36871_inst ( .DIN1(_33982), .DIN2(_37016), .Q(_37015) );
  xor2s1 _36872_inst ( .DIN1(_26523), .DIN2(_36989), .Q(_37016) );
  nnd2s1 _36873_inst ( .DIN1(_37017), .DIN2(_37018), .Q(_36989) );
  nnd2s1 _36874_inst ( .DIN1(_37019), .DIN2(_26651), .Q(_37018) );
  nnd2s1 _36875_inst ( .DIN1(_33333), .DIN2(_37020), .Q(_37019) );
  xnr2s1 _36876_inst ( .DIN1(_30674), .DIN2(_37021), .Q(_37017) );
  nor2s1 _36877_inst ( .DIN1(_33333), .DIN2(_37020), .Q(_37021) );
  xor2s1 _36878_inst ( .DIN1(_36994), .DIN2(_37022), .Q(_33982) );
  xor2s1 _36879_inst ( .DIN1(_53374), .DIN2(_53377), .Q(_37022) );
  nnd2s1 _36880_inst ( .DIN1(_37023), .DIN2(_37024), .Q(_36994) );
  nnd2s1 _36881_inst ( .DIN1(_53372), .DIN2(_37025), .Q(_37024) );
  or2s1 _36882_inst ( .DIN1(_37026), .DIN2(_53379), .Q(_37025) );
  nnd2s1 _36883_inst ( .DIN1(_53379), .DIN2(_37026), .Q(_37023) );
  nor2s1 _36884_inst ( .DIN1(_36899), .DIN2(_37027), .Q(_37013) );
  nor2s1 _36885_inst ( .DIN1(_53213), .DIN2(_27614), .Q(_37027) );
  hi1s1 _36886_inst ( .DIN(_36885), .Q(_36899) );
  nnd2s1 _36887_inst ( .DIN1(_37028), .DIN2(_37029), .Q(_36885) );
  nor2s1 _36888_inst ( .DIN1(_35114), .DIN2(_37030), .Q(_37029) );
  nor2s1 _36889_inst ( .DIN1(_36209), .DIN2(_35888), .Q(_37028) );
  nnd2s1 _36890_inst ( .DIN1(_37031), .DIN2(_36950), .Q(_35888) );
  nor2s1 _36891_inst ( .DIN1(_37032), .DIN2(_36067), .Q(_36950) );
  nnd2s1 _36892_inst ( .DIN1(_35930), .DIN2(_35271), .Q(_37032) );
  nor2s1 _36893_inst ( .DIN1(_37033), .DIN2(_35253), .Q(_37031) );
  hi1s1 _36894_inst ( .DIN(_37034), .Q(_35253) );
  nor2s1 _36895_inst ( .DIN1(_27994), .DIN2(_26349), .Q(_37007) );
  nnd2s1 _36896_inst ( .DIN1(_37035), .DIN2(_37036), .Q(
        _____________________________171________) );
  nnd2s1 _36897_inst ( .DIN1(_37037), .DIN2(_28178), .Q(_37036) );
  nor2s1 _36898_inst ( .DIN1(_37038), .DIN2(_27291), .Q(_37037) );
  xor2s1 _36899_inst ( .DIN1(_26600), .DIN2(_53405), .Q(_37038) );
  nnd2s1 _36900_inst ( .DIN1(_28010), .DIN2(_37039), .Q(_37035) );
  nnd2s1 _36901_inst ( .DIN1(_37040), .DIN2(_37041), .Q(_37039) );
  nnd2s1 _36902_inst ( .DIN1(_37042), .DIN2(_37043), .Q(_37041) );
  xor2s1 _36903_inst ( .DIN1(_33333), .DIN2(_37044), .Q(_37043) );
  xor2s1 _36904_inst ( .DIN1(_26651), .DIN2(_37020), .Q(_37044) );
  nnd2s1 _36905_inst ( .DIN1(_37045), .DIN2(_37046), .Q(_37020) );
  nnd2s1 _36906_inst ( .DIN1(_37047), .DIN2(_26566), .Q(_37046) );
  nnd2s1 _36907_inst ( .DIN1(_33349), .DIN2(_37048), .Q(_37047) );
  or2s1 _36908_inst ( .DIN1(_37048), .DIN2(_26801), .Q(_37045) );
  hi1s1 _36909_inst ( .DIN(_33344), .Q(_33333) );
  xor2s1 _36910_inst ( .DIN1(_37026), .DIN2(_37049), .Q(_33344) );
  xor2s1 _36911_inst ( .DIN1(_53372), .DIN2(_53379), .Q(_37049) );
  nnd2s1 _36912_inst ( .DIN1(_37050), .DIN2(_37051), .Q(_37026) );
  nnd2s1 _36913_inst ( .DIN1(_53338), .DIN2(_37052), .Q(_37051) );
  or2s1 _36914_inst ( .DIN1(_37053), .DIN2(_53346), .Q(_37052) );
  nnd2s1 _36915_inst ( .DIN1(_53346), .DIN2(_37053), .Q(_37050) );
  nnd2s1 _36916_inst ( .DIN1(_53206), .DIN2(_37054), .Q(_37040) );
  nnd2s1 _36917_inst ( .DIN1(_37055), .DIN2(_37056), .Q(
        _____________________________170________) );
  nnd2s1 _36918_inst ( .DIN1(_37057), .DIN2(_27915), .Q(_37056) );
  nor2s1 _36919_inst ( .DIN1(_37042), .DIN2(_37058), .Q(_37057) );
  nor2s1 _36920_inst ( .DIN1(_37059), .DIN2(_37060), .Q(_37058) );
  nnd2s1 _36921_inst ( .DIN1(_37061), .DIN2(_37054), .Q(_37060) );
  or2s1 _36922_inst ( .DIN1(_37001), .DIN2(_53158), .Q(_37061) );
  nor2s1 _36923_inst ( .DIN1(_26407), .DIN2(_26265), .Q(_37001) );
  nor2s1 _36924_inst ( .DIN1(_26407), .DIN2(_37002), .Q(_37059) );
  nnd2s1 _36925_inst ( .DIN1(_53158), .DIN2(_53206), .Q(_37002) );
  nor2s1 _36926_inst ( .DIN1(_37062), .DIN2(_37063), .Q(_37055) );
  nor2s1 _36927_inst ( .DIN1(_53264), .DIN2(_37064), .Q(_37063) );
  nor2s1 _36928_inst ( .DIN1(_37065), .DIN2(_37066), .Q(_37064) );
  nor2s1 _36929_inst ( .DIN1(_27913), .DIN2(_37067), .Q(_37066) );
  hi1s1 _36930_inst ( .DIN(_37068), .Q(_37067) );
  nor2s1 _36931_inst ( .DIN1(_37069), .DIN2(_37070), .Q(_37065) );
  nor2s1 _36932_inst ( .DIN1(_37071), .DIN2(_26566), .Q(_37062) );
  nor2s1 _36933_inst ( .DIN1(_37072), .DIN2(_37073), .Q(_37071) );
  nor2s1 _36934_inst ( .DIN1(_27913), .DIN2(_37068), .Q(_37073) );
  and2s1 _36935_inst ( .DIN1(_37069), .DIN2(_37074), .Q(_37072) );
  xnr2s1 _36936_inst ( .DIN1(_37048), .DIN2(_34034), .Q(_37069) );
  hi1s1 _36937_inst ( .DIN(_33349), .Q(_34034) );
  xor2s1 _36938_inst ( .DIN1(_37053), .DIN2(_37075), .Q(_33349) );
  xor2s1 _36939_inst ( .DIN1(_53338), .DIN2(_53346), .Q(_37075) );
  nnd2s1 _36940_inst ( .DIN1(_37076), .DIN2(_37077), .Q(_37053) );
  nnd2s1 _36941_inst ( .DIN1(_37078), .DIN2(_34787), .Q(_37077) );
  or2s1 _36942_inst ( .DIN1(_37079), .DIN2(_53381), .Q(_37078) );
  nnd2s1 _36943_inst ( .DIN1(_53381), .DIN2(_37079), .Q(_37076) );
  nnd2s1 _36944_inst ( .DIN1(_37080), .DIN2(_37081), .Q(_37048) );
  nnd2s1 _36945_inst ( .DIN1(_53260), .DIN2(_37082), .Q(_37081) );
  or2s1 _36946_inst ( .DIN1(_37083), .DIN2(_33388), .Q(_37082) );
  nnd2s1 _36947_inst ( .DIN1(_33388), .DIN2(_37083), .Q(_37080) );
  hi1s1 _36948_inst ( .DIN(_33393), .Q(_33388) );
  nnd2s1 _36949_inst ( .DIN1(_37084), .DIN2(_37085), .Q(
        _____________________________16________) );
  nnd2s1 _36950_inst ( .DIN1(_37086), .DIN2(_37087), .Q(_37085) );
  xnr2s1 _36951_inst ( .DIN1(_32833), .DIN2(_53209), .Q(_37087) );
  and2s1 _36952_inst ( .DIN1(______[20]), .DIN2(_33039), .Q(_37086) );
  nnd2s1 _36953_inst ( .DIN1(_32837), .DIN2(_37088), .Q(_37084) );
  nnd2s1 _36954_inst ( .DIN1(_37089), .DIN2(_37090), .Q(_37088) );
  nnd2s1 _36955_inst ( .DIN1(_36804), .DIN2(_37091), .Q(_37090) );
  nnd2s1 _36956_inst ( .DIN1(______[26]), .DIN2(_26379), .Q(_37091) );
  nor2s1 _36957_inst ( .DIN1(_36808), .DIN2(_37092), .Q(_37089) );
  nor2s1 _36958_inst ( .DIN1(_37093), .DIN2(_36810), .Q(_37092) );
  xor2s1 _36959_inst ( .DIN1(_35338), .DIN2(_37094), .Q(_37093) );
  xor2s1 _36960_inst ( .DIN1(_26534), .DIN2(_36816), .Q(_37094) );
  nnd2s1 _36961_inst ( .DIN1(_37095), .DIN2(_37096), .Q(_36816) );
  nnd2s1 _36962_inst ( .DIN1(_53229), .DIN2(_37097), .Q(_37096) );
  or2s1 _36963_inst ( .DIN1(_37098), .DIN2(_35356), .Q(_37097) );
  nnd2s1 _36964_inst ( .DIN1(_35356), .DIN2(_37098), .Q(_37095) );
  hi1s1 _36965_inst ( .DIN(_35353), .Q(_35356) );
  xnr2s1 _36966_inst ( .DIN1(_37099), .DIN2(_36822), .Q(_35338) );
  xor2s1 _36967_inst ( .DIN1(_26323), .DIN2(_36821), .Q(_37099) );
  nnd2s1 _36968_inst ( .DIN1(_37100), .DIN2(_37101), .Q(_36821) );
  nnd2s1 _36969_inst ( .DIN1(_37102), .DIN2(_27731), .Q(_37101) );
  or2s1 _36970_inst ( .DIN1(_37103), .DIN2(_37104), .Q(_37102) );
  nnd2s1 _36971_inst ( .DIN1(_37104), .DIN2(_37103), .Q(_37100) );
  hi1s1 _36972_inst ( .DIN(_37105), .Q(_36808) );
  nnd2s1 _36973_inst ( .DIN1(_37106), .DIN2(_27256), .Q(
        _____________________________169________) );
  nnd2s1 _36974_inst ( .DIN1(_27123), .DIN2(_27122), .Q(_27256) );
  nor2s1 _36975_inst ( .DIN1(_37107), .DIN2(_37108), .Q(_37106) );
  nor2s1 _36976_inst ( .DIN1(_27122), .DIN2(_37109), .Q(_37108) );
  nnd2s1 _36977_inst ( .DIN1(_37110), .DIN2(_37111), .Q(_37109) );
  nnd2s1 _36978_inst ( .DIN1(_37112), .DIN2(_37042), .Q(_37111) );
  xor2s1 _36979_inst ( .DIN1(_33393), .DIN2(_37113), .Q(_37112) );
  xor2s1 _36980_inst ( .DIN1(_26610), .DIN2(_37083), .Q(_37113) );
  nnd2s1 _36981_inst ( .DIN1(_37114), .DIN2(_37115), .Q(_37083) );
  nnd2s1 _36982_inst ( .DIN1(_53265), .DIN2(_37116), .Q(_37115) );
  or2s1 _36983_inst ( .DIN1(_37117), .DIN2(_26802), .Q(_37116) );
  nnd2s1 _36984_inst ( .DIN1(_26802), .DIN2(_37117), .Q(_37114) );
  xnr2s1 _36985_inst ( .DIN1(_37118), .DIN2(_37079), .Q(_33393) );
  nnd2s1 _36986_inst ( .DIN1(_37119), .DIN2(_37120), .Q(_37079) );
  nnd2s1 _36987_inst ( .DIN1(_53377), .DIN2(_37121), .Q(_37120) );
  or2s1 _36988_inst ( .DIN1(_37122), .DIN2(_53380), .Q(_37121) );
  nnd2s1 _36989_inst ( .DIN1(_53380), .DIN2(_37122), .Q(_37119) );
  xor2s1 _36990_inst ( .DIN1(_34787), .DIN2(_53381), .Q(_37118) );
  nnd2s1 _36991_inst ( .DIN1(_37123), .DIN2(_37124), .Q(_37110) );
  nor2s1 _36992_inst ( .DIN1(_37125), .DIN2(_37126), .Q(_37124) );
  nor2s1 _36993_inst ( .DIN1(_53256), .DIN2(_26351), .Q(_37126) );
  nor2s1 _36994_inst ( .DIN1(_27774), .DIN2(_37127), .Q(_37123) );
  hi1s1 _36995_inst ( .DIN(_27116), .Q(_27122) );
  nor2s1 _36996_inst ( .DIN1(_27116), .DIN2(_37128), .Q(_37107) );
  nor2s1 _36997_inst ( .DIN1(_53057), .DIN2(_27241), .Q(_37128) );
  nor2s1 _36998_inst ( .DIN1(_27663), .DIN2(_37129), .Q(_27116) );
  nnd2s1 _36999_inst ( .DIN1(_37130), .DIN2(_37131), .Q(
        _____________________________168________) );
  nnd2s1 _37000_inst ( .DIN1(_37132), .DIN2(_37133), .Q(_37131) );
  xor2s1 _37001_inst ( .DIN1(_33396), .DIN2(_37134), .Q(_37133) );
  xor2s1 _37002_inst ( .DIN1(_26255), .DIN2(_37117), .Q(_37134) );
  nnd2s1 _37003_inst ( .DIN1(_37135), .DIN2(_37136), .Q(_37117) );
  nnd2s1 _37004_inst ( .DIN1(_53257), .DIN2(_37137), .Q(_37136) );
  or2s1 _37005_inst ( .DIN1(_37138), .DIN2(_33419), .Q(_37137) );
  nnd2s1 _37006_inst ( .DIN1(_33419), .DIN2(_37138), .Q(_37135) );
  hi1s1 _37007_inst ( .DIN(_33398), .Q(_33396) );
  xor2s1 _37008_inst ( .DIN1(_37122), .DIN2(_37139), .Q(_33398) );
  xor2s1 _37009_inst ( .DIN1(_53377), .DIN2(_53380), .Q(_37139) );
  nnd2s1 _37010_inst ( .DIN1(_37140), .DIN2(_37141), .Q(_37122) );
  nnd2s1 _37011_inst ( .DIN1(_53350), .DIN2(_37142), .Q(_37141) );
  or2s1 _37012_inst ( .DIN1(_37143), .DIN2(_53379), .Q(_37142) );
  nnd2s1 _37013_inst ( .DIN1(_53379), .DIN2(_37143), .Q(_37140) );
  hi1s1 _37014_inst ( .DIN(_37144), .Q(_37132) );
  nor2s1 _37015_inst ( .DIN1(_37145), .DIN2(_37146), .Q(_37130) );
  nor2s1 _37016_inst ( .DIN1(_37147), .DIN2(_37148), .Q(_37146) );
  nnd2s1 _37017_inst ( .DIN1(_37149), .DIN2(_53210), .Q(_37148) );
  nor2s1 _37018_inst ( .DIN1(_37125), .DIN2(_37042), .Q(_37149) );
  nor2s1 _37019_inst ( .DIN1(_35829), .DIN2(_37150), .Q(_37145) );
  nor2s1 _37020_inst ( .DIN1(_26774), .DIN2(_37151), .Q(_37150) );
  nnd2s1 _37021_inst ( .DIN1(_37152), .DIN2(_37153), .Q(_37151) );
  xor2s1 _37022_inst ( .DIN1(_26372), .DIN2(_37154), .Q(_37152) );
  nnd2s1 _37023_inst ( .DIN1(_53214), .DIN2(_53212), .Q(_37154) );
  nnd2s1 _37024_inst ( .DIN1(_37155), .DIN2(_37156), .Q(
        _____________________________167________) );
  nnd2s1 _37025_inst ( .DIN1(_37157), .DIN2(_37147), .Q(_37156) );
  nnd2s1 _37026_inst ( .DIN1(_37158), .DIN2(_53212), .Q(_37157) );
  nor2s1 _37027_inst ( .DIN1(_36927), .DIN2(_27393), .Q(_37158) );
  nor2s1 _37028_inst ( .DIN1(_37159), .DIN2(_37160), .Q(_37155) );
  nor2s1 _37029_inst ( .DIN1(_37161), .DIN2(_37144), .Q(_37160) );
  nnd2s1 _37030_inst ( .DIN1(_37042), .DIN2(_35829), .Q(_37144) );
  xor2s1 _37031_inst ( .DIN1(_33419), .DIN2(_37162), .Q(_37161) );
  xnr2s1 _37032_inst ( .DIN1(_53257), .DIN2(_37138), .Q(_37162) );
  nnd2s1 _37033_inst ( .DIN1(_37163), .DIN2(_37164), .Q(_37138) );
  nnd2s1 _37034_inst ( .DIN1(_53268), .DIN2(_37165), .Q(_37164) );
  or2s1 _37035_inst ( .DIN1(_37166), .DIN2(_26831), .Q(_37165) );
  nnd2s1 _37036_inst ( .DIN1(_26831), .DIN2(_37166), .Q(_37163) );
  xnr2s1 _37037_inst ( .DIN1(_37167), .DIN2(_37143), .Q(_33419) );
  nnd2s1 _37038_inst ( .DIN1(_37168), .DIN2(_37169), .Q(_37143) );
  nnd2s1 _37039_inst ( .DIN1(_53346), .DIN2(_37170), .Q(_37169) );
  or2s1 _37040_inst ( .DIN1(_37171), .DIN2(_53352), .Q(_37170) );
  nnd2s1 _37041_inst ( .DIN1(_53352), .DIN2(_37171), .Q(_37168) );
  xor2s1 _37042_inst ( .DIN1(_26320), .DIN2(_53379), .Q(_37167) );
  nor2s1 _37043_inst ( .DIN1(_37042), .DIN2(_37172), .Q(_37159) );
  nnd2s1 _37044_inst ( .DIN1(_37054), .DIN2(_26351), .Q(_37172) );
  hi1s1 _37045_inst ( .DIN(_37125), .Q(_37054) );
  nnd2s1 _37046_inst ( .DIN1(_37173), .DIN2(_37174), .Q(
        _____________________________166________) );
  nnd2s1 _37047_inst ( .DIN1(_37074), .DIN2(_37175), .Q(_37174) );
  xnr2s1 _37048_inst ( .DIN1(_26831), .DIN2(_37176), .Q(_37175) );
  xnr2s1 _37049_inst ( .DIN1(_53268), .DIN2(_37166), .Q(_37176) );
  nnd2s1 _37050_inst ( .DIN1(_37177), .DIN2(_37178), .Q(_37166) );
  nnd2s1 _37051_inst ( .DIN1(_37179), .DIN2(_26664), .Q(_37178) );
  nnd2s1 _37052_inst ( .DIN1(_37180), .DIN2(_34138), .Q(_37179) );
  xor2s1 _37053_inst ( .DIN1(_30163), .DIN2(_37181), .Q(_37177) );
  nor2s1 _37054_inst ( .DIN1(_37180), .DIN2(_34138), .Q(_37181) );
  xor2s1 _37055_inst ( .DIN1(_53346), .DIN2(_53352), .Q(_37182) );
  nnd2s1 _37056_inst ( .DIN1(_37183), .DIN2(_37184), .Q(_37171) );
  nnd2s1 _37057_inst ( .DIN1(_53357), .DIN2(_37185), .Q(_37184) );
  or2s1 _37058_inst ( .DIN1(_37186), .DIN2(_53381), .Q(_37185) );
  nnd2s1 _37059_inst ( .DIN1(_53381), .DIN2(_37186), .Q(_37183) );
  hi1s1 _37060_inst ( .DIN(_37070), .Q(_37074) );
  nnd2s1 _37061_inst ( .DIN1(_37042), .DIN2(_27915), .Q(_37070) );
  and2s1 _37062_inst ( .DIN1(_37187), .DIN2(_37188), .Q(_37042) );
  nor2s1 _37063_inst ( .DIN1(_37189), .DIN2(_37190), .Q(_37188) );
  nnd2s1 _37064_inst ( .DIN1(_35271), .DIN2(_37034), .Q(_37190) );
  nor2s1 _37065_inst ( .DIN1(_36228), .DIN2(_35933), .Q(_37187) );
  nnd2s1 _37066_inst ( .DIN1(_37191), .DIN2(_37192), .Q(_36228) );
  nor2s1 _37067_inst ( .DIN1(_37193), .DIN2(_37194), .Q(_37192) );
  nor2s1 _37068_inst ( .DIN1(_36209), .DIN2(_36067), .Q(_37191) );
  xnr2s1 _37069_inst ( .DIN1(_37195), .DIN2(_37196), .Q(_36067) );
  nor2s1 _37070_inst ( .DIN1(_37197), .DIN2(_37198), .Q(_37196) );
  nnd2s1 _37071_inst ( .DIN1(_36066), .DIN2(_37199), .Q(_36209) );
  nnd2s1 _37072_inst ( .DIN1(______[18]), .DIN2(_37200), .Q(_37173) );
  nnd2s1 _37073_inst ( .DIN1(_37201), .DIN2(_37202), .Q(_37200) );
  nnd2s1 _37074_inst ( .DIN1(_37203), .DIN2(_27915), .Q(_37202) );
  nor2s1 _37075_inst ( .DIN1(_37125), .DIN2(_37204), .Q(_37203) );
  nor2s1 _37076_inst ( .DIN1(_37205), .DIN2(_37127), .Q(_37204) );
  nnd2s1 _37077_inst ( .DIN1(_37206), .DIN2(_37207), .Q(_37127) );
  nnd2s1 _37078_inst ( .DIN1(_26272), .DIN2(_26716), .Q(_37207) );
  nnd2s1 _37079_inst ( .DIN1(_37208), .DIN2(_53214), .Q(_37206) );
  nor2s1 _37080_inst ( .DIN1(_53212), .DIN2(_26272), .Q(_37208) );
  nor2s1 _37081_inst ( .DIN1(_53214), .DIN2(_26351), .Q(_37205) );
  nor2s1 _37082_inst ( .DIN1(_36059), .DIN2(_37030), .Q(_37125) );
  nnd2s1 _37083_inst ( .DIN1(_37209), .DIN2(_37210), .Q(_36059) );
  and2s1 _37084_inst ( .DIN1(_36066), .DIN2(_37211), .Q(_37210) );
  nor2s1 _37085_inst ( .DIN1(_37189), .DIN2(_37198), .Q(_37209) );
  or2s1 _37086_inst ( .DIN1(_35113), .DIN2(_35929), .Q(_37198) );
  nnd2s1 _37087_inst ( .DIN1(_37212), .DIN2(_37213), .Q(_37201) );
  xor2s1 _37088_inst ( .DIN1(_37068), .DIN2(_53207), .Q(_37212) );
  nnd2s1 _37089_inst ( .DIN1(_37214), .DIN2(_37215), .Q(
        _____________________________165________) );
  nnd2s1 _37090_inst ( .DIN1(_37216), .DIN2(_37217), .Q(_37215) );
  nnd2s1 _37091_inst ( .DIN1(_37218), .DIN2(______[6]), .Q(_37217) );
  nor2s1 _37092_inst ( .DIN1(_37219), .DIN2(_37220), .Q(_37218) );
  xor2s1 _37093_inst ( .DIN1(_37221), .DIN2(_37222), .Q(_37220) );
  xor2s1 _37094_inst ( .DIN1(_53218), .DIN2(_53220), .Q(_37222) );
  nnd2s1 _37095_inst ( .DIN1(_26533), .DIN2(_26268), .Q(_37221) );
  nor2s1 _37096_inst ( .DIN1(_37223), .DIN2(_37224), .Q(_37214) );
  nor2s1 _37097_inst ( .DIN1(_37225), .DIN2(_37004), .Q(_37224) );
  xor2s1 _37098_inst ( .DIN1(_26372), .DIN2(_53214), .Q(_37225) );
  nor2s1 _37099_inst ( .DIN1(_37226), .DIN2(_37227), .Q(_37223) );
  xor2s1 _37100_inst ( .DIN1(_34138), .DIN2(_37228), .Q(_37227) );
  xor2s1 _37101_inst ( .DIN1(_26664), .DIN2(_37180), .Q(_37228) );
  and2s1 _37102_inst ( .DIN1(_37229), .DIN2(_37230), .Q(_37180) );
  nnd2s1 _37103_inst ( .DIN1(_37231), .DIN2(_26385), .Q(_37230) );
  or2s1 _37104_inst ( .DIN1(_37232), .DIN2(_26833), .Q(_37231) );
  nnd2s1 _37105_inst ( .DIN1(_26833), .DIN2(_37232), .Q(_37229) );
  xor2s1 _37106_inst ( .DIN1(_37233), .DIN2(_37234), .Q(_34138) );
  xor2s1 _37107_inst ( .DIN1(_29518), .DIN2(_37186), .Q(_37234) );
  nnd2s1 _37108_inst ( .DIN1(_37235), .DIN2(_37236), .Q(_37186) );
  nnd2s1 _37109_inst ( .DIN1(_53358), .DIN2(_37237), .Q(_37236) );
  or2s1 _37110_inst ( .DIN1(_37238), .DIN2(_53380), .Q(_37237) );
  nnd2s1 _37111_inst ( .DIN1(_53380), .DIN2(_37238), .Q(_37235) );
  xor2s1 _37112_inst ( .DIN1(_26396), .DIN2(_53381), .Q(_37233) );
  nnd2s1 _37113_inst ( .DIN1(_37239), .DIN2(_28298), .Q(
        _____________________________164________) );
  nnd2s1 _37114_inst ( .DIN1(_37240), .DIN2(_28302), .Q(_28298) );
  nor2s1 _37115_inst ( .DIN1(_37241), .DIN2(_37242), .Q(_37239) );
  nor2s1 _37116_inst ( .DIN1(_28302), .DIN2(_37243), .Q(_37242) );
  nor2s1 _37117_inst ( .DIN1(_37244), .DIN2(_37245), .Q(_37243) );
  nor2s1 _37118_inst ( .DIN1(_35771), .DIN2(_37246), .Q(_37245) );
  nnd2s1 _37119_inst ( .DIN1(_37247), .DIN2(______[14]), .Q(_37246) );
  nor2s1 _37120_inst ( .DIN1(_53216), .DIN2(_37219), .Q(_37247) );
  nor2s1 _37121_inst ( .DIN1(_35764), .DIN2(_37248), .Q(_37244) );
  xnr2s1 _37122_inst ( .DIN1(_26833), .DIN2(_37249), .Q(_37248) );
  xor2s1 _37123_inst ( .DIN1(_26385), .DIN2(_37232), .Q(_37249) );
  nnd2s1 _37124_inst ( .DIN1(_37250), .DIN2(_37251), .Q(_37232) );
  nnd2s1 _37125_inst ( .DIN1(_37252), .DIN2(_26375), .Q(_37251) );
  or2s1 _37126_inst ( .DIN1(_37253), .DIN2(_33504), .Q(_37252) );
  nnd2s1 _37127_inst ( .DIN1(_33504), .DIN2(_37253), .Q(_37250) );
  xor2s1 _37128_inst ( .DIN1(_53358), .DIN2(_53380), .Q(_37254) );
  nnd2s1 _37129_inst ( .DIN1(_37255), .DIN2(_37256), .Q(_37238) );
  nnd2s1 _37130_inst ( .DIN1(_53350), .DIN2(_37257), .Q(_37256) );
  or2s1 _37131_inst ( .DIN1(_37258), .DIN2(_53467), .Q(_37257) );
  nnd2s1 _37132_inst ( .DIN1(_53467), .DIN2(_37258), .Q(_37255) );
  nor2s1 _37133_inst ( .DIN1(_28308), .DIN2(_37259), .Q(_37241) );
  nor2s1 _37134_inst ( .DIN1(_28100), .DIN2(_37260), .Q(_37259) );
  xor2s1 _37135_inst ( .DIN1(_53215), .DIN2(_37261), .Q(_37260) );
  nor2s1 _37136_inst ( .DIN1(_53510), .DIN2(_53489), .Q(_37261) );
  nnd2s1 _37137_inst ( .DIN1(_37262), .DIN2(_27994), .Q(
        _____________________________163________) );
  nor2s1 _37138_inst ( .DIN1(_37263), .DIN2(_37264), .Q(_37262) );
  nor2s1 _37139_inst ( .DIN1(_35764), .DIN2(_37265), .Q(_37264) );
  xor2s1 _37140_inst ( .DIN1(_37253), .DIN2(_37266), .Q(_37265) );
  xor2s1 _37141_inst ( .DIN1(_26375), .DIN2(_33504), .Q(_37266) );
  xnr2s1 _37142_inst ( .DIN1(_37267), .DIN2(_37258), .Q(_33504) );
  nnd2s1 _37143_inst ( .DIN1(_37268), .DIN2(_37269), .Q(_37258) );
  nnd2s1 _37144_inst ( .DIN1(_53352), .DIN2(_37270), .Q(_37269) );
  or2s1 _37145_inst ( .DIN1(_37271), .DIN2(_26329), .Q(_37270) );
  nnd2s1 _37146_inst ( .DIN1(_37271), .DIN2(_26329), .Q(_37268) );
  xor2s1 _37147_inst ( .DIN1(_26341), .DIN2(_53350), .Q(_37267) );
  xnr2s1 _37148_inst ( .DIN1(_37272), .DIN2(_36328), .Q(_37253) );
  hi1s1 _37149_inst ( .DIN(_31282), .Q(_36328) );
  nnd2s1 _37150_inst ( .DIN1(_37273), .DIN2(_37274), .Q(_37272) );
  or2s1 _37151_inst ( .DIN1(_33534), .DIN2(_53093), .Q(_37274) );
  nnd2s1 _37152_inst ( .DIN1(_37275), .DIN2(_37276), .Q(_37273) );
  nnd2s1 _37153_inst ( .DIN1(_53093), .DIN2(_33534), .Q(_37276) );
  hi1s1 _37154_inst ( .DIN(_34172), .Q(_33534) );
  xor2s1 _37155_inst ( .DIN1(_33214), .DIN2(_33517), .Q(_34172) );
  nor2s1 _37156_inst ( .DIN1(_35771), .DIN2(_37277), .Q(_37263) );
  nor2s1 _37157_inst ( .DIN1(_37219), .DIN2(_26594), .Q(_37277) );
  hi1s1 _37158_inst ( .DIN(_35775), .Q(_37219) );
  nnd2s1 _37159_inst ( .DIN1(_37278), .DIN2(_37279), .Q(
        _____________________________162________) );
  nnd2s1 _37160_inst ( .DIN1(_37280), .DIN2(_37281), .Q(_37279) );
  hi1s1 _37161_inst ( .DIN(_37226), .Q(_37281) );
  nnd2s1 _37162_inst ( .DIN1(_35829), .DIN2(_35771), .Q(_37226) );
  hi1s1 _37163_inst ( .DIN(_37147), .Q(_35829) );
  xor2s1 _37164_inst ( .DIN1(_37282), .DIN2(_33517), .Q(_37280) );
  xnr2s1 _37165_inst ( .DIN1(_37271), .DIN2(_37283), .Q(_33517) );
  xor2s1 _37166_inst ( .DIN1(_53352), .DIN2(_53353), .Q(_37283) );
  nnd2s1 _37167_inst ( .DIN1(_37284), .DIN2(_37285), .Q(_37271) );
  nnd2s1 _37168_inst ( .DIN1(_53357), .DIN2(_37286), .Q(_37285) );
  nnd2s1 _37169_inst ( .DIN1(_53366), .DIN2(_37287), .Q(_37286) );
  nnd2s1 _37170_inst ( .DIN1(_37288), .DIN2(_26698), .Q(_37284) );
  hi1s1 _37171_inst ( .DIN(_37287), .Q(_37288) );
  xnr2s1 _37172_inst ( .DIN1(_37275), .DIN2(_53093), .Q(_37282) );
  nor2s1 _37173_inst ( .DIN1(_37289), .DIN2(_37290), .Q(_37278) );
  nor2s1 _37174_inst ( .DIN1(_37004), .DIN2(_37291), .Q(_37290) );
  nnd2s1 _37175_inst ( .DIN1(_26859), .DIN2(_37292), .Q(_37291) );
  xor2s1 _37176_inst ( .DIN1(_37293), .DIN2(_37294), .Q(_37292) );
  xor2s1 _37177_inst ( .DIN1(_53098), .DIN2(_53217), .Q(_37294) );
  nor2s1 _37178_inst ( .DIN1(_26263), .DIN2(_26595), .Q(_37293) );
  nnd2s1 _37179_inst ( .DIN1(_37147), .DIN2(_37153), .Q(_37004) );
  nor2s1 _37180_inst ( .DIN1(_37295), .DIN2(_37296), .Q(_37289) );
  nnd2s1 _37181_inst ( .DIN1(_37297), .DIN2(_37216), .Q(_37296) );
  nor2s1 _37182_inst ( .DIN1(_37147), .DIN2(_35771), .Q(_37216) );
  nnd2s1 _37183_inst ( .DIN1(_37298), .DIN2(_37299), .Q(_37147) );
  xor2s1 _37184_inst ( .DIN1(_26268), .DIN2(_53220), .Q(_37297) );
  nnd2s1 _37185_inst ( .DIN1(______[16]), .DIN2(_35775), .Q(_37295) );
  nnd2s1 _37186_inst ( .DIN1(_37300), .DIN2(_37301), .Q(
        _____________________________161________) );
  nnd2s1 _37187_inst ( .DIN1(_37302), .DIN2(_53222), .Q(_37301) );
  hi1s1 _37188_inst ( .DIN(_36929), .Q(_37302) );
  nnd2s1 _37189_inst ( .DIN1(_37303), .DIN2(_53221), .Q(_36929) );
  and2s1 _37190_inst ( .DIN1(_33149), .DIN2(_53223), .Q(_37303) );
  nor2s1 _37191_inst ( .DIN1(_37304), .DIN2(_37305), .Q(_37300) );
  nor2s1 _37192_inst ( .DIN1(_33149), .DIN2(_37306), .Q(_37305) );
  nor2s1 _37193_inst ( .DIN1(_37307), .DIN2(_37308), .Q(_37306) );
  nor2s1 _37194_inst ( .DIN1(_37309), .DIN2(_35764), .Q(_37308) );
  nor2s1 _37195_inst ( .DIN1(_37310), .DIN2(_37275), .Q(_37309) );
  and2s1 _37196_inst ( .DIN1(_33515), .DIN2(_26569), .Q(_37275) );
  nor2s1 _37197_inst ( .DIN1(_33515), .DIN2(_26569), .Q(_37310) );
  xor2s1 _37198_inst ( .DIN1(_37287), .DIN2(_37311), .Q(_33515) );
  xor2s1 _37199_inst ( .DIN1(_53357), .DIN2(_53366), .Q(_37311) );
  nnd2s1 _37200_inst ( .DIN1(_53358), .DIN2(_53369), .Q(_37287) );
  nor2s1 _37201_inst ( .DIN1(_35771), .DIN2(_37312), .Q(_37307) );
  nor2s1 _37202_inst ( .DIN1(_37313), .DIN2(_37314), .Q(_37312) );
  nnd2s1 _37203_inst ( .DIN1(______[0]), .DIN2(_35775), .Q(_37314) );
  nnd2s1 _37204_inst ( .DIN1(_37315), .DIN2(_37316), .Q(_35775) );
  nor2s1 _37205_inst ( .DIN1(_36456), .DIN2(_37317), .Q(_37316) );
  nnd2s1 _37206_inst ( .DIN1(_37318), .DIN2(_37034), .Q(_37317) );
  nor2s1 _37207_inst ( .DIN1(_35115), .DIN2(_37319), .Q(_37315) );
  nnd2s1 _37208_inst ( .DIN1(_37320), .DIN2(_37211), .Q(_37319) );
  nnd2s1 _37209_inst ( .DIN1(_37321), .DIN2(_37322), .Q(_35115) );
  nor2s1 _37210_inst ( .DIN1(_37197), .DIN2(_36199), .Q(_37322) );
  nor2s1 _37211_inst ( .DIN1(_35887), .DIN2(_37030), .Q(_37321) );
  nnd2s1 _37212_inst ( .DIN1(_37323), .DIN2(_36949), .Q(_37030) );
  nnd2s1 _37213_inst ( .DIN1(_35269), .DIN2(_36207), .Q(_35887) );
  xor2s1 _37214_inst ( .DIN1(_26455), .DIN2(_35824), .Q(_37313) );
  nnd2s1 _37215_inst ( .DIN1(_53225), .DIN2(_53224), .Q(_35824) );
  hi1s1 _37216_inst ( .DIN(_35764), .Q(_35771) );
  nnd2s1 _37217_inst ( .DIN1(_37324), .DIN2(_37325), .Q(_35764) );
  nor2s1 _37218_inst ( .DIN1(_36456), .DIN2(_37326), .Q(_37325) );
  nnd2s1 _37219_inst ( .DIN1(_37034), .DIN2(_35104), .Q(_37326) );
  nor2s1 _37220_inst ( .DIN1(_35273), .DIN2(_35931), .Q(_37324) );
  nnd2s1 _37221_inst ( .DIN1(_37320), .DIN2(_35271), .Q(_35931) );
  nnd2s1 _37222_inst ( .DIN1(_37327), .DIN2(_37328), .Q(_35271) );
  nor2s1 _37223_inst ( .DIN1(_53425), .DIN2(_37329), .Q(_37327) );
  nnd2s1 _37224_inst ( .DIN1(_37330), .DIN2(_37331), .Q(_35273) );
  nor2s1 _37225_inst ( .DIN1(_37332), .DIN2(_37193), .Q(_37331) );
  nor2s1 _37226_inst ( .DIN1(_35256), .DIN2(_35933), .Q(_37330) );
  nnd2s1 _37227_inst ( .DIN1(_37333), .DIN2(_37211), .Q(_35933) );
  nor2s1 _37228_inst ( .DIN1(_37012), .DIN2(_35114), .Q(_37333) );
  or2s1 _37229_inst ( .DIN1(_37334), .DIN2(_36203), .Q(_35256) );
  nor2s1 _37230_inst ( .DIN1(_33132), .DIN2(_37335), .Q(_37304) );
  nor2s1 _37231_inst ( .DIN1(_36952), .DIN2(_37336), .Q(_37335) );
  nnd2s1 _37232_inst ( .DIN1(______[22]), .DIN2(_37337), .Q(_37336) );
  or2s1 _37233_inst ( .DIN1(_53222), .DIN2(_53221), .Q(_37337) );
  nnd2s1 _37234_inst ( .DIN1(_33152), .DIN2(_37338), .Q(_36952) );
  or2s1 _37235_inst ( .DIN1(_53223), .DIN2(_53221), .Q(_37338) );
  nnd2s1 _37236_inst ( .DIN1(_37339), .DIN2(_37340), .Q(
        _____________________________160________) );
  nnd2s1 _37237_inst ( .DIN1(_37341), .DIN2(_37342), .Q(_37340) );
  xor2s1 _37238_inst ( .DIN1(_53355), .DIN2(_53356), .Q(_37342) );
  nnd2s1 _37239_inst ( .DIN1(_27655), .DIN2(_37343), .Q(_37339) );
  nnd2s1 _37240_inst ( .DIN1(_37344), .DIN2(_37345), .Q(_37343) );
  nnd2s1 _37241_inst ( .DIN1(_53136), .DIN2(_32920), .Q(_37345) );
  nor2s1 _37242_inst ( .DIN1(_37346), .DIN2(_37347), .Q(_37344) );
  nor2s1 _37243_inst ( .DIN1(_26300), .DIN2(_37348), .Q(_37347) );
  nor2s1 _37244_inst ( .DIN1(_37349), .DIN2(_37350), .Q(_37348) );
  nor2s1 _37245_inst ( .DIN1(_33578), .DIN2(_37351), .Q(_37350) );
  nor2s1 _37246_inst ( .DIN1(_37352), .DIN2(_33577), .Q(_37349) );
  nor2s1 _37247_inst ( .DIN1(_53226), .DIN2(_37353), .Q(_37346) );
  nor2s1 _37248_inst ( .DIN1(_37354), .DIN2(_37355), .Q(_37353) );
  nor2s1 _37249_inst ( .DIN1(_33577), .DIN2(_37351), .Q(_37355) );
  nor2s1 _37250_inst ( .DIN1(_37352), .DIN2(_33578), .Q(_37354) );
  hi1s1 _37251_inst ( .DIN(_37351), .Q(_37352) );
  nnd2s1 _37252_inst ( .DIN1(_37356), .DIN2(_37357), .Q(_37351) );
  nnd2s1 _37253_inst ( .DIN1(_37358), .DIN2(_26213), .Q(_37357) );
  nnd2s1 _37254_inst ( .DIN1(_37359), .DIN2(_37360), .Q(_37358) );
  or2s1 _37255_inst ( .DIN1(_37360), .DIN2(_37359), .Q(_37356) );
  nnd2s1 _37256_inst ( .DIN1(_37361), .DIN2(_37362), .Q(
        _____________________________15________) );
  nor2s1 _37257_inst ( .DIN1(_37363), .DIN2(_37364), .Q(_37362) );
  nor2s1 _37258_inst ( .DIN1(_28016), .DIN2(_37365), .Q(_37364) );
  nnd2s1 _37259_inst ( .DIN1(_37366), .DIN2(_37367), .Q(_37365) );
  nnd2s1 _37260_inst ( .DIN1(_36530), .DIN2(_37368), .Q(_37367) );
  xor2s1 _37261_inst ( .DIN1(_53227), .DIN2(_53228), .Q(_37368) );
  nnd2s1 _37262_inst ( .DIN1(_37369), .DIN2(_36533), .Q(_37366) );
  xor2s1 _37263_inst ( .DIN1(_35353), .DIN2(_37370), .Q(_37369) );
  xnr2s1 _37264_inst ( .DIN1(_53229), .DIN2(_37098), .Q(_37370) );
  nnd2s1 _37265_inst ( .DIN1(_37371), .DIN2(_37372), .Q(_37098) );
  nnd2s1 _37266_inst ( .DIN1(_53241), .DIN2(_37373), .Q(_37372) );
  or2s1 _37267_inst ( .DIN1(_37374), .DIN2(_35407), .Q(_37373) );
  xor2s1 _37268_inst ( .DIN1(_31842), .DIN2(_37375), .Q(_37371) );
  nnd2s1 _37269_inst ( .DIN1(_35407), .DIN2(_37374), .Q(_37375) );
  hi1s1 _37270_inst ( .DIN(_37376), .Q(_35407) );
  xnr2s1 _37271_inst ( .DIN1(_37377), .DIN2(_37104), .Q(_35353) );
  xor2s1 _37272_inst ( .DIN1(_27731), .DIN2(_37103), .Q(_37377) );
  nnd2s1 _37273_inst ( .DIN1(_37378), .DIN2(_37379), .Q(_37103) );
  nnd2s1 _37274_inst ( .DIN1(_53373), .DIN2(_37380), .Q(_37379) );
  or2s1 _37275_inst ( .DIN1(_37381), .DIN2(_37382), .Q(_37380) );
  nnd2s1 _37276_inst ( .DIN1(_37382), .DIN2(_37381), .Q(_37378) );
  nor2s1 _37277_inst ( .DIN1(_28024), .DIN2(_37383), .Q(_37363) );
  nor2s1 _37278_inst ( .DIN1(_37384), .DIN2(_28684), .Q(_37383) );
  nor2s1 _37279_inst ( .DIN1(_37385), .DIN2(_26683), .Q(_37384) );
  nor2s1 _37280_inst ( .DIN1(_35064), .DIN2(_37386), .Q(_37361) );
  nor2s1 _37281_inst ( .DIN1(_53230), .DIN2(_28027), .Q(_37386) );
  nnd2s1 _37282_inst ( .DIN1(_37385), .DIN2(_28016), .Q(_28027) );
  hi1s1 _37283_inst ( .DIN(_35063), .Q(_37385) );
  nnd2s1 _37284_inst ( .DIN1(_53231), .DIN2(_53232), .Q(_35063) );
  hi1s1 _37285_inst ( .DIN(_28026), .Q(_35064) );
  nnd2s1 _37286_inst ( .DIN1(_37387), .DIN2(_37388), .Q(
        _____________________________159________) );
  nnd2s1 _37287_inst ( .DIN1(_37389), .DIN2(_28923), .Q(_37388) );
  nor2s1 _37288_inst ( .DIN1(_28308), .DIN2(_37240), .Q(_28923) );
  nor2s1 _37289_inst ( .DIN1(_37390), .DIN2(_27393), .Q(_37389) );
  xor2s1 _37290_inst ( .DIN1(_26551), .DIN2(_53489), .Q(_37390) );
  nnd2s1 _37291_inst ( .DIN1(_28308), .DIN2(_37391), .Q(_37387) );
  xor2s1 _37292_inst ( .DIN1(_32330), .DIN2(_37392), .Q(_37391) );
  nnd2s1 _37293_inst ( .DIN1(_37393), .DIN2(_37394), .Q(_37392) );
  nor2s1 _37294_inst ( .DIN1(_37395), .DIN2(_37396), .Q(_37393) );
  nor2s1 _37295_inst ( .DIN1(_32855), .DIN2(_37397), .Q(_37396) );
  xnr2s1 _37296_inst ( .DIN1(_37359), .DIN2(_37398), .Q(_37397) );
  xor2s1 _37297_inst ( .DIN1(_26213), .DIN2(_37360), .Q(_37398) );
  nnd2s1 _37298_inst ( .DIN1(_37399), .DIN2(_37400), .Q(_37360) );
  nnd2s1 _37299_inst ( .DIN1(_37401), .DIN2(_26436), .Q(_37400) );
  xor2s1 _37300_inst ( .DIN1(_31282), .DIN2(_37402), .Q(_37401) );
  nnd2s1 _37301_inst ( .DIN1(_37403), .DIN2(_37404), .Q(_31282) );
  nnd2s1 _37302_inst ( .DIN1(_34289), .DIN2(_53500), .Q(_37404) );
  nor2s1 _37303_inst ( .DIN1(_32878), .DIN2(_37405), .Q(_37395) );
  nor2s1 _37304_inst ( .DIN1(_26772), .DIN2(_37406), .Q(_37405) );
  nnd2s1 _37305_inst ( .DIN1(_37407), .DIN2(_37408), .Q(_37406) );
  or2s1 _37306_inst ( .DIN1(_32857), .DIN2(_53275), .Q(_37408) );
  nor2s1 _37307_inst ( .DIN1(_26518), .DIN2(_53344), .Q(_32857) );
  nnd2s1 _37308_inst ( .DIN1(_32856), .DIN2(_53215), .Q(_37407) );
  and2s1 _37309_inst ( .DIN1(_53275), .DIN2(_26613), .Q(_32856) );
  hi1s1 _37310_inst ( .DIN(_28302), .Q(_28308) );
  nnd2s1 _37311_inst ( .DIN1(_37409), .DIN2(_37410), .Q(_28302) );
  nor2s1 _37312_inst ( .DIN1(_37411), .DIN2(_37412), .Q(_37410) );
  nnd2s1 _37313_inst ( .DIN1(_37413), .DIN2(_34485), .Q(_37412) );
  nor2s1 _37314_inst ( .DIN1(_37414), .DIN2(_29184), .Q(_37409) );
  nnd2s1 _37315_inst ( .DIN1(_37415), .DIN2(_27660), .Q(
        _____________________________158________) );
  nnd2s1 _37316_inst ( .DIN1(_37416), .DIN2(_28380), .Q(_27660) );
  nor2s1 _37317_inst ( .DIN1(_37417), .DIN2(_37418), .Q(_28380) );
  nor2s1 _37318_inst ( .DIN1(_27672), .DIN2(_37419), .Q(_37416) );
  nor2s1 _37319_inst ( .DIN1(_37420), .DIN2(_37421), .Q(_37415) );
  nor2s1 _37320_inst ( .DIN1(_27663), .DIN2(_37422), .Q(_37421) );
  nor2s1 _37321_inst ( .DIN1(_37423), .DIN2(_37424), .Q(_37422) );
  nor2s1 _37322_inst ( .DIN1(_32855), .DIN2(_37425), .Q(_37424) );
  xnr2s1 _37323_inst ( .DIN1(_37426), .DIN2(_37427), .Q(_37425) );
  xor2s1 _37324_inst ( .DIN1(_26436), .DIN2(_37428), .Q(_37427) );
  nnd2s1 _37325_inst ( .DIN1(_37399), .DIN2(_37402), .Q(_37428) );
  nnd2s1 _37326_inst ( .DIN1(_37429), .DIN2(_37430), .Q(_37402) );
  nor2s1 _37327_inst ( .DIN1(_37431), .DIN2(_37432), .Q(_37429) );
  nor2s1 _37328_inst ( .DIN1(_53297), .DIN2(_37433), .Q(_37431) );
  nnd2s1 _37329_inst ( .DIN1(_37434), .DIN2(_37435), .Q(_37399) );
  nor2s1 _37330_inst ( .DIN1(_37436), .DIN2(_37433), .Q(_37434) );
  nor2s1 _37331_inst ( .DIN1(_37437), .DIN2(_37438), .Q(_37433) );
  nor2s1 _37332_inst ( .DIN1(_37432), .DIN2(_26266), .Q(_37436) );
  nor2s1 _37333_inst ( .DIN1(_37439), .DIN2(_37440), .Q(_37432) );
  hi1s1 _37334_inst ( .DIN(_37438), .Q(_37439) );
  nor2s1 _37335_inst ( .DIN1(_32878), .DIN2(_37441), .Q(_37423) );
  nor2s1 _37336_inst ( .DIN1(_37442), .DIN2(_37443), .Q(_37441) );
  nnd2s1 _37337_inst ( .DIN1(______[22]), .DIN2(_37444), .Q(_37443) );
  nnd2s1 _37338_inst ( .DIN1(_36688), .DIN2(_37445), .Q(_37444) );
  xor2s1 _37339_inst ( .DIN1(_26476), .DIN2(_37446), .Q(_37442) );
  nnd2s1 _37340_inst ( .DIN1(_53323), .DIN2(_53234), .Q(_37446) );
  nor2s1 _37341_inst ( .DIN1(_27672), .DIN2(_37447), .Q(_37420) );
  xor2s1 _37342_inst ( .DIN1(_27674), .DIN2(_53233), .Q(_37447) );
  nnd2s1 _37343_inst ( .DIN1(_53267), .DIN2(_53268), .Q(_27674) );
  hi1s1 _37344_inst ( .DIN(_27663), .Q(_27672) );
  nnd2s1 _37345_inst ( .DIN1(_37448), .DIN2(_27154), .Q(_27663) );
  nnd2s1 _37346_inst ( .DIN1(_37449), .DIN2(_30228), .Q(
        _____________________________157________) );
  nnd2s1 _37347_inst ( .DIN1(_33489), .DIN2(_29555), .Q(_30228) );
  nor2s1 _37348_inst ( .DIN1(_37450), .DIN2(_37451), .Q(_37449) );
  nor2s1 _37349_inst ( .DIN1(_37452), .DIN2(_29555), .Q(_37451) );
  nor2s1 _37350_inst ( .DIN1(_32861), .DIN2(_37453), .Q(_37452) );
  nnd2s1 _37351_inst ( .DIN1(_37454), .DIN2(_37455), .Q(_37453) );
  nnd2s1 _37352_inst ( .DIN1(_37456), .DIN2(_32855), .Q(_37455) );
  xor2s1 _37353_inst ( .DIN1(_26260), .DIN2(_53267), .Q(_37456) );
  nnd2s1 _37354_inst ( .DIN1(_37457), .DIN2(_32878), .Q(_37454) );
  xor2s1 _37355_inst ( .DIN1(_37440), .DIN2(_37458), .Q(_37457) );
  xor2s1 _37356_inst ( .DIN1(_26266), .DIN2(_37438), .Q(_37458) );
  nnd2s1 _37357_inst ( .DIN1(_37459), .DIN2(_37460), .Q(_37438) );
  nnd2s1 _37358_inst ( .DIN1(_53285), .DIN2(_37461), .Q(_37460) );
  or2s1 _37359_inst ( .DIN1(_37462), .DIN2(_37463), .Q(_37461) );
  nnd2s1 _37360_inst ( .DIN1(_37463), .DIN2(_37462), .Q(_37459) );
  hi1s1 _37361_inst ( .DIN(_37437), .Q(_37440) );
  hi1s1 _37362_inst ( .DIN(_37394), .Q(_32861) );
  nnd2s1 _37363_inst ( .DIN1(_37464), .DIN2(_36688), .Q(_37394) );
  hi1s1 _37364_inst ( .DIN(_36662), .Q(_36688) );
  nnd2s1 _37365_inst ( .DIN1(_37465), .DIN2(_37466), .Q(_36662) );
  nor2s1 _37366_inst ( .DIN1(_37467), .DIN2(_36695), .Q(_37465) );
  nor2s1 _37367_inst ( .DIN1(_32878), .DIN2(_37468), .Q(_37464) );
  hi1s1 _37368_inst ( .DIN(_32855), .Q(_32878) );
  nnd2s1 _37369_inst ( .DIN1(_36748), .DIN2(_37445), .Q(_32855) );
  hi1s1 _37370_inst ( .DIN(_36736), .Q(_36748) );
  nnd2s1 _37371_inst ( .DIN1(_37469), .DIN2(_37470), .Q(_36736) );
  nor2s1 _37372_inst ( .DIN1(_37467), .DIN2(_37471), .Q(_37469) );
  nor2s1 _37373_inst ( .DIN1(_53347), .DIN2(_29560), .Q(_37450) );
  nnd2s1 _37374_inst ( .DIN1(_37472), .DIN2(_37473), .Q(
        _____________________________156________) );
  nnd2s1 _37375_inst ( .DIN1(_37474), .DIN2(_33149), .Q(_37473) );
  nor2s1 _37376_inst ( .DIN1(_26400), .DIN2(_37475), .Q(_37474) );
  nnd2s1 _37377_inst ( .DIN1(______[22]), .DIN2(_33152), .Q(_37475) );
  nnd2s1 _37378_inst ( .DIN1(_37476), .DIN2(_33132), .Q(_37472) );
  nor2s1 _37379_inst ( .DIN1(_37477), .DIN2(_37478), .Q(_37476) );
  xor2s1 _37380_inst ( .DIN1(_37463), .DIN2(_37479), .Q(_37477) );
  xor2s1 _37381_inst ( .DIN1(_26394), .DIN2(_37462), .Q(_37479) );
  nnd2s1 _37382_inst ( .DIN1(_37480), .DIN2(_37481), .Q(_37462) );
  nnd2s1 _37383_inst ( .DIN1(_37482), .DIN2(_26682), .Q(_37481) );
  xor2s1 _37384_inst ( .DIN1(_30674), .DIN2(_37483), .Q(_37482) );
  nnd2s1 _37385_inst ( .DIN1(_37484), .DIN2(_37485), .Q(
        _____________________________155________) );
  nnd2s1 _37386_inst ( .DIN1(_37486), .DIN2(_33403), .Q(_37485) );
  nor2s1 _37387_inst ( .DIN1(_37487), .DIN2(_27365), .Q(_37486) );
  xor2s1 _37388_inst ( .DIN1(_37488), .DIN2(_53335), .Q(_37487) );
  nnd2s1 _37389_inst ( .DIN1(_53255), .DIN2(_53271), .Q(_37488) );
  nnd2s1 _37390_inst ( .DIN1(_28470), .DIN2(_37489), .Q(_37484) );
  nnd2s1 _37391_inst ( .DIN1(_37490), .DIN2(_37491), .Q(_37489) );
  xor2s1 _37392_inst ( .DIN1(_37492), .DIN2(_53235), .Q(_37490) );
  nnd2s1 _37393_inst ( .DIN1(_37483), .DIN2(_37480), .Q(_37492) );
  nnd2s1 _37394_inst ( .DIN1(_37493), .DIN2(_37494), .Q(_37480) );
  or2s1 _37395_inst ( .DIN1(_37494), .DIN2(_37493), .Q(_37483) );
  nnd2s1 _37396_inst ( .DIN1(_37495), .DIN2(_37496), .Q(_37494) );
  nnd2s1 _37397_inst ( .DIN1(_37497), .DIN2(_26510), .Q(_37496) );
  or2s1 _37398_inst ( .DIN1(_37498), .DIN2(_37499), .Q(_37497) );
  nnd2s1 _37399_inst ( .DIN1(_37499), .DIN2(_37498), .Q(_37495) );
  nnd2s1 _37400_inst ( .DIN1(_37500), .DIN2(_37501), .Q(
        _____________________________154________) );
  nnd2s1 _37401_inst ( .DIN1(_37491), .DIN2(_37502), .Q(_37501) );
  xor2s1 _37402_inst ( .DIN1(_37499), .DIN2(_37503), .Q(_37502) );
  xor2s1 _37403_inst ( .DIN1(_26510), .DIN2(_37498), .Q(_37503) );
  nnd2s1 _37404_inst ( .DIN1(_37504), .DIN2(_37505), .Q(_37498) );
  nnd2s1 _37405_inst ( .DIN1(_53236), .DIN2(_37506), .Q(_37505) );
  or2s1 _37406_inst ( .DIN1(_37507), .DIN2(_37508), .Q(_37506) );
  nnd2s1 _37407_inst ( .DIN1(_37508), .DIN2(_37507), .Q(_37504) );
  hi1s1 _37408_inst ( .DIN(_37478), .Q(_37491) );
  nor2s1 _37409_inst ( .DIN1(_37509), .DIN2(_32873), .Q(
        _____________________________153________) );
  nor2s1 _37410_inst ( .DIN1(_37478), .DIN2(_37510), .Q(_37509) );
  xor2s1 _37411_inst ( .DIN1(_37508), .DIN2(_37511), .Q(_37510) );
  xnr2s1 _37412_inst ( .DIN1(_53236), .DIN2(_37507), .Q(_37511) );
  nnd2s1 _37413_inst ( .DIN1(_37512), .DIN2(_37513), .Q(_37507) );
  nnd2s1 _37414_inst ( .DIN1(_37514), .DIN2(_26445), .Q(_37513) );
  or2s1 _37415_inst ( .DIN1(_37515), .DIN2(_37516), .Q(_37514) );
  nnd2s1 _37416_inst ( .DIN1(_37516), .DIN2(_37515), .Q(_37512) );
  nnd2s1 _37417_inst ( .DIN1(_37517), .DIN2(_37518), .Q(
        _____________________________152________) );
  nnd2s1 _37418_inst ( .DIN1(_37519), .DIN2(_37520), .Q(_37518) );
  xor2s1 _37419_inst ( .DIN1(_37521), .DIN2(_37522), .Q(_37520) );
  xnr2s1 _37420_inst ( .DIN1(_37515), .DIN2(_37516), .Q(_37522) );
  nnd2s1 _37421_inst ( .DIN1(_37523), .DIN2(_37524), .Q(_37515) );
  nnd2s1 _37422_inst ( .DIN1(_53282), .DIN2(_37525), .Q(_37524) );
  or2s1 _37423_inst ( .DIN1(_37526), .DIN2(_37527), .Q(_37525) );
  nnd2s1 _37424_inst ( .DIN1(_37527), .DIN2(_37526), .Q(_37523) );
  xor2s1 _37425_inst ( .DIN1(_30186), .DIN2(_53281), .Q(_37521) );
  nor2s1 _37426_inst ( .DIN1(_37528), .DIN2(_37478), .Q(_37519) );
  nnd2s1 _37427_inst ( .DIN1(_37529), .DIN2(_53300), .Q(_37517) );
  and2s1 _37428_inst ( .DIN1(_26865), .DIN2(_28968), .Q(_37529) );
  nnd2s1 _37429_inst ( .DIN1(_37530), .DIN2(_30774), .Q(
        _____________________________151________) );
  nnd2s1 _37430_inst ( .DIN1(_34809), .DIN2(_30777), .Q(_30774) );
  nor2s1 _37431_inst ( .DIN1(_33616), .DIN2(_35699), .Q(_34809) );
  nnd2s1 _37432_inst ( .DIN1(_37531), .DIN2(_37532), .Q(_33616) );
  and2s1 _37433_inst ( .DIN1(_37533), .DIN2(_35784), .Q(_37531) );
  nor2s1 _37434_inst ( .DIN1(_37534), .DIN2(_37535), .Q(_37530) );
  nor2s1 _37435_inst ( .DIN1(_37536), .DIN2(_30777), .Q(_37535) );
  nor2s1 _37436_inst ( .DIN1(_37478), .DIN2(_37537), .Q(_37536) );
  xor2s1 _37437_inst ( .DIN1(_37527), .DIN2(_37538), .Q(_37537) );
  xnr2s1 _37438_inst ( .DIN1(_53282), .DIN2(_37526), .Q(_37538) );
  nnd2s1 _37439_inst ( .DIN1(_37539), .DIN2(_37540), .Q(_37526) );
  nnd2s1 _37440_inst ( .DIN1(_53239), .DIN2(_37541), .Q(_37540) );
  nnd2s1 _37441_inst ( .DIN1(_37542), .DIN2(_37543), .Q(_37541) );
  or2s1 _37442_inst ( .DIN1(_37543), .DIN2(_37542), .Q(_37539) );
  nnd2s1 _37443_inst ( .DIN1(_36488), .DIN2(_37466), .Q(_37478) );
  nor2s1 _37444_inst ( .DIN1(_27227), .DIN2(_37544), .Q(_37534) );
  nor2s1 _37445_inst ( .DIN1(_37545), .DIN2(_27448), .Q(_37544) );
  xnr2s1 _37446_inst ( .DIN1(_53238), .DIN2(_53237), .Q(_37545) );
  hi1s1 _37447_inst ( .DIN(_30777), .Q(_27227) );
  nnd2s1 _37448_inst ( .DIN1(_37546), .DIN2(_37547), .Q(_30777) );
  nor2s1 _37449_inst ( .DIN1(_37548), .DIN2(_37549), .Q(_37547) );
  nnd2s1 _37450_inst ( .DIN1(_37550), .DIN2(_35757), .Q(_37549) );
  nnd2s1 _37451_inst ( .DIN1(_35707), .DIN2(_37551), .Q(_37548) );
  nor2s1 _37452_inst ( .DIN1(_37552), .DIN2(_37553), .Q(_37546) );
  or2s1 _37453_inst ( .DIN1(_36612), .DIN2(_34397), .Q(_37553) );
  hi1s1 _37454_inst ( .DIN(_35708), .Q(_36612) );
  nor2s1 _37455_inst ( .DIN1(_27936), .DIN2(_34673), .Q(_35708) );
  nnd2s1 _37456_inst ( .DIN1(_37554), .DIN2(_37555), .Q(_27936) );
  nor2s1 _37457_inst ( .DIN1(_34678), .DIN2(_37556), .Q(_37554) );
  nnd2s1 _37458_inst ( .DIN1(_37533), .DIN2(_37557), .Q(_37552) );
  nnd2s1 _37459_inst ( .DIN1(_37500), .DIN2(_37558), .Q(
        _____________________________150________) );
  nnd2s1 _37460_inst ( .DIN1(_37559), .DIN2(_37560), .Q(_37558) );
  nnd2s1 _37461_inst ( .DIN1(_37561), .DIN2(_37562), .Q(_37560) );
  nnd2s1 _37462_inst ( .DIN1(_37563), .DIN2(_37564), .Q(_37562) );
  xor2s1 _37463_inst ( .DIN1(_37565), .DIN2(_37566), .Q(_37563) );
  xor2s1 _37464_inst ( .DIN1(_53197), .DIN2(_53240), .Q(_37566) );
  nor2s1 _37465_inst ( .DIN1(_53245), .DIN2(_53242), .Q(_37565) );
  nnd2s1 _37466_inst ( .DIN1(_37567), .DIN2(_37568), .Q(_37559) );
  xor2s1 _37467_inst ( .DIN1(_37542), .DIN2(_37569), .Q(_37568) );
  xnr2s1 _37468_inst ( .DIN1(_53239), .DIN2(_37543), .Q(_37569) );
  xnr2s1 _37469_inst ( .DIN1(_37570), .DIN2(_2064), .Q(_37543) );
  nnd2s1 _37470_inst ( .DIN1(_37571), .DIN2(_37572), .Q(_37570) );
  nnd2s1 _37471_inst ( .DIN1(_53300), .DIN2(_37573), .Q(_37572) );
  or2s1 _37472_inst ( .DIN1(_37574), .DIN2(_37575), .Q(_37573) );
  nnd2s1 _37473_inst ( .DIN1(_37575), .DIN2(_37574), .Q(_37571) );
  nnd2s1 _37474_inst ( .DIN1(_28253), .DIN2(_37576), .Q(
        _____________________________14________) );
  xor2s1 _37475_inst ( .DIN1(_37577), .DIN2(_37578), .Q(_37576) );
  nnd2s1 _37476_inst ( .DIN1(_37579), .DIN2(_37580), .Q(_37578) );
  nnd2s1 _37477_inst ( .DIN1(_37581), .DIN2(_36533), .Q(_37580) );
  xor2s1 _37478_inst ( .DIN1(_37376), .DIN2(_37582), .Q(_37581) );
  xnr2s1 _37479_inst ( .DIN1(_53241), .DIN2(_37374), .Q(_37582) );
  nnd2s1 _37480_inst ( .DIN1(_37583), .DIN2(_37584), .Q(_37374) );
  nnd2s1 _37481_inst ( .DIN1(_53254), .DIN2(_37585), .Q(_37584) );
  or2s1 _37482_inst ( .DIN1(_37586), .DIN2(_35427), .Q(_37585) );
  nnd2s1 _37483_inst ( .DIN1(_35427), .DIN2(_37586), .Q(_37583) );
  xor2s1 _37484_inst ( .DIN1(_37382), .DIN2(_37587), .Q(_37376) );
  xor2s1 _37485_inst ( .DIN1(_26333), .DIN2(_37381), .Q(_37587) );
  nnd2s1 _37486_inst ( .DIN1(_37588), .DIN2(_37589), .Q(_37381) );
  nnd2s1 _37487_inst ( .DIN1(_53374), .DIN2(_37590), .Q(_37589) );
  or2s1 _37488_inst ( .DIN1(_37591), .DIN2(_37592), .Q(_37590) );
  nnd2s1 _37489_inst ( .DIN1(_37592), .DIN2(_37591), .Q(_37588) );
  nnd2s1 _37490_inst ( .DIN1(_36530), .DIN2(_37593), .Q(_37579) );
  xor2s1 _37491_inst ( .DIN1(_37594), .DIN2(_37595), .Q(_37593) );
  xor2s1 _37492_inst ( .DIN1(_53035), .DIN2(_53252), .Q(_37595) );
  and2s1 _37493_inst ( .DIN1(_26290), .DIN2(_53034), .Q(_37594) );
  nnd2s1 _37494_inst ( .DIN1(_37596), .DIN2(_37597), .Q(
        _____________________________149________) );
  nnd2s1 _37495_inst ( .DIN1(_34160), .DIN2(_37598), .Q(_37597) );
  xor2s1 _37496_inst ( .DIN1(_53243), .DIN2(_53285), .Q(_37598) );
  nnd2s1 _37497_inst ( .DIN1(_37599), .DIN2(_30856), .Q(_37596) );
  nor2s1 _37498_inst ( .DIN1(_37600), .DIN2(_37601), .Q(_37599) );
  nor2s1 _37499_inst ( .DIN1(_37602), .DIN2(_37603), .Q(_37601) );
  xor2s1 _37500_inst ( .DIN1(_37575), .DIN2(_37604), .Q(_37603) );
  xnr2s1 _37501_inst ( .DIN1(_53300), .DIN2(_37574), .Q(_37604) );
  nnd2s1 _37502_inst ( .DIN1(_37605), .DIN2(_37606), .Q(_37574) );
  nnd2s1 _37503_inst ( .DIN1(_53303), .DIN2(_37607), .Q(_37606) );
  or2s1 _37504_inst ( .DIN1(_37608), .DIN2(_37609), .Q(_37607) );
  nnd2s1 _37505_inst ( .DIN1(_37609), .DIN2(_37608), .Q(_37605) );
  nor2s1 _37506_inst ( .DIN1(_37567), .DIN2(_37610), .Q(_37600) );
  nnd2s1 _37507_inst ( .DIN1(_37564), .DIN2(_26557), .Q(_37610) );
  nor2s1 _37508_inst ( .DIN1(_27749), .DIN2(_37611), .Q(
        _____________________________148________) );
  nnd2s1 _37509_inst ( .DIN1(_37612), .DIN2(_37613), .Q(_37611) );
  nnd2s1 _37510_inst ( .DIN1(_37614), .DIN2(_37602), .Q(_37613) );
  nnd2s1 _37511_inst ( .DIN1(_53240), .DIN2(_37564), .Q(_37614) );
  nnd2s1 _37512_inst ( .DIN1(_37615), .DIN2(_37567), .Q(_37612) );
  xor2s1 _37513_inst ( .DIN1(_37609), .DIN2(_37616), .Q(_37615) );
  xor2s1 _37514_inst ( .DIN1(_26601), .DIN2(_37608), .Q(_37616) );
  nnd2s1 _37515_inst ( .DIN1(_37617), .DIN2(_37618), .Q(_37608) );
  nnd2s1 _37516_inst ( .DIN1(_37619), .DIN2(_26309), .Q(_37618) );
  or2s1 _37517_inst ( .DIN1(_37620), .DIN2(_37621), .Q(_37619) );
  nnd2s1 _37518_inst ( .DIN1(_37621), .DIN2(_37620), .Q(_37617) );
  nnd2s1 _37519_inst ( .DIN1(_37622), .DIN2(_33050), .Q(
        _____________________________147________) );
  nnd2s1 _37520_inst ( .DIN1(_37623), .DIN2(_53244), .Q(_33050) );
  nor2s1 _37521_inst ( .DIN1(_33069), .DIN2(_26503), .Q(_37623) );
  nor2s1 _37522_inst ( .DIN1(_37624), .DIN2(_37625), .Q(_37622) );
  nor2s1 _37523_inst ( .DIN1(_33053), .DIN2(_37626), .Q(_37625) );
  nor2s1 _37524_inst ( .DIN1(_37627), .DIN2(_37628), .Q(_37626) );
  nor2s1 _37525_inst ( .DIN1(_37602), .DIN2(_37629), .Q(_37628) );
  xor2s1 _37526_inst ( .DIN1(_37621), .DIN2(_37630), .Q(_37629) );
  xor2s1 _37527_inst ( .DIN1(_26309), .DIN2(_37620), .Q(_37630) );
  nnd2s1 _37528_inst ( .DIN1(_37631), .DIN2(_37632), .Q(_37620) );
  nnd2s1 _37529_inst ( .DIN1(_37633), .DIN2(_26750), .Q(_37632) );
  or2s1 _37530_inst ( .DIN1(_37634), .DIN2(_37635), .Q(_37633) );
  nnd2s1 _37531_inst ( .DIN1(_37635), .DIN2(_37634), .Q(_37631) );
  nor2s1 _37532_inst ( .DIN1(_37567), .DIN2(_37636), .Q(_37627) );
  nor2s1 _37533_inst ( .DIN1(_37470), .DIN2(_37637), .Q(_37636) );
  xor2s1 _37534_inst ( .DIN1(_53240), .DIN2(_53245), .Q(_37637) );
  nor2s1 _37535_inst ( .DIN1(_33069), .DIN2(_37638), .Q(_37624) );
  nor2s1 _37536_inst ( .DIN1(_27448), .DIN2(_33071), .Q(_37638) );
  nnd2s1 _37537_inst ( .DIN1(_29039), .DIN2(_37639), .Q(_33071) );
  nnd2s1 _37538_inst ( .DIN1(_26503), .DIN2(_26287), .Q(_37639) );
  nnd2s1 _37539_inst ( .DIN1(_37640), .DIN2(_37641), .Q(
        _____________________________146________) );
  nnd2s1 _37540_inst ( .DIN1(_37642), .DIN2(_37500), .Q(_37641) );
  nor2s1 _37541_inst ( .DIN1(_37567), .DIN2(_37643), .Q(_37642) );
  nor2s1 _37542_inst ( .DIN1(_37470), .DIN2(_37644), .Q(_37643) );
  xor2s1 _37543_inst ( .DIN1(_37645), .DIN2(_37646), .Q(_37644) );
  nnd2s1 _37544_inst ( .DIN1(_37647), .DIN2(_37648), .Q(_37645) );
  or2s1 _37545_inst ( .DIN1(_26342), .DIN2(_53251), .Q(_37648) );
  nnd2s1 _37546_inst ( .DIN1(_37649), .DIN2(_37650), .Q(_37640) );
  xor2s1 _37547_inst ( .DIN1(_37651), .DIN2(_37652), .Q(_37650) );
  xor2s1 _37548_inst ( .DIN1(_37634), .DIN2(_37635), .Q(_37652) );
  nnd2s1 _37549_inst ( .DIN1(_37653), .DIN2(_37654), .Q(_37634) );
  nnd2s1 _37550_inst ( .DIN1(_37655), .DIN2(_26757), .Q(_37654) );
  or2s1 _37551_inst ( .DIN1(_37656), .DIN2(_37657), .Q(_37655) );
  nnd2s1 _37552_inst ( .DIN1(_37657), .DIN2(_37656), .Q(_37653) );
  xor2s1 _37553_inst ( .DIN1(_31947), .DIN2(_53247), .Q(_37651) );
  hi1s1 _37554_inst ( .DIN(_37561), .Q(_37649) );
  nnd2s1 _37555_inst ( .DIN1(_37567), .DIN2(_37500), .Q(_37561) );
  nnd2s1 _37556_inst ( .DIN1(_37658), .DIN2(_37500), .Q(
        _____________________________145________) );
  hi1s1 _37557_inst ( .DIN(_32873), .Q(_37500) );
  nnd2s1 _37558_inst ( .DIN1(_33359), .DIN2(_27828), .Q(_32873) );
  nor2s1 _37559_inst ( .DIN1(_37659), .DIN2(_37660), .Q(_37658) );
  nor2s1 _37560_inst ( .DIN1(_37602), .DIN2(_37661), .Q(_37660) );
  xor2s1 _37561_inst ( .DIN1(_37657), .DIN2(_37662), .Q(_37661) );
  xor2s1 _37562_inst ( .DIN1(_37656), .DIN2(_53248), .Q(_37662) );
  nnd2s1 _37563_inst ( .DIN1(_37663), .DIN2(_37664), .Q(_37656) );
  nnd2s1 _37564_inst ( .DIN1(_53310), .DIN2(_37665), .Q(_37664) );
  or2s1 _37565_inst ( .DIN1(_37666), .DIN2(_37667), .Q(_37665) );
  nnd2s1 _37566_inst ( .DIN1(_37667), .DIN2(_37666), .Q(_37663) );
  nor2s1 _37567_inst ( .DIN1(_37567), .DIN2(_37668), .Q(_37659) );
  nnd2s1 _37568_inst ( .DIN1(_37669), .DIN2(______[18]), .Q(_37668) );
  nor2s1 _37569_inst ( .DIN1(_53249), .DIN2(_37470), .Q(_37669) );
  hi1s1 _37570_inst ( .DIN(_37564), .Q(_37470) );
  nnd2s1 _37571_inst ( .DIN1(_37466), .DIN2(_37670), .Q(_37564) );
  hi1s1 _37572_inst ( .DIN(_37671), .Q(_37466) );
  hi1s1 _37573_inst ( .DIN(_37602), .Q(_37567) );
  nnd2s1 _37574_inst ( .DIN1(_37672), .DIN2(_36693), .Q(_37602) );
  nor2s1 _37575_inst ( .DIN1(_37467), .DIN2(_37673), .Q(_37672) );
  nnd2s1 _37576_inst ( .DIN1(_37674), .DIN2(_28284), .Q(
        _____________________________144________) );
  nnd2s1 _37577_inst ( .DIN1(_27606), .DIN2(_27144), .Q(_28284) );
  nor2s1 _37578_inst ( .DIN1(_37675), .DIN2(_37676), .Q(_37674) );
  nor2s1 _37579_inst ( .DIN1(_27144), .DIN2(_37677), .Q(_37676) );
  nnd2s1 _37580_inst ( .DIN1(_37678), .DIN2(_37679), .Q(_37677) );
  nnd2s1 _37581_inst ( .DIN1(_53251), .DIN2(_37680), .Q(_37679) );
  nnd2s1 _37582_inst ( .DIN1(_37681), .DIN2(_37682), .Q(_37678) );
  xor2s1 _37583_inst ( .DIN1(_37683), .DIN2(_37684), .Q(_37682) );
  xnr2s1 _37584_inst ( .DIN1(_53310), .DIN2(_37666), .Q(_37684) );
  nnd2s1 _37585_inst ( .DIN1(_37685), .DIN2(_37686), .Q(_37666) );
  nnd2s1 _37586_inst ( .DIN1(_37687), .DIN2(_26555), .Q(_37686) );
  or2s1 _37587_inst ( .DIN1(_37688), .DIN2(_37689), .Q(_37687) );
  nnd2s1 _37588_inst ( .DIN1(_37689), .DIN2(_37688), .Q(_37685) );
  hi1s1 _37589_inst ( .DIN(_37667), .Q(_37683) );
  nor2s1 _37590_inst ( .DIN1(_27146), .DIN2(_37690), .Q(_37675) );
  nor2s1 _37591_inst ( .DIN1(_27241), .DIN2(_37691), .Q(_37690) );
  xor2s1 _37592_inst ( .DIN1(_52879), .DIN2(_53250), .Q(_37691) );
  hi1s1 _37593_inst ( .DIN(_27144), .Q(_27146) );
  nnd2s1 _37594_inst ( .DIN1(_37692), .DIN2(_28253), .Q(_27144) );
  nor2s1 _37595_inst ( .DIN1(_35510), .DIN2(_35342), .Q(_37692) );
  nnd2s1 _37596_inst ( .DIN1(_37693), .DIN2(_37694), .Q(
        _____________________________143________) );
  nnd2s1 _37597_inst ( .DIN1(_37695), .DIN2(_33149), .Q(_37694) );
  nnd2s1 _37598_inst ( .DIN1(_37696), .DIN2(_37697), .Q(_37695) );
  nnd2s1 _37599_inst ( .DIN1(_26400), .DIN2(_26260), .Q(_37697) );
  nor2s1 _37600_inst ( .DIN1(_33714), .DIN2(_33683), .Q(_37696) );
  nnd2s1 _37601_inst ( .DIN1(_37698), .DIN2(_33132), .Q(_37693) );
  hi1s1 _37602_inst ( .DIN(_33149), .Q(_33132) );
  nnd2s1 _37603_inst ( .DIN1(_37699), .DIN2(_37700), .Q(_33149) );
  nor2s1 _37604_inst ( .DIN1(_31809), .DIN2(_37701), .Q(_37700) );
  nor2s1 _37605_inst ( .DIN1(_33182), .DIN2(_37702), .Q(_37699) );
  nor2s1 _37606_inst ( .DIN1(_37703), .DIN2(_37704), .Q(_37698) );
  nor2s1 _37607_inst ( .DIN1(_37705), .DIN2(_37706), .Q(_37704) );
  nnd2s1 _37608_inst ( .DIN1(______[26]), .DIN2(_37707), .Q(_37706) );
  nnd2s1 _37609_inst ( .DIN1(_37646), .DIN2(_26342), .Q(_37707) );
  and2s1 _37610_inst ( .DIN1(_53251), .DIN2(_53246), .Q(_37646) );
  nnd2s1 _37611_inst ( .DIN1(_37708), .DIN2(_37680), .Q(_37705) );
  nnd2s1 _37612_inst ( .DIN1(_37647), .DIN2(_26549), .Q(_37708) );
  nnd2s1 _37613_inst ( .DIN1(_53251), .DIN2(_26342), .Q(_37647) );
  nor2s1 _37614_inst ( .DIN1(_37709), .DIN2(_37710), .Q(_37703) );
  hi1s1 _37615_inst ( .DIN(_37681), .Q(_37710) );
  xnr2s1 _37616_inst ( .DIN1(_37689), .DIN2(_37711), .Q(_37709) );
  xor2s1 _37617_inst ( .DIN1(_26555), .DIN2(_37688), .Q(_37711) );
  nnd2s1 _37618_inst ( .DIN1(_37712), .DIN2(_37713), .Q(_37688) );
  nnd2s1 _37619_inst ( .DIN1(_53325), .DIN2(_37714), .Q(_37713) );
  or2s1 _37620_inst ( .DIN1(_37715), .DIN2(_37716), .Q(_37714) );
  nnd2s1 _37621_inst ( .DIN1(_37716), .DIN2(_37715), .Q(_37712) );
  nnd2s1 _37622_inst ( .DIN1(_37717), .DIN2(_37718), .Q(
        _____________________________142________) );
  nor2s1 _37623_inst ( .DIN1(_37719), .DIN2(_37720), .Q(_37718) );
  nor2s1 _37624_inst ( .DIN1(_37721), .DIN2(_37722), .Q(_37720) );
  xor2s1 _37625_inst ( .DIN1(_53271), .DIN2(_37723), .Q(_37722) );
  nor2s1 _37626_inst ( .DIN1(_37724), .DIN2(_37725), .Q(_37717) );
  nor2s1 _37627_inst ( .DIN1(_37726), .DIN2(_37727), .Q(_37725) );
  xor2s1 _37628_inst ( .DIN1(_37716), .DIN2(_37728), .Q(_37727) );
  xnr2s1 _37629_inst ( .DIN1(_53325), .DIN2(_37715), .Q(_37728) );
  nnd2s1 _37630_inst ( .DIN1(_37729), .DIN2(_37730), .Q(_37715) );
  nnd2s1 _37631_inst ( .DIN1(_53324), .DIN2(_37731), .Q(_37730) );
  or2s1 _37632_inst ( .DIN1(_37732), .DIN2(_37733), .Q(_37731) );
  nnd2s1 _37633_inst ( .DIN1(_37733), .DIN2(_37732), .Q(_37729) );
  nor2s1 _37634_inst ( .DIN1(_37734), .DIN2(_37735), .Q(_37724) );
  xor2s1 _37635_inst ( .DIN1(_37736), .DIN2(_53257), .Q(_37735) );
  nnd2s1 _37636_inst ( .DIN1(_37737), .DIN2(_37738), .Q(
        _____________________________141________) );
  nor2s1 _37637_inst ( .DIN1(_37739), .DIN2(_37740), .Q(_37738) );
  nor2s1 _37638_inst ( .DIN1(_53204), .DIN2(_37741), .Q(_37740) );
  nor2s1 _37639_inst ( .DIN1(_37742), .DIN2(_37743), .Q(_37741) );
  nor2s1 _37640_inst ( .DIN1(_37734), .DIN2(_37736), .Q(_37743) );
  nor2s1 _37641_inst ( .DIN1(_53263), .DIN2(_37721), .Q(_37742) );
  nor2s1 _37642_inst ( .DIN1(_37744), .DIN2(_26597), .Q(_37739) );
  nor2s1 _37643_inst ( .DIN1(_37745), .DIN2(_37746), .Q(_37744) );
  nor2s1 _37644_inst ( .DIN1(_37747), .DIN2(_37734), .Q(_37746) );
  nor2s1 _37645_inst ( .DIN1(_26523), .DIN2(_37721), .Q(_37745) );
  nnd2s1 _37646_inst ( .DIN1(_37734), .DIN2(_37680), .Q(_37721) );
  nor2s1 _37647_inst ( .DIN1(_37719), .DIN2(_37748), .Q(_37737) );
  nor2s1 _37648_inst ( .DIN1(_37749), .DIN2(_37726), .Q(_37748) );
  xor2s1 _37649_inst ( .DIN1(_37733), .DIN2(_37750), .Q(_37749) );
  xor2s1 _37650_inst ( .DIN1(_26456), .DIN2(_37732), .Q(_37750) );
  nnd2s1 _37651_inst ( .DIN1(_37751), .DIN2(_37752), .Q(_37732) );
  nnd2s1 _37652_inst ( .DIN1(_53326), .DIN2(_37753), .Q(_37752) );
  or2s1 _37653_inst ( .DIN1(_37754), .DIN2(_37755), .Q(_37753) );
  nnd2s1 _37654_inst ( .DIN1(_37755), .DIN2(_37754), .Q(_37751) );
  nnd2s1 _37655_inst ( .DIN1(_37756), .DIN2(_37757), .Q(
        _____________________________140________) );
  nor2s1 _37656_inst ( .DIN1(_37719), .DIN2(_37758), .Q(_37757) );
  nor2s1 _37657_inst ( .DIN1(_53262), .DIN2(_37759), .Q(_37758) );
  nor2s1 _37658_inst ( .DIN1(_37680), .DIN2(_37760), .Q(_37759) );
  nor2s1 _37659_inst ( .DIN1(_37761), .DIN2(_37762), .Q(_37756) );
  nor2s1 _37660_inst ( .DIN1(______[0]), .DIN2(_37734), .Q(_37762) );
  nor2s1 _37661_inst ( .DIN1(_37763), .DIN2(_37726), .Q(_37761) );
  nnd2s1 _37662_inst ( .DIN1(_37734), .DIN2(_37681), .Q(_37726) );
  xor2s1 _37663_inst ( .DIN1(_37755), .DIN2(_37764), .Q(_37763) );
  xor2s1 _37664_inst ( .DIN1(_26400), .DIN2(_37754), .Q(_37764) );
  nnd2s1 _37665_inst ( .DIN1(_37765), .DIN2(_37766), .Q(_37754) );
  nnd2s1 _37666_inst ( .DIN1(_37767), .DIN2(_26284), .Q(_37766) );
  or2s1 _37667_inst ( .DIN1(_37768), .DIN2(_37769), .Q(_37767) );
  nnd2s1 _37668_inst ( .DIN1(_37769), .DIN2(_37768), .Q(_37765) );
  nnd2s1 _37669_inst ( .DIN1(_37770), .DIN2(_37771), .Q(
        _____________________________13________) );
  nnd2s1 _37670_inst ( .DIN1(_37772), .DIN2(_32830), .Q(_37771) );
  nnd2s1 _37671_inst ( .DIN1(_37773), .DIN2(_36777), .Q(_37772) );
  xnr2s1 _37672_inst ( .DIN1(_32833), .DIN2(_53228), .Q(_37773) );
  nor2s1 _37673_inst ( .DIN1(_26521), .DIN2(_26290), .Q(_32833) );
  nnd2s1 _37674_inst ( .DIN1(_37774), .DIN2(_32837), .Q(_37770) );
  nor2s1 _37675_inst ( .DIN1(_37775), .DIN2(_37776), .Q(_37774) );
  nnd2s1 _37676_inst ( .DIN1(_37777), .DIN2(_37105), .Q(_37776) );
  nnd2s1 _37677_inst ( .DIN1(_36810), .DIN2(_37778), .Q(_37105) );
  nnd2s1 _37678_inst ( .DIN1(_37779), .DIN2(_37780), .Q(_37777) );
  hi1s1 _37679_inst ( .DIN(_36810), .Q(_37780) );
  xor2s1 _37680_inst ( .DIN1(_35427), .DIN2(_37781), .Q(_37779) );
  xnr2s1 _37681_inst ( .DIN1(_53254), .DIN2(_37586), .Q(_37781) );
  nnd2s1 _37682_inst ( .DIN1(_37782), .DIN2(_37783), .Q(_37586) );
  nnd2s1 _37683_inst ( .DIN1(_37784), .DIN2(_26488), .Q(_37783) );
  or2s1 _37684_inst ( .DIN1(_37785), .DIN2(_35443), .Q(_37784) );
  nnd2s1 _37685_inst ( .DIN1(_35443), .DIN2(_37785), .Q(_37782) );
  xnr2s1 _37686_inst ( .DIN1(_37592), .DIN2(_26813), .Q(_35427) );
  nnd2s1 _37687_inst ( .DIN1(_37787), .DIN2(_37788), .Q(_37591) );
  nnd2s1 _37688_inst ( .DIN1(_53372), .DIN2(_37789), .Q(_37788) );
  or2s1 _37689_inst ( .DIN1(_37790), .DIN2(_37791), .Q(_37789) );
  nnd2s1 _37690_inst ( .DIN1(_37791), .DIN2(_37790), .Q(_37787) );
  nor2s1 _37691_inst ( .DIN1(_53034), .DIN2(_36533), .Q(_37775) );
  hi1s1 _37692_inst ( .DIN(_36804), .Q(_36533) );
  xnr2s1 _37693_inst ( .DIN1(_36810), .DIN2(_37792), .Q(_36804) );
  nnd2s1 _37694_inst ( .DIN1(_37793), .DIN2(_27721), .Q(_36810) );
  xor2s1 _37695_inst ( .DIN1(_37794), .DIN2(_32005), .Q(_27721) );
  nnd2s1 _37696_inst ( .DIN1(_34913), .DIN2(_37778), .Q(_37794) );
  and2s1 _37697_inst ( .DIN1(_36308), .DIN2(_36336), .Q(_37793) );
  nnd2s1 _37698_inst ( .DIN1(_37795), .DIN2(_37796), .Q(
        _____________________________139________) );
  nnd2s1 _37699_inst ( .DIN1(_28470), .DIN2(_37797), .Q(_37796) );
  nnd2s1 _37700_inst ( .DIN1(_37798), .DIN2(_37799), .Q(_37797) );
  nnd2s1 _37701_inst ( .DIN1(_37800), .DIN2(_37801), .Q(_37799) );
  and2s1 _37702_inst ( .DIN1(_37736), .DIN2(_37680), .Q(_37801) );
  nor2s1 _37703_inst ( .DIN1(_37723), .DIN2(_28646), .Q(_37800) );
  nnd2s1 _37704_inst ( .DIN1(_37681), .DIN2(_37802), .Q(_37798) );
  xor2s1 _37705_inst ( .DIN1(_37769), .DIN2(_37803), .Q(_37802) );
  xor2s1 _37706_inst ( .DIN1(_26284), .DIN2(_37768), .Q(_37803) );
  nnd2s1 _37707_inst ( .DIN1(_37804), .DIN2(_37805), .Q(_37768) );
  nnd2s1 _37708_inst ( .DIN1(_37806), .DIN2(_26447), .Q(_37805) );
  or2s1 _37709_inst ( .DIN1(_37807), .DIN2(_37808), .Q(_37806) );
  nnd2s1 _37710_inst ( .DIN1(_37808), .DIN2(_37807), .Q(_37804) );
  nor2s1 _37711_inst ( .DIN1(_37680), .DIN2(_37471), .Q(_37681) );
  nnd2s1 _37712_inst ( .DIN1(_37809), .DIN2(_37810), .Q(_37680) );
  nor2s1 _37713_inst ( .DIN1(_37467), .DIN2(_37468), .Q(_37809) );
  nnd2s1 _37714_inst ( .DIN1(_37811), .DIN2(_28467), .Q(_37795) );
  nnd2s1 _37715_inst ( .DIN1(_37812), .DIN2(_53255), .Q(_37811) );
  nor2s1 _37716_inst ( .DIN1(_28182), .DIN2(_27651), .Q(_37812) );
  nnd2s1 _37717_inst ( .DIN1(_37813), .DIN2(_33335), .Q(
        _____________________________138________) );
  nnd2s1 _37718_inst ( .DIN1(_33338), .DIN2(_30174), .Q(_33335) );
  nor2s1 _37719_inst ( .DIN1(_37814), .DIN2(_37815), .Q(_37813) );
  nor2s1 _37720_inst ( .DIN1(_30175), .DIN2(_37816), .Q(_37815) );
  nor2s1 _37721_inst ( .DIN1(_27082), .DIN2(_37817), .Q(_37816) );
  nnd2s1 _37722_inst ( .DIN1(_37818), .DIN2(_37068), .Q(_37817) );
  nnd2s1 _37723_inst ( .DIN1(_53256), .DIN2(_53211), .Q(_37068) );
  nnd2s1 _37724_inst ( .DIN1(_26272), .DIN2(_26718), .Q(_37818) );
  nor2s1 _37725_inst ( .DIN1(_37819), .DIN2(_33338), .Q(_37814) );
  nor2s1 _37726_inst ( .DIN1(_37820), .DIN2(_37821), .Q(_37819) );
  nor2s1 _37727_inst ( .DIN1(_37822), .DIN2(_37445), .Q(_37821) );
  xor2s1 _37728_inst ( .DIN1(_26255), .DIN2(_53257), .Q(_37822) );
  nor2s1 _37729_inst ( .DIN1(_37823), .DIN2(_37824), .Q(_37820) );
  xnr2s1 _37730_inst ( .DIN1(_37808), .DIN2(_37825), .Q(_37823) );
  xor2s1 _37731_inst ( .DIN1(_26447), .DIN2(_37807), .Q(_37825) );
  nnd2s1 _37732_inst ( .DIN1(_37826), .DIN2(_37827), .Q(_37807) );
  nnd2s1 _37733_inst ( .DIN1(_37828), .DIN2(_26553), .Q(_37827) );
  or2s1 _37734_inst ( .DIN1(_37829), .DIN2(_37830), .Q(_37828) );
  xor2s1 _37735_inst ( .DIN1(_37831), .DIN2(_37832), .Q(_37826) );
  xor2s1 _37736_inst ( .DIN1(_31456), .DIN2(_37577), .Q(_37832) );
  nnd2s1 _37737_inst ( .DIN1(_37830), .DIN2(_37829), .Q(_37831) );
  nnd2s1 _37738_inst ( .DIN1(_37833), .DIN2(_37834), .Q(
        _____________________________137________) );
  nnd2s1 _37739_inst ( .DIN1(_27007), .DIN2(_37835), .Q(_37834) );
  nnd2s1 _37740_inst ( .DIN1(_37836), .DIN2(_37837), .Q(_37835) );
  nor2s1 _37741_inst ( .DIN1(_37838), .DIN2(_37839), .Q(_37837) );
  nor2s1 _37742_inst ( .DIN1(_37824), .DIN2(_37840), .Q(_37839) );
  xor2s1 _37743_inst ( .DIN1(_37830), .DIN2(_37841), .Q(_37840) );
  xor2s1 _37744_inst ( .DIN1(_26553), .DIN2(_37829), .Q(_37841) );
  nnd2s1 _37745_inst ( .DIN1(_37842), .DIN2(_37843), .Q(_37829) );
  nnd2s1 _37746_inst ( .DIN1(_53261), .DIN2(_37844), .Q(_37843) );
  or2s1 _37747_inst ( .DIN1(_37845), .DIN2(_37846), .Q(_37844) );
  nnd2s1 _37748_inst ( .DIN1(_37846), .DIN2(_37845), .Q(_37842) );
  nor2s1 _37749_inst ( .DIN1(_36693), .DIN2(_37847), .Q(_37838) );
  nor2s1 _37750_inst ( .DIN1(_37848), .DIN2(_27039), .Q(_37847) );
  nor2s1 _37751_inst ( .DIN1(_53260), .DIN2(_53264), .Q(_37848) );
  nor2s1 _37752_inst ( .DIN1(_37849), .DIN2(_37850), .Q(_37836) );
  nor2s1 _37753_inst ( .DIN1(_26610), .DIN2(_37851), .Q(_37850) );
  hi1s1 _37754_inst ( .DIN(_37852), .Q(_37849) );
  hi1s1 _37755_inst ( .DIN(_26996), .Q(_27007) );
  nnd2s1 _37756_inst ( .DIN1(_37853), .DIN2(_26996), .Q(_37833) );
  nnd2s1 _37757_inst ( .DIN1(_33683), .DIN2(_37854), .Q(_26996) );
  hi1s1 _37758_inst ( .DIN(_33152), .Q(_33683) );
  nor2s1 _37759_inst ( .DIN1(_35961), .DIN2(_37855), .Q(_37853) );
  xor2s1 _37760_inst ( .DIN1(_26236), .DIN2(_37856), .Q(_37855) );
  nnd2s1 _37761_inst ( .DIN1(_53259), .DIN2(_53258), .Q(_37856) );
  and2s1 _37762_inst ( .DIN1(_37857), .DIN2(_37240), .Q(_35961) );
  nor2s1 _37763_inst ( .DIN1(_36302), .DIN2(_31809), .Q(_37240) );
  nor2s1 _37764_inst ( .DIN1(_34490), .DIN2(_33182), .Q(_37857) );
  nnd2s1 _37765_inst ( .DIN1(_37858), .DIN2(_27994), .Q(
        _____________________________136________) );
  nor2s1 _37766_inst ( .DIN1(_37859), .DIN2(_37860), .Q(_37858) );
  nor2s1 _37767_inst ( .DIN1(_37861), .DIN2(_37824), .Q(_37860) );
  xor2s1 _37768_inst ( .DIN1(_37846), .DIN2(_37862), .Q(_37861) );
  xor2s1 _37769_inst ( .DIN1(_26503), .DIN2(_37845), .Q(_37862) );
  nnd2s1 _37770_inst ( .DIN1(_37863), .DIN2(_37864), .Q(_37845) );
  nnd2s1 _37771_inst ( .DIN1(_37865), .DIN2(_26357), .Q(_37864) );
  or2s1 _37772_inst ( .DIN1(_37866), .DIN2(_37867), .Q(_37865) );
  nnd2s1 _37773_inst ( .DIN1(_37867), .DIN2(_37866), .Q(_37863) );
  nor2s1 _37774_inst ( .DIN1(_37445), .DIN2(_37868), .Q(_37859) );
  nnd2s1 _37775_inst ( .DIN1(_53260), .DIN2(______[28]), .Q(_37868) );
  nnd2s1 _37776_inst ( .DIN1(_37869), .DIN2(_37870), .Q(
        _____________________________135________) );
  nnd2s1 _37777_inst ( .DIN1(_37734), .DIN2(_37871), .Q(_37870) );
  nnd2s1 _37778_inst ( .DIN1(_37852), .DIN2(_37851), .Q(_37871) );
  nnd2s1 _37779_inst ( .DIN1(_37872), .DIN2(_53264), .Q(_37851) );
  nor2s1 _37780_inst ( .DIN1(_36693), .DIN2(_26255), .Q(_37872) );
  nnd2s1 _37781_inst ( .DIN1(_37873), .DIN2(_37824), .Q(_37852) );
  nnd2s1 _37782_inst ( .DIN1(_37468), .DIN2(_37874), .Q(_37873) );
  nnd2s1 _37783_inst ( .DIN1(_26255), .DIN2(_26566), .Q(_37874) );
  nor2s1 _37784_inst ( .DIN1(_37875), .DIN2(_37876), .Q(_37869) );
  nor2s1 _37785_inst ( .DIN1(_37877), .DIN2(_37878), .Q(_37876) );
  xor2s1 _37786_inst ( .DIN1(_37867), .DIN2(_37879), .Q(_37877) );
  xor2s1 _37787_inst ( .DIN1(_26357), .DIN2(_37866), .Q(_37879) );
  nnd2s1 _37788_inst ( .DIN1(_37880), .DIN2(_37881), .Q(_37866) );
  nnd2s1 _37789_inst ( .DIN1(_37882), .DIN2(_26344), .Q(_37881) );
  or2s1 _37790_inst ( .DIN1(_37883), .DIN2(_37884), .Q(_37882) );
  nnd2s1 _37791_inst ( .DIN1(_37884), .DIN2(_37883), .Q(_37880) );
  nor2s1 _37792_inst ( .DIN1(_37885), .DIN2(_37886), .Q(_37875) );
  nnd2s1 _37793_inst ( .DIN1(_37887), .DIN2(______[22]), .Q(_37886) );
  or2s1 _37794_inst ( .DIN1(_37723), .DIN2(_37747), .Q(_37885) );
  hi1s1 _37795_inst ( .DIN(_37736), .Q(_37747) );
  nnd2s1 _37796_inst ( .DIN1(_53263), .DIN2(_53262), .Q(_37736) );
  nor2s1 _37797_inst ( .DIN1(_53262), .DIN2(_53263), .Q(_37723) );
  nnd2s1 _37798_inst ( .DIN1(_37888), .DIN2(_28238), .Q(
        _____________________________134________) );
  nor2s1 _37799_inst ( .DIN1(_37889), .DIN2(_37890), .Q(_37888) );
  nor2s1 _37800_inst ( .DIN1(_28241), .DIN2(_37891), .Q(_37890) );
  nnd2s1 _37801_inst ( .DIN1(_37892), .DIN2(_37893), .Q(_37891) );
  nnd2s1 _37802_inst ( .DIN1(_37894), .DIN2(_37468), .Q(_37893) );
  xor2s1 _37803_inst ( .DIN1(_26375), .DIN2(_37895), .Q(_37894) );
  nor2s1 _37804_inst ( .DIN1(_53269), .DIN2(_53266), .Q(_37895) );
  xor2s1 _37805_inst ( .DIN1(_27329), .DIN2(_37896), .Q(_37892) );
  nnd2s1 _37806_inst ( .DIN1(_37897), .DIN2(_36693), .Q(_37896) );
  xor2s1 _37807_inst ( .DIN1(_37884), .DIN2(_37898), .Q(_37897) );
  xor2s1 _37808_inst ( .DIN1(_26344), .DIN2(_37883), .Q(_37898) );
  nnd2s1 _37809_inst ( .DIN1(_37899), .DIN2(_37900), .Q(_37883) );
  nnd2s1 _37810_inst ( .DIN1(_53340), .DIN2(_37901), .Q(_37900) );
  or2s1 _37811_inst ( .DIN1(_37902), .DIN2(_37903), .Q(_37901) );
  nnd2s1 _37812_inst ( .DIN1(_37903), .DIN2(_37902), .Q(_37899) );
  nor2s1 _37813_inst ( .DIN1(_28250), .DIN2(_37904), .Q(_37889) );
  and2s1 _37814_inst ( .DIN1(______[0]), .DIN2(_53267), .Q(_37904) );
  nnd2s1 _37815_inst ( .DIN1(_37905), .DIN2(_37906), .Q(
        _____________________________133________) );
  nor2s1 _37816_inst ( .DIN1(_37907), .DIN2(_37908), .Q(_37906) );
  nor2s1 _37817_inst ( .DIN1(_37760), .DIN2(_37909), .Q(_37908) );
  nnd2s1 _37818_inst ( .DIN1(_37468), .DIN2(_37910), .Q(_37909) );
  xor2s1 _37819_inst ( .DIN1(_53268), .DIN2(_26385), .Q(_37910) );
  nor2s1 _37820_inst ( .DIN1(_37734), .DIN2(_37911), .Q(_37907) );
  xor2s1 _37821_inst ( .DIN1(_37912), .DIN2(_53191), .Q(_37911) );
  nnd2s1 _37822_inst ( .DIN1(_53269), .DIN2(_53270), .Q(_37912) );
  nor2s1 _37823_inst ( .DIN1(_37719), .DIN2(_37913), .Q(_37905) );
  nor2s1 _37824_inst ( .DIN1(_37878), .DIN2(_37914), .Q(_37913) );
  xor2s1 _37825_inst ( .DIN1(_37903), .DIN2(_37915), .Q(_37914) );
  xnr2s1 _37826_inst ( .DIN1(_53340), .DIN2(_37902), .Q(_37915) );
  nnd2s1 _37827_inst ( .DIN1(_37916), .DIN2(_37917), .Q(_37902) );
  nnd2s1 _37828_inst ( .DIN1(_53349), .DIN2(_37918), .Q(_37917) );
  or2s1 _37829_inst ( .DIN1(_37919), .DIN2(_37920), .Q(_37918) );
  xor2s1 _37830_inst ( .DIN1(_31947), .DIN2(_37921), .Q(_37916) );
  nnd2s1 _37831_inst ( .DIN1(_37920), .DIN2(_37919), .Q(_37921) );
  nnd2s1 _37832_inst ( .DIN1(_31802), .DIN2(_37922), .Q(_31947) );
  nnd2s1 _37833_inst ( .DIN1(_37734), .DIN2(_36693), .Q(_37878) );
  hi1s1 _37834_inst ( .DIN(_37824), .Q(_36693) );
  nnd2s1 _37835_inst ( .DIN1(_37923), .DIN2(_37445), .Q(_37824) );
  and2s1 _37836_inst ( .DIN1(_37924), .DIN2(_31109), .Q(_37719) );
  nor2s1 _37837_inst ( .DIN1(_36829), .DIN2(_37734), .Q(_37924) );
  nnd2s1 _37838_inst ( .DIN1(_37925), .DIN2(_37926), .Q(
        _____________________________132________) );
  nnd2s1 _37839_inst ( .DIN1(_37887), .DIN2(_37927), .Q(_37926) );
  xor2s1 _37840_inst ( .DIN1(_53266), .DIN2(_53270), .Q(_37927) );
  and2s1 _37841_inst ( .DIN1(_37760), .DIN2(_37928), .Q(_37887) );
  nnd2s1 _37842_inst ( .DIN1(_31109), .DIN2(_36832), .Q(_37928) );
  hi1s1 _37843_inst ( .DIN(_31173), .Q(_31109) );
  nnd2s1 _37844_inst ( .DIN1(_37929), .DIN2(_37930), .Q(_31173) );
  nor2s1 _37845_inst ( .DIN1(_31196), .DIN2(_37931), .Q(_37929) );
  nnd2s1 _37846_inst ( .DIN1(_37734), .DIN2(_37932), .Q(_37925) );
  nnd2s1 _37847_inst ( .DIN1(_36488), .DIN2(_37933), .Q(_37932) );
  xor2s1 _37848_inst ( .DIN1(_37920), .DIN2(_37934), .Q(_37933) );
  xor2s1 _37849_inst ( .DIN1(_53349), .DIN2(_37919), .Q(_37934) );
  xor2s1 _37850_inst ( .DIN1(_37935), .DIN2(_31975), .Q(_37919) );
  nnd2s1 _37851_inst ( .DIN1(_37936), .DIN2(_37937), .Q(_37935) );
  nnd2s1 _37852_inst ( .DIN1(_37938), .DIN2(_26678), .Q(_37937) );
  or2s1 _37853_inst ( .DIN1(_37939), .DIN2(_32867), .Q(_37938) );
  nnd2s1 _37854_inst ( .DIN1(_32867), .DIN2(_37939), .Q(_37936) );
  hi1s1 _37855_inst ( .DIN(_37760), .Q(_37734) );
  nnd2s1 _37856_inst ( .DIN1(_27827), .DIN2(_36832), .Q(_37760) );
  nor2s1 _37857_inst ( .DIN1(_37940), .DIN2(_37941), .Q(_27827) );
  nnd2s1 _37858_inst ( .DIN1(_37942), .DIN2(_37299), .Q(_37940) );
  nnd2s1 _37859_inst ( .DIN1(_37943), .DIN2(_37944), .Q(
        _____________________________131________) );
  nnd2s1 _37860_inst ( .DIN1(_33403), .DIN2(_37945), .Q(_37944) );
  xor2s1 _37861_inst ( .DIN1(_53271), .DIN2(_53335), .Q(_37945) );
  nor2s1 _37862_inst ( .DIN1(_28182), .DIN2(_28470), .Q(_33403) );
  nnd2s1 _37863_inst ( .DIN1(_28470), .DIN2(_37946), .Q(_37943) );
  nnd2s1 _37864_inst ( .DIN1(_37947), .DIN2(_36488), .Q(_37946) );
  xor2s1 _37865_inst ( .DIN1(_32867), .DIN2(_37948), .Q(_37947) );
  xor2s1 _37866_inst ( .DIN1(_26678), .DIN2(_37939), .Q(_37948) );
  nnd2s1 _37867_inst ( .DIN1(_37949), .DIN2(_37950), .Q(_37939) );
  nnd2s1 _37868_inst ( .DIN1(_37951), .DIN2(_26613), .Q(_37950) );
  nnd2s1 _37869_inst ( .DIN1(_37952), .DIN2(_37953), .Q(_37951) );
  nnd2s1 _37870_inst ( .DIN1(_37954), .DIN2(_32880), .Q(_37949) );
  hi1s1 _37871_inst ( .DIN(_28467), .Q(_28470) );
  nnd2s1 _37872_inst ( .DIN1(_37955), .DIN2(_34090), .Q(_28467) );
  nnd2s1 _37873_inst ( .DIN1(_37956), .DIN2(_37957), .Q(
        _____________________________130________) );
  nnd2s1 _37874_inst ( .DIN1(_29096), .DIN2(_37958), .Q(_37957) );
  nnd2s1 _37875_inst ( .DIN1(_37959), .DIN2(_36488), .Q(_37958) );
  xor2s1 _37876_inst ( .DIN1(_37960), .DIN2(_32880), .Q(_37959) );
  xor2s1 _37877_inst ( .DIN1(_37953), .DIN2(_53344), .Q(_37960) );
  nnd2s1 _37878_inst ( .DIN1(_29094), .DIN2(_52875), .Q(_37956) );
  nor2s1 _37879_inst ( .DIN1(_29096), .DIN2(_27123), .Q(_29094) );
  nor2s1 _37880_inst ( .DIN1(_37961), .DIN2(_27161), .Q(_27123) );
  hi1s1 _37881_inst ( .DIN(_34707), .Q(_29096) );
  nnd2s1 _37882_inst ( .DIN1(_37962), .DIN2(_37963), .Q(_34707) );
  nor2s1 _37883_inst ( .DIN1(_37961), .DIN2(_37129), .Q(_37962) );
  nnd2s1 _37884_inst ( .DIN1(_37964), .DIN2(_37965), .Q(
        _____________________________12________) );
  nnd2s1 _37885_inst ( .DIN1(_32837), .DIN2(_37966), .Q(_37965) );
  nnd2s1 _37886_inst ( .DIN1(_37967), .DIN2(_33044), .Q(_37966) );
  xor2s1 _37887_inst ( .DIN1(_35443), .DIN2(_37968), .Q(_37967) );
  xor2s1 _37888_inst ( .DIN1(_26488), .DIN2(_37785), .Q(_37968) );
  nnd2s1 _37889_inst ( .DIN1(_37969), .DIN2(_37970), .Q(_37785) );
  nnd2s1 _37890_inst ( .DIN1(_53295), .DIN2(_37971), .Q(_37970) );
  nnd2s1 _37891_inst ( .DIN1(_37972), .DIN2(_35482), .Q(_37971) );
  nnd2s1 _37892_inst ( .DIN1(_35459), .DIN2(_37973), .Q(_37969) );
  hi1s1 _37893_inst ( .DIN(_35482), .Q(_35459) );
  xor2s1 _37894_inst ( .DIN1(_37974), .DIN2(_37975), .Q(_35443) );
  xor2s1 _37895_inst ( .DIN1(_26336), .DIN2(_37790), .Q(_37975) );
  nnd2s1 _37896_inst ( .DIN1(_37976), .DIN2(_37977), .Q(_37790) );
  nnd2s1 _37897_inst ( .DIN1(_53338), .DIN2(_37978), .Q(_37977) );
  or2s1 _37898_inst ( .DIN1(_37979), .DIN2(_37980), .Q(_37978) );
  nnd2s1 _37899_inst ( .DIN1(_37980), .DIN2(_37979), .Q(_37976) );
  nnd2s1 _37900_inst ( .DIN1(_33039), .DIN2(_53252), .Q(_37964) );
  nor2s1 _37901_inst ( .DIN1(_32834), .DIN2(_32837), .Q(_33039) );
  hi1s1 _37902_inst ( .DIN(_32830), .Q(_32837) );
  nnd2s1 _37903_inst ( .DIN1(_31193), .DIN2(_37981), .Q(_32830) );
  nor2s1 _37904_inst ( .DIN1(_27821), .DIN2(_36828), .Q(_37981) );
  nor2s1 _37905_inst ( .DIN1(_37941), .DIN2(_37153), .Q(_31193) );
  hi1s1 _37906_inst ( .DIN(_36927), .Q(_37153) );
  nor2s1 _37907_inst ( .DIN1(_33295), .DIN2(_37931), .Q(_36927) );
  nnd2s1 _37908_inst ( .DIN1(_37982), .DIN2(_37983), .Q(_33295) );
  nnd2s1 _37909_inst ( .DIN1(_37984), .DIN2(_33293), .Q(_37941) );
  hi1s1 _37910_inst ( .DIN(_36777), .Q(_32834) );
  nnd2s1 _37911_inst ( .DIN1(_37985), .DIN2(_37986), .Q(_36777) );
  nor2s1 _37912_inst ( .DIN1(_37987), .DIN2(_36828), .Q(_37985) );
  nnd2s1 _37913_inst ( .DIN1(_37988), .DIN2(_37989), .Q(
        _____________________________129________) );
  nnd2s1 _37914_inst ( .DIN1(_37990), .DIN2(_30298), .Q(_37989) );
  hi1s1 _37915_inst ( .DIN(_27182), .Q(_30298) );
  nnd2s1 _37916_inst ( .DIN1(_30129), .DIN2(_28084), .Q(_27182) );
  nor2s1 _37917_inst ( .DIN1(_37991), .DIN2(_26988), .Q(_37990) );
  xor2s1 _37918_inst ( .DIN1(_26377), .DIN2(_53273), .Q(_37991) );
  nnd2s1 _37919_inst ( .DIN1(_27183), .DIN2(_37992), .Q(_37988) );
  nnd2s1 _37920_inst ( .DIN1(_37993), .DIN2(_36488), .Q(_37992) );
  hi1s1 _37921_inst ( .DIN(_36513), .Q(_36488) );
  nnd2s1 _37922_inst ( .DIN1(_37994), .DIN2(_37995), .Q(_36513) );
  nor2s1 _37923_inst ( .DIN1(_37471), .DIN2(_37673), .Q(_37994) );
  nor2s1 _37924_inst ( .DIN1(_37954), .DIN2(_37996), .Q(_37993) );
  nor2s1 _37925_inst ( .DIN1(_53275), .DIN2(_37997), .Q(_37996) );
  hi1s1 _37926_inst ( .DIN(_37953), .Q(_37954) );
  nnd2s1 _37927_inst ( .DIN1(_53275), .DIN2(_37997), .Q(_37953) );
  nnd2s1 _37928_inst ( .DIN1(_37998), .DIN2(_28811), .Q(
        _____________________________128________) );
  nnd2s1 _37929_inst ( .DIN1(_33992), .DIN2(_28814), .Q(_28811) );
  hi1s1 _37930_inst ( .DIN(_28364), .Q(_33992) );
  nnd2s1 _37931_inst ( .DIN1(_34580), .DIN2(_37532), .Q(_28364) );
  hi1s1 _37932_inst ( .DIN(_37999), .Q(_37532) );
  nor2s1 _37933_inst ( .DIN1(_38000), .DIN2(_38001), .Q(_37998) );
  nor2s1 _37934_inst ( .DIN1(_28814), .DIN2(_38002), .Q(_38001) );
  nnd2s1 _37935_inst ( .DIN1(_38003), .DIN2(_38004), .Q(_38002) );
  nnd2s1 _37936_inst ( .DIN1(_38005), .DIN2(_53277), .Q(_38004) );
  nor2s1 _37937_inst ( .DIN1(_33571), .DIN2(_28100), .Q(_38005) );
  nor2s1 _37938_inst ( .DIN1(_38006), .DIN2(_38007), .Q(_38003) );
  nor2s1 _37939_inst ( .DIN1(_26743), .DIN2(_38008), .Q(_38007) );
  nor2s1 _37940_inst ( .DIN1(_38009), .DIN2(_38010), .Q(_38008) );
  nor2s1 _37941_inst ( .DIN1(_33578), .DIN2(_38011), .Q(_38010) );
  nor2s1 _37942_inst ( .DIN1(_38012), .DIN2(_33577), .Q(_38009) );
  nor2s1 _37943_inst ( .DIN1(_53276), .DIN2(_38013), .Q(_38006) );
  nor2s1 _37944_inst ( .DIN1(_38014), .DIN2(_38015), .Q(_38013) );
  nor2s1 _37945_inst ( .DIN1(_33577), .DIN2(_38011), .Q(_38015) );
  nnd2s1 _37946_inst ( .DIN1(_32916), .DIN2(_26850), .Q(_33577) );
  nor2s1 _37947_inst ( .DIN1(_38012), .DIN2(_33578), .Q(_38014) );
  nnd2s1 _37948_inst ( .DIN1(_32916), .DIN2(_26849), .Q(_33578) );
  hi1s1 _37949_inst ( .DIN(_34223), .Q(_32916) );
  nnd2s1 _37950_inst ( .DIN1(_38016), .DIN2(_33571), .Q(_34223) );
  nor2s1 _37951_inst ( .DIN1(_38017), .DIN2(_38018), .Q(_38016) );
  hi1s1 _37952_inst ( .DIN(_38011), .Q(_38012) );
  nnd2s1 _37953_inst ( .DIN1(_38019), .DIN2(_38020), .Q(_38011) );
  nnd2s1 _37954_inst ( .DIN1(_38021), .DIN2(_26367), .Q(_38020) );
  nnd2s1 _37955_inst ( .DIN1(_37359), .DIN2(_38022), .Q(_38021) );
  or2s1 _37956_inst ( .DIN1(_38022), .DIN2(_37359), .Q(_38019) );
  nor2s1 _37957_inst ( .DIN1(_28356), .DIN2(_38023), .Q(_38000) );
  xor2s1 _37958_inst ( .DIN1(_38024), .DIN2(_52971), .Q(_38023) );
  nnd2s1 _37959_inst ( .DIN1(_53279), .DIN2(_53278), .Q(_38024) );
  hi1s1 _37960_inst ( .DIN(_28814), .Q(_28356) );
  nnd2s1 _37961_inst ( .DIN1(_38025), .DIN2(_38026), .Q(_28814) );
  nor2s1 _37962_inst ( .DIN1(_33617), .DIN2(_34602), .Q(_38026) );
  hi1s1 _37963_inst ( .DIN(_36585), .Q(_33617) );
  nnd2s1 _37964_inst ( .DIN1(_38027), .DIN2(_38028), .Q(_36585) );
  nor2s1 _37965_inst ( .DIN1(_37999), .DIN2(_36613), .Q(_38025) );
  nnd2s1 _37966_inst ( .DIN1(_37557), .DIN2(_35694), .Q(_37999) );
  nnd2s1 _37967_inst ( .DIN1(_38029), .DIN2(_28794), .Q(
        _____________________________127________) );
  or2s1 _37968_inst ( .DIN1(_32985), .DIN2(_28797), .Q(_28794) );
  nnd2s1 _37969_inst ( .DIN1(_38030), .DIN2(_28182), .Q(_32985) );
  nor2s1 _37970_inst ( .DIN1(_38031), .DIN2(_35998), .Q(_38030) );
  nor2s1 _37971_inst ( .DIN1(_38032), .DIN2(_38033), .Q(_38029) );
  nor2s1 _37972_inst ( .DIN1(_28801), .DIN2(_38034), .Q(_38033) );
  nnd2s1 _37973_inst ( .DIN1(_38035), .DIN2(_38036), .Q(_38034) );
  nnd2s1 _37974_inst ( .DIN1(_38037), .DIN2(_33536), .Q(_38036) );
  xnr2s1 _37975_inst ( .DIN1(_37359), .DIN2(_38038), .Q(_38037) );
  xor2s1 _37976_inst ( .DIN1(_26367), .DIN2(_38022), .Q(_38038) );
  nnd2s1 _37977_inst ( .DIN1(_38039), .DIN2(_38040), .Q(_38022) );
  nnd2s1 _37978_inst ( .DIN1(_38041), .DIN2(_26740), .Q(_38040) );
  nnd2s1 _37979_inst ( .DIN1(_37430), .DIN2(_38042), .Q(_38041) );
  or2s1 _37980_inst ( .DIN1(_38042), .DIN2(_37430), .Q(_38039) );
  xor2s1 _37981_inst ( .DIN1(_38043), .DIN2(_35087), .Q(_37359) );
  xor2s1 _37982_inst ( .DIN1(_35082), .DIN2(_38044), .Q(_35087) );
  nor2s1 _37983_inst ( .DIN1(_38045), .DIN2(_38046), .Q(_38044) );
  nor2s1 _37984_inst ( .DIN1(_26850), .DIN2(_38047), .Q(_38046) );
  nor2s1 _37985_inst ( .DIN1(_53364), .DIN2(_38048), .Q(_38045) );
  and2s1 _37986_inst ( .DIN1(_38047), .DIN2(_26850), .Q(_38048) );
  nnd2s1 _37987_inst ( .DIN1(_35059), .DIN2(_35056), .Q(_35082) );
  nnd2s1 _37988_inst ( .DIN1(_26849), .DIN2(_53363), .Q(_35056) );
  nnd2s1 _37989_inst ( .DIN1(_26335), .DIN2(_26850), .Q(_35059) );
  xor2s1 _37990_inst ( .DIN1(_38049), .DIN2(_53384), .Q(_38043) );
  nnd2s1 _37991_inst ( .DIN1(_38050), .DIN2(_38051), .Q(_38049) );
  nnd2s1 _37992_inst ( .DIN1(_26849), .DIN2(_38052), .Q(_38051) );
  nnd2s1 _37993_inst ( .DIN1(_38053), .DIN2(_38054), .Q(_38052) );
  or2s1 _37994_inst ( .DIN1(_38054), .DIN2(_38053), .Q(_38050) );
  hi1s1 _37995_inst ( .DIN(_35129), .Q(_38053) );
  nnd2s1 _37996_inst ( .DIN1(_38055), .DIN2(_38056), .Q(_38035) );
  hi1s1 _37997_inst ( .DIN(_33550), .Q(_38056) );
  nnd2s1 _37998_inst ( .DIN1(_33531), .DIN2(_38057), .Q(_33550) );
  nnd2s1 _37999_inst ( .DIN1(_38058), .DIN2(_33519), .Q(_38057) );
  nor2s1 _38000_inst ( .DIN1(_38059), .DIN2(_27291), .Q(_38055) );
  xnr2s1 _38001_inst ( .DIN1(_38060), .DIN2(_38061), .Q(_38059) );
  nnd2s1 _38002_inst ( .DIN1(_38062), .DIN2(_38063), .Q(_38060) );
  nnd2s1 _38003_inst ( .DIN1(_53286), .DIN2(_26394), .Q(_38063) );
  nor2s1 _38004_inst ( .DIN1(_28797), .DIN2(_38064), .Q(_38032) );
  nor2s1 _38005_inst ( .DIN1(_36509), .DIN2(_38065), .Q(_38064) );
  nnd2s1 _38006_inst ( .DIN1(_38066), .DIN2(_38067), .Q(_38065) );
  nnd2s1 _38007_inst ( .DIN1(_26213), .DIN2(_26224), .Q(_38067) );
  nnd2s1 _38008_inst ( .DIN1(_38068), .DIN2(_53284), .Q(_38066) );
  nor2s1 _38009_inst ( .DIN1(_26445), .DIN2(_26213), .Q(_38068) );
  nnd2s1 _38010_inst ( .DIN1(______[4]), .DIN2(_38069), .Q(_36509) );
  nnd2s1 _38011_inst ( .DIN1(_26224), .DIN2(_26445), .Q(_38069) );
  hi1s1 _38012_inst ( .DIN(_28801), .Q(_28797) );
  nnd2s1 _38013_inst ( .DIN1(_32292), .DIN2(_28792), .Q(_28801) );
  hi1s1 _38014_inst ( .DIN(_28786), .Q(_28792) );
  nnd2s1 _38015_inst ( .DIN1(_38070), .DIN2(_34090), .Q(_28786) );
  nor2s1 _38016_inst ( .DIN1(_36492), .DIN2(_38071), .Q(_38070) );
  nor2s1 _38017_inst ( .DIN1(_38072), .DIN2(_38031), .Q(_32292) );
  nnd2s1 _38018_inst ( .DIN1(_38073), .DIN2(_38074), .Q(
        _____________________________126________) );
  nnd2s1 _38019_inst ( .DIN1(_38075), .DIN2(_38076), .Q(_38074) );
  xor2s1 _38020_inst ( .DIN1(_38077), .DIN2(_38078), .Q(_38076) );
  xor2s1 _38021_inst ( .DIN1(_38042), .DIN2(_37435), .Q(_38078) );
  hi1s1 _38022_inst ( .DIN(_37430), .Q(_37435) );
  xor2s1 _38023_inst ( .DIN1(_35129), .DIN2(_38079), .Q(_37430) );
  xor2s1 _38024_inst ( .DIN1(_26850), .DIN2(_38054), .Q(_38079) );
  nnd2s1 _38025_inst ( .DIN1(_38080), .DIN2(_38081), .Q(_38054) );
  nnd2s1 _38026_inst ( .DIN1(_38082), .DIN2(_26850), .Q(_38081) );
  or2s1 _38027_inst ( .DIN1(_38083), .DIN2(_35169), .Q(_38082) );
  nnd2s1 _38028_inst ( .DIN1(_35169), .DIN2(_38083), .Q(_38080) );
  xnr2s1 _38029_inst ( .DIN1(_36565), .DIN2(_38047), .Q(_35129) );
  nnd2s1 _38030_inst ( .DIN1(_38084), .DIN2(_38085), .Q(_38047) );
  nnd2s1 _38031_inst ( .DIN1(_38086), .DIN2(_26338), .Q(_38085) );
  or2s1 _38032_inst ( .DIN1(_38087), .DIN2(_26335), .Q(_38086) );
  nnd2s1 _38033_inst ( .DIN1(_38087), .DIN2(_26335), .Q(_38084) );
  xor2s1 _38034_inst ( .DIN1(_27620), .DIN2(_53384), .Q(_36565) );
  nnd2s1 _38035_inst ( .DIN1(_38088), .DIN2(_38089), .Q(_38042) );
  nnd2s1 _38036_inst ( .DIN1(_53283), .DIN2(_38090), .Q(_38089) );
  nnd2s1 _38037_inst ( .DIN1(_37437), .DIN2(_38091), .Q(_38090) );
  or2s1 _38038_inst ( .DIN1(_38091), .DIN2(_37437), .Q(_38088) );
  xor2s1 _38039_inst ( .DIN1(_35291), .DIN2(_53462), .Q(_38077) );
  hi1s1 _38040_inst ( .DIN(_38092), .Q(_38075) );
  nor2s1 _38041_inst ( .DIN1(_38093), .DIN2(_38094), .Q(_38073) );
  nor2s1 _38042_inst ( .DIN1(_38095), .DIN2(_33356), .Q(_38094) );
  nor2s1 _38043_inst ( .DIN1(_38096), .DIN2(_38097), .Q(_38095) );
  hi1s1 _38044_inst ( .DIN(_33528), .Q(_38097) );
  nor2s1 _38045_inst ( .DIN1(_33536), .DIN2(_38098), .Q(_38096) );
  nor2s1 _38046_inst ( .DIN1(_27365), .DIN2(_26213), .Q(_38098) );
  nor2s1 _38047_inst ( .DIN1(_38099), .DIN2(_38100), .Q(_38093) );
  nnd2s1 _38048_inst ( .DIN1(_33422), .DIN2(______[2]), .Q(_38100) );
  hi1s1 _38049_inst ( .DIN(_38101), .Q(_33422) );
  xor2s1 _38050_inst ( .DIN1(_53282), .DIN2(_38102), .Q(_38099) );
  nnd2s1 _38051_inst ( .DIN1(_38103), .DIN2(_38104), .Q(
        _____________________________125________) );
  nnd2s1 _38052_inst ( .DIN1(_33359), .DIN2(_38105), .Q(_38104) );
  nnd2s1 _38053_inst ( .DIN1(_33528), .DIN2(_38106), .Q(_38105) );
  nnd2s1 _38054_inst ( .DIN1(_53286), .DIN2(_33531), .Q(_38106) );
  nor2s1 _38055_inst ( .DIN1(_38107), .DIN2(_38108), .Q(_38103) );
  nor2s1 _38056_inst ( .DIN1(_38109), .DIN2(_38092), .Q(_38108) );
  nnd2s1 _38057_inst ( .DIN1(_33536), .DIN2(_33359), .Q(_38092) );
  xor2s1 _38058_inst ( .DIN1(_37437), .DIN2(_38110), .Q(_38109) );
  xor2s1 _38059_inst ( .DIN1(_26420), .DIN2(_38091), .Q(_38110) );
  nnd2s1 _38060_inst ( .DIN1(_38111), .DIN2(_38112), .Q(_38091) );
  nnd2s1 _38061_inst ( .DIN1(_38113), .DIN2(_26224), .Q(_38112) );
  or2s1 _38062_inst ( .DIN1(_38114), .DIN2(_37463), .Q(_38113) );
  nnd2s1 _38063_inst ( .DIN1(_37463), .DIN2(_38114), .Q(_38111) );
  xor2s1 _38064_inst ( .DIN1(_35169), .DIN2(_38115), .Q(_37437) );
  xor2s1 _38065_inst ( .DIN1(_26850), .DIN2(_38083), .Q(_38115) );
  nnd2s1 _38066_inst ( .DIN1(_38116), .DIN2(_38117), .Q(_38083) );
  nnd2s1 _38067_inst ( .DIN1(_38118), .DIN2(_26850), .Q(_38117) );
  or2s1 _38068_inst ( .DIN1(_38119), .DIN2(_35189), .Q(_38118) );
  nnd2s1 _38069_inst ( .DIN1(_38119), .DIN2(_35189), .Q(_38116) );
  xor2s1 _38070_inst ( .DIN1(_38087), .DIN2(_38120), .Q(_35169) );
  nnd2s1 _38071_inst ( .DIN1(_38121), .DIN2(_38122), .Q(_38087) );
  nnd2s1 _38072_inst ( .DIN1(_38123), .DIN2(_34515), .Q(_38122) );
  nnd2s1 _38073_inst ( .DIN1(_38124), .DIN2(_53364), .Q(_38123) );
  nor2s1 _38074_inst ( .DIN1(_38101), .DIN2(_38125), .Q(_38107) );
  nnd2s1 _38075_inst ( .DIN1(______[12]), .DIN2(_38126), .Q(_38125) );
  xor2s1 _38076_inst ( .DIN1(_53286), .DIN2(_53298), .Q(_38126) );
  nnd2s1 _38077_inst ( .DIN1(_38127), .DIN2(_38128), .Q(
        _____________________________124________) );
  nnd2s1 _38078_inst ( .DIN1(_30856), .DIN2(_38129), .Q(_38128) );
  nnd2s1 _38079_inst ( .DIN1(_38130), .DIN2(_33528), .Q(_38129) );
  nnd2s1 _38080_inst ( .DIN1(_38131), .DIN2(_38058), .Q(_33528) );
  nor2s1 _38081_inst ( .DIN1(_38132), .DIN2(_38133), .Q(_38058) );
  nor2s1 _38082_inst ( .DIN1(_33536), .DIN2(_33281), .Q(_38131) );
  nor2s1 _38083_inst ( .DIN1(_38134), .DIN2(_38135), .Q(_38130) );
  nor2s1 _38084_inst ( .DIN1(_33531), .DIN2(_38136), .Q(_38135) );
  xor2s1 _38085_inst ( .DIN1(_37463), .DIN2(_38137), .Q(_38136) );
  xor2s1 _38086_inst ( .DIN1(_26224), .DIN2(_38114), .Q(_38137) );
  nnd2s1 _38087_inst ( .DIN1(_38138), .DIN2(_38139), .Q(_38114) );
  nnd2s1 _38088_inst ( .DIN1(_38140), .DIN2(_26281), .Q(_38139) );
  or2s1 _38089_inst ( .DIN1(_38141), .DIN2(_37493), .Q(_38140) );
  nnd2s1 _38090_inst ( .DIN1(_37493), .DIN2(_38141), .Q(_38138) );
  xnr2s1 _38091_inst ( .DIN1(_38142), .DIN2(_38119), .Q(_37463) );
  nnd2s1 _38092_inst ( .DIN1(_38143), .DIN2(_38144), .Q(_38119) );
  nnd2s1 _38093_inst ( .DIN1(_38145), .DIN2(_26850), .Q(_38144) );
  nnd2s1 _38094_inst ( .DIN1(_38146), .DIN2(_35598), .Q(_38145) );
  hi1s1 _38095_inst ( .DIN(_35386), .Q(_35598) );
  nnd2s1 _38096_inst ( .DIN1(_35386), .DIN2(_38147), .Q(_38143) );
  xor2s1 _38097_inst ( .DIN1(_26850), .DIN2(_35381), .Q(_38142) );
  hi1s1 _38098_inst ( .DIN(_35189), .Q(_35381) );
  nnd2s1 _38099_inst ( .DIN1(_38148), .DIN2(_38149), .Q(_35189) );
  nnd2s1 _38100_inst ( .DIN1(_38150), .DIN2(_38124), .Q(_38149) );
  nor2s1 _38101_inst ( .DIN1(_38151), .DIN2(_38152), .Q(_38148) );
  nor2s1 _38102_inst ( .DIN1(_34515), .DIN2(_38153), .Q(_38152) );
  xor2s1 _38103_inst ( .DIN1(_27620), .DIN2(_38124), .Q(_38153) );
  hi1s1 _38104_inst ( .DIN(_38154), .Q(_38124) );
  nor2s1 _38105_inst ( .DIN1(_53361), .DIN2(_38121), .Q(_38151) );
  nnd2s1 _38106_inst ( .DIN1(_38154), .DIN2(_27620), .Q(_38121) );
  nnd2s1 _38107_inst ( .DIN1(_38155), .DIN2(_38156), .Q(_38154) );
  nnd2s1 _38108_inst ( .DIN1(_53362), .DIN2(_38157), .Q(_38156) );
  or2s1 _38109_inst ( .DIN1(_38158), .DIN2(_53365), .Q(_38157) );
  nnd2s1 _38110_inst ( .DIN1(_53365), .DIN2(_38158), .Q(_38155) );
  nor2s1 _38111_inst ( .DIN1(_33536), .DIN2(_38159), .Q(_38134) );
  nor2s1 _38112_inst ( .DIN1(_38160), .DIN2(_38161), .Q(_38159) );
  nor2s1 _38113_inst ( .DIN1(_26394), .DIN2(_38061), .Q(_38161) );
  nnd2s1 _38114_inst ( .DIN1(_26436), .DIN2(_26266), .Q(_38061) );
  and2s1 _38115_inst ( .DIN1(_38062), .DIN2(_53297), .Q(_38160) );
  nnd2s1 _38116_inst ( .DIN1(_53285), .DIN2(_26436), .Q(_38062) );
  nnd2s1 _38117_inst ( .DIN1(_34160), .DIN2(_26658), .Q(_38127) );
  nor2s1 _38118_inst ( .DIN1(_30856), .DIN2(_33743), .Q(_34160) );
  hi1s1 _38119_inst ( .DIN(_30854), .Q(_33743) );
  nnd2s1 _38120_inst ( .DIN1(_38162), .DIN2(_38163), .Q(_30854) );
  hi1s1 _38121_inst ( .DIN(_30853), .Q(_30856) );
  nnd2s1 _38122_inst ( .DIN1(_38164), .DIN2(_36388), .Q(_30853) );
  nor2s1 _38123_inst ( .DIN1(_38165), .DIN2(_38166), .Q(_38164) );
  nnd2s1 _38124_inst ( .DIN1(_38167), .DIN2(_38168), .Q(
        _____________________________123________) );
  nnd2s1 _38125_inst ( .DIN1(_38169), .DIN2(_38170), .Q(_38168) );
  xor2s1 _38126_inst ( .DIN1(_37493), .DIN2(_38171), .Q(_38170) );
  xor2s1 _38127_inst ( .DIN1(_26281), .DIN2(_38141), .Q(_38171) );
  nnd2s1 _38128_inst ( .DIN1(_38172), .DIN2(_38173), .Q(_38141) );
  nnd2s1 _38129_inst ( .DIN1(_38174), .DIN2(_26423), .Q(_38173) );
  or2s1 _38130_inst ( .DIN1(_38175), .DIN2(_37499), .Q(_38174) );
  nnd2s1 _38131_inst ( .DIN1(_37499), .DIN2(_38175), .Q(_38172) );
  xor2s1 _38132_inst ( .DIN1(_35386), .DIN2(_38176), .Q(_37493) );
  xor2s1 _38133_inst ( .DIN1(_53384), .DIN2(_38146), .Q(_38176) );
  hi1s1 _38134_inst ( .DIN(_38147), .Q(_38146) );
  nnd2s1 _38135_inst ( .DIN1(_38177), .DIN2(_38178), .Q(_38147) );
  nnd2s1 _38136_inst ( .DIN1(_38179), .DIN2(_26850), .Q(_38178) );
  or2s1 _38137_inst ( .DIN1(_38180), .DIN2(_35603), .Q(_38179) );
  nnd2s1 _38138_inst ( .DIN1(_35603), .DIN2(_38180), .Q(_38177) );
  xor2s1 _38139_inst ( .DIN1(_38158), .DIN2(_38181), .Q(_35386) );
  xor2s1 _38140_inst ( .DIN1(_53362), .DIN2(_53365), .Q(_38181) );
  nnd2s1 _38141_inst ( .DIN1(_38182), .DIN2(_38183), .Q(_38158) );
  nnd2s1 _38142_inst ( .DIN1(_53361), .DIN2(_38184), .Q(_38183) );
  nnd2s1 _38143_inst ( .DIN1(_38185), .DIN2(_26780), .Q(_38184) );
  nnd2s1 _38144_inst ( .DIN1(_26781), .DIN2(_38186), .Q(_38182) );
  nor2s1 _38145_inst ( .DIN1(_29555), .DIN2(_38187), .Q(_38169) );
  nnd2s1 _38146_inst ( .DIN1(_38188), .DIN2(_29039), .Q(_38167) );
  nor2s1 _38147_inst ( .DIN1(_38189), .DIN2(_27241), .Q(_38188) );
  xor2s1 _38148_inst ( .DIN1(_26497), .DIN2(_53289), .Q(_38189) );
  nnd2s1 _38149_inst ( .DIN1(_38190), .DIN2(_38191), .Q(
        _____________________________122________) );
  nnd2s1 _38150_inst ( .DIN1(_38192), .DIN2(_53297), .Q(_38191) );
  nor2s1 _38151_inst ( .DIN1(_26772), .DIN2(_38101), .Q(_38192) );
  nnd2s1 _38152_inst ( .DIN1(_33357), .DIN2(_33356), .Q(_38101) );
  nnd2s1 _38153_inst ( .DIN1(_33359), .DIN2(_38193), .Q(_38190) );
  nnd2s1 _38154_inst ( .DIN1(_38194), .DIN2(_38195), .Q(_38193) );
  xor2s1 _38155_inst ( .DIN1(_37499), .DIN2(_38196), .Q(_38195) );
  xor2s1 _38156_inst ( .DIN1(_26423), .DIN2(_38175), .Q(_38196) );
  nnd2s1 _38157_inst ( .DIN1(_38197), .DIN2(_38198), .Q(_38175) );
  nnd2s1 _38158_inst ( .DIN1(_53293), .DIN2(_38199), .Q(_38198) );
  or2s1 _38159_inst ( .DIN1(_38200), .DIN2(_37508), .Q(_38199) );
  nnd2s1 _38160_inst ( .DIN1(_37508), .DIN2(_38200), .Q(_38197) );
  xor2s1 _38161_inst ( .DIN1(_35603), .DIN2(_38201), .Q(_37499) );
  xor2s1 _38162_inst ( .DIN1(_26803), .DIN2(_38180), .Q(_38201) );
  nnd2s1 _38163_inst ( .DIN1(_38202), .DIN2(_38203), .Q(_38180) );
  nnd2s1 _38164_inst ( .DIN1(_38204), .DIN2(_26850), .Q(_38203) );
  or2s1 _38165_inst ( .DIN1(_38205), .DIN2(_35861), .Q(_38204) );
  nnd2s1 _38166_inst ( .DIN1(_35861), .DIN2(_38205), .Q(_38202) );
  xnr2s1 _38167_inst ( .DIN1(_38206), .DIN2(_26776), .Q(_35603) );
  hi1s1 _38168_inst ( .DIN(_38186), .Q(_38185) );
  nnd2s1 _38169_inst ( .DIN1(_38208), .DIN2(_38209), .Q(_38186) );
  nnd2s1 _38170_inst ( .DIN1(_38210), .DIN2(_26331), .Q(_38209) );
  or2s1 _38171_inst ( .DIN1(_38211), .DIN2(_53367), .Q(_38210) );
  nnd2s1 _38172_inst ( .DIN1(_53367), .DIN2(_38211), .Q(_38208) );
  hi1s1 _38173_inst ( .DIN(_38212), .Q(_29231) );
  xor2s1 _38174_inst ( .DIN1(_34515), .DIN2(_53368), .Q(_38206) );
  nnd2s1 _38175_inst ( .DIN1(_38213), .DIN2(_38214), .Q(
        _____________________________121________) );
  nor2s1 _38176_inst ( .DIN1(_38215), .DIN2(_38216), .Q(_38213) );
  nor2s1 _38177_inst ( .DIN1(_38217), .DIN2(_37528), .Q(_38216) );
  nor2s1 _38178_inst ( .DIN1(_38187), .DIN2(_38218), .Q(_38217) );
  xor2s1 _38179_inst ( .DIN1(_37508), .DIN2(_38219), .Q(_38218) );
  xor2s1 _38180_inst ( .DIN1(_26570), .DIN2(_38200), .Q(_38219) );
  nnd2s1 _38181_inst ( .DIN1(_38220), .DIN2(_38221), .Q(_38200) );
  nnd2s1 _38182_inst ( .DIN1(_38222), .DIN2(_26412), .Q(_38221) );
  or2s1 _38183_inst ( .DIN1(_38223), .DIN2(_37516), .Q(_38222) );
  nnd2s1 _38184_inst ( .DIN1(_37516), .DIN2(_38223), .Q(_38220) );
  xor2s1 _38185_inst ( .DIN1(_35861), .DIN2(_38224), .Q(_37508) );
  xor2s1 _38186_inst ( .DIN1(_26803), .DIN2(_38205), .Q(_38224) );
  nnd2s1 _38187_inst ( .DIN1(_38225), .DIN2(_38226), .Q(_38205) );
  nnd2s1 _38188_inst ( .DIN1(_38227), .DIN2(_26850), .Q(_38226) );
  or2s1 _38189_inst ( .DIN1(_38228), .DIN2(_36111), .Q(_38227) );
  nnd2s1 _38190_inst ( .DIN1(_36111), .DIN2(_38228), .Q(_38225) );
  hi1s1 _38191_inst ( .DIN(_36110), .Q(_36111) );
  xnr2s1 _38192_inst ( .DIN1(_38211), .DIN2(_38229), .Q(_35861) );
  nnd2s1 _38193_inst ( .DIN1(_38230), .DIN2(_38231), .Q(_38211) );
  nnd2s1 _38194_inst ( .DIN1(_53309), .DIN2(_38232), .Q(_38231) );
  or2s1 _38195_inst ( .DIN1(_38233), .DIN2(_26780), .Q(_38232) );
  nnd2s1 _38196_inst ( .DIN1(_38233), .DIN2(_26780), .Q(_38230) );
  nor2s1 _38197_inst ( .DIN1(_28971), .DIN2(_38234), .Q(_38215) );
  nor2s1 _38198_inst ( .DIN1(_38235), .DIN2(_27291), .Q(_38234) );
  xnr2s1 _38199_inst ( .DIN1(_53292), .DIN2(_53036), .Q(_38235) );
  nnd2s1 _38200_inst ( .DIN1(_38236), .DIN2(_36504), .Q(
        _____________________________120________) );
  nor2s1 _38201_inst ( .DIN1(_38237), .DIN2(_38238), .Q(_38236) );
  nor2s1 _38202_inst ( .DIN1(_36511), .DIN2(_38239), .Q(_38238) );
  nnd2s1 _38203_inst ( .DIN1(_38194), .DIN2(_38240), .Q(_38239) );
  xor2s1 _38204_inst ( .DIN1(_37516), .DIN2(_38241), .Q(_38240) );
  xor2s1 _38205_inst ( .DIN1(_26412), .DIN2(_38223), .Q(_38241) );
  nnd2s1 _38206_inst ( .DIN1(_38242), .DIN2(_38243), .Q(_38223) );
  nnd2s1 _38207_inst ( .DIN1(_53296), .DIN2(_38244), .Q(_38243) );
  or2s1 _38208_inst ( .DIN1(_38245), .DIN2(_37527), .Q(_38244) );
  nnd2s1 _38209_inst ( .DIN1(_37527), .DIN2(_38245), .Q(_38242) );
  hi1s1 _38210_inst ( .DIN(_38246), .Q(_37527) );
  xnr2s1 _38211_inst ( .DIN1(_36110), .DIN2(_38247), .Q(_37516) );
  xor2s1 _38212_inst ( .DIN1(_26803), .DIN2(_38228), .Q(_38247) );
  nnd2s1 _38213_inst ( .DIN1(_38248), .DIN2(_38249), .Q(_38228) );
  nnd2s1 _38214_inst ( .DIN1(_38250), .DIN2(_26335), .Q(_38249) );
  or2s1 _38215_inst ( .DIN1(_38251), .DIN2(_36333), .Q(_38250) );
  nnd2s1 _38216_inst ( .DIN1(_36333), .DIN2(_38251), .Q(_38248) );
  xnr2s1 _38217_inst ( .DIN1(_38252), .DIN2(_38233), .Q(_36110) );
  nnd2s1 _38218_inst ( .DIN1(_38253), .DIN2(_38254), .Q(_38233) );
  nnd2s1 _38219_inst ( .DIN1(_53314), .DIN2(_38255), .Q(_38254) );
  or2s1 _38220_inst ( .DIN1(_38256), .DIN2(_26209), .Q(_38255) );
  nnd2s1 _38221_inst ( .DIN1(_38256), .DIN2(_26209), .Q(_38253) );
  xor2s1 _38222_inst ( .DIN1(_26526), .DIN2(_26781), .Q(_38252) );
  nor2s1 _38223_inst ( .DIN1(_35940), .DIN2(_38257), .Q(_38237) );
  nor2s1 _38224_inst ( .DIN1(_27082), .DIN2(_26213), .Q(_38257) );
  nnd2s1 _38225_inst ( .DIN1(_38258), .DIN2(_33379), .Q(
        _____________________________11________) );
  nnd2s1 _38226_inst ( .DIN1(_33771), .DIN2(_33399), .Q(_33379) );
  and2s1 _38227_inst ( .DIN1(_38259), .DIN2(_30992), .Q(_33771) );
  hi1s1 _38228_inst ( .DIN(_36023), .Q(_30992) );
  nnd2s1 _38229_inst ( .DIN1(_38260), .DIN2(_38261), .Q(_36023) );
  nor2s1 _38230_inst ( .DIN1(_36493), .DIN2(_38031), .Q(_38260) );
  nor2s1 _38231_inst ( .DIN1(_36976), .DIN2(_38072), .Q(_38259) );
  nor2s1 _38232_inst ( .DIN1(_38262), .DIN2(_38263), .Q(_38258) );
  nor2s1 _38233_inst ( .DIN1(_33399), .DIN2(_38264), .Q(_38263) );
  nnd2s1 _38234_inst ( .DIN1(_33044), .DIN2(_38265), .Q(_38264) );
  xor2s1 _38235_inst ( .DIN1(_38266), .DIN2(_38267), .Q(_38265) );
  xor2s1 _38236_inst ( .DIN1(_35482), .DIN2(_37972), .Q(_38267) );
  hi1s1 _38237_inst ( .DIN(_37973), .Q(_37972) );
  nnd2s1 _38238_inst ( .DIN1(_38268), .DIN2(_38269), .Q(_37973) );
  nnd2s1 _38239_inst ( .DIN1(_53316), .DIN2(_38270), .Q(_38269) );
  or2s1 _38240_inst ( .DIN1(_38271), .DIN2(_35488), .Q(_38270) );
  nnd2s1 _38241_inst ( .DIN1(_35488), .DIN2(_38271), .Q(_38268) );
  xor2s1 _38242_inst ( .DIN1(_37980), .DIN2(_26810), .Q(_35482) );
  nnd2s1 _38243_inst ( .DIN1(_38273), .DIN2(_38274), .Q(_37979) );
  nnd2s1 _38244_inst ( .DIN1(_38275), .DIN2(_34787), .Q(_38274) );
  or2s1 _38245_inst ( .DIN1(_38276), .DIN2(_38277), .Q(_38275) );
  nnd2s1 _38246_inst ( .DIN1(_38277), .DIN2(_38276), .Q(_38273) );
  xor2s1 _38247_inst ( .DIN1(_53295), .DIN2(_32753), .Q(_38266) );
  hi1s1 _38248_inst ( .DIN(_32839), .Q(_33044) );
  hi1s1 _38249_inst ( .DIN(_33305), .Q(_33399) );
  nor2s1 _38250_inst ( .DIN1(_53470), .DIN2(_33305), .Q(_38262) );
  nor2s1 _38251_inst ( .DIN1(_27967), .DIN2(_35998), .Q(_33305) );
  nnd2s1 _38252_inst ( .DIN1(_38278), .DIN2(_38279), .Q(_35998) );
  nor2s1 _38253_inst ( .DIN1(_36493), .DIN2(_38071), .Q(_38278) );
  hi1s1 _38254_inst ( .DIN(_38280), .Q(_36493) );
  hi1s1 _38255_inst ( .DIN(_28755), .Q(_27967) );
  nor2s1 _38256_inst ( .DIN1(_38281), .DIN2(_38282), .Q(_28755) );
  nnd2s1 _38257_inst ( .DIN1(_38283), .DIN2(_38284), .Q(_38281) );
  nnd2s1 _38258_inst ( .DIN1(_38285), .DIN2(_38286), .Q(
        _____________________________119________) );
  nnd2s1 _38259_inst ( .DIN1(_38287), .DIN2(_33356), .Q(_38286) );
  nnd2s1 _38260_inst ( .DIN1(_38288), .DIN2(_38289), .Q(_38287) );
  nor2s1 _38261_inst ( .DIN1(_38290), .DIN2(_38102), .Q(_38289) );
  nor2s1 _38262_inst ( .DIN1(_26510), .DIN2(_26266), .Q(_38102) );
  hi1s1 _38263_inst ( .DIN(_33357), .Q(_38290) );
  nnd2s1 _38264_inst ( .DIN1(_37986), .DIN2(_37930), .Q(_33357) );
  nor2s1 _38265_inst ( .DIN1(_38291), .DIN2(_27651), .Q(_38288) );
  nor2s1 _38266_inst ( .DIN1(_53297), .DIN2(_53298), .Q(_38291) );
  nnd2s1 _38267_inst ( .DIN1(_38292), .DIN2(_33359), .Q(_38285) );
  hi1s1 _38268_inst ( .DIN(_33356), .Q(_33359) );
  nnd2s1 _38269_inst ( .DIN1(_36926), .DIN2(_34126), .Q(_33356) );
  and2s1 _38270_inst ( .DIN1(_37930), .DIN2(_37983), .Q(_34126) );
  nor2s1 _38271_inst ( .DIN1(_31195), .DIN2(_36826), .Q(_37930) );
  hi1s1 _38272_inst ( .DIN(_37299), .Q(_36826) );
  nor2s1 _38273_inst ( .DIN1(_27822), .DIN2(_36827), .Q(_36926) );
  nor2s1 _38274_inst ( .DIN1(_38293), .DIN2(_38187), .Q(_38292) );
  xor2s1 _38275_inst ( .DIN1(_38246), .DIN2(_38294), .Q(_38293) );
  xor2s1 _38276_inst ( .DIN1(_53296), .DIN2(_38245), .Q(_38294) );
  nnd2s1 _38277_inst ( .DIN1(_38295), .DIN2(_38296), .Q(_38245) );
  nnd2s1 _38278_inst ( .DIN1(_38297), .DIN2(_26269), .Q(_38296) );
  or2s1 _38279_inst ( .DIN1(_38298), .DIN2(_38299), .Q(_38297) );
  nnd2s1 _38280_inst ( .DIN1(_38299), .DIN2(_38298), .Q(_38295) );
  hi1s1 _38281_inst ( .DIN(_37542), .Q(_38299) );
  xnr2s1 _38282_inst ( .DIN1(_38300), .DIN2(_36333), .Q(_38246) );
  xor2s1 _38283_inst ( .DIN1(_26335), .DIN2(_38251), .Q(_38300) );
  nnd2s1 _38284_inst ( .DIN1(_38301), .DIN2(_38302), .Q(_38251) );
  nnd2s1 _38285_inst ( .DIN1(_38303), .DIN2(_27620), .Q(_38302) );
  or2s1 _38286_inst ( .DIN1(_38304), .DIN2(_36543), .Q(_38303) );
  nnd2s1 _38287_inst ( .DIN1(_36543), .DIN2(_38304), .Q(_38301) );
  xnr2s1 _38288_inst ( .DIN1(_38256), .DIN2(_38305), .Q(_36333) );
  xor2s1 _38289_inst ( .DIN1(_53314), .DIN2(_53367), .Q(_38305) );
  nnd2s1 _38290_inst ( .DIN1(_38306), .DIN2(_38307), .Q(_38256) );
  nnd2s1 _38291_inst ( .DIN1(_38308), .DIN2(_26526), .Q(_38307) );
  or2s1 _38292_inst ( .DIN1(_38309), .DIN2(_53371), .Q(_38308) );
  nnd2s1 _38293_inst ( .DIN1(_53371), .DIN2(_38309), .Q(_38306) );
  nnd2s1 _38294_inst ( .DIN1(_38310), .DIN2(_38311), .Q(
        _____________________________118________) );
  nnd2s1 _38295_inst ( .DIN1(_38312), .DIN2(_38194), .Q(_38311) );
  hi1s1 _38296_inst ( .DIN(_38187), .Q(_38194) );
  nnd2s1 _38297_inst ( .DIN1(_33285), .DIN2(_33520), .Q(_38187) );
  hi1s1 _38298_inst ( .DIN(_33365), .Q(_33285) );
  nnd2s1 _38299_inst ( .DIN1(_38313), .DIN2(_33519), .Q(_33365) );
  nor2s1 _38300_inst ( .DIN1(_38132), .DIN2(_38314), .Q(_38313) );
  nor2s1 _38301_inst ( .DIN1(_38315), .DIN2(_37528), .Q(_38312) );
  xor2s1 _38302_inst ( .DIN1(_37542), .DIN2(_38316), .Q(_38315) );
  xor2s1 _38303_inst ( .DIN1(_26269), .DIN2(_38298), .Q(_38316) );
  nnd2s1 _38304_inst ( .DIN1(_38317), .DIN2(_38318), .Q(_38298) );
  nnd2s1 _38305_inst ( .DIN1(_53221), .DIN2(_38319), .Q(_38318) );
  nnd2s1 _38306_inst ( .DIN1(_38320), .DIN2(_38321), .Q(_38319) );
  or2s1 _38307_inst ( .DIN1(_38320), .DIN2(_38321), .Q(_38317) );
  hi1s1 _38308_inst ( .DIN(_37575), .Q(_38321) );
  xnr2s1 _38309_inst ( .DIN1(_36543), .DIN2(_26760), .Q(_37542) );
  nnd2s1 _38310_inst ( .DIN1(_38322), .DIN2(_38323), .Q(_38304) );
  nnd2s1 _38311_inst ( .DIN1(_53362), .DIN2(_38324), .Q(_38323) );
  or2s1 _38312_inst ( .DIN1(_38325), .DIN2(_36822), .Q(_38324) );
  nnd2s1 _38313_inst ( .DIN1(_36822), .DIN2(_38325), .Q(_38322) );
  xor2s1 _38314_inst ( .DIN1(_38326), .DIN2(_38309), .Q(_36543) );
  nnd2s1 _38315_inst ( .DIN1(_38327), .DIN2(_38328), .Q(_38309) );
  nnd2s1 _38316_inst ( .DIN1(_38329), .DIN2(_26343), .Q(_38328) );
  or2s1 _38317_inst ( .DIN1(_38330), .DIN2(_53370), .Q(_38329) );
  nnd2s1 _38318_inst ( .DIN1(_53370), .DIN2(_38330), .Q(_38327) );
  xor2s1 _38319_inst ( .DIN1(_26526), .DIN2(_53371), .Q(_38326) );
  nnd2s1 _38320_inst ( .DIN1(_28968), .DIN2(_38331), .Q(_38310) );
  xor2s1 _38321_inst ( .DIN1(_52989), .DIN2(_53301), .Q(_38331) );
  nor2s1 _38322_inst ( .DIN1(_28971), .DIN2(_38332), .Q(_28968) );
  nnd2s1 _38323_inst ( .DIN1(_38333), .DIN2(_38214), .Q(
        _____________________________117________) );
  nor2s1 _38324_inst ( .DIN1(_38334), .DIN2(_38335), .Q(_38333) );
  nor2s1 _38325_inst ( .DIN1(_28971), .DIN2(_38336), .Q(_38335) );
  xnr2s1 _38326_inst ( .DIN1(_53239), .DIN2(_38337), .Q(_38336) );
  nnd2s1 _38327_inst ( .DIN1(_53300), .DIN2(_53301), .Q(_38337) );
  nor2s1 _38328_inst ( .DIN1(_38338), .DIN2(_37528), .Q(_38334) );
  nor2s1 _38329_inst ( .DIN1(_38339), .DIN2(_38340), .Q(_38338) );
  xor2s1 _38330_inst ( .DIN1(_38341), .DIN2(_38320), .Q(_38339) );
  xor2s1 _38331_inst ( .DIN1(_38342), .DIN2(_30674), .Q(_38320) );
  nnd2s1 _38332_inst ( .DIN1(_38343), .DIN2(_35037), .Q(_30674) );
  hi1s1 _38333_inst ( .DIN(_31456), .Q(_35037) );
  nor2s1 _38334_inst ( .DIN1(_38344), .DIN2(_38345), .Q(_38343) );
  nnd2s1 _38335_inst ( .DIN1(_38346), .DIN2(_38347), .Q(_38342) );
  nnd2s1 _38336_inst ( .DIN1(_53302), .DIN2(_38348), .Q(_38347) );
  nnd2s1 _38337_inst ( .DIN1(_37609), .DIN2(_38349), .Q(_38348) );
  or2s1 _38338_inst ( .DIN1(_38349), .DIN2(_37609), .Q(_38346) );
  xor2s1 _38339_inst ( .DIN1(_53221), .DIN2(_37575), .Q(_38341) );
  xnr2s1 _38340_inst ( .DIN1(_36822), .DIN2(_38350), .Q(_37575) );
  xor2s1 _38341_inst ( .DIN1(_26338), .DIN2(_38325), .Q(_38350) );
  nnd2s1 _38342_inst ( .DIN1(_38351), .DIN2(_38352), .Q(_38325) );
  nnd2s1 _38343_inst ( .DIN1(_53361), .DIN2(_38353), .Q(_38352) );
  or2s1 _38344_inst ( .DIN1(_38354), .DIN2(_37104), .Q(_38353) );
  nnd2s1 _38345_inst ( .DIN1(_37104), .DIN2(_38354), .Q(_38351) );
  xnr2s1 _38346_inst ( .DIN1(_38330), .DIN2(_38355), .Q(_36822) );
  xor2s1 _38347_inst ( .DIN1(_53314), .DIN2(_53370), .Q(_38355) );
  nnd2s1 _38348_inst ( .DIN1(_38356), .DIN2(_38357), .Q(_38330) );
  nnd2s1 _38349_inst ( .DIN1(_38358), .DIN2(_36332), .Q(_38357) );
  or2s1 _38350_inst ( .DIN1(_38359), .DIN2(_53517), .Q(_38358) );
  nnd2s1 _38351_inst ( .DIN1(_53517), .DIN2(_38359), .Q(_38356) );
  nnd2s1 _38352_inst ( .DIN1(_38360), .DIN2(_38361), .Q(
        _____________________________116________) );
  nor2s1 _38353_inst ( .DIN1(_38362), .DIN2(_38363), .Q(_38361) );
  nor2s1 _38354_inst ( .DIN1(_26456), .DIN2(_38364), .Q(_38363) );
  nor2s1 _38355_inst ( .DIN1(_53324), .DIN2(_38365), .Q(_38362) );
  nor2s1 _38356_inst ( .DIN1(_38366), .DIN2(_38367), .Q(_38360) );
  nor2s1 _38357_inst ( .DIN1(_38368), .DIN2(_38369), .Q(_38367) );
  xnr2s1 _38358_inst ( .DIN1(_37609), .DIN2(_38370), .Q(_38369) );
  xnr2s1 _38359_inst ( .DIN1(_53302), .DIN2(_38349), .Q(_38370) );
  nnd2s1 _38360_inst ( .DIN1(_38371), .DIN2(_38372), .Q(_38349) );
  nnd2s1 _38361_inst ( .DIN1(_38373), .DIN2(_26378), .Q(_38372) );
  or2s1 _38362_inst ( .DIN1(_38374), .DIN2(_37621), .Q(_38373) );
  nnd2s1 _38363_inst ( .DIN1(_37621), .DIN2(_38374), .Q(_38371) );
  xnr2s1 _38364_inst ( .DIN1(_37104), .DIN2(_26759), .Q(_37609) );
  nnd2s1 _38365_inst ( .DIN1(_38375), .DIN2(_38376), .Q(_38354) );
  nnd2s1 _38366_inst ( .DIN1(_38377), .DIN2(_26331), .Q(_38376) );
  or2s1 _38367_inst ( .DIN1(_38378), .DIN2(_37382), .Q(_38377) );
  nnd2s1 _38368_inst ( .DIN1(_37382), .DIN2(_38378), .Q(_38375) );
  xnr2s1 _38369_inst ( .DIN1(_38379), .DIN2(_38359), .Q(_37104) );
  nnd2s1 _38370_inst ( .DIN1(_38380), .DIN2(_38381), .Q(_38359) );
  nnd2s1 _38371_inst ( .DIN1(_38382), .DIN2(_26778), .Q(_38381) );
  or2s1 _38372_inst ( .DIN1(_38383), .DIN2(_27731), .Q(_38382) );
  nnd2s1 _38373_inst ( .DIN1(_38383), .DIN2(_27731), .Q(_38380) );
  nnd2s1 _38374_inst ( .DIN1(_38384), .DIN2(_38385), .Q(
        _____________________________115________) );
  nor2s1 _38375_inst ( .DIN1(_38386), .DIN2(_38387), .Q(_38385) );
  nor2s1 _38376_inst ( .DIN1(_26601), .DIN2(_38364), .Q(_38387) );
  nnd2s1 _38377_inst ( .DIN1(_32847), .DIN2(_38388), .Q(_38364) );
  nor2s1 _38378_inst ( .DIN1(_53303), .DIN2(_38365), .Q(_38386) );
  hi1s1 _38379_inst ( .DIN(_38389), .Q(_38365) );
  nor2s1 _38380_inst ( .DIN1(_38366), .DIN2(_38390), .Q(_38384) );
  nor2s1 _38381_inst ( .DIN1(_38368), .DIN2(_38391), .Q(_38390) );
  xnr2s1 _38382_inst ( .DIN1(_37621), .DIN2(_38392), .Q(_38391) );
  xor2s1 _38383_inst ( .DIN1(_26378), .DIN2(_38374), .Q(_38392) );
  nnd2s1 _38384_inst ( .DIN1(_38393), .DIN2(_38394), .Q(_38374) );
  nnd2s1 _38385_inst ( .DIN1(_38395), .DIN2(_26403), .Q(_38394) );
  or2s1 _38386_inst ( .DIN1(_38396), .DIN2(_37635), .Q(_38395) );
  nnd2s1 _38387_inst ( .DIN1(_37635), .DIN2(_38396), .Q(_38393) );
  hi1s1 _38388_inst ( .DIN(_38397), .Q(_37635) );
  xnr2s1 _38389_inst ( .DIN1(_37382), .DIN2(_38398), .Q(_37621) );
  xor2s1 _38390_inst ( .DIN1(_38383), .DIN2(_38399), .Q(_37382) );
  xor2s1 _38391_inst ( .DIN1(_53370), .DIN2(_53375), .Q(_38399) );
  nnd2s1 _38392_inst ( .DIN1(_38400), .DIN2(_38401), .Q(_38383) );
  nnd2s1 _38393_inst ( .DIN1(_53373), .DIN2(_38402), .Q(_38401) );
  or2s1 _38394_inst ( .DIN1(_38403), .DIN2(_26323), .Q(_38402) );
  nnd2s1 _38395_inst ( .DIN1(_38403), .DIN2(_26323), .Q(_38400) );
  xor2s1 _38396_inst ( .DIN1(_38378), .DIN2(_53365), .Q(_38398) );
  nnd2s1 _38397_inst ( .DIN1(_38404), .DIN2(_38405), .Q(_38378) );
  nnd2s1 _38398_inst ( .DIN1(_38406), .DIN2(_26780), .Q(_38405) );
  or2s1 _38399_inst ( .DIN1(_38407), .DIN2(_37592), .Q(_38406) );
  xor2s1 _38400_inst ( .DIN1(_38212), .DIN2(_38408), .Q(_38404) );
  nnd2s1 _38401_inst ( .DIN1(_37592), .DIN2(_38407), .Q(_38408) );
  nnd2s1 _38402_inst ( .DIN1(_37403), .DIN2(_31459), .Q(_38212) );
  nnd2s1 _38403_inst ( .DIN1(_38409), .DIN2(_32868), .Q(_38368) );
  nnd2s1 _38404_inst ( .DIN1(_38410), .DIN2(_27198), .Q(
        _____________________________114________) );
  nnd2s1 _38405_inst ( .DIN1(_36552), .DIN2(_27204), .Q(_27198) );
  nor2s1 _38406_inst ( .DIN1(_38411), .DIN2(_38412), .Q(_38410) );
  nor2s1 _38407_inst ( .DIN1(_38413), .DIN2(_27204), .Q(_38412) );
  nor2s1 _38408_inst ( .DIN1(_38414), .DIN2(_38340), .Q(_38413) );
  xor2s1 _38409_inst ( .DIN1(_38397), .DIN2(_38415), .Q(_38414) );
  xor2s1 _38410_inst ( .DIN1(_26403), .DIN2(_38396), .Q(_38415) );
  nnd2s1 _38411_inst ( .DIN1(_38416), .DIN2(_38417), .Q(_38396) );
  nnd2s1 _38412_inst ( .DIN1(_53308), .DIN2(_38418), .Q(_38417) );
  or2s1 _38413_inst ( .DIN1(_38419), .DIN2(_37657), .Q(_38418) );
  nnd2s1 _38414_inst ( .DIN1(_37657), .DIN2(_38419), .Q(_38416) );
  xnr2s1 _38415_inst ( .DIN1(_37592), .DIN2(_26786), .Q(_38397) );
  nnd2s1 _38416_inst ( .DIN1(_38421), .DIN2(_38422), .Q(_38407) );
  nnd2s1 _38417_inst ( .DIN1(_38423), .DIN2(_26209), .Q(_38422) );
  xor2s1 _38418_inst ( .DIN1(_33328), .DIN2(_38424), .Q(_38423) );
  xor2s1 _38419_inst ( .DIN1(_38425), .DIN2(_38403), .Q(_37592) );
  nnd2s1 _38420_inst ( .DIN1(_38426), .DIN2(_38427), .Q(_38403) );
  nnd2s1 _38421_inst ( .DIN1(_53374), .DIN2(_38428), .Q(_38427) );
  or2s1 _38422_inst ( .DIN1(_38429), .DIN2(_53375), .Q(_38428) );
  nnd2s1 _38423_inst ( .DIN1(_53375), .DIN2(_38429), .Q(_38426) );
  xor2s1 _38424_inst ( .DIN1(_26333), .DIN2(_53517), .Q(_38425) );
  nor2s1 _38425_inst ( .DIN1(_27201), .DIN2(_38430), .Q(_38411) );
  nor2s1 _38426_inst ( .DIN1(_27393), .DIN2(_38431), .Q(_38430) );
  nnd2s1 _38427_inst ( .DIN1(_38432), .DIN2(_28991), .Q(_38431) );
  or2s1 _38428_inst ( .DIN1(_53311), .DIN2(_53310), .Q(_38432) );
  nnd2s1 _38429_inst ( .DIN1(_38433), .DIN2(_38434), .Q(
        _____________________________113________) );
  nnd2s1 _38430_inst ( .DIN1(_38435), .DIN2(_38436), .Q(_38434) );
  xor2s1 _38431_inst ( .DIN1(_37657), .DIN2(_38437), .Q(_38436) );
  xor2s1 _38432_inst ( .DIN1(_38419), .DIN2(_53308), .Q(_38437) );
  nnd2s1 _38433_inst ( .DIN1(_38438), .DIN2(_38439), .Q(_38419) );
  nnd2s1 _38434_inst ( .DIN1(_53331), .DIN2(_38440), .Q(_38439) );
  or2s1 _38435_inst ( .DIN1(_38441), .DIN2(_37667), .Q(_38440) );
  nnd2s1 _38436_inst ( .DIN1(_37667), .DIN2(_38441), .Q(_38438) );
  nnd2s1 _38437_inst ( .DIN1(_38442), .DIN2(_38443), .Q(_37657) );
  nnd2s1 _38438_inst ( .DIN1(_38444), .DIN2(_26209), .Q(_38443) );
  nnd2s1 _38439_inst ( .DIN1(_38424), .DIN2(_38421), .Q(_38444) );
  nnd2s1 _38440_inst ( .DIN1(_37791), .DIN2(_38445), .Q(_38421) );
  hi1s1 _38441_inst ( .DIN(_37974), .Q(_37791) );
  nnd2s1 _38442_inst ( .DIN1(_38446), .DIN2(_37974), .Q(_38424) );
  nnd2s1 _38443_inst ( .DIN1(_38447), .DIN2(_53367), .Q(_38442) );
  xor2s1 _38444_inst ( .DIN1(_37974), .DIN2(_38446), .Q(_38447) );
  hi1s1 _38445_inst ( .DIN(_38445), .Q(_38446) );
  nnd2s1 _38446_inst ( .DIN1(_38448), .DIN2(_38449), .Q(_38445) );
  nnd2s1 _38447_inst ( .DIN1(_38450), .DIN2(_26526), .Q(_38449) );
  or2s1 _38448_inst ( .DIN1(_38451), .DIN2(_37980), .Q(_38450) );
  nnd2s1 _38449_inst ( .DIN1(_37980), .DIN2(_38451), .Q(_38448) );
  xor2s1 _38450_inst ( .DIN1(_38429), .DIN2(_38452), .Q(_37974) );
  nnd2s1 _38451_inst ( .DIN1(_38453), .DIN2(_38454), .Q(_38429) );
  nnd2s1 _38452_inst ( .DIN1(_53372), .DIN2(_38455), .Q(_38454) );
  or2s1 _38453_inst ( .DIN1(_38456), .DIN2(_26333), .Q(_38455) );
  nnd2s1 _38454_inst ( .DIN1(_38456), .DIN2(_26333), .Q(_38453) );
  nor2s1 _38455_inst ( .DIN1(_27132), .DIN2(_38340), .Q(_38435) );
  nnd2s1 _38456_inst ( .DIN1(_38457), .DIN2(_38458), .Q(_38433) );
  xnr2s1 _38457_inst ( .DIN1(_52878), .DIN2(_29787), .Q(_38458) );
  nor2s1 _38458_inst ( .DIN1(_26679), .DIN2(_53307), .Q(_29787) );
  nor2s1 _38459_inst ( .DIN1(_28100), .DIN2(_29789), .Q(_38457) );
  nnd2s1 _38460_inst ( .DIN1(_27132), .DIN2(_38459), .Q(_29789) );
  nnd2s1 _38461_inst ( .DIN1(_34826), .DIN2(_38460), .Q(_38459) );
  nnd2s1 _38462_inst ( .DIN1(_36552), .DIN2(_34827), .Q(_27132) );
  nnd2s1 _38463_inst ( .DIN1(_38461), .DIN2(_38462), .Q(
        _____________________________112________) );
  nnd2s1 _38464_inst ( .DIN1(_38463), .DIN2(_38409), .Q(_38462) );
  hi1s1 _38465_inst ( .DIN(_38340), .Q(_38409) );
  nnd2s1 _38466_inst ( .DIN1(_38464), .DIN2(_33519), .Q(_38340) );
  hi1s1 _38467_inst ( .DIN(_33281), .Q(_33519) );
  nnd2s1 _38468_inst ( .DIN1(_38465), .DIN2(_38466), .Q(_33281) );
  nor2s1 _38469_inst ( .DIN1(_38467), .DIN2(_27204), .Q(_38463) );
  xor2s1 _38470_inst ( .DIN1(_37667), .DIN2(_38468), .Q(_38467) );
  xnr2s1 _38471_inst ( .DIN1(_53331), .DIN2(_38441), .Q(_38468) );
  nnd2s1 _38472_inst ( .DIN1(_38469), .DIN2(_38470), .Q(_38441) );
  nnd2s1 _38473_inst ( .DIN1(_38471), .DIN2(_26531), .Q(_38470) );
  or2s1 _38474_inst ( .DIN1(_38472), .DIN2(_37689), .Q(_38471) );
  nnd2s1 _38475_inst ( .DIN1(_37689), .DIN2(_38472), .Q(_38469) );
  xor2s1 _38476_inst ( .DIN1(_37980), .DIN2(_38473), .Q(_37667) );
  xor2s1 _38477_inst ( .DIN1(_26526), .DIN2(_38451), .Q(_38473) );
  nnd2s1 _38478_inst ( .DIN1(_38474), .DIN2(_38475), .Q(_38451) );
  nnd2s1 _38479_inst ( .DIN1(_38476), .DIN2(_26343), .Q(_38475) );
  or2s1 _38480_inst ( .DIN1(_38477), .DIN2(_38277), .Q(_38476) );
  nnd2s1 _38481_inst ( .DIN1(_38277), .DIN2(_38477), .Q(_38474) );
  xor2s1 _38482_inst ( .DIN1(_38478), .DIN2(_38456), .Q(_37980) );
  xnr2s1 _38483_inst ( .DIN1(_38479), .DIN2(_27338), .Q(_38456) );
  nnd2s1 _38484_inst ( .DIN1(_38480), .DIN2(_38481), .Q(_38479) );
  nnd2s1 _38485_inst ( .DIN1(_53338), .DIN2(_38482), .Q(_38481) );
  or2s1 _38486_inst ( .DIN1(_38483), .DIN2(_26322), .Q(_38482) );
  nnd2s1 _38487_inst ( .DIN1(_38483), .DIN2(_26322), .Q(_38480) );
  xor2s1 _38488_inst ( .DIN1(_26336), .DIN2(_53373), .Q(_38478) );
  nnd2s1 _38489_inst ( .DIN1(_38484), .DIN2(_28992), .Q(_38461) );
  nor2s1 _38490_inst ( .DIN1(_27201), .DIN2(_36552), .Q(_28992) );
  hi1s1 _38491_inst ( .DIN(_27204), .Q(_27201) );
  nnd2s1 _38492_inst ( .DIN1(_38485), .DIN2(_34828), .Q(_27204) );
  nor2s1 _38493_inst ( .DIN1(_38486), .DIN2(_35617), .Q(_38485) );
  xor2s1 _38494_inst ( .DIN1(_28991), .DIN2(_52994), .Q(_38484) );
  nnd2s1 _38495_inst ( .DIN1(_53310), .DIN2(_53311), .Q(_28991) );
  nnd2s1 _38496_inst ( .DIN1(_38487), .DIN2(_32844), .Q(
        _____________________________111________) );
  hi1s1 _38497_inst ( .DIN(_38366), .Q(_32844) );
  nor2s1 _38498_inst ( .DIN1(_38488), .DIN2(_38489), .Q(_38487) );
  nor2s1 _38499_inst ( .DIN1(_38490), .DIN2(_32847), .Q(_38489) );
  nor2s1 _38500_inst ( .DIN1(_38491), .DIN2(_38492), .Q(_38490) );
  nor2s1 _38501_inst ( .DIN1(_38493), .DIN2(_38494), .Q(_38492) );
  xor2s1 _38502_inst ( .DIN1(_38495), .DIN2(_38496), .Q(_38494) );
  xor2s1 _38503_inst ( .DIN1(_53325), .DIN2(_53326), .Q(_38496) );
  nnd2s1 _38504_inst ( .DIN1(_53324), .DIN2(_53325), .Q(_38495) );
  nor2s1 _38505_inst ( .DIN1(_38497), .DIN2(_33531), .Q(_38491) );
  xnr2s1 _38506_inst ( .DIN1(_37689), .DIN2(_38498), .Q(_38497) );
  xor2s1 _38507_inst ( .DIN1(_26531), .DIN2(_38472), .Q(_38498) );
  nnd2s1 _38508_inst ( .DIN1(_38499), .DIN2(_38500), .Q(_38472) );
  nnd2s1 _38509_inst ( .DIN1(_38501), .DIN2(_26545), .Q(_38500) );
  or2s1 _38510_inst ( .DIN1(_38502), .DIN2(_37716), .Q(_38501) );
  nnd2s1 _38511_inst ( .DIN1(_37716), .DIN2(_38502), .Q(_38499) );
  xor2s1 _38512_inst ( .DIN1(_38277), .DIN2(_38503), .Q(_37689) );
  xor2s1 _38513_inst ( .DIN1(_26343), .DIN2(_38477), .Q(_38503) );
  nnd2s1 _38514_inst ( .DIN1(_38504), .DIN2(_38505), .Q(_38477) );
  nnd2s1 _38515_inst ( .DIN1(_38506), .DIN2(_36332), .Q(_38505) );
  or2s1 _38516_inst ( .DIN1(_38507), .DIN2(_38508), .Q(_38506) );
  nnd2s1 _38517_inst ( .DIN1(_38508), .DIN2(_38507), .Q(_38504) );
  nor2s1 _38518_inst ( .DIN1(_53321), .DIN2(_32868), .Q(_38488) );
  nnd2s1 _38519_inst ( .DIN1(_38509), .DIN2(_28530), .Q(
        _____________________________110________) );
  nnd2s1 _38520_inst ( .DIN1(_29215), .DIN2(_28533), .Q(_28530) );
  hi1s1 _38521_inst ( .DIN(_36302), .Q(_29215) );
  nor2s1 _38522_inst ( .DIN1(_38510), .DIN2(_38511), .Q(_38509) );
  nor2s1 _38523_inst ( .DIN1(_28533), .DIN2(_38512), .Q(_38511) );
  nnd2s1 _38524_inst ( .DIN1(_38513), .DIN2(_38514), .Q(_38512) );
  nnd2s1 _38525_inst ( .DIN1(_33536), .DIN2(_38515), .Q(_38514) );
  xor2s1 _38526_inst ( .DIN1(_37716), .DIN2(_38516), .Q(_38515) );
  xor2s1 _38527_inst ( .DIN1(_26545), .DIN2(_38502), .Q(_38516) );
  nnd2s1 _38528_inst ( .DIN1(_38517), .DIN2(_38518), .Q(_38502) );
  nnd2s1 _38529_inst ( .DIN1(_38519), .DIN2(_26267), .Q(_38518) );
  or2s1 _38530_inst ( .DIN1(_38520), .DIN2(_37733), .Q(_38519) );
  nnd2s1 _38531_inst ( .DIN1(_37733), .DIN2(_38520), .Q(_38517) );
  xnr2s1 _38532_inst ( .DIN1(_38521), .DIN2(_38522), .Q(_37716) );
  xor2s1 _38533_inst ( .DIN1(_38507), .DIN2(_38508), .Q(_38522) );
  nnd2s1 _38534_inst ( .DIN1(_38523), .DIN2(_38524), .Q(_38507) );
  nnd2s1 _38535_inst ( .DIN1(_38525), .DIN2(_26778), .Q(_38524) );
  or2s1 _38536_inst ( .DIN1(_38526), .DIN2(_38527), .Q(_38525) );
  nnd2s1 _38537_inst ( .DIN1(_38526), .DIN2(_38527), .Q(_38523) );
  xor2s1 _38538_inst ( .DIN1(_36332), .DIN2(_31802), .Q(_38521) );
  hi1s1 _38539_inst ( .DIN(_31585), .Q(_31802) );
  nnd2s1 _38540_inst ( .DIN1(_32762), .DIN2(_38528), .Q(_31585) );
  hi1s1 _38541_inst ( .DIN(_29544), .Q(_32762) );
  nnd2s1 _38542_inst ( .DIN1(_38529), .DIN2(______[4]), .Q(_38513) );
  nor2s1 _38543_inst ( .DIN1(_53304), .DIN2(_38493), .Q(_38529) );
  nor2s1 _38544_inst ( .DIN1(_28542), .DIN2(_38530), .Q(_38510) );
  nor2s1 _38545_inst ( .DIN1(_27651), .DIN2(_26602), .Q(_38530) );
  nnd2s1 _38546_inst ( .DIN1(_38531), .DIN2(_38214), .Q(
        _____________________________10________) );
  nnd2s1 _38547_inst ( .DIN1(_38332), .DIN2(_37528), .Q(_38214) );
  nor2s1 _38548_inst ( .DIN1(_38532), .DIN2(_38533), .Q(_38531) );
  nor2s1 _38549_inst ( .DIN1(_28971), .DIN2(_38534), .Q(_38533) );
  and2s1 _38550_inst ( .DIN1(______[12]), .DIN2(_53229), .Q(_38534) );
  hi1s1 _38551_inst ( .DIN(_37528), .Q(_28971) );
  nor2s1 _38552_inst ( .DIN1(_38535), .DIN2(_37528), .Q(_38532) );
  nnd2s1 _38553_inst ( .DIN1(_38536), .DIN2(_34826), .Q(_37528) );
  hi1s1 _38554_inst ( .DIN(_30129), .Q(_34826) );
  nnd2s1 _38555_inst ( .DIN1(_32015), .DIN2(_31103), .Q(_30129) );
  nor2s1 _38556_inst ( .DIN1(_38486), .DIN2(_38537), .Q(_38536) );
  nor2s1 _38557_inst ( .DIN1(_32839), .DIN2(_38538), .Q(_38535) );
  xor2s1 _38558_inst ( .DIN1(_35488), .DIN2(_38539), .Q(_38538) );
  xor2s1 _38559_inst ( .DIN1(_26462), .DIN2(_38271), .Q(_38539) );
  nnd2s1 _38560_inst ( .DIN1(_38540), .DIN2(_38541), .Q(_38271) );
  nnd2s1 _38561_inst ( .DIN1(_53008), .DIN2(_38542), .Q(_38541) );
  or2s1 _38562_inst ( .DIN1(_32840), .DIN2(_32842), .Q(_38542) );
  nnd2s1 _38563_inst ( .DIN1(_32840), .DIN2(_32842), .Q(_38540) );
  nnd2s1 _38564_inst ( .DIN1(_33047), .DIN2(_38543), .Q(_32842) );
  nnd2s1 _38565_inst ( .DIN1(_38544), .DIN2(_26528), .Q(_38543) );
  xor2s1 _38566_inst ( .DIN1(_33046), .DIN2(_38545), .Q(_38544) );
  xor2s1 _38567_inst ( .DIN1(_33328), .DIN2(_28613), .Q(_38545) );
  nnd2s1 _38568_inst ( .DIN1(_32612), .DIN2(_37922), .Q(_33328) );
  or2s1 _38569_inst ( .DIN1(_38546), .DIN2(_35520), .Q(_33046) );
  nnd2s1 _38570_inst ( .DIN1(_35520), .DIN2(_38546), .Q(_33047) );
  nnd2s1 _38571_inst ( .DIN1(_38547), .DIN2(_38548), .Q(_38546) );
  nnd2s1 _38572_inst ( .DIN1(_53011), .DIN2(_38549), .Q(_38548) );
  or2s1 _38573_inst ( .DIN1(_33255), .DIN2(_33253), .Q(_38549) );
  nnd2s1 _38574_inst ( .DIN1(_33253), .DIN2(_33255), .Q(_38547) );
  nnd2s1 _38575_inst ( .DIN1(_38550), .DIN2(_38551), .Q(_33255) );
  nnd2s1 _38576_inst ( .DIN1(_53012), .DIN2(_38552), .Q(_38551) );
  or2s1 _38577_inst ( .DIN1(_33463), .DIN2(_33461), .Q(_38552) );
  nnd2s1 _38578_inst ( .DIN1(_33461), .DIN2(_33463), .Q(_38550) );
  nnd2s1 _38579_inst ( .DIN1(_38553), .DIN2(_38554), .Q(_33463) );
  nnd2s1 _38580_inst ( .DIN1(_53023), .DIN2(_38555), .Q(_38554) );
  or2s1 _38581_inst ( .DIN1(_33674), .DIN2(_33675), .Q(_38555) );
  nnd2s1 _38582_inst ( .DIN1(_33675), .DIN2(_33674), .Q(_38553) );
  nnd2s1 _38583_inst ( .DIN1(_38556), .DIN2(_38557), .Q(_33674) );
  nnd2s1 _38584_inst ( .DIN1(_38558), .DIN2(_26479), .Q(_38557) );
  or2s1 _38585_inst ( .DIN1(_33874), .DIN2(_33872), .Q(_38558) );
  nnd2s1 _38586_inst ( .DIN1(_33872), .DIN2(_33874), .Q(_38556) );
  nnd2s1 _38587_inst ( .DIN1(_38559), .DIN2(_38560), .Q(_33874) );
  nnd2s1 _38588_inst ( .DIN1(_38561), .DIN2(_26399), .Q(_38560) );
  or2s1 _38589_inst ( .DIN1(_34086), .DIN2(_34084), .Q(_38561) );
  nnd2s1 _38590_inst ( .DIN1(_34084), .DIN2(_34086), .Q(_38559) );
  nnd2s1 _38591_inst ( .DIN1(_38562), .DIN2(_38563), .Q(_34086) );
  nnd2s1 _38592_inst ( .DIN1(_38564), .DIN2(_53319), .Q(_38563) );
  nor2s1 _38593_inst ( .DIN1(_38565), .DIN2(_36306), .Q(_38564) );
  hi1s1 _38594_inst ( .DIN(_34288), .Q(_36306) );
  nnd2s1 _38595_inst ( .DIN1(_38566), .DIN2(_38567), .Q(_34288) );
  nnd2s1 _38596_inst ( .DIN1(_53358), .DIN2(_38568), .Q(_38567) );
  nnd2s1 _38597_inst ( .DIN1(_38569), .DIN2(_38570), .Q(_38568) );
  nnd2s1 _38598_inst ( .DIN1(_38571), .DIN2(_26448), .Q(_38566) );
  xor2s1 _38599_inst ( .DIN1(_38572), .DIN2(_38573), .Q(_38571) );
  nor2s1 _38600_inst ( .DIN1(_53053), .DIN2(_34287), .Q(_38565) );
  nnd2s1 _38601_inst ( .DIN1(_34287), .DIN2(_53053), .Q(_38562) );
  xnr2s1 _38602_inst ( .DIN1(_38574), .DIN2(_38575), .Q(_34287) );
  xor2s1 _38603_inst ( .DIN1(_26396), .DIN2(_38576), .Q(_38575) );
  hi1s1 _38604_inst ( .DIN(_35665), .Q(_34084) );
  xnr2s1 _38605_inst ( .DIN1(_38577), .DIN2(_38578), .Q(_35665) );
  xor2s1 _38606_inst ( .DIN1(_38579), .DIN2(_53352), .Q(_38577) );
  xnr2s1 _38607_inst ( .DIN1(_38581), .DIN2(_38580), .Q(_33872) );
  xor2s1 _38608_inst ( .DIN1(_26320), .DIN2(_38582), .Q(_38581) );
  xnr2s1 _38609_inst ( .DIN1(_38583), .DIN2(_38584), .Q(_33675) );
  xnr2s1 _38610_inst ( .DIN1(_38585), .DIN2(_38586), .Q(_38584) );
  xor2s1 _38611_inst ( .DIN1(_26330), .DIN2(_32005), .Q(_38583) );
  xor2s1 _38612_inst ( .DIN1(_38587), .DIN2(_38588), .Q(_33461) );
  xor2s1 _38613_inst ( .DIN1(_38589), .DIN2(_38590), .Q(_38588) );
  xnr2s1 _38614_inst ( .DIN1(_38591), .DIN2(_38592), .Q(_33253) );
  xor2s1 _38615_inst ( .DIN1(_27558), .DIN2(_38593), .Q(_38592) );
  xnr2s1 _38616_inst ( .DIN1(_38527), .DIN2(_26811), .Q(_35520) );
  xnr2s1 _38617_inst ( .DIN1(_38508), .DIN2(_26815), .Q(_32840) );
  xor2s1 _38618_inst ( .DIN1(_38277), .DIN2(_26785), .Q(_35488) );
  nnd2s1 _38619_inst ( .DIN1(_38599), .DIN2(_38600), .Q(_38276) );
  nnd2s1 _38620_inst ( .DIN1(_53377), .DIN2(_38601), .Q(_38600) );
  or2s1 _38621_inst ( .DIN1(_38597), .DIN2(_38508), .Q(_38601) );
  nnd2s1 _38622_inst ( .DIN1(_38508), .DIN2(_38597), .Q(_38599) );
  nnd2s1 _38623_inst ( .DIN1(_38602), .DIN2(_38603), .Q(_38597) );
  nnd2s1 _38624_inst ( .DIN1(_53379), .DIN2(_38604), .Q(_38603) );
  or2s1 _38625_inst ( .DIN1(_38595), .DIN2(_38527), .Q(_38604) );
  nnd2s1 _38626_inst ( .DIN1(_38527), .DIN2(_38595), .Q(_38602) );
  nnd2s1 _38627_inst ( .DIN1(_38605), .DIN2(_38606), .Q(_38595) );
  nnd2s1 _38628_inst ( .DIN1(_53346), .DIN2(_38607), .Q(_38606) );
  or2s1 _38629_inst ( .DIN1(_38593), .DIN2(_38591), .Q(_38607) );
  nnd2s1 _38630_inst ( .DIN1(_38591), .DIN2(_38593), .Q(_38605) );
  nnd2s1 _38631_inst ( .DIN1(_38608), .DIN2(_38609), .Q(_38593) );
  nnd2s1 _38632_inst ( .DIN1(_53381), .DIN2(_38610), .Q(_38609) );
  or2s1 _38633_inst ( .DIN1(_38590), .DIN2(_38611), .Q(_38610) );
  nnd2s1 _38634_inst ( .DIN1(_38611), .DIN2(_38590), .Q(_38608) );
  nnd2s1 _38635_inst ( .DIN1(_38612), .DIN2(_38613), .Q(_38590) );
  nnd2s1 _38636_inst ( .DIN1(_53380), .DIN2(_38614), .Q(_38613) );
  or2s1 _38637_inst ( .DIN1(_38585), .DIN2(_38586), .Q(_38614) );
  nnd2s1 _38638_inst ( .DIN1(_38586), .DIN2(_38585), .Q(_38612) );
  nnd2s1 _38639_inst ( .DIN1(_38615), .DIN2(_38616), .Q(_38585) );
  nnd2s1 _38640_inst ( .DIN1(_53350), .DIN2(_38617), .Q(_38616) );
  or2s1 _38641_inst ( .DIN1(_38582), .DIN2(_38580), .Q(_38617) );
  nnd2s1 _38642_inst ( .DIN1(_38580), .DIN2(_38582), .Q(_38615) );
  nnd2s1 _38643_inst ( .DIN1(_38618), .DIN2(_38619), .Q(_38582) );
  nnd2s1 _38644_inst ( .DIN1(_53352), .DIN2(_38620), .Q(_38619) );
  or2s1 _38645_inst ( .DIN1(_38579), .DIN2(_38578), .Q(_38620) );
  nnd2s1 _38646_inst ( .DIN1(_38578), .DIN2(_38579), .Q(_38618) );
  nnd2s1 _38647_inst ( .DIN1(_38621), .DIN2(_38622), .Q(_38578) );
  nnd2s1 _38648_inst ( .DIN1(_53357), .DIN2(_38623), .Q(_38622) );
  or2s1 _38649_inst ( .DIN1(_38576), .DIN2(_38574), .Q(_38623) );
  nnd2s1 _38650_inst ( .DIN1(_38574), .DIN2(_38576), .Q(_38621) );
  nnd2s1 _38651_inst ( .DIN1(_38570), .DIN2(_38624), .Q(_38576) );
  nnd2s1 _38652_inst ( .DIN1(_53358), .DIN2(_38625), .Q(_38624) );
  xor2s1 _38653_inst ( .DIN1(_34026), .DIN2(_38569), .Q(_38625) );
  or2s1 _38654_inst ( .DIN1(_38572), .DIN2(_38573), .Q(_38569) );
  nnd2s1 _38655_inst ( .DIN1(_38573), .DIN2(_38572), .Q(_38570) );
  nnd2s1 _38656_inst ( .DIN1(_38626), .DIN2(_38627), .Q(_38572) );
  nnd2s1 _38657_inst ( .DIN1(_53467), .DIN2(_38628), .Q(_38627) );
  nnd2s1 _38658_inst ( .DIN1(_38629), .DIN2(_38630), .Q(_38626) );
  nnd2s1 _38659_inst ( .DIN1(_38631), .DIN2(_26341), .Q(_38630) );
  nor2s1 _38660_inst ( .DIN1(_38632), .DIN2(_38633), .Q(_38629) );
  nor2s1 _38661_inst ( .DIN1(_38634), .DIN2(_38635), .Q(_38633) );
  nor2s1 _38662_inst ( .DIN1(_38636), .DIN2(_26329), .Q(_38632) );
  and2s1 _38663_inst ( .DIN1(_38635), .DIN2(_38634), .Q(_38636) );
  nnd2s1 _38664_inst ( .DIN1(_38637), .DIN2(_38638), .Q(_38635) );
  nnd2s1 _38665_inst ( .DIN1(_38639), .DIN2(_53369), .Q(_38638) );
  nor2s1 _38666_inst ( .DIN1(_38640), .DIN2(_38641), .Q(_38639) );
  nor2s1 _38667_inst ( .DIN1(_38642), .DIN2(_26698), .Q(_38640) );
  nnd2s1 _38668_inst ( .DIN1(_38642), .DIN2(_26698), .Q(_38637) );
  xnr2s1 _38669_inst ( .DIN1(_38643), .DIN2(_38644), .Q(_38508) );
  xor2s1 _38670_inst ( .DIN1(_26336), .DIN2(_53376), .Q(_38643) );
  xnr2s1 _38671_inst ( .DIN1(_38483), .DIN2(_38645), .Q(_38277) );
  xor2s1 _38672_inst ( .DIN1(_53338), .DIN2(_53374), .Q(_38645) );
  nnd2s1 _38673_inst ( .DIN1(_38646), .DIN2(_38647), .Q(_38483) );
  nnd2s1 _38674_inst ( .DIN1(_38648), .DIN2(_26336), .Q(_38647) );
  or2s1 _38675_inst ( .DIN1(_38644), .DIN2(_34787), .Q(_38648) );
  nnd2s1 _38676_inst ( .DIN1(_38644), .DIN2(_34787), .Q(_38646) );
  nnd2s1 _38677_inst ( .DIN1(_38649), .DIN2(_38650), .Q(_38644) );
  nnd2s1 _38678_inst ( .DIN1(_38651), .DIN2(_26319), .Q(_38650) );
  or2s1 _38679_inst ( .DIN1(_38652), .DIN2(_53377), .Q(_38651) );
  nnd2s1 _38680_inst ( .DIN1(_53377), .DIN2(_38652), .Q(_38649) );
  nnd2s1 _38681_inst ( .DIN1(_27567), .DIN2(_36336), .Q(_32839) );
  hi1s1 _38682_inst ( .DIN(_27557), .Q(_27567) );
  nnd2s1 _38683_inst ( .DIN1(_27555), .DIN2(_34913), .Q(_27557) );
  hi1s1 _38684_inst ( .DIN(_27683), .Q(_27555) );
  xor2s1 _38685_inst ( .DIN1(_31222), .DIN2(_27585), .Q(_27683) );
  nnd2s1 _38686_inst ( .DIN1(_38653), .DIN2(_38654), .Q(
        _____________________________109________) );
  nor2s1 _38687_inst ( .DIN1(_38655), .DIN2(_38656), .Q(_38654) );
  nor2s1 _38688_inst ( .DIN1(_32847), .DIN2(_38657), .Q(_38656) );
  xor2s1 _38689_inst ( .DIN1(_26998), .DIN2(_38658), .Q(_38657) );
  nnd2s1 _38690_inst ( .DIN1(_38659), .DIN2(_38660), .Q(_38658) );
  nnd2s1 _38691_inst ( .DIN1(_38661), .DIN2(_33531), .Q(_38660) );
  nnd2s1 _38692_inst ( .DIN1(_53325), .DIN2(_38662), .Q(_38661) );
  nnd2s1 _38693_inst ( .DIN1(_38663), .DIN2(_33536), .Q(_38659) );
  xnr2s1 _38694_inst ( .DIN1(_37733), .DIN2(_38664), .Q(_38663) );
  xor2s1 _38695_inst ( .DIN1(_26267), .DIN2(_38520), .Q(_38664) );
  nnd2s1 _38696_inst ( .DIN1(_38665), .DIN2(_38666), .Q(_38520) );
  nnd2s1 _38697_inst ( .DIN1(_38667), .DIN2(_26520), .Q(_38666) );
  xor2s1 _38698_inst ( .DIN1(_27413), .DIN2(_38668), .Q(_38667) );
  xor2s1 _38699_inst ( .DIN1(_38669), .DIN2(_38526), .Q(_37733) );
  xnr2s1 _38700_inst ( .DIN1(_34026), .DIN2(_38670), .Q(_38526) );
  nor2s1 _38701_inst ( .DIN1(_38671), .DIN2(_38672), .Q(_38670) );
  and2s1 _38702_inst ( .DIN1(_38673), .DIN2(_38591), .Q(_38672) );
  nor2s1 _38703_inst ( .DIN1(_53517), .DIN2(_38674), .Q(_38671) );
  nor2s1 _38704_inst ( .DIN1(_38591), .DIN2(_38673), .Q(_38674) );
  xor2s1 _38705_inst ( .DIN1(_26778), .DIN2(_38527), .Q(_38669) );
  xor2s1 _38706_inst ( .DIN1(_38675), .DIN2(_38652), .Q(_38527) );
  nnd2s1 _38707_inst ( .DIN1(_38676), .DIN2(_38677), .Q(_38652) );
  nnd2s1 _38708_inst ( .DIN1(_53376), .DIN2(_38678), .Q(_38677) );
  or2s1 _38709_inst ( .DIN1(_38679), .DIN2(_53379), .Q(_38678) );
  nnd2s1 _38710_inst ( .DIN1(_53379), .DIN2(_38679), .Q(_38676) );
  xor2s1 _38711_inst ( .DIN1(_26319), .DIN2(_53377), .Q(_38675) );
  nor2s1 _38712_inst ( .DIN1(_32868), .DIN2(_38680), .Q(_38655) );
  nnd2s1 _38713_inst ( .DIN1(_26309), .DIN2(_26555), .Q(_38680) );
  nor2s1 _38714_inst ( .DIN1(_38366), .DIN2(_38389), .Q(_38653) );
  nor2s1 _38715_inst ( .DIN1(_38388), .DIN2(_32868), .Q(_38389) );
  nnd2s1 _38716_inst ( .DIN1(_53304), .DIN2(_53321), .Q(_38388) );
  nor2s1 _38717_inst ( .DIN1(_38681), .DIN2(_33294), .Q(_38366) );
  nnd2s1 _38718_inst ( .DIN1(_38682), .DIN2(_32847), .Q(_38681) );
  nnd2s1 _38719_inst ( .DIN1(_38683), .DIN2(_38684), .Q(
        _____________________________108________) );
  nnd2s1 _38720_inst ( .DIN1(_38685), .DIN2(_38686), .Q(_38684) );
  xor2s1 _38721_inst ( .DIN1(_33714), .DIN2(_26376), .Q(_38686) );
  nor2s1 _38722_inst ( .DIN1(_26260), .DIN2(_26400), .Q(_33714) );
  nor2s1 _38723_inst ( .DIN1(_27039), .DIN2(_36633), .Q(_38685) );
  nnd2s1 _38724_inst ( .DIN1(_29184), .DIN2(_33696), .Q(_36633) );
  nnd2s1 _38725_inst ( .DIN1(_29206), .DIN2(_38687), .Q(_38683) );
  nnd2s1 _38726_inst ( .DIN1(_38688), .DIN2(_38689), .Q(_38687) );
  nnd2s1 _38727_inst ( .DIN1(_38690), .DIN2(_33536), .Q(_38689) );
  xor2s1 _38728_inst ( .DIN1(_38691), .DIN2(_53327), .Q(_38690) );
  nnd2s1 _38729_inst ( .DIN1(_38668), .DIN2(_38665), .Q(_38691) );
  nnd2s1 _38730_inst ( .DIN1(_37755), .DIN2(_38692), .Q(_38665) );
  or2s1 _38731_inst ( .DIN1(_38692), .DIN2(_37755), .Q(_38668) );
  xor2s1 _38732_inst ( .DIN1(_38591), .DIN2(_38693), .Q(_37755) );
  xor2s1 _38733_inst ( .DIN1(_26323), .DIN2(_38673), .Q(_38693) );
  nnd2s1 _38734_inst ( .DIN1(_38694), .DIN2(_38695), .Q(_38673) );
  nnd2s1 _38735_inst ( .DIN1(_53375), .DIN2(_38696), .Q(_38695) );
  nnd2s1 _38736_inst ( .DIN1(_38587), .DIN2(_38697), .Q(_38696) );
  xor2s1 _38737_inst ( .DIN1(_32612), .DIN2(_38698), .Q(_38694) );
  nor2s1 _38738_inst ( .DIN1(_38587), .DIN2(_38697), .Q(_38698) );
  xor2s1 _38739_inst ( .DIN1(_38679), .DIN2(_38699), .Q(_38591) );
  nnd2s1 _38740_inst ( .DIN1(_38700), .DIN2(_38701), .Q(_38679) );
  nnd2s1 _38741_inst ( .DIN1(_53346), .DIN2(_38702), .Q(_38701) );
  or2s1 _38742_inst ( .DIN1(_38703), .DIN2(_26318), .Q(_38702) );
  nnd2s1 _38743_inst ( .DIN1(_38703), .DIN2(_26318), .Q(_38700) );
  nnd2s1 _38744_inst ( .DIN1(_38704), .DIN2(_38705), .Q(_38692) );
  nnd2s1 _38745_inst ( .DIN1(_53328), .DIN2(_38706), .Q(_38705) );
  or2s1 _38746_inst ( .DIN1(_38707), .DIN2(_37769), .Q(_38706) );
  nnd2s1 _38747_inst ( .DIN1(_37769), .DIN2(_38707), .Q(_38704) );
  hi1s1 _38748_inst ( .DIN(_38708), .Q(_37769) );
  nnd2s1 _38749_inst ( .DIN1(_38709), .DIN2(_38662), .Q(_38688) );
  xor2s1 _38750_inst ( .DIN1(_26456), .DIN2(_38710), .Q(_38709) );
  nnd2s1 _38751_inst ( .DIN1(_53326), .DIN2(_53325), .Q(_38710) );
  hi1s1 _38752_inst ( .DIN(_29184), .Q(_29206) );
  nnd2s1 _38753_inst ( .DIN1(_38711), .DIN2(_37854), .Q(_29184) );
  and2s1 _38754_inst ( .DIN1(_38712), .DIN2(_38713), .Q(_37854) );
  nor2s1 _38755_inst ( .DIN1(_31809), .DIN2(_34489), .Q(_38712) );
  nor2s1 _38756_inst ( .DIN1(_38714), .DIN2(_33182), .Q(_38711) );
  nnd2s1 _38757_inst ( .DIN1(_38715), .DIN2(_33229), .Q(
        _____________________________107________) );
  nnd2s1 _38758_inst ( .DIN1(_35873), .DIN2(_27509), .Q(_33229) );
  nor2s1 _38759_inst ( .DIN1(_38716), .DIN2(_38717), .Q(_38715) );
  nor2s1 _38760_inst ( .DIN1(_27509), .DIN2(_38718), .Q(_38717) );
  nnd2s1 _38761_inst ( .DIN1(_38719), .DIN2(_38720), .Q(_38718) );
  nnd2s1 _38762_inst ( .DIN1(_38721), .DIN2(_38722), .Q(_38720) );
  xor2s1 _38763_inst ( .DIN1(_38723), .DIN2(_38724), .Q(_38722) );
  xor2s1 _38764_inst ( .DIN1(_53261), .DIN2(_53329), .Q(_38724) );
  nnd2s1 _38765_inst ( .DIN1(_26284), .DIN2(_26553), .Q(_38723) );
  nor2s1 _38766_inst ( .DIN1(_38493), .DIN2(_26771), .Q(_38721) );
  xor2s1 _38767_inst ( .DIN1(_29579), .DIN2(_38725), .Q(_38719) );
  nnd2s1 _38768_inst ( .DIN1(_33536), .DIN2(_38726), .Q(_38725) );
  xor2s1 _38769_inst ( .DIN1(_38727), .DIN2(_38728), .Q(_38726) );
  xor2s1 _38770_inst ( .DIN1(_38707), .DIN2(_38708), .Q(_38728) );
  xor2s1 _38771_inst ( .DIN1(_38729), .DIN2(_38611), .Q(_38708) );
  hi1s1 _38772_inst ( .DIN(_38587), .Q(_38611) );
  xor2s1 _38773_inst ( .DIN1(_38703), .DIN2(_38730), .Q(_38587) );
  xor2s1 _38774_inst ( .DIN1(_53346), .DIN2(_53377), .Q(_38730) );
  nnd2s1 _38775_inst ( .DIN1(_38731), .DIN2(_38732), .Q(_38703) );
  nnd2s1 _38776_inst ( .DIN1(_38733), .DIN2(_26332), .Q(_38732) );
  nnd2s1 _38777_inst ( .DIN1(_38734), .DIN2(_38589), .Q(_38733) );
  or2s1 _38778_inst ( .DIN1(_38734), .DIN2(_38589), .Q(_38731) );
  xor2s1 _38779_inst ( .DIN1(_38697), .DIN2(_53375), .Q(_38729) );
  nnd2s1 _38780_inst ( .DIN1(_38735), .DIN2(_38736), .Q(_38697) );
  nnd2s1 _38781_inst ( .DIN1(_53373), .DIN2(_38737), .Q(_38736) );
  nnd2s1 _38782_inst ( .DIN1(_38586), .DIN2(_38738), .Q(_38737) );
  or2s1 _38783_inst ( .DIN1(_38738), .DIN2(_38586), .Q(_38735) );
  nnd2s1 _38784_inst ( .DIN1(_38739), .DIN2(_38740), .Q(_38707) );
  nnd2s1 _38785_inst ( .DIN1(_38741), .DIN2(_26550), .Q(_38740) );
  or2s1 _38786_inst ( .DIN1(_38742), .DIN2(_37808), .Q(_38741) );
  nnd2s1 _38787_inst ( .DIN1(_37808), .DIN2(_38742), .Q(_38739) );
  xor2s1 _38788_inst ( .DIN1(_26605), .DIN2(_29544), .Q(_38727) );
  nor2s1 _38789_inst ( .DIN1(_27512), .DIN2(_38743), .Q(_38716) );
  nor2s1 _38790_inst ( .DIN1(_38744), .DIN2(_28100), .Q(_38743) );
  xnr2s1 _38791_inst ( .DIN1(_53331), .DIN2(_53330), .Q(_38744) );
  nnd2s1 _38792_inst ( .DIN1(_38745), .DIN2(_31861), .Q(
        _____________________________106________) );
  nor2s1 _38793_inst ( .DIN1(_38746), .DIN2(_38747), .Q(_38745) );
  nor2s1 _38794_inst ( .DIN1(_31864), .DIN2(_38748), .Q(_38747) );
  nnd2s1 _38795_inst ( .DIN1(_38749), .DIN2(_38750), .Q(_38748) );
  nnd2s1 _38796_inst ( .DIN1(_33536), .DIN2(_38751), .Q(_38750) );
  xor2s1 _38797_inst ( .DIN1(_37808), .DIN2(_38752), .Q(_38751) );
  xor2s1 _38798_inst ( .DIN1(_26550), .DIN2(_38742), .Q(_38752) );
  nnd2s1 _38799_inst ( .DIN1(_38753), .DIN2(_38754), .Q(_38742) );
  nnd2s1 _38800_inst ( .DIN1(_53334), .DIN2(_38755), .Q(_38754) );
  or2s1 _38801_inst ( .DIN1(_38756), .DIN2(_37830), .Q(_38755) );
  nnd2s1 _38802_inst ( .DIN1(_37830), .DIN2(_38756), .Q(_38753) );
  xor2s1 _38803_inst ( .DIN1(_38586), .DIN2(_38757), .Q(_37808) );
  xor2s1 _38804_inst ( .DIN1(_26333), .DIN2(_38738), .Q(_38757) );
  nnd2s1 _38805_inst ( .DIN1(_38758), .DIN2(_38759), .Q(_38738) );
  nnd2s1 _38806_inst ( .DIN1(_38760), .DIN2(_26322), .Q(_38759) );
  or2s1 _38807_inst ( .DIN1(_38761), .DIN2(_38580), .Q(_38760) );
  nnd2s1 _38808_inst ( .DIN1(_38580), .DIN2(_38761), .Q(_38758) );
  xnr2s1 _38809_inst ( .DIN1(_38762), .DIN2(_38734), .Q(_38586) );
  xnr2s1 _38810_inst ( .DIN1(_32657), .DIN2(_38763), .Q(_38734) );
  nor2s1 _38811_inst ( .DIN1(_38764), .DIN2(_38765), .Q(_38763) );
  nor2s1 _38812_inst ( .DIN1(_53380), .DIN2(_38766), .Q(_38765) );
  nor2s1 _38813_inst ( .DIN1(_38767), .DIN2(_27558), .Q(_38764) );
  and2s1 _38814_inst ( .DIN1(_38766), .DIN2(_53380), .Q(_38767) );
  xor2s1 _38815_inst ( .DIN1(_26332), .DIN2(_53381), .Q(_38762) );
  hi1s1 _38816_inst ( .DIN(_33531), .Q(_33536) );
  nnd2s1 _38817_inst ( .DIN1(_38768), .DIN2(_33520), .Q(_33531) );
  nnd2s1 _38818_inst ( .DIN1(_38662), .DIN2(_26284), .Q(_38749) );
  nor2s1 _38819_inst ( .DIN1(_53332), .DIN2(_31907), .Q(_38746) );
  nor2s1 _38820_inst ( .DIN1(_38769), .DIN2(_27500), .Q(
        _____________________________105________) );
  nor2s1 _38821_inst ( .DIN1(_38770), .DIN2(_38771), .Q(_38769) );
  and2s1 _38822_inst ( .DIN1(_26447), .DIN2(_38772), .Q(_38771) );
  nor2s1 _38823_inst ( .DIN1(_38773), .DIN2(_38774), .Q(_38770) );
  xor2s1 _38824_inst ( .DIN1(_37830), .DIN2(_38775), .Q(_38774) );
  xor2s1 _38825_inst ( .DIN1(_26582), .DIN2(_38756), .Q(_38775) );
  nnd2s1 _38826_inst ( .DIN1(_38776), .DIN2(_38777), .Q(_38756) );
  nnd2s1 _38827_inst ( .DIN1(_38778), .DIN2(_26474), .Q(_38777) );
  nnd2s1 _38828_inst ( .DIN1(_38779), .DIN2(_38780), .Q(_38778) );
  hi1s1 _38829_inst ( .DIN(_37846), .Q(_38780) );
  nnd2s1 _38830_inst ( .DIN1(_37846), .DIN2(_38781), .Q(_38776) );
  xor2s1 _38831_inst ( .DIN1(_38580), .DIN2(_38782), .Q(_37830) );
  xor2s1 _38832_inst ( .DIN1(_26322), .DIN2(_38761), .Q(_38782) );
  nnd2s1 _38833_inst ( .DIN1(_38783), .DIN2(_38784), .Q(_38761) );
  nnd2s1 _38834_inst ( .DIN1(_38785), .DIN2(_26336), .Q(_38784) );
  or2s1 _38835_inst ( .DIN1(_38786), .DIN2(_38579), .Q(_38785) );
  nnd2s1 _38836_inst ( .DIN1(_38786), .DIN2(_38579), .Q(_38783) );
  xnr2s1 _38837_inst ( .DIN1(_38787), .DIN2(_38766), .Q(_38580) );
  nnd2s1 _38838_inst ( .DIN1(_38788), .DIN2(_38789), .Q(_38766) );
  nnd2s1 _38839_inst ( .DIN1(_53350), .DIN2(_38790), .Q(_38789) );
  nnd2s1 _38840_inst ( .DIN1(_38791), .DIN2(_53381), .Q(_38790) );
  nnd2s1 _38841_inst ( .DIN1(_38792), .DIN2(_38793), .Q(
        _____________________________104________) );
  nnd2s1 _38842_inst ( .DIN1(_38794), .DIN2(_33053), .Q(_38793) );
  nnd2s1 _38843_inst ( .DIN1(_33951), .DIN2(_53293), .Q(_38794) );
  nor2s1 _38844_inst ( .DIN1(_33489), .DIN2(_27066), .Q(_33951) );
  nnd2s1 _38845_inst ( .DIN1(_38795), .DIN2(_33069), .Q(_38792) );
  hi1s1 _38846_inst ( .DIN(_33053), .Q(_33069) );
  nnd2s1 _38847_inst ( .DIN1(_28738), .DIN2(_38163), .Q(_33053) );
  hi1s1 _38848_inst ( .DIN(_28733), .Q(_28738) );
  nnd2s1 _38849_inst ( .DIN1(_33489), .DIN2(_35368), .Q(_28733) );
  nor2s1 _38850_inst ( .DIN1(_38796), .DIN2(_38797), .Q(_38795) );
  nor2s1 _38851_inst ( .DIN1(_27448), .DIN2(_38798), .Q(_38797) );
  nnd2s1 _38852_inst ( .DIN1(_38799), .DIN2(_38662), .Q(_38798) );
  xor2s1 _38853_inst ( .DIN1(_53329), .DIN2(_53336), .Q(_38799) );
  nor2s1 _38854_inst ( .DIN1(_38773), .DIN2(_38800), .Q(_38796) );
  xor2s1 _38855_inst ( .DIN1(_37846), .DIN2(_38801), .Q(_38800) );
  xor2s1 _38856_inst ( .DIN1(_26474), .DIN2(_38779), .Q(_38801) );
  hi1s1 _38857_inst ( .DIN(_38781), .Q(_38779) );
  nnd2s1 _38858_inst ( .DIN1(_38802), .DIN2(_38803), .Q(_38781) );
  nnd2s1 _38859_inst ( .DIN1(_53337), .DIN2(_38804), .Q(_38803) );
  or2s1 _38860_inst ( .DIN1(_38805), .DIN2(_37867), .Q(_38804) );
  nnd2s1 _38861_inst ( .DIN1(_37867), .DIN2(_38805), .Q(_38802) );
  xnr2s1 _38862_inst ( .DIN1(_38806), .DIN2(_38786), .Q(_37846) );
  nnd2s1 _38863_inst ( .DIN1(_38807), .DIN2(_38808), .Q(_38786) );
  nnd2s1 _38864_inst ( .DIN1(_38809), .DIN2(_26319), .Q(_38808) );
  or2s1 _38865_inst ( .DIN1(_38810), .DIN2(_38574), .Q(_38809) );
  nnd2s1 _38866_inst ( .DIN1(_38574), .DIN2(_38810), .Q(_38807) );
  xor2s1 _38867_inst ( .DIN1(_38579), .DIN2(_53372), .Q(_38806) );
  nnd2s1 _38868_inst ( .DIN1(_38811), .DIN2(_38812), .Q(_38579) );
  nnd2s1 _38869_inst ( .DIN1(_38813), .DIN2(_38791), .Q(_38812) );
  hi1s1 _38870_inst ( .DIN(_38814), .Q(_38791) );
  nor2s1 _38871_inst ( .DIN1(_38815), .DIN2(_38816), .Q(_38811) );
  nor2s1 _38872_inst ( .DIN1(_53350), .DIN2(_38817), .Q(_38816) );
  xor2s1 _38873_inst ( .DIN1(_38814), .DIN2(_53381), .Q(_38817) );
  nor2s1 _38874_inst ( .DIN1(_26320), .DIN2(_38788), .Q(_38815) );
  nnd2s1 _38875_inst ( .DIN1(_38814), .DIN2(_38589), .Q(_38788) );
  nnd2s1 _38876_inst ( .DIN1(_38818), .DIN2(_38819), .Q(_38814) );
  nnd2s1 _38877_inst ( .DIN1(_53352), .DIN2(_38820), .Q(_38819) );
  or2s1 _38878_inst ( .DIN1(_38821), .DIN2(_26330), .Q(_38820) );
  nnd2s1 _38879_inst ( .DIN1(_38821), .DIN2(_26330), .Q(_38818) );
  nnd2s1 _38880_inst ( .DIN1(_38822), .DIN2(_38823), .Q(
        _____________________________103________) );
  nnd2s1 _38881_inst ( .DIN1(_29849), .DIN2(_38824), .Q(_38823) );
  nnd2s1 _38882_inst ( .DIN1(_38825), .DIN2(_38826), .Q(_38824) );
  nnd2s1 _38883_inst ( .DIN1(_38827), .DIN2(_38772), .Q(_38826) );
  xor2s1 _38884_inst ( .DIN1(_38828), .DIN2(_38829), .Q(_38827) );
  xor2s1 _38885_inst ( .DIN1(_53348), .DIN2(_53349), .Q(_38829) );
  nnd2s1 _38886_inst ( .DIN1(_53340), .DIN2(_26357), .Q(_38828) );
  nnd2s1 _38887_inst ( .DIN1(_38768), .DIN2(_38830), .Q(_38825) );
  xnr2s1 _38888_inst ( .DIN1(_37867), .DIN2(_38831), .Q(_38830) );
  xnr2s1 _38889_inst ( .DIN1(_53337), .DIN2(_38805), .Q(_38831) );
  nnd2s1 _38890_inst ( .DIN1(_38832), .DIN2(_38833), .Q(_38805) );
  nnd2s1 _38891_inst ( .DIN1(_53259), .DIN2(_38834), .Q(_38833) );
  or2s1 _38892_inst ( .DIN1(_38835), .DIN2(_37884), .Q(_38834) );
  nnd2s1 _38893_inst ( .DIN1(_37884), .DIN2(_38835), .Q(_38832) );
  xor2s1 _38894_inst ( .DIN1(_38836), .DIN2(_38837), .Q(_37867) );
  xnr2s1 _38895_inst ( .DIN1(_38574), .DIN2(_38810), .Q(_38837) );
  xor2s1 _38896_inst ( .DIN1(_38838), .DIN2(_38821), .Q(_38574) );
  nnd2s1 _38897_inst ( .DIN1(_38839), .DIN2(_38840), .Q(_38821) );
  nnd2s1 _38898_inst ( .DIN1(_38841), .DIN2(_26320), .Q(_38840) );
  or2s1 _38899_inst ( .DIN1(_38842), .DIN2(_53357), .Q(_38841) );
  nnd2s1 _38900_inst ( .DIN1(_53357), .DIN2(_38842), .Q(_38839) );
  xor2s1 _38901_inst ( .DIN1(_26221), .DIN2(_53380), .Q(_38838) );
  nnd2s1 _38902_inst ( .DIN1(_38843), .DIN2(_38844), .Q(_38810) );
  nnd2s1 _38903_inst ( .DIN1(_53376), .DIN2(_38845), .Q(_38844) );
  or2s1 _38904_inst ( .DIN1(_38846), .DIN2(_38573), .Q(_38845) );
  nnd2s1 _38905_inst ( .DIN1(_38573), .DIN2(_38846), .Q(_38843) );
  hi1s1 _38906_inst ( .DIN(_38847), .Q(_38573) );
  xor2s1 _38907_inst ( .DIN1(_38848), .DIN2(_53338), .Q(_38836) );
  nnd2s1 _38908_inst ( .DIN1(_38849), .DIN2(_29828), .Q(_38822) );
  nor2s1 _38909_inst ( .DIN1(_28381), .DIN2(_38850), .Q(_38849) );
  xor2s1 _38910_inst ( .DIN1(_26401), .DIN2(_28835), .Q(_38850) );
  nnd2s1 _38911_inst ( .DIN1(_38851), .DIN2(_31861), .Q(
        _____________________________102________) );
  nnd2s1 _38912_inst ( .DIN1(_38852), .DIN2(_36676), .Q(_31861) );
  nor2s1 _38913_inst ( .DIN1(_38853), .DIN2(_38714), .Q(_36676) );
  nor2s1 _38914_inst ( .DIN1(_31907), .DIN2(_33152), .Q(_38852) );
  nnd2s1 _38915_inst ( .DIN1(_38854), .DIN2(_38855), .Q(_33152) );
  nor2s1 _38916_inst ( .DIN1(_34490), .DIN2(_37411), .Q(_38855) );
  nor2s1 _38917_inst ( .DIN1(_37701), .DIN2(_33182), .Q(_38854) );
  nor2s1 _38918_inst ( .DIN1(_38856), .DIN2(_38857), .Q(_38851) );
  nor2s1 _38919_inst ( .DIN1(_31864), .DIN2(_38858), .Q(_38857) );
  nnd2s1 _38920_inst ( .DIN1(_38859), .DIN2(_38860), .Q(_38858) );
  nnd2s1 _38921_inst ( .DIN1(_38861), .DIN2(_38768), .Q(_38860) );
  xor2s1 _38922_inst ( .DIN1(_38862), .DIN2(_38835), .Q(_38861) );
  xnr2s1 _38923_inst ( .DIN1(_38863), .DIN2(_32615), .Q(_38835) );
  nor2s1 _38924_inst ( .DIN1(_29544), .DIN2(_38344), .Q(_32615) );
  nnd2s1 _38925_inst ( .DIN1(_38864), .DIN2(_38865), .Q(_29544) );
  nnd2s1 _38926_inst ( .DIN1(_38866), .DIN2(_38867), .Q(_38863) );
  nnd2s1 _38927_inst ( .DIN1(_38868), .DIN2(_26490), .Q(_38867) );
  or2s1 _38928_inst ( .DIN1(_38869), .DIN2(_37903), .Q(_38868) );
  nnd2s1 _38929_inst ( .DIN1(_37903), .DIN2(_38869), .Q(_38866) );
  hi1s1 _38930_inst ( .DIN(_38870), .Q(_37903) );
  xor2s1 _38931_inst ( .DIN1(_53259), .DIN2(_37884), .Q(_38862) );
  xor2s1 _38932_inst ( .DIN1(_38847), .DIN2(_26812), .Q(_37884) );
  nnd2s1 _38933_inst ( .DIN1(_38872), .DIN2(_38873), .Q(_38846) );
  nnd2s1 _38934_inst ( .DIN1(_38874), .DIN2(_26318), .Q(_38873) );
  or2s1 _38935_inst ( .DIN1(_38875), .DIN2(_38628), .Q(_38874) );
  nnd2s1 _38936_inst ( .DIN1(_38628), .DIN2(_38875), .Q(_38872) );
  hi1s1 _38937_inst ( .DIN(_38631), .Q(_38628) );
  hi1s1 _38938_inst ( .DIN(_53376), .Q(_34787) );
  xor2s1 _38939_inst ( .DIN1(_38842), .DIN2(_38876), .Q(_38847) );
  xor2s1 _38940_inst ( .DIN1(_53350), .DIN2(_53357), .Q(_38876) );
  nnd2s1 _38941_inst ( .DIN1(_38877), .DIN2(_38878), .Q(_38842) );
  nnd2s1 _38942_inst ( .DIN1(_38879), .DIN2(_26221), .Q(_38878) );
  or2s1 _38943_inst ( .DIN1(_38880), .DIN2(_53358), .Q(_38879) );
  nnd2s1 _38944_inst ( .DIN1(_53358), .DIN2(_38880), .Q(_38877) );
  nnd2s1 _38945_inst ( .DIN1(_38772), .DIN2(_26357), .Q(_38859) );
  nor2s1 _38946_inst ( .DIN1(_27082), .DIN2(_38493), .Q(_38772) );
  nor2s1 _38947_inst ( .DIN1(_31907), .DIN2(_38881), .Q(_38856) );
  and2s1 _38948_inst ( .DIN1(______[0]), .DIN2(_53342), .Q(_38881) );
  hi1s1 _38949_inst ( .DIN(_31864), .Q(_31907) );
  nnd2s1 _38950_inst ( .DIN1(_38882), .DIN2(_38883), .Q(_31864) );
  nor2s1 _38951_inst ( .DIN1(_38884), .DIN2(_37411), .Q(_38883) );
  nor2s1 _38952_inst ( .DIN1(_38853), .DIN2(_38885), .Q(_38882) );
  nnd2s1 _38953_inst ( .DIN1(_38886), .DIN2(_38887), .Q(
        _____________________________101________) );
  nnd2s1 _38954_inst ( .DIN1(_38888), .DIN2(_32847), .Q(_38887) );
  nor2s1 _38955_inst ( .DIN1(_38889), .DIN2(_38890), .Q(_38888) );
  xnr2s1 _38956_inst ( .DIN1(_53187), .DIN2(_32871), .Q(_38890) );
  nnd2s1 _38957_inst ( .DIN1(_53343), .DIN2(_53344), .Q(_32871) );
  nor2s1 _38958_inst ( .DIN1(_31196), .DIN2(_33294), .Q(_38889) );
  nnd2s1 _38959_inst ( .DIN1(_38891), .DIN2(_36832), .Q(_33294) );
  nor2s1 _38960_inst ( .DIN1(_27822), .DIN2(_37987), .Q(_38891) );
  hi1s1 _38961_inst ( .DIN(_38682), .Q(_31196) );
  nnd2s1 _38962_inst ( .DIN1(_38892), .DIN2(_32868), .Q(_38886) );
  hi1s1 _38963_inst ( .DIN(_32847), .Q(_32868) );
  nnd2s1 _38964_inst ( .DIN1(_38893), .DIN2(_37298), .Q(_32847) );
  and2s1 _38965_inst ( .DIN1(_38894), .DIN2(_37986), .Q(_37298) );
  and2s1 _38966_inst ( .DIN1(_38895), .DIN2(_38682), .Q(_37986) );
  nor2s1 _38967_inst ( .DIN1(_27822), .DIN2(_36833), .Q(_38895) );
  hi1s1 _38968_inst ( .DIN(_37983), .Q(_36833) );
  nor2s1 _38969_inst ( .DIN1(_27821), .DIN2(_36827), .Q(_38894) );
  hi1s1 _38970_inst ( .DIN(_37984), .Q(_36827) );
  nor2s1 _38971_inst ( .DIN1(_37931), .DIN2(_36829), .Q(_38893) );
  nnd2s1 _38972_inst ( .DIN1(_38896), .DIN2(_38897), .Q(_38892) );
  nnd2s1 _38973_inst ( .DIN1(_38898), .DIN2(_38773), .Q(_38897) );
  nnd2s1 _38974_inst ( .DIN1(_26344), .DIN2(_38662), .Q(_38898) );
  nnd2s1 _38975_inst ( .DIN1(_38899), .DIN2(_38768), .Q(_38896) );
  xor2s1 _38976_inst ( .DIN1(_38870), .DIN2(_38900), .Q(_38899) );
  xor2s1 _38977_inst ( .DIN1(_26490), .DIN2(_38869), .Q(_38900) );
  nnd2s1 _38978_inst ( .DIN1(_38901), .DIN2(_38902), .Q(_38869) );
  nnd2s1 _38979_inst ( .DIN1(_53347), .DIN2(_38903), .Q(_38902) );
  nnd2s1 _38980_inst ( .DIN1(_38904), .DIN2(_38905), .Q(_38903) );
  or2s1 _38981_inst ( .DIN1(_38905), .DIN2(_38904), .Q(_38901) );
  hi1s1 _38982_inst ( .DIN(_37920), .Q(_38904) );
  xor2s1 _38983_inst ( .DIN1(_38631), .DIN2(_26784), .Q(_38870) );
  nnd2s1 _38984_inst ( .DIN1(_38907), .DIN2(_38908), .Q(_38875) );
  nnd2s1 _38985_inst ( .DIN1(_38909), .DIN2(_26332), .Q(_38908) );
  xor2s1 _38986_inst ( .DIN1(_38910), .DIN2(_37426), .Q(_38909) );
  xnr2s1 _38987_inst ( .DIN1(_30081), .DIN2(_32612), .Q(_37426) );
  hi1s1 _38988_inst ( .DIN(_32427), .Q(_32612) );
  nnd2s1 _38989_inst ( .DIN1(_38911), .DIN2(_38528), .Q(_32427) );
  and2s1 _38990_inst ( .DIN1(_36898), .DIN2(_38912), .Q(_38911) );
  xnr2s1 _38991_inst ( .DIN1(_38913), .DIN2(_38880), .Q(_38631) );
  nnd2s1 _38992_inst ( .DIN1(_38914), .DIN2(_38915), .Q(_38880) );
  nnd2s1 _38993_inst ( .DIN1(_38916), .DIN2(_26396), .Q(_38915) );
  or2s1 _38994_inst ( .DIN1(_38917), .DIN2(_53467), .Q(_38916) );
  nnd2s1 _38995_inst ( .DIN1(_53467), .DIN2(_38917), .Q(_38914) );
  xor2s1 _38996_inst ( .DIN1(_26448), .DIN2(_53352), .Q(_38913) );
  nnd2s1 _38997_inst ( .DIN1(_38918), .DIN2(_28238), .Q(
        _____________________________100________) );
  nnd2s1 _38998_inst ( .DIN1(_38919), .DIN2(_28241), .Q(_28238) );
  nor2s1 _38999_inst ( .DIN1(_38920), .DIN2(_38921), .Q(_38918) );
  nor2s1 _39000_inst ( .DIN1(_28241), .DIN2(_38922), .Q(_38921) );
  nnd2s1 _39001_inst ( .DIN1(_38923), .DIN2(_38924), .Q(_38922) );
  nnd2s1 _39002_inst ( .DIN1(_38925), .DIN2(_38768), .Q(_38924) );
  hi1s1 _39003_inst ( .DIN(_38773), .Q(_38768) );
  nnd2s1 _39004_inst ( .DIN1(_38464), .DIN2(_38493), .Q(_38773) );
  nor2s1 _39005_inst ( .DIN1(_38314), .DIN2(_38133), .Q(_38464) );
  xor2s1 _39006_inst ( .DIN1(_38926), .DIN2(_38927), .Q(_38925) );
  xor2s1 _39007_inst ( .DIN1(_38905), .DIN2(_37920), .Q(_38927) );
  nnd2s1 _39008_inst ( .DIN1(_38928), .DIN2(_38929), .Q(_37920) );
  nnd2s1 _39009_inst ( .DIN1(_38930), .DIN2(_26332), .Q(_38929) );
  nnd2s1 _39010_inst ( .DIN1(_38910), .DIN2(_38907), .Q(_38930) );
  nnd2s1 _39011_inst ( .DIN1(_38931), .DIN2(_38634), .Q(_38907) );
  hi1s1 _39012_inst ( .DIN(_38932), .Q(_38634) );
  nnd2s1 _39013_inst ( .DIN1(_38932), .DIN2(_38933), .Q(_38910) );
  nnd2s1 _39014_inst ( .DIN1(_38934), .DIN2(_53379), .Q(_38928) );
  xor2s1 _39015_inst ( .DIN1(_38932), .DIN2(_38933), .Q(_38934) );
  hi1s1 _39016_inst ( .DIN(_38931), .Q(_38933) );
  xor2s1 _39017_inst ( .DIN1(_38935), .DIN2(_2064), .Q(_38931) );
  nnd2s1 _39018_inst ( .DIN1(_38936), .DIN2(_38937), .Q(_38935) );
  nnd2s1 _39019_inst ( .DIN1(_38938), .DIN2(_27558), .Q(_38937) );
  or2s1 _39020_inst ( .DIN1(_38939), .DIN2(_38642), .Q(_38938) );
  nnd2s1 _39021_inst ( .DIN1(_38642), .DIN2(_38939), .Q(_38936) );
  xor2s1 _39022_inst ( .DIN1(_38917), .DIN2(_38940), .Q(_38932) );
  xor2s1 _39023_inst ( .DIN1(_53357), .DIN2(_53467), .Q(_38940) );
  nnd2s1 _39024_inst ( .DIN1(_38941), .DIN2(_38942), .Q(_38917) );
  nnd2s1 _39025_inst ( .DIN1(_38943), .DIN2(_26329), .Q(_38942) );
  or2s1 _39026_inst ( .DIN1(_26448), .DIN2(_38944), .Q(_38943) );
  nnd2s1 _39027_inst ( .DIN1(_38944), .DIN2(_26448), .Q(_38941) );
  nnd2s1 _39028_inst ( .DIN1(_38945), .DIN2(_38946), .Q(_38905) );
  nnd2s1 _39029_inst ( .DIN1(_38947), .DIN2(_26220), .Q(_38946) );
  nnd2s1 _39030_inst ( .DIN1(_32867), .DIN2(_32866), .Q(_38947) );
  or2s1 _39031_inst ( .DIN1(_32866), .DIN2(_32867), .Q(_38945) );
  xor2s1 _39032_inst ( .DIN1(_38642), .DIN2(_38948), .Q(_32867) );
  xor2s1 _39033_inst ( .DIN1(_27558), .DIN2(_38939), .Q(_38948) );
  nnd2s1 _39034_inst ( .DIN1(_38949), .DIN2(_38950), .Q(_38939) );
  nnd2s1 _39035_inst ( .DIN1(_38951), .DIN2(_38589), .Q(_38950) );
  or2s1 _39036_inst ( .DIN1(_38952), .DIN2(_38953), .Q(_38951) );
  nnd2s1 _39037_inst ( .DIN1(_38953), .DIN2(_38952), .Q(_38949) );
  hi1s1 _39038_inst ( .DIN(_38641), .Q(_38953) );
  xnr2s1 _39039_inst ( .DIN1(_38954), .DIN2(_38944), .Q(_38642) );
  nnd2s1 _39040_inst ( .DIN1(_38955), .DIN2(_38956), .Q(_38944) );
  nnd2s1 _39041_inst ( .DIN1(_38957), .DIN2(_26698), .Q(_38956) );
  nnd2s1 _39042_inst ( .DIN1(_53467), .DIN2(_38958), .Q(_38957) );
  or2s1 _39043_inst ( .DIN1(_38958), .DIN2(_53467), .Q(_38955) );
  nnd2s1 _39044_inst ( .DIN1(_38959), .DIN2(_38960), .Q(_32866) );
  nnd2s1 _39045_inst ( .DIN1(_53015), .DIN2(_38961), .Q(_38960) );
  nnd2s1 _39046_inst ( .DIN1(_37952), .DIN2(_32881), .Q(_38961) );
  nnd2s1 _39047_inst ( .DIN1(_38962), .DIN2(_32880), .Q(_38959) );
  hi1s1 _39048_inst ( .DIN(_37952), .Q(_32880) );
  xor2s1 _39049_inst ( .DIN1(_38641), .DIN2(_38963), .Q(_37952) );
  xor2s1 _39050_inst ( .DIN1(_38589), .DIN2(_38952), .Q(_38963) );
  nnd2s1 _39051_inst ( .DIN1(_38964), .DIN2(_38965), .Q(_38952) );
  nnd2s1 _39052_inst ( .DIN1(_38966), .DIN2(_26330), .Q(_38965) );
  nnd2s1 _39053_inst ( .DIN1(_38967), .DIN2(_38968), .Q(_38966) );
  nnd2s1 _39054_inst ( .DIN1(_38969), .DIN2(_38970), .Q(_38964) );
  hi1s1 _39055_inst ( .DIN(_38968), .Q(_38969) );
  xnr2s1 _39056_inst ( .DIN1(_38971), .DIN2(_38958), .Q(_38641) );
  nnd2s1 _39057_inst ( .DIN1(_53353), .DIN2(_38972), .Q(_38958) );
  nnd2s1 _39058_inst ( .DIN1(_26242), .DIN2(_26698), .Q(_38972) );
  xor2s1 _39059_inst ( .DIN1(_26341), .DIN2(_53366), .Q(_38971) );
  hi1s1 _39060_inst ( .DIN(_32881), .Q(_38962) );
  nnd2s1 _39061_inst ( .DIN1(_37997), .DIN2(_26441), .Q(_32881) );
  hi1s1 _39062_inst ( .DIN(_32891), .Q(_37997) );
  xor2s1 _39063_inst ( .DIN1(_38968), .DIN2(_38973), .Q(_32891) );
  xor2s1 _39064_inst ( .DIN1(_53380), .DIN2(_38967), .Q(_38973) );
  hi1s1 _39065_inst ( .DIN(_38970), .Q(_38967) );
  nnd2s1 _39066_inst ( .DIN1(_38974), .DIN2(_38975), .Q(_38970) );
  nnd2s1 _39067_inst ( .DIN1(_38976), .DIN2(_53366), .Q(_38975) );
  nor2s1 _39068_inst ( .DIN1(_53352), .DIN2(_26242), .Q(_38976) );
  nnd2s1 _39069_inst ( .DIN1(_38977), .DIN2(_26320), .Q(_38974) );
  nnd2s1 _39070_inst ( .DIN1(_38978), .DIN2(_38979), .Q(_38977) );
  nnd2s1 _39071_inst ( .DIN1(_38980), .DIN2(_38981), .Q(_38979) );
  nor2s1 _39072_inst ( .DIN1(_53358), .DIN2(_38982), .Q(_38981) );
  nnd2s1 _39073_inst ( .DIN1(_26396), .DIN2(_26221), .Q(_38982) );
  nor2s1 _39074_inst ( .DIN1(_53467), .DIN2(_26329), .Q(_38980) );
  nor2s1 _39075_inst ( .DIN1(_38983), .DIN2(_38984), .Q(_38978) );
  nor2s1 _39076_inst ( .DIN1(_38985), .DIN2(_26242), .Q(_38984) );
  nor2s1 _39077_inst ( .DIN1(_53366), .DIN2(_26221), .Q(_38985) );
  nor2s1 _39078_inst ( .DIN1(_53366), .DIN2(_53369), .Q(_38983) );
  xor2s1 _39079_inst ( .DIN1(_38986), .DIN2(_38987), .Q(_38968) );
  xor2s1 _39080_inst ( .DIN1(_53353), .DIN2(_53369), .Q(_38987) );
  nnd2s1 _39081_inst ( .DIN1(_53366), .DIN2(_26242), .Q(_38986) );
  xor2s1 _39082_inst ( .DIN1(_26519), .DIN2(_31456), .Q(_38926) );
  nnd2s1 _39083_inst ( .DIN1(_38864), .DIN2(_36898), .Q(_31456) );
  nnd2s1 _39084_inst ( .DIN1(_38988), .DIN2(_38989), .Q(_38923) );
  xor2s1 _39085_inst ( .DIN1(_53340), .DIN2(_26344), .Q(_38989) );
  nor2s1 _39086_inst ( .DIN1(_38493), .DIN2(_28100), .Q(_38988) );
  hi1s1 _39087_inst ( .DIN(_38662), .Q(_38493) );
  nnd2s1 _39088_inst ( .DIN1(_38466), .DIN2(_38990), .Q(_38662) );
  nor2s1 _39089_inst ( .DIN1(_28250), .DIN2(_38991), .Q(_38920) );
  nor2s1 _39090_inst ( .DIN1(_26772), .DIN2(_38992), .Q(_38991) );
  xor2s1 _39091_inst ( .DIN1(_38993), .DIN2(_38994), .Q(_38992) );
  xor2s1 _39092_inst ( .DIN1(_52850), .DIN2(_53409), .Q(_38994) );
  nor2s1 _39093_inst ( .DIN1(_26668), .DIN2(_26305), .Q(_38993) );
  nor2s1 _39094_inst ( .DIN1(_38995), .DIN2(_38996), .Q(
        _______9____2________________9____________________) );
  nor2s1 _39095_inst ( .DIN1(_38997), .DIN2(_38998), .Q(_38995) );
  nnd2s1 _39096_inst ( .DIN1(_38999), .DIN2(_39000), .Q(_38998) );
  nnd2s1 _39097_inst ( .DIN1(_39001), .DIN2(_39002), .Q(_39000) );
  nnd2s1 _39098_inst ( .DIN1(_39003), .DIN2(_26330), .Q(_38999) );
  nor2s1 _39099_inst ( .DIN1(_39004), .DIN2(_38996), .Q(
        _______8____2________________8____________________) );
  nor2s1 _39100_inst ( .DIN1(_39005), .DIN2(_39006), .Q(_39004) );
  nnd2s1 _39101_inst ( .DIN1(_39007), .DIN2(_39008), .Q(_39006) );
  nnd2s1 _39102_inst ( .DIN1(_34947), .DIN2(_26854), .Q(_39008) );
  nnd2s1 _39103_inst ( .DIN1(_39009), .DIN2(_34943), .Q(_39007) );
  nnd2s1 _39104_inst ( .DIN1(_53350), .DIN2(______[20]), .Q(_39009) );
  hi1s1 _39105_inst ( .DIN(_34935), .Q(_39005) );
  nnd2s1 _39106_inst ( .DIN1(_39010), .DIN2(_36436), .Q(
        _______7____2________________7____________________) );
  nor2s1 _39107_inst ( .DIN1(_39011), .DIN2(_39012), .Q(_39010) );
  nor2s1 _39108_inst ( .DIN1(_39013), .DIN2(_39014), .Q(_39012) );
  xnr2s1 _39109_inst ( .DIN1(_38813), .DIN2(_38787), .Q(_39013) );
  xor2s1 _39110_inst ( .DIN1(_27558), .DIN2(_26330), .Q(_38787) );
  nor2s1 _39111_inst ( .DIN1(_26320), .DIN2(_38589), .Q(_38813) );
  nor2s1 _39112_inst ( .DIN1(_34943), .DIN2(_39015), .Q(_39011) );
  nnd2s1 _39113_inst ( .DIN1(_39016), .DIN2(_27994), .Q(
        _______6____2________________6____________________) );
  nor2s1 _39114_inst ( .DIN1(_39017), .DIN2(_39018), .Q(_39016) );
  nor2s1 _39115_inst ( .DIN1(_39019), .DIN2(_39014), .Q(_39018) );
  nnd2s1 _39116_inst ( .DIN1(_34935), .DIN2(_34943), .Q(_39014) );
  nnd2s1 _39117_inst ( .DIN1(_39020), .DIN2(_39021), .Q(_34935) );
  nor2s1 _39118_inst ( .DIN1(_34960), .DIN2(_34947), .Q(_39021) );
  xor2s1 _39119_inst ( .DIN1(_34925), .DIN2(_26406), .Q(_39019) );
  nor2s1 _39120_inst ( .DIN1(_26221), .DIN2(_53090), .Q(_34925) );
  nor2s1 _39121_inst ( .DIN1(_28646), .DIN2(_34943), .Q(_39017) );
  hi1s1 _39122_inst ( .DIN(_34947), .Q(_34943) );
  nor2s1 _39123_inst ( .DIN1(_39022), .DIN2(_34712), .Q(_34947) );
  nnd2s1 _39124_inst ( .DIN1(_39023), .DIN2(_39024), .Q(_34712) );
  nor2s1 _39125_inst ( .DIN1(_34891), .DIN2(_39025), .Q(_39024) );
  nnd2s1 _39126_inst ( .DIN1(_39026), .DIN2(_39027), .Q(_39025) );
  nor2s1 _39127_inst ( .DIN1(_39028), .DIN2(_39029), .Q(_39023) );
  xor2s1 _39128_inst ( .DIN1(_27338), .DIN2(_39030), .Q(_39029) );
  nor2s1 _39129_inst ( .DIN1(_39031), .DIN2(_34531), .Q(_39030) );
  nnd2s1 _39130_inst ( .DIN1(_39032), .DIN2(_34638), .Q(_39022) );
  nnd2s1 _39131_inst ( .DIN1(_39033), .DIN2(_39034), .Q(
        _______5____2________________5____________________) );
  and2s1 _39132_inst ( .DIN1(_39035), .DIN2(_39036), .Q(_39033) );
  nnd2s1 _39133_inst ( .DIN1(_38954), .DIN2(_35685), .Q(_39036) );
  xor2s1 _39134_inst ( .DIN1(_26329), .DIN2(_53358), .Q(_38954) );
  nnd2s1 _39135_inst ( .DIN1(______[5]), .DIN2(_28317), .Q(_39035) );
  hi1s1 _39136_inst ( .DIN(_35735), .Q(_28317) );
  nnd2s1 _39137_inst ( .DIN1(_39037), .DIN2(_36266), .Q(
        _______4____2________________4____________________) );
  nor2s1 _39138_inst ( .DIN1(_39038), .DIN2(_39039), .Q(_39037) );
  nor2s1 _39139_inst ( .DIN1(_28321), .DIN2(_26341), .Q(_39039) );
  hi1s1 _39140_inst ( .DIN(_35685), .Q(_28321) );
  nnd2s1 _39141_inst ( .DIN1(_39040), .DIN2(_35688), .Q(_35685) );
  nor2s1 _39142_inst ( .DIN1(_28684), .DIN2(_35735), .Q(_39038) );
  nnd2s1 _39143_inst ( .DIN1(_39041), .DIN2(_35684), .Q(_35735) );
  and2s1 _39144_inst ( .DIN1(_28622), .DIN2(_39042), .Q(_35684) );
  nor2s1 _39145_inst ( .DIN1(_28599), .DIN2(_38017), .Q(_28622) );
  nor2s1 _39146_inst ( .DIN1(_28526), .DIN2(_28389), .Q(_39041) );
  nnd2s1 _39147_inst ( .DIN1(_39043), .DIN2(_39044), .Q(_28389) );
  nor2s1 _39148_inst ( .DIN1(_38018), .DIN2(_35433), .Q(_39044) );
  nor2s1 _39149_inst ( .DIN1(_28525), .DIN2(_28595), .Q(_39043) );
  nnd2s1 _39150_inst ( .DIN1(_39045), .DIN2(_39046), .Q(
        _______3____2________________3____________________) );
  nnd2s1 _39151_inst ( .DIN1(_39047), .DIN2(______[10]), .Q(_39046) );
  nor2s1 _39152_inst ( .DIN1(_53471), .DIN2(_27522), .Q(_39047) );
  nnd2s1 _39153_inst ( .DIN1(_39048), .DIN2(_27524), .Q(_39045) );
  nor2s1 _39154_inst ( .DIN1(_39049), .DIN2(_39050), .Q(_39048) );
  and2s1 _39155_inst ( .DIN1(______[3]), .DIN2(_28333), .Q(_39050) );
  nor2s1 _39156_inst ( .DIN1(_28333), .DIN2(_39051), .Q(_39049) );
  nnd2s1 _39157_inst ( .DIN1(_39052), .DIN2(______[24]), .Q(_39051) );
  nor2s1 _39158_inst ( .DIN1(_28336), .DIN2(_39053), .Q(_39052) );
  xor2s1 _39159_inst ( .DIN1(_26329), .DIN2(_39054), .Q(_39053) );
  nnd2s1 _39160_inst ( .DIN1(_53358), .DIN2(_53467), .Q(_39054) );
  hi1s1 _39161_inst ( .DIN(_39055), .Q(_28336) );
  nnd2s1 _39162_inst ( .DIN1(_39056), .DIN2(_28091), .Q(
        _______31____2________________31____________________) );
  nor2s1 _39163_inst ( .DIN1(_39057), .DIN2(_39058), .Q(_39056) );
  nor2s1 _39164_inst ( .DIN1(_28095), .DIN2(_39059), .Q(_39058) );
  nor2s1 _39165_inst ( .DIN1(_39060), .DIN2(_39061), .Q(_39059) );
  nor2s1 _39166_inst ( .DIN1(_27135), .DIN2(_39062), .Q(_39061) );
  nor2s1 _39167_inst ( .DIN1(_27160), .DIN2(_39063), .Q(_39062) );
  xor2s1 _39168_inst ( .DIN1(_53208), .DIN2(_53354), .Q(_39063) );
  hi1s1 _39169_inst ( .DIN(_27361), .Q(_27160) );
  nnd2s1 _39170_inst ( .DIN1(_39064), .DIN2(_39065), .Q(_27361) );
  nor2s1 _39171_inst ( .DIN1(_27342), .DIN2(_29801), .Q(_39065) );
  and2s1 _39172_inst ( .DIN1(_27473), .DIN2(_29345), .Q(_39064) );
  hi1s1 _39173_inst ( .DIN(_27158), .Q(_27135) );
  nor2s1 _39174_inst ( .DIN1(______[31]), .DIN2(_27158), .Q(_39060) );
  nnd2s1 _39175_inst ( .DIN1(_39066), .DIN2(_39067), .Q(_27158) );
  nor2s1 _39176_inst ( .DIN1(_39068), .DIN2(_27376), .Q(_39067) );
  nnd2s1 _39177_inst ( .DIN1(_27471), .DIN2(_29481), .Q(_27376) );
  and2s1 _39178_inst ( .DIN1(_27348), .DIN2(_39069), .Q(_27471) );
  nor2s1 _39179_inst ( .DIN1(_29483), .DIN2(_29656), .Q(_39066) );
  nnd2s1 _39180_inst ( .DIN1(_39070), .DIN2(_29345), .Q(_29656) );
  nor2s1 _39181_inst ( .DIN1(_29325), .DIN2(_29820), .Q(_29345) );
  nor2s1 _39182_inst ( .DIN1(_27296), .DIN2(_27343), .Q(_39070) );
  nnd2s1 _39183_inst ( .DIN1(_27497), .DIN2(_27466), .Q(_27343) );
  nnd2s1 _39184_inst ( .DIN1(_27359), .DIN2(_29351), .Q(_29483) );
  nor2s1 _39185_inst ( .DIN1(_28098), .DIN2(_39071), .Q(_39057) );
  nor2s1 _39186_inst ( .DIN1(_53383), .DIN2(_27365), .Q(_39071) );
  nnd2s1 _39187_inst ( .DIN1(_39072), .DIN2(_39073), .Q(
        _______30____2________________30____________________) );
  nnd2s1 _39188_inst ( .DIN1(_37341), .DIN2(_39074), .Q(_39073) );
  xor2s1 _39189_inst ( .DIN1(_26449), .DIN2(_39075), .Q(_39074) );
  nnd2s1 _39190_inst ( .DIN1(_53356), .DIN2(_53363), .Q(_39075) );
  and2s1 _39191_inst ( .DIN1(_27648), .DIN2(_36407), .Q(_37341) );
  nnd2s1 _39192_inst ( .DIN1(_39076), .DIN2(_39077), .Q(_36407) );
  nor2s1 _39193_inst ( .DIN1(_39078), .DIN2(_39079), .Q(_39077) );
  nnd2s1 _39194_inst ( .DIN1(_34672), .DIN2(_37551), .Q(_39079) );
  nor2s1 _39195_inst ( .DIN1(_36587), .DIN2(_35699), .Q(_39076) );
  nnd2s1 _39196_inst ( .DIN1(_35707), .DIN2(_37555), .Q(_35699) );
  nnd2s1 _39197_inst ( .DIN1(_27655), .DIN2(_39080), .Q(_39072) );
  nnd2s1 _39198_inst ( .DIN1(_39081), .DIN2(_39082), .Q(_39080) );
  nnd2s1 _39199_inst ( .DIN1(_39083), .DIN2(_27797), .Q(_39082) );
  xor2s1 _39200_inst ( .DIN1(_26338), .DIN2(_53364), .Q(_39083) );
  nnd2s1 _39201_inst ( .DIN1(______[30]), .DIN2(_27795), .Q(_39081) );
  hi1s1 _39202_inst ( .DIN(_27648), .Q(_27655) );
  nnd2s1 _39203_inst ( .DIN1(_39084), .DIN2(_39085), .Q(_27648) );
  nor2s1 _39204_inst ( .DIN1(_39086), .DIN2(_39087), .Q(_39085) );
  nnd2s1 _39205_inst ( .DIN1(_35784), .DIN2(_37533), .Q(_39087) );
  nnd2s1 _39206_inst ( .DIN1(_35707), .DIN2(_35781), .Q(_39086) );
  hi1s1 _39207_inst ( .DIN(_34676), .Q(_35707) );
  nor2s1 _39208_inst ( .DIN1(_36613), .DIN2(_39088), .Q(_39084) );
  or2s1 _39209_inst ( .DIN1(_27934), .DIN2(_34394), .Q(_39088) );
  nnd2s1 _39210_inst ( .DIN1(_39089), .DIN2(_39090), .Q(_34394) );
  nor2s1 _39211_inst ( .DIN1(_34399), .DIN2(_39091), .Q(_39090) );
  nor2s1 _39212_inst ( .DIN1(_33611), .DIN2(_34602), .Q(_39089) );
  nnd2s1 _39213_inst ( .DIN1(_35695), .DIN2(_35785), .Q(_34602) );
  nnd2s1 _39214_inst ( .DIN1(_34671), .DIN2(_39092), .Q(_27934) );
  nnd2s1 _39215_inst ( .DIN1(_39093), .DIN2(_34580), .Q(_36613) );
  and2s1 _39216_inst ( .DIN1(_39094), .DIN2(_39095), .Q(_34580) );
  nor2s1 _39217_inst ( .DIN1(_35706), .DIN2(_39096), .Q(_39094) );
  nor2s1 _39218_inst ( .DIN1(_39078), .DIN2(_34397), .Q(_39093) );
  nnd2s1 _39219_inst ( .DIN1(_33614), .DIN2(_39097), .Q(_34397) );
  nnd2s1 _39220_inst ( .DIN1(_39098), .DIN2(_36266), .Q(
        _______2____2________________2____________________) );
  nor2s1 _39221_inst ( .DIN1(_39099), .DIN2(_39100), .Q(_39098) );
  nor2s1 _39222_inst ( .DIN1(_28333), .DIN2(_39101), .Q(_39100) );
  nor2s1 _39223_inst ( .DIN1(_26772), .DIN2(_39102), .Q(_39101) );
  nnd2s1 _39224_inst ( .DIN1(_39103), .DIN2(_39055), .Q(_39102) );
  xor2s1 _39225_inst ( .DIN1(_53357), .DIN2(_53358), .Q(_39103) );
  nor2s1 _39226_inst ( .DIN1(______[2]), .DIN2(_28337), .Q(_39099) );
  nnd2s1 _39227_inst ( .DIN1(_39104), .DIN2(_39105), .Q(
        _______29____2________________29____________________) );
  nnd2s1 _39228_inst ( .DIN1(_39106), .DIN2(_39107), .Q(_39105) );
  xor2s1 _39229_inst ( .DIN1(_27880), .DIN2(_53359), .Q(_39107) );
  nnd2s1 _39230_inst ( .DIN1(_53485), .DIN2(_53360), .Q(_27880) );
  nor2s1 _39231_inst ( .DIN1(_27365), .DIN2(_27881), .Q(_39106) );
  nnd2s1 _39232_inst ( .DIN1(_28139), .DIN2(_28137), .Q(_27881) );
  nnd2s1 _39233_inst ( .DIN1(_39108), .DIN2(_34869), .Q(_28139) );
  and2s1 _39234_inst ( .DIN1(_39109), .DIN2(_39110), .Q(_34869) );
  nor2s1 _39235_inst ( .DIN1(_34415), .DIN2(_30925), .Q(_39109) );
  hi1s1 _39236_inst ( .DIN(_39111), .Q(_34415) );
  nor2s1 _39237_inst ( .DIN1(_30771), .DIN2(_30030), .Q(_39108) );
  nnd2s1 _39238_inst ( .DIN1(_39112), .DIN2(_27882), .Q(_39104) );
  hi1s1 _39239_inst ( .DIN(_28137), .Q(_27882) );
  nnd2s1 _39240_inst ( .DIN1(_39113), .DIN2(_28930), .Q(_28137) );
  hi1s1 _39241_inst ( .DIN(_30640), .Q(_28930) );
  nnd2s1 _39242_inst ( .DIN1(_39114), .DIN2(_32091), .Q(_30640) );
  nor2s1 _39243_inst ( .DIN1(_30029), .DIN2(_30432), .Q(_39113) );
  nnd2s1 _39244_inst ( .DIN1(_39115), .DIN2(_30407), .Q(_30432) );
  and2s1 _39245_inst ( .DIN1(_39116), .DIN2(_39111), .Q(_30407) );
  nor2s1 _39246_inst ( .DIN1(_30027), .DIN2(_30030), .Q(_39116) );
  hi1s1 _39247_inst ( .DIN(_30939), .Q(_30030) );
  hi1s1 _39248_inst ( .DIN(_39117), .Q(_30027) );
  nor2s1 _39249_inst ( .DIN1(_30771), .DIN2(_29940), .Q(_39115) );
  hi1s1 _39250_inst ( .DIN(_30940), .Q(_30029) );
  nor2s1 _39251_inst ( .DIN1(_39118), .DIN2(_39119), .Q(_39112) );
  nor2s1 _39252_inst ( .DIN1(_27786), .DIN2(_39120), .Q(_39119) );
  nor2s1 _39253_inst ( .DIN1(_27795), .DIN2(_39121), .Q(_39118) );
  nnd2s1 _39254_inst ( .DIN1(_39122), .DIN2(______[22]), .Q(_39121) );
  nor2s1 _39255_inst ( .DIN1(_53362), .DIN2(_27787), .Q(_39122) );
  hi1s1 _39256_inst ( .DIN(_27797), .Q(_27787) );
  nnd2s1 _39257_inst ( .DIN1(_39123), .DIN2(_36266), .Q(
        _______28____2________________28____________________) );
  nor2s1 _39258_inst ( .DIN1(_39124), .DIN2(_39125), .Q(_39123) );
  nor2s1 _39259_inst ( .DIN1(_26774), .DIN2(_27786), .Q(_39125) );
  nor2s1 _39260_inst ( .DIN1(_39126), .DIN2(_39127), .Q(_39124) );
  nnd2s1 _39261_inst ( .DIN1(______[8]), .DIN2(_34515), .Q(_39127) );
  nnd2s1 _39262_inst ( .DIN1(_39128), .DIN2(_36266), .Q(
        _______27____2________________27____________________) );
  nor2s1 _39263_inst ( .DIN1(_39129), .DIN2(_39130), .Q(_39128) );
  and2s1 _39264_inst ( .DIN1(______[27]), .DIN2(_27795), .Q(_39130) );
  nor2s1 _39265_inst ( .DIN1(_39126), .DIN2(_39131), .Q(_39129) );
  xor2s1 _39266_inst ( .DIN1(_38150), .DIN2(_38120), .Q(_39131) );
  xor2s1 _39267_inst ( .DIN1(_53363), .DIN2(_53362), .Q(_38120) );
  nor2s1 _39268_inst ( .DIN1(_27620), .DIN2(_53361), .Q(_38150) );
  nnd2s1 _39269_inst ( .DIN1(_27797), .DIN2(_27786), .Q(_39126) );
  hi1s1 _39270_inst ( .DIN(_27795), .Q(_27786) );
  nor2s1 _39271_inst ( .DIN1(_39132), .DIN2(_34530), .Q(_27795) );
  nnd2s1 _39272_inst ( .DIN1(_27630), .DIN2(_39133), .Q(_39132) );
  nnd2s1 _39273_inst ( .DIN1(_39134), .DIN2(_39133), .Q(_27797) );
  nor2s1 _39274_inst ( .DIN1(_34960), .DIN2(_39135), .Q(_39134) );
  nnd2s1 _39275_inst ( .DIN1(_39136), .DIN2(_39137), .Q(
        _______26____2________________26____________________) );
  nnd2s1 _39276_inst ( .DIN1(_39138), .DIN2(______[26]), .Q(_39137) );
  nor2s1 _39277_inst ( .DIN1(_39139), .DIN2(_39140), .Q(_39136) );
  nor2s1 _39278_inst ( .DIN1(_26781), .DIN2(_39141), .Q(_39140) );
  nnd2s1 _39279_inst ( .DIN1(_39142), .DIN2(_39143), .Q(_39141) );
  hi1s1 _39280_inst ( .DIN(_39144), .Q(_39142) );
  nor2s1 _39281_inst ( .DIN1(_39145), .DIN2(_26780), .Q(_39139) );
  nor2s1 _39282_inst ( .DIN1(_39146), .DIN2(_39147), .Q(_39145) );
  nor2s1 _39283_inst ( .DIN1(_39143), .DIN2(_39144), .Q(_39147) );
  nor2s1 _39284_inst ( .DIN1(_26209), .DIN2(_26331), .Q(_39143) );
  nor2s1 _39285_inst ( .DIN1(_27241), .DIN2(_39148), .Q(_39146) );
  nnd2s1 _39286_inst ( .DIN1(_39149), .DIN2(_39150), .Q(
        _______25____2________________25____________________) );
  nnd2s1 _39287_inst ( .DIN1(______[25]), .DIN2(_39138), .Q(_39150) );
  nor2s1 _39288_inst ( .DIN1(_39151), .DIN2(_39152), .Q(_39149) );
  nor2s1 _39289_inst ( .DIN1(_26526), .DIN2(_39148), .Q(_39152) );
  nor2s1 _39290_inst ( .DIN1(_39144), .DIN2(_39153), .Q(_39151) );
  nnd2s1 _39291_inst ( .DIN1(_53367), .DIN2(______[22]), .Q(_39153) );
  nor2s1 _39292_inst ( .DIN1(_27593), .DIN2(_39154), .Q(
        _______24____2________________24____________________) );
  nnd2s1 _39293_inst ( .DIN1(_39155), .DIN2(_39156), .Q(_39154) );
  nnd2s1 _39294_inst ( .DIN1(_39157), .DIN2(_39158), .Q(_39156) );
  nor2s1 _39295_inst ( .DIN1(_26526), .DIN2(_39159), .Q(_39157) );
  nnd2s1 _39296_inst ( .DIN1(______[12]), .DIN2(_39160), .Q(_39159) );
  nnd2s1 _39297_inst ( .DIN1(_39161), .DIN2(______[24]), .Q(_39155) );
  nnd2s1 _39298_inst ( .DIN1(_39162), .DIN2(_39163), .Q(
        _______23____2________________23____________________) );
  nor2s1 _39299_inst ( .DIN1(_39164), .DIN2(_39165), .Q(_39162) );
  nor2s1 _39300_inst ( .DIN1(_39166), .DIN2(_39167), .Q(_39165) );
  nnd2s1 _39301_inst ( .DIN1(_39168), .DIN2(_39169), .Q(_39167) );
  nnd2s1 _39302_inst ( .DIN1(_39170), .DIN2(_39160), .Q(_39169) );
  xor2s1 _39303_inst ( .DIN1(_39171), .DIN2(_38229), .Q(_39170) );
  xor2s1 _39304_inst ( .DIN1(_53365), .DIN2(_53367), .Q(_38229) );
  nor2s1 _39305_inst ( .DIN1(_26780), .DIN2(_26209), .Q(_39171) );
  nnd2s1 _39306_inst ( .DIN1(______[23]), .DIN2(_39161), .Q(_39168) );
  nor2s1 _39307_inst ( .DIN1(_36436), .DIN2(_39172), .Q(_39164) );
  nor2s1 _39308_inst ( .DIN1(_27066), .DIN2(_39173), .Q(_39172) );
  xnr2s1 _39309_inst ( .DIN1(_39174), .DIN2(_39175), .Q(_39173) );
  xor2s1 _39310_inst ( .DIN1(_26698), .DIN2(_26781), .Q(_39175) );
  nnd2s1 _39311_inst ( .DIN1(_39176), .DIN2(_39177), .Q(
        _______22____2________________22____________________) );
  nnd2s1 _39312_inst ( .DIN1(_39138), .DIN2(______[22]), .Q(_39177) );
  nor2s1 _39313_inst ( .DIN1(_39158), .DIN2(_39166), .Q(_39138) );
  nor2s1 _39314_inst ( .DIN1(_39178), .DIN2(_39179), .Q(_39176) );
  nor2s1 _39315_inst ( .DIN1(_36889), .DIN2(_39148), .Q(_39179) );
  or2s1 _39316_inst ( .DIN1(_36386), .DIN2(_36436), .Q(_39148) );
  xor2s1 _39317_inst ( .DIN1(_53371), .DIN2(_26333), .Q(_36889) );
  nor2s1 _39318_inst ( .DIN1(_39180), .DIN2(_39144), .Q(_39178) );
  nnd2s1 _39319_inst ( .DIN1(_36436), .DIN2(_39160), .Q(_39144) );
  xor2s1 _39320_inst ( .DIN1(_36332), .DIN2(_53370), .Q(_39180) );
  nnd2s1 _39321_inst ( .DIN1(_39181), .DIN2(_39163), .Q(
        _______21____2________________21____________________) );
  nor2s1 _39322_inst ( .DIN1(_39182), .DIN2(_39183), .Q(_39181) );
  nor2s1 _39323_inst ( .DIN1(_39166), .DIN2(_39184), .Q(_39183) );
  nnd2s1 _39324_inst ( .DIN1(_39185), .DIN2(_39186), .Q(_39184) );
  nnd2s1 _39325_inst ( .DIN1(______[21]), .DIN2(_39161), .Q(_39186) );
  hi1s1 _39326_inst ( .DIN(_39158), .Q(_39161) );
  nnd2s1 _39327_inst ( .DIN1(_39187), .DIN2(_34641), .Q(_39158) );
  nnd2s1 _39328_inst ( .DIN1(_39188), .DIN2(_53370), .Q(_39185) );
  nor2s1 _39329_inst ( .DIN1(_34637), .DIN2(_27241), .Q(_39188) );
  hi1s1 _39330_inst ( .DIN(_39160), .Q(_34637) );
  nnd2s1 _39331_inst ( .DIN1(_39189), .DIN2(_34866), .Q(_39160) );
  hi1s1 _39332_inst ( .DIN(_27707), .Q(_34866) );
  nnd2s1 _39333_inst ( .DIN1(_39190), .DIN2(_39191), .Q(_27707) );
  xor2s1 _39334_inst ( .DIN1(_2064), .DIN2(_39192), .Q(_39191) );
  nor2s1 _39335_inst ( .DIN1(_39031), .DIN2(_39193), .Q(_39192) );
  nor2s1 _39336_inst ( .DIN1(_27653), .DIN2(_39135), .Q(_39190) );
  hi1s1 _39337_inst ( .DIN(_34890), .Q(_39135) );
  nor2s1 _39338_inst ( .DIN1(_34765), .DIN2(_34891), .Q(_39189) );
  nor2s1 _39339_inst ( .DIN1(_36436), .DIN2(_39194), .Q(_39182) );
  nor2s1 _39340_inst ( .DIN1(_53370), .DIN2(_28684), .Q(_39194) );
  nnd2s1 _39341_inst ( .DIN1(_39195), .DIN2(_39034), .Q(
        _______20____2________________20____________________) );
  nor2s1 _39342_inst ( .DIN1(_39196), .DIN2(_39197), .Q(_39195) );
  nor2s1 _39343_inst ( .DIN1(_27448), .DIN2(_39198), .Q(_39197) );
  nor2s1 _39344_inst ( .DIN1(_39199), .DIN2(_39200), .Q(_39196) );
  nnd2s1 _39345_inst ( .DIN1(______[28]), .DIN2(_38379), .Q(_39200) );
  xor2s1 _39346_inst ( .DIN1(_36332), .DIN2(_26323), .Q(_38379) );
  hi1s1 _39347_inst ( .DIN(_53371), .Q(_36332) );
  nnd2s1 _39348_inst ( .DIN1(_39201), .DIN2(_39163), .Q(
        _______1____2________________1____________________) );
  nnd2s1 _39349_inst ( .DIN1(_36386), .DIN2(_39166), .Q(_39163) );
  nor2s1 _39350_inst ( .DIN1(_28420), .DIN2(_39202), .Q(_36386) );
  hi1s1 _39351_inst ( .DIN(_35720), .Q(_39202) );
  nor2s1 _39352_inst ( .DIN1(_39203), .DIN2(_39204), .Q(_39201) );
  nor2s1 _39353_inst ( .DIN1(_39166), .DIN2(_39205), .Q(_39204) );
  nor2s1 _39354_inst ( .DIN1(_39206), .DIN2(_39207), .Q(_39205) );
  nor2s1 _39355_inst ( .DIN1(_28333), .DIN2(_39208), .Q(_39207) );
  nor2s1 _39356_inst ( .DIN1(_27393), .DIN2(_39209), .Q(_39208) );
  nnd2s1 _39357_inst ( .DIN1(_39210), .DIN2(_39055), .Q(_39209) );
  xor2s1 _39358_inst ( .DIN1(_52851), .DIN2(_53369), .Q(_39210) );
  nor2s1 _39359_inst ( .DIN1(______[1]), .DIN2(_28337), .Q(_39206) );
  nor2s1 _39360_inst ( .DIN1(_36436), .DIN2(_39211), .Q(_39203) );
  nor2s1 _39361_inst ( .DIN1(_27774), .DIN2(_39212), .Q(_39211) );
  nnd2s1 _39362_inst ( .DIN1(_39213), .DIN2(_39214), .Q(_39212) );
  nnd2s1 _39363_inst ( .DIN1(_39215), .DIN2(_26331), .Q(_39214) );
  nnd2s1 _39364_inst ( .DIN1(_26781), .DIN2(_26698), .Q(_39215) );
  nnd2s1 _39365_inst ( .DIN1(_39174), .DIN2(_26698), .Q(_39213) );
  nor2s1 _39366_inst ( .DIN1(_26780), .DIN2(_26331), .Q(_39174) );
  nnd2s1 _39367_inst ( .DIN1(_39216), .DIN2(_39217), .Q(
        _______19____2________________19____________________) );
  nnd2s1 _39368_inst ( .DIN1(_39218), .DIN2(______[12]), .Q(_39217) );
  nor2s1 _39369_inst ( .DIN1(_27522), .DIN2(_39219), .Q(_39218) );
  xor2s1 _39370_inst ( .DIN1(_26341), .DIN2(_53471), .Q(_39219) );
  nnd2s1 _39371_inst ( .DIN1(_39220), .DIN2(_27524), .Q(_39216) );
  nor2s1 _39372_inst ( .DIN1(_39221), .DIN2(_39222), .Q(_39220) );
  nor2s1 _39373_inst ( .DIN1(_39187), .DIN2(_39223), .Q(_39222) );
  nor2s1 _39374_inst ( .DIN1(_27448), .DIN2(_39224), .Q(_39223) );
  nnd2s1 _39375_inst ( .DIN1(_39225), .DIN2(_39226), .Q(_39224) );
  xor2s1 _39376_inst ( .DIN1(_26343), .DIN2(_39227), .Q(_39225) );
  nnd2s1 _39377_inst ( .DIN1(_53370), .DIN2(_53371), .Q(_39227) );
  hi1s1 _39378_inst ( .DIN(_39198), .Q(_39187) );
  nor2s1 _39379_inst ( .DIN1(______[19]), .DIN2(_39198), .Q(_39221) );
  nnd2s1 _39380_inst ( .DIN1(_39228), .DIN2(_36266), .Q(
        _______18____2________________18____________________) );
  hi1s1 _39381_inst ( .DIN(_39229), .Q(_36266) );
  nor2s1 _39382_inst ( .DIN1(_39230), .DIN2(_39231), .Q(_39228) );
  nor2s1 _39383_inst ( .DIN1(_27291), .DIN2(_39198), .Q(_39231) );
  nor2s1 _39384_inst ( .DIN1(_39199), .DIN2(_39232), .Q(_39230) );
  nnd2s1 _39385_inst ( .DIN1(_26858), .DIN2(_39233), .Q(_39232) );
  xor2s1 _39386_inst ( .DIN1(_53373), .DIN2(_39234), .Q(_39233) );
  nor2s1 _39387_inst ( .DIN1(_38996), .DIN2(_39235), .Q(
        _______17____2________________17____________________) );
  nnd2s1 _39388_inst ( .DIN1(_39236), .DIN2(_39237), .Q(_39235) );
  or2s1 _39389_inst ( .DIN1(______[17]), .DIN2(_39198), .Q(_39237) );
  nnd2s1 _39390_inst ( .DIN1(_39238), .DIN2(_39198), .Q(_39236) );
  nnd2s1 _39391_inst ( .DIN1(_39239), .DIN2(_53374), .Q(_39238) );
  nor2s1 _39392_inst ( .DIN1(_39240), .DIN2(_27291), .Q(_39239) );
  hi1s1 _39393_inst ( .DIN(_39034), .Q(_38996) );
  nnd2s1 _39394_inst ( .DIN1(_39241), .DIN2(_39034), .Q(
        _______16____2________________16____________________) );
  nor2s1 _39395_inst ( .DIN1(_28420), .DIN2(_35302), .Q(_39034) );
  nor2s1 _39396_inst ( .DIN1(_39242), .DIN2(_39243), .Q(_39241) );
  nor2s1 _39397_inst ( .DIN1(_26771), .DIN2(_39198), .Q(_39243) );
  nor2s1 _39398_inst ( .DIN1(_39199), .DIN2(_39244), .Q(_39242) );
  nnd2s1 _39399_inst ( .DIN1(_53372), .DIN2(______[20]), .Q(_39244) );
  nnd2s1 _39400_inst ( .DIN1(_39245), .DIN2(_36436), .Q(
        _______15____2________________15____________________) );
  nor2s1 _39401_inst ( .DIN1(_39246), .DIN2(_39247), .Q(_39245) );
  nor2s1 _39402_inst ( .DIN1(_39198), .DIN2(_39248), .Q(_39247) );
  nor2s1 _39403_inst ( .DIN1(_39249), .DIN2(_39199), .Q(_39246) );
  nnd2s1 _39404_inst ( .DIN1(_39226), .DIN2(_39198), .Q(_39199) );
  nnd2s1 _39405_inst ( .DIN1(_39250), .DIN2(_39251), .Q(_39198) );
  nor2s1 _39406_inst ( .DIN1(_27653), .DIN2(_39193), .Q(_39251) );
  nor2s1 _39407_inst ( .DIN1(_34891), .DIN2(_34530), .Q(_39250) );
  nnd2s1 _39408_inst ( .DIN1(_39252), .DIN2(_34959), .Q(_34530) );
  nor2s1 _39409_inst ( .DIN1(_34960), .DIN2(_34894), .Q(_39252) );
  hi1s1 _39410_inst ( .DIN(_39240), .Q(_39226) );
  nor2s1 _39411_inst ( .DIN1(_27810), .DIN2(_39193), .Q(_39240) );
  nnd2s1 _39412_inst ( .DIN1(_39020), .DIN2(_39253), .Q(_27810) );
  nor2s1 _39413_inst ( .DIN1(_27653), .DIN2(_34891), .Q(_39253) );
  nor2s1 _39414_inst ( .DIN1(_34766), .DIN2(_39028), .Q(_39020) );
  hi1s1 _39415_inst ( .DIN(_34959), .Q(_39028) );
  xor2s1 _39416_inst ( .DIN1(_31842), .DIN2(_39254), .Q(_34959) );
  nor2s1 _39417_inst ( .DIN1(_39255), .DIN2(_39256), .Q(_39254) );
  nnd2s1 _39418_inst ( .DIN1(_34890), .DIN2(_39257), .Q(_39256) );
  xor2s1 _39419_inst ( .DIN1(_39258), .DIN2(_38452), .Q(_39249) );
  nor2s1 _39420_inst ( .DIN1(_39234), .DIN2(_39259), .Q(_38452) );
  nor2s1 _39421_inst ( .DIN1(_27731), .DIN2(_53374), .Q(_39259) );
  hi1s1 _39422_inst ( .DIN(_53375), .Q(_27731) );
  nor2s1 _39423_inst ( .DIN1(_26322), .DIN2(_53375), .Q(_39234) );
  nnd2s1 _39424_inst ( .DIN1(_53374), .DIN2(_53373), .Q(_39258) );
  nnd2s1 _39425_inst ( .DIN1(_39260), .DIN2(_39261), .Q(
        _______14____2________________14____________________) );
  nnd2s1 _39426_inst ( .DIN1(_39262), .DIN2(_39263), .Q(_39261) );
  nor2s1 _39427_inst ( .DIN1(_39264), .DIN2(_39265), .Q(_39262) );
  nor2s1 _39428_inst ( .DIN1(_39001), .DIN2(_39266), .Q(_39265) );
  nor2s1 _39429_inst ( .DIN1(_27365), .DIN2(_39267), .Q(_39266) );
  xor2s1 _39430_inst ( .DIN1(_53376), .DIN2(_53377), .Q(_39267) );
  nor2s1 _39431_inst ( .DIN1(______[14]), .DIN2(_39003), .Q(_39264) );
  nnd2s1 _39432_inst ( .DIN1(_36436), .DIN2(_39268), .Q(
        _______13____2________________13____________________) );
  nnd2s1 _39433_inst ( .DIN1(_39269), .DIN2(_39263), .Q(_39268) );
  nor2s1 _39434_inst ( .DIN1(_39270), .DIN2(_39271), .Q(_39269) );
  nor2s1 _39435_inst ( .DIN1(_53377), .DIN2(_39001), .Q(_39271) );
  nor2s1 _39436_inst ( .DIN1(______[13]), .DIN2(_39003), .Q(_39270) );
  nnd2s1 _39437_inst ( .DIN1(_39272), .DIN2(_28091), .Q(
        _______12____2________________12____________________) );
  nor2s1 _39438_inst ( .DIN1(_39273), .DIN2(_39274), .Q(_39272) );
  nor2s1 _39439_inst ( .DIN1(_28095), .DIN2(_39275), .Q(_39274) );
  nnd2s1 _39440_inst ( .DIN1(_39276), .DIN2(_39263), .Q(_39275) );
  nor2s1 _39441_inst ( .DIN1(_39277), .DIN2(_39278), .Q(_39276) );
  nor2s1 _39442_inst ( .DIN1(_39001), .DIN2(_39279), .Q(_39278) );
  nor2s1 _39443_inst ( .DIN1(_27291), .DIN2(_38699), .Q(_39279) );
  xor2s1 _39444_inst ( .DIN1(_53379), .DIN2(_53376), .Q(_38699) );
  nor2s1 _39445_inst ( .DIN1(______[12]), .DIN2(_39003), .Q(_39277) );
  nor2s1 _39446_inst ( .DIN1(_28098), .DIN2(_39280), .Q(_39273) );
  xor2s1 _39447_inst ( .DIN1(_26237), .DIN2(_53384), .Q(_39280) );
  nnd2s1 _39448_inst ( .DIN1(_39281), .DIN2(_28310), .Q(
        _______11____2________________11____________________) );
  hi1s1 _39449_inst ( .DIN(_28384), .Q(_28310) );
  nor2s1 _39450_inst ( .DIN1(_28420), .DIN2(_28322), .Q(_28384) );
  nnd2s1 _39451_inst ( .DIN1(_39282), .DIN2(_35300), .Q(_28420) );
  nor2s1 _39452_inst ( .DIN1(_39283), .DIN2(_39284), .Q(_39281) );
  nor2s1 _39453_inst ( .DIN1(_28313), .DIN2(_39285), .Q(_39284) );
  nnd2s1 _39454_inst ( .DIN1(_39286), .DIN2(_39287), .Q(_39285) );
  nnd2s1 _39455_inst ( .DIN1(______[11]), .DIN2(_39001), .Q(_39287) );
  nnd2s1 _39456_inst ( .DIN1(_39288), .DIN2(______[10]), .Q(_39286) );
  nor2s1 _39457_inst ( .DIN1(_39289), .DIN2(_39290), .Q(_39288) );
  xor2s1 _39458_inst ( .DIN1(_26319), .DIN2(_39291), .Q(_39290) );
  nor2s1 _39459_inst ( .DIN1(_53376), .DIN2(_26318), .Q(_39291) );
  nor2s1 _39460_inst ( .DIN1(_28322), .DIN2(_39292), .Q(_39283) );
  nor2s1 _39461_inst ( .DIN1(_27448), .DIN2(_39293), .Q(_39292) );
  xor2s1 _39462_inst ( .DIN1(_53378), .DIN2(_28324), .Q(_39293) );
  nor2s1 _39463_inst ( .DIN1(_26332), .DIN2(_53367), .Q(_28324) );
  hi1s1 _39464_inst ( .DIN(_28313), .Q(_28322) );
  nnd2s1 _39465_inst ( .DIN1(_39260), .DIN2(_35720), .Q(_28313) );
  hi1s1 _39466_inst ( .DIN(_27593), .Q(_39260) );
  nor2s1 _39467_inst ( .DIN1(_39294), .DIN2(_39166), .Q(
        _______10____2________________10____________________) );
  nor2s1 _39468_inst ( .DIN1(_38997), .DIN2(_39295), .Q(_39294) );
  nnd2s1 _39469_inst ( .DIN1(_39296), .DIN2(_39297), .Q(_39295) );
  nnd2s1 _39470_inst ( .DIN1(_39001), .DIN2(_27614), .Q(_39297) );
  hi1s1 _39471_inst ( .DIN(_39003), .Q(_39001) );
  nnd2s1 _39472_inst ( .DIN1(_39298), .DIN2(_39003), .Q(_39296) );
  xor2s1 _39473_inst ( .DIN1(_38589), .DIN2(_53380), .Q(_39298) );
  hi1s1 _39474_inst ( .DIN(_53381), .Q(_38589) );
  hi1s1 _39475_inst ( .DIN(_39263), .Q(_38997) );
  nnd2s1 _39476_inst ( .DIN1(_39289), .DIN2(_39003), .Q(_39263) );
  nnd2s1 _39477_inst ( .DIN1(_39299), .DIN2(_34764), .Q(_39003) );
  nor2s1 _39478_inst ( .DIN1(_34894), .DIN2(_39193), .Q(_34764) );
  nor2s1 _39479_inst ( .DIN1(_27843), .DIN2(_39300), .Q(_39299) );
  nnd2s1 _39480_inst ( .DIN1(_39301), .DIN2(_39027), .Q(_27843) );
  hi1s1 _39481_inst ( .DIN(_39300), .Q(_39289) );
  nnd2s1 _39482_inst ( .DIN1(_39302), .DIN2(_34641), .Q(_39300) );
  nor2s1 _39483_inst ( .DIN1(_34766), .DIN2(_39031), .Q(_34641) );
  nor2s1 _39484_inst ( .DIN1(_34891), .DIN2(_39255), .Q(_39302) );
  nor2s1 _39485_inst ( .DIN1(_39229), .DIN2(_39303), .Q(
        _______0____2________________0____________________) );
  nnd2s1 _39486_inst ( .DIN1(_39304), .DIN2(_39305), .Q(_39303) );
  nnd2s1 _39487_inst ( .DIN1(_39306), .DIN2(_28337), .Q(_39305) );
  nor2s1 _39488_inst ( .DIN1(_26774), .DIN2(_39307), .Q(_39306) );
  nnd2s1 _39489_inst ( .DIN1(_52851), .DIN2(_39055), .Q(_39307) );
  nnd2s1 _39490_inst ( .DIN1(_39308), .DIN2(_33571), .Q(_39055) );
  hi1s1 _39491_inst ( .DIN(_32920), .Q(_33571) );
  nnd2s1 _39492_inst ( .DIN1(_39309), .DIN2(_39310), .Q(_32920) );
  xnr2s1 _39493_inst ( .DIN1(_28527), .DIN2(_29994), .Q(_39310) );
  nnd2s1 _39494_inst ( .DIN1(_39311), .DIN2(_39312), .Q(_28527) );
  nor2s1 _39495_inst ( .DIN1(_28597), .DIN2(_28603), .Q(_39309) );
  nnd2s1 _39496_inst ( .DIN1(_39313), .DIN2(_39314), .Q(_28603) );
  nor2s1 _39497_inst ( .DIN1(_28599), .DIN2(_38018), .Q(_39308) );
  nnd2s1 _39498_inst ( .DIN1(_28333), .DIN2(______[0]), .Q(_39304) );
  hi1s1 _39499_inst ( .DIN(_28337), .Q(_28333) );
  nnd2s1 _39500_inst ( .DIN1(_39315), .DIN2(_35432), .Q(_28337) );
  and2s1 _39501_inst ( .DIN1(_39316), .DIN2(_28442), .Q(_35432) );
  hi1s1 _39502_inst ( .DIN(_28598), .Q(_28442) );
  nnd2s1 _39503_inst ( .DIN1(_39040), .DIN2(_35533), .Q(_28598) );
  nor2s1 _39504_inst ( .DIN1(_38017), .DIN2(_39317), .Q(_39316) );
  nor2s1 _39505_inst ( .DIN1(_28599), .DIN2(_28596), .Q(_39315) );
  nnd2s1 _39506_inst ( .DIN1(_39318), .DIN2(_35723), .Q(_39229) );
  nor2s1 _39507_inst ( .DIN1(_39319), .DIN2(_35302), .Q(_39318) );
  hi1s1 _39508_inst ( .DIN(_35721), .Q(_35302) );
  nnd2s1 _39509_inst ( .DIN1(_36436), .DIN2(_39320), .Q(
        ____3____________9_____) );
  nnd2s1 _39510_inst ( .DIN1(_39321), .DIN2(_39322), .Q(_39320) );
  nor2s1 _39511_inst ( .DIN1(_39323), .DIN2(_39324), .Q(_39322) );
  nnd2s1 _39512_inst ( .DIN1(_39325), .DIN2(_39326), .Q(_39324) );
  hi1s1 _39513_inst ( .DIN(_39327), .Q(_39326) );
  nor2s1 _39514_inst ( .DIN1(_39328), .DIN2(_39329), .Q(_39325) );
  nor2s1 _39515_inst ( .DIN1(_39330), .DIN2(_39331), .Q(_39329) );
  nor2s1 _39516_inst ( .DIN1(_39332), .DIN2(_39333), .Q(_39328) );
  nor2s1 _39517_inst ( .DIN1(_39334), .DIN2(_39335), .Q(_39332) );
  nnd2s1 _39518_inst ( .DIN1(_39336), .DIN2(_39337), .Q(_39323) );
  nor2s1 _39519_inst ( .DIN1(_39338), .DIN2(_39339), .Q(_39337) );
  nor2s1 _39520_inst ( .DIN1(_39340), .DIN2(_39341), .Q(_39336) );
  nor2s1 _39521_inst ( .DIN1(_39342), .DIN2(_39343), .Q(_39341) );
  nor2s1 _39522_inst ( .DIN1(_39344), .DIN2(_39345), .Q(_39342) );
  hi1s1 _39523_inst ( .DIN(_39346), .Q(_39340) );
  nor2s1 _39524_inst ( .DIN1(_39347), .DIN2(_39348), .Q(_39321) );
  nnd2s1 _39525_inst ( .DIN1(_39349), .DIN2(_39350), .Q(_39348) );
  nor2s1 _39526_inst ( .DIN1(_39351), .DIN2(_39352), .Q(_39349) );
  nnd2s1 _39527_inst ( .DIN1(_39353), .DIN2(_39354), .Q(_39347) );
  nor2s1 _39528_inst ( .DIN1(_39355), .DIN2(_39356), .Q(_39354) );
  nor2s1 _39529_inst ( .DIN1(_39357), .DIN2(_39358), .Q(_39353) );
  hi1s1 _39530_inst ( .DIN(_39166), .Q(_36436) );
  nnd2s1 _39531_inst ( .DIN1(_39359), .DIN2(_39360), .Q(
        ____3____________8_____) );
  nnd2s1 _39532_inst ( .DIN1(_27397), .DIN2(_39361), .Q(_39360) );
  nnd2s1 _39533_inst ( .DIN1(_39362), .DIN2(_39363), .Q(_39361) );
  nor2s1 _39534_inst ( .DIN1(_39364), .DIN2(_39365), .Q(_39363) );
  nnd2s1 _39535_inst ( .DIN1(_39366), .DIN2(_39367), .Q(_39365) );
  or2s1 _39536_inst ( .DIN1(_39368), .DIN2(_39369), .Q(_39367) );
  nor2s1 _39537_inst ( .DIN1(_39370), .DIN2(_39371), .Q(_39366) );
  nor2s1 _39538_inst ( .DIN1(_39372), .DIN2(_39373), .Q(_39371) );
  nor2s1 _39539_inst ( .DIN1(_39343), .DIN2(_39374), .Q(_39370) );
  nnd2s1 _39540_inst ( .DIN1(_39375), .DIN2(_39376), .Q(_39364) );
  nor2s1 _39541_inst ( .DIN1(_39377), .DIN2(_39378), .Q(_39376) );
  nor2s1 _39542_inst ( .DIN1(_39379), .DIN2(_39380), .Q(_39378) );
  nor2s1 _39543_inst ( .DIN1(_39381), .DIN2(_39382), .Q(_39379) );
  nor2s1 _39544_inst ( .DIN1(_39383), .DIN2(_39384), .Q(_39377) );
  and2s1 _39545_inst ( .DIN1(_39385), .DIN2(_39386), .Q(_39384) );
  nor2s1 _39546_inst ( .DIN1(_39387), .DIN2(_39388), .Q(_39375) );
  nor2s1 _39547_inst ( .DIN1(_39389), .DIN2(_39390), .Q(_39387) );
  and2s1 _39548_inst ( .DIN1(_39391), .DIN2(_39392), .Q(_39389) );
  nor2s1 _39549_inst ( .DIN1(_39393), .DIN2(_39394), .Q(_39362) );
  nnd2s1 _39550_inst ( .DIN1(_39395), .DIN2(_39396), .Q(_39394) );
  xor2s1 _39551_inst ( .DIN1(_39397), .DIN2(_27840), .Q(_39396) );
  or2s1 _39552_inst ( .DIN1(_39398), .DIN2(_39356), .Q(_39397) );
  nnd2s1 _39553_inst ( .DIN1(_39399), .DIN2(_39400), .Q(_39356) );
  nor2s1 _39554_inst ( .DIN1(_39401), .DIN2(_39402), .Q(_39400) );
  nnd2s1 _39555_inst ( .DIN1(_39403), .DIN2(_39404), .Q(_39402) );
  nor2s1 _39556_inst ( .DIN1(_39405), .DIN2(_39406), .Q(_39399) );
  nor2s1 _39557_inst ( .DIN1(_39383), .DIN2(_39407), .Q(_39405) );
  nor2s1 _39558_inst ( .DIN1(_39408), .DIN2(_39409), .Q(_39395) );
  nnd2s1 _39559_inst ( .DIN1(_39410), .DIN2(_39411), .Q(_39393) );
  nor2s1 _39560_inst ( .DIN1(_39412), .DIN2(_39413), .Q(_39410) );
  hi1s1 _39561_inst ( .DIN(_27392), .Q(_27397) );
  nnd2s1 _39562_inst ( .DIN1(_39414), .DIN2(_27392), .Q(_39359) );
  nnd2s1 _39563_inst ( .DIN1(_27183), .DIN2(_38460), .Q(_27392) );
  hi1s1 _39564_inst ( .DIN(_28084), .Q(_27183) );
  nnd2s1 _39565_inst ( .DIN1(_38332), .DIN2(_34827), .Q(_28084) );
  and2s1 _39566_inst ( .DIN1(_39415), .DIN2(_34828), .Q(_38332) );
  nor2s1 _39567_inst ( .DIN1(_38537), .DIN2(_27903), .Q(_39415) );
  hi1s1 _39568_inst ( .DIN(_32015), .Q(_27903) );
  nor2s1 _39569_inst ( .DIN1(_36552), .DIN2(_26493), .Q(_39414) );
  hi1s1 _39570_inst ( .DIN(_27396), .Q(_36552) );
  nnd2s1 _39571_inst ( .DIN1(_39416), .DIN2(_31103), .Q(_27396) );
  nor2s1 _39572_inst ( .DIN1(_38537), .DIN2(_35617), .Q(_39416) );
  hi1s1 _39573_inst ( .DIN(_39417), .Q(_38537) );
  nnd2s1 _39574_inst ( .DIN1(_39418), .DIN2(_39419), .Q(
        ____3____________7_____) );
  nnd2s1 _39575_inst ( .DIN1(_29849), .DIN2(_39420), .Q(_39419) );
  nnd2s1 _39576_inst ( .DIN1(_39421), .DIN2(_39422), .Q(_39420) );
  nor2s1 _39577_inst ( .DIN1(_39423), .DIN2(_39424), .Q(_39422) );
  nnd2s1 _39578_inst ( .DIN1(_39425), .DIN2(_39426), .Q(_39424) );
  hi1s1 _39579_inst ( .DIN(_39427), .Q(_39426) );
  nor2s1 _39580_inst ( .DIN1(_39428), .DIN2(_39429), .Q(_39425) );
  nor2s1 _39581_inst ( .DIN1(_39430), .DIN2(_39431), .Q(_39428) );
  nnd2s1 _39582_inst ( .DIN1(_39432), .DIN2(_39433), .Q(_39423) );
  nor2s1 _39583_inst ( .DIN1(_39434), .DIN2(_39435), .Q(_39433) );
  nor2s1 _39584_inst ( .DIN1(_39436), .DIN2(_39437), .Q(_39435) );
  nor2s1 _39585_inst ( .DIN1(_39438), .DIN2(_39343), .Q(_39434) );
  and2s1 _39586_inst ( .DIN1(_39373), .DIN2(_39374), .Q(_39438) );
  nor2s1 _39587_inst ( .DIN1(_39439), .DIN2(_39440), .Q(_39432) );
  nor2s1 _39588_inst ( .DIN1(_39441), .DIN2(_39368), .Q(_39440) );
  nor2s1 _39589_inst ( .DIN1(_39380), .DIN2(_39442), .Q(_39439) );
  nor2s1 _39590_inst ( .DIN1(_39443), .DIN2(_39444), .Q(_39421) );
  nnd2s1 _39591_inst ( .DIN1(_39445), .DIN2(_39446), .Q(_39444) );
  hi1s1 _39592_inst ( .DIN(_39447), .Q(_39446) );
  nor2s1 _39593_inst ( .DIN1(_39448), .DIN2(_39449), .Q(_39445) );
  nnd2s1 _39594_inst ( .DIN1(_39450), .DIN2(_39451), .Q(_39443) );
  nor2s1 _39595_inst ( .DIN1(_39452), .DIN2(_39453), .Q(_39450) );
  nnd2s1 _39596_inst ( .DIN1(_39454), .DIN2(_29828), .Q(_39418) );
  hi1s1 _39597_inst ( .DIN(_29849), .Q(_29828) );
  nor2s1 _39598_inst ( .DIN1(_39455), .DIN2(_39456), .Q(_29849) );
  or2s1 _39599_inst ( .DIN1(_37129), .DIN2(_39457), .Q(_39455) );
  nor2s1 _39600_inst ( .DIN1(_28381), .DIN2(_39458), .Q(_39454) );
  xor2s1 _39601_inst ( .DIN1(_26357), .DIN2(_28835), .Q(_39458) );
  nnd2s1 _39602_inst ( .DIN1(_53410), .DIN2(_53437), .Q(_28835) );
  hi1s1 _39603_inst ( .DIN(_37419), .Q(_28381) );
  nnd2s1 _39604_inst ( .DIN1(_39459), .DIN2(_39460), .Q(_37419) );
  nor2s1 _39605_inst ( .DIN1(_27161), .DIN2(_37129), .Q(_39460) );
  nor2s1 _39606_inst ( .DIN1(_39461), .DIN2(_39457), .Q(_39459) );
  hi1s1 _39607_inst ( .DIN(_39462), .Q(_39457) );
  nnd2s1 _39608_inst ( .DIN1(_39463), .DIN2(_28091), .Q(
        ____3____________6_____) );
  or2s1 _39609_inst ( .DIN1(_28857), .DIN2(_28098), .Q(_28091) );
  nor2s1 _39610_inst ( .DIN1(_39464), .DIN2(_39465), .Q(_39463) );
  nor2s1 _39611_inst ( .DIN1(_28095), .DIN2(_39466), .Q(_39465) );
  nnd2s1 _39612_inst ( .DIN1(_39467), .DIN2(_39468), .Q(_39466) );
  nor2s1 _39613_inst ( .DIN1(_39469), .DIN2(_39470), .Q(_39468) );
  nnd2s1 _39614_inst ( .DIN1(_39471), .DIN2(_39472), .Q(_39470) );
  nor2s1 _39615_inst ( .DIN1(_39473), .DIN2(_39474), .Q(_39472) );
  nor2s1 _39616_inst ( .DIN1(_39372), .DIN2(_39475), .Q(_39474) );
  nor2s1 _39617_inst ( .DIN1(_39476), .DIN2(_39477), .Q(_39473) );
  nor2s1 _39618_inst ( .DIN1(_39478), .DIN2(_39479), .Q(_39471) );
  nnd2s1 _39619_inst ( .DIN1(_39480), .DIN2(_39481), .Q(_39469) );
  and2s1 _39620_inst ( .DIN1(_39482), .DIN2(_39403), .Q(_39481) );
  nor2s1 _39621_inst ( .DIN1(_39483), .DIN2(_39484), .Q(_39480) );
  nor2s1 _39622_inst ( .DIN1(_39485), .DIN2(_39486), .Q(_39484) );
  nor2s1 _39623_inst ( .DIN1(_39487), .DIN2(_39488), .Q(_39467) );
  nnd2s1 _39624_inst ( .DIN1(_39489), .DIN2(_39490), .Q(_39488) );
  nor2s1 _39625_inst ( .DIN1(_39491), .DIN2(_39492), .Q(_39490) );
  nor2s1 _39626_inst ( .DIN1(_39493), .DIN2(_39494), .Q(_39489) );
  nnd2s1 _39627_inst ( .DIN1(_39495), .DIN2(_39496), .Q(_39487) );
  nor2s1 _39628_inst ( .DIN1(_39497), .DIN2(_39498), .Q(_39496) );
  nor2s1 _39629_inst ( .DIN1(_39413), .DIN2(_39499), .Q(_39495) );
  nnd2s1 _39630_inst ( .DIN1(_39500), .DIN2(_39501), .Q(_39413) );
  nor2s1 _39631_inst ( .DIN1(_39502), .DIN2(_39503), .Q(_39501) );
  nnd2s1 _39632_inst ( .DIN1(_39504), .DIN2(_39505), .Q(_39503) );
  nor2s1 _39633_inst ( .DIN1(_39506), .DIN2(_39507), .Q(_39500) );
  nor2s1 _39634_inst ( .DIN1(_28098), .DIN2(_39508), .Q(_39464) );
  nor2s1 _39635_inst ( .DIN1(_39509), .DIN2(_27614), .Q(_39508) );
  xor2s1 _39636_inst ( .DIN1(_39510), .DIN2(_39511), .Q(_39509) );
  xor2s1 _39637_inst ( .DIN1(_53377), .DIN2(_53383), .Q(_39511) );
  nnd2s1 _39638_inst ( .DIN1(_26849), .DIN2(_26211), .Q(_39510) );
  hi1s1 _39639_inst ( .DIN(_28095), .Q(_28098) );
  nnd2s1 _39640_inst ( .DIN1(_39512), .DIN2(_39513), .Q(_28095) );
  nor2s1 _39641_inst ( .DIN1(_39514), .DIN2(_39515), .Q(_39513) );
  nnd2s1 _39642_inst ( .DIN1(_39516), .DIN2(_39517), .Q(_39515) );
  nor2s1 _39643_inst ( .DIN1(_39518), .DIN2(_27745), .Q(_39512) );
  nnd2s1 _39644_inst ( .DIN1(_39519), .DIN2(_39520), .Q(_27745) );
  nor2s1 _39645_inst ( .DIN1(_39521), .DIN2(_39522), .Q(_39520) );
  nor2s1 _39646_inst ( .DIN1(_39523), .DIN2(_27747), .Q(_39519) );
  nnd2s1 _39647_inst ( .DIN1(_39524), .DIN2(_30112), .Q(
        ____3____________5_____) );
  nor2s1 _39648_inst ( .DIN1(_39525), .DIN2(_39526), .Q(_39524) );
  nor2s1 _39649_inst ( .DIN1(_28032), .DIN2(_39527), .Q(_39526) );
  nnd2s1 _39650_inst ( .DIN1(_39528), .DIN2(_39529), .Q(_39527) );
  nor2s1 _39651_inst ( .DIN1(_39530), .DIN2(_39531), .Q(_39529) );
  nnd2s1 _39652_inst ( .DIN1(_39532), .DIN2(_39533), .Q(_39531) );
  nor2s1 _39653_inst ( .DIN1(_39534), .DIN2(_39535), .Q(_39532) );
  xor2s1 _39654_inst ( .DIN1(_39536), .DIN2(_35821), .Q(_39535) );
  nnd2s1 _39655_inst ( .DIN1(_39537), .DIN2(_39538), .Q(_39536) );
  nnd2s1 _39656_inst ( .DIN1(_39539), .DIN2(_39540), .Q(_39538) );
  nor2s1 _39657_inst ( .DIN1(_39541), .DIN2(_39542), .Q(_39540) );
  nnd2s1 _39658_inst ( .DIN1(_39543), .DIN2(_39544), .Q(_39542) );
  nor2s1 _39659_inst ( .DIN1(_39545), .DIN2(_39546), .Q(_39544) );
  nor2s1 _39660_inst ( .DIN1(_39547), .DIN2(_39548), .Q(_39543) );
  nor2s1 _39661_inst ( .DIN1(_39549), .DIN2(_39550), .Q(_39548) );
  nor2s1 _39662_inst ( .DIN1(_39551), .DIN2(_39381), .Q(_39550) );
  nnd2s1 _39663_inst ( .DIN1(_39552), .DIN2(_39553), .Q(_39541) );
  nor2s1 _39664_inst ( .DIN1(_39554), .DIN2(_39555), .Q(_39553) );
  and2s1 _39665_inst ( .DIN1(_39556), .DIN2(_39557), .Q(_39552) );
  nor2s1 _39666_inst ( .DIN1(_39558), .DIN2(_39559), .Q(_39539) );
  nnd2s1 _39667_inst ( .DIN1(_39560), .DIN2(_39561), .Q(_39559) );
  nor2s1 _39668_inst ( .DIN1(_39562), .DIN2(_39563), .Q(_39561) );
  nnd2s1 _39669_inst ( .DIN1(_39564), .DIN2(_39565), .Q(_39563) );
  nnd2s1 _39670_inst ( .DIN1(_39566), .DIN2(_39567), .Q(_39565) );
  nnd2s1 _39671_inst ( .DIN1(_39568), .DIN2(_39569), .Q(_39564) );
  nnd2s1 _39672_inst ( .DIN1(_39570), .DIN2(_39571), .Q(_39569) );
  nnd2s1 _39673_inst ( .DIN1(_39572), .DIN2(_39573), .Q(_39571) );
  nor2s1 _39674_inst ( .DIN1(_39574), .DIN2(_39575), .Q(_39570) );
  nnd2s1 _39675_inst ( .DIN1(_39576), .DIN2(_39577), .Q(_39562) );
  nnd2s1 _39676_inst ( .DIN1(_39578), .DIN2(_39579), .Q(_39577) );
  nnd2s1 _39677_inst ( .DIN1(_39580), .DIN2(_39581), .Q(_39576) );
  nnd2s1 _39678_inst ( .DIN1(_39582), .DIN2(_39583), .Q(_39581) );
  hi1s1 _39679_inst ( .DIN(_39584), .Q(_39583) );
  nor2s1 _39680_inst ( .DIN1(_39585), .DIN2(_39586), .Q(_39582) );
  nor2s1 _39681_inst ( .DIN1(_39587), .DIN2(_39588), .Q(_39586) );
  nor2s1 _39682_inst ( .DIN1(_39589), .DIN2(_39590), .Q(_39560) );
  nnd2s1 _39683_inst ( .DIN1(_39591), .DIN2(_39592), .Q(_39590) );
  nnd2s1 _39684_inst ( .DIN1(_39593), .DIN2(_39594), .Q(_39592) );
  nnd2s1 _39685_inst ( .DIN1(_39486), .DIN2(_39407), .Q(_39593) );
  nnd2s1 _39686_inst ( .DIN1(_39595), .DIN2(_39596), .Q(_39591) );
  nnd2s1 _39687_inst ( .DIN1(_39597), .DIN2(_39598), .Q(_39596) );
  nnd2s1 _39688_inst ( .DIN1(_39599), .DIN2(_39600), .Q(_39589) );
  nnd2s1 _39689_inst ( .DIN1(_39335), .DIN2(_39601), .Q(_39600) );
  hi1s1 _39690_inst ( .DIN(_39602), .Q(_39335) );
  nnd2s1 _39691_inst ( .DIN1(_39603), .DIN2(_39604), .Q(_39599) );
  nnd2s1 _39692_inst ( .DIN1(_39605), .DIN2(_39606), .Q(_39558) );
  nor2s1 _39693_inst ( .DIN1(_37195), .DIN2(_39607), .Q(_39606) );
  nnd2s1 _39694_inst ( .DIN1(_39608), .DIN2(_39609), .Q(_39607) );
  nnd2s1 _39695_inst ( .DIN1(_39610), .DIN2(_39611), .Q(_39609) );
  nnd2s1 _39696_inst ( .DIN1(_39612), .DIN2(_39613), .Q(_39608) );
  nnd2s1 _39697_inst ( .DIN1(_39392), .DIN2(_39614), .Q(_39613) );
  nor2s1 _39698_inst ( .DIN1(_39615), .DIN2(_39616), .Q(_39605) );
  nnd2s1 _39699_inst ( .DIN1(_39617), .DIN2(_39618), .Q(_39616) );
  nnd2s1 _39700_inst ( .DIN1(_39619), .DIN2(_39620), .Q(_39618) );
  nnd2s1 _39701_inst ( .DIN1(_39621), .DIN2(_39475), .Q(_39620) );
  nor2s1 _39702_inst ( .DIN1(_39622), .DIN2(_39623), .Q(_39621) );
  nnd2s1 _39703_inst ( .DIN1(_39624), .DIN2(_39625), .Q(_39617) );
  nnd2s1 _39704_inst ( .DIN1(_39626), .DIN2(_39627), .Q(_39624) );
  nnd2s1 _39705_inst ( .DIN1(_39628), .DIN2(_39629), .Q(_39615) );
  or2s1 _39706_inst ( .DIN1(_39331), .DIN2(_39630), .Q(_39629) );
  nnd2s1 _39707_inst ( .DIN1(_39630), .DIN2(_39631), .Q(_39628) );
  nnd2s1 _39708_inst ( .DIN1(_39632), .DIN2(_39633), .Q(_39631) );
  nor2s1 _39709_inst ( .DIN1(_39634), .DIN2(_39635), .Q(_39632) );
  hi1s1 _39710_inst ( .DIN(_39636), .Q(_39634) );
  and2s1 _39711_inst ( .DIN1(_39637), .DIN2(_39638), .Q(_39534) );
  nnd2s1 _39712_inst ( .DIN1(_39639), .DIN2(_39640), .Q(_39530) );
  and2s1 _39713_inst ( .DIN1(_39641), .DIN2(_39404), .Q(_39639) );
  nor2s1 _39714_inst ( .DIN1(_39642), .DIN2(_39643), .Q(_39528) );
  nnd2s1 _39715_inst ( .DIN1(_39644), .DIN2(_39645), .Q(_39643) );
  hi1s1 _39716_inst ( .DIN(_39646), .Q(_39645) );
  nnd2s1 _39717_inst ( .DIN1(_39647), .DIN2(_39648), .Q(_39642) );
  hi1s1 _39718_inst ( .DIN(_39649), .Q(_39648) );
  nor2s1 _39719_inst ( .DIN1(_39352), .DIN2(_39499), .Q(_39647) );
  nor2s1 _39720_inst ( .DIN1(_28037), .DIN2(_39650), .Q(_39525) );
  nor2s1 _39721_inst ( .DIN1(_39651), .DIN2(_27082), .Q(_39650) );
  xor2s1 _39722_inst ( .DIN1(_39652), .DIN2(_39653), .Q(_39651) );
  xor2s1 _39723_inst ( .DIN1(_53085), .DIN2(_53385), .Q(_39653) );
  nnd2s1 _39724_inst ( .DIN1(_53085), .DIN2(_53076), .Q(_39652) );
  nnd2s1 _39725_inst ( .DIN1(_39654), .DIN2(_39655), .Q(
        ____3____________4_____) );
  nnd2s1 _39726_inst ( .DIN1(_39656), .DIN2(_36302), .Q(_39655) );
  xor2s1 _39727_inst ( .DIN1(_26591), .DIN2(_28545), .Q(_39656) );
  nor2s1 _39728_inst ( .DIN1(_53387), .DIN2(_53388), .Q(_28545) );
  nnd2s1 _39729_inst ( .DIN1(_28542), .DIN2(_39657), .Q(_39654) );
  nnd2s1 _39730_inst ( .DIN1(_39658), .DIN2(_39659), .Q(_39657) );
  nor2s1 _39731_inst ( .DIN1(_39660), .DIN2(_39661), .Q(_39659) );
  nnd2s1 _39732_inst ( .DIN1(_39662), .DIN2(_39663), .Q(_39661) );
  nor2s1 _39733_inst ( .DIN1(_39664), .DIN2(_39665), .Q(_39663) );
  nor2s1 _39734_inst ( .DIN1(_39436), .DIN2(_39386), .Q(_39665) );
  nor2s1 _39735_inst ( .DIN1(_39485), .DIN2(_39666), .Q(_39664) );
  nor2s1 _39736_inst ( .DIN1(_39478), .DIN2(_39667), .Q(_39662) );
  nnd2s1 _39737_inst ( .DIN1(_39668), .DIN2(_39669), .Q(_39660) );
  nor2s1 _39738_inst ( .DIN1(_39670), .DIN2(_39671), .Q(_39669) );
  nnd2s1 _39739_inst ( .DIN1(_39672), .DIN2(_39673), .Q(_39671) );
  nor2s1 _39740_inst ( .DIN1(_39674), .DIN2(_39675), .Q(_39668) );
  nor2s1 _39741_inst ( .DIN1(_39383), .DIN2(_39676), .Q(_39675) );
  nor2s1 _39742_inst ( .DIN1(_39677), .DIN2(_39678), .Q(_39676) );
  nor2s1 _39743_inst ( .DIN1(_39679), .DIN2(_39372), .Q(_39674) );
  nor2s1 _39744_inst ( .DIN1(_39554), .DIN2(_39680), .Q(_39679) );
  nor2s1 _39745_inst ( .DIN1(_39681), .DIN2(_39682), .Q(_39658) );
  nnd2s1 _39746_inst ( .DIN1(_39683), .DIN2(_39684), .Q(_39682) );
  nor2s1 _39747_inst ( .DIN1(_39685), .DIN2(_39492), .Q(_39684) );
  nnd2s1 _39748_inst ( .DIN1(_39686), .DIN2(_39687), .Q(_39492) );
  nor2s1 _39749_inst ( .DIN1(_39688), .DIN2(_39689), .Q(_39687) );
  nnd2s1 _39750_inst ( .DIN1(_39690), .DIN2(_39691), .Q(_39689) );
  nnd2s1 _39751_inst ( .DIN1(_39692), .DIN2(_39693), .Q(_39688) );
  nnd2s1 _39752_inst ( .DIN1(_39694), .DIN2(_39695), .Q(_39693) );
  nor2s1 _39753_inst ( .DIN1(_39696), .DIN2(_39697), .Q(_39692) );
  nor2s1 _39754_inst ( .DIN1(_39383), .DIN2(_39698), .Q(_39697) );
  nor2s1 _39755_inst ( .DIN1(_39699), .DIN2(_39700), .Q(_39698) );
  nnd2s1 _39756_inst ( .DIN1(_39368), .DIN2(_39556), .Q(_39700) );
  nor2s1 _39757_inst ( .DIN1(_39701), .DIN2(_39702), .Q(_39686) );
  or2s1 _39758_inst ( .DIN1(_39703), .DIN2(_39412), .Q(_39702) );
  or2s1 _39759_inst ( .DIN1(_39704), .DIN2(_39705), .Q(_39412) );
  and2s1 _39760_inst ( .DIN1(_39547), .DIN2(_39706), .Q(_39705) );
  nnd2s1 _39761_inst ( .DIN1(_39707), .DIN2(_39708), .Q(_39701) );
  nnd2s1 _39762_inst ( .DIN1(_39709), .DIN2(_39710), .Q(_39708) );
  or2s1 _39763_inst ( .DIN1(_39374), .DIN2(_39372), .Q(_39707) );
  nor2s1 _39764_inst ( .DIN1(_39646), .DIN2(_39711), .Q(_39683) );
  nnd2s1 _39765_inst ( .DIN1(_39712), .DIN2(_39713), .Q(_39646) );
  nnd2s1 _39766_inst ( .DIN1(_39714), .DIN2(_39715), .Q(_39681) );
  nor2s1 _39767_inst ( .DIN1(_39716), .DIN2(_39408), .Q(_39715) );
  nnd2s1 _39768_inst ( .DIN1(_39717), .DIN2(_39718), .Q(_39408) );
  nor2s1 _39769_inst ( .DIN1(_39719), .DIN2(_39720), .Q(_39718) );
  nor2s1 _39770_inst ( .DIN1(_39441), .DIN2(_39721), .Q(_39720) );
  nor2s1 _39771_inst ( .DIN1(_39722), .DIN2(_39723), .Q(_39717) );
  nor2s1 _39772_inst ( .DIN1(_39724), .DIN2(_39448), .Q(_39714) );
  nnd2s1 _39773_inst ( .DIN1(_39725), .DIN2(_39726), .Q(_39448) );
  nor2s1 _39774_inst ( .DIN1(_39483), .DIN2(_39727), .Q(_39726) );
  nnd2s1 _39775_inst ( .DIN1(_39728), .DIN2(_39729), .Q(_39727) );
  hi1s1 _39776_inst ( .DIN(_39730), .Q(_39483) );
  nor2s1 _39777_inst ( .DIN1(_39731), .DIN2(_39732), .Q(_39725) );
  nnd2s1 _39778_inst ( .DIN1(_39733), .DIN2(_39734), .Q(_39732) );
  or2s1 _39779_inst ( .DIN1(_39407), .DIN2(_39735), .Q(_39734) );
  nnd2s1 _39780_inst ( .DIN1(_39334), .DIN2(_39736), .Q(_39733) );
  nor2s1 _39781_inst ( .DIN1(_39737), .DIN2(_39391), .Q(_39731) );
  hi1s1 _39782_inst ( .DIN(_28533), .Q(_28542) );
  nnd2s1 _39783_inst ( .DIN1(_39738), .DIN2(_39739), .Q(_28533) );
  nor2s1 _39784_inst ( .DIN1(_39740), .DIN2(_39741), .Q(_39739) );
  nnd2s1 _39785_inst ( .DIN1(_39742), .DIN2(_34485), .Q(_39741) );
  nor2s1 _39786_inst ( .DIN1(_37414), .DIN2(_33338), .Q(_39738) );
  hi1s1 _39787_inst ( .DIN(_30175), .Q(_33338) );
  nor2s1 _39788_inst ( .DIN1(_39743), .DIN2(_38885), .Q(_30175) );
  nnd2s1 _39789_inst ( .DIN1(_39744), .DIN2(_37413), .Q(_38885) );
  nor2s1 _39790_inst ( .DIN1(_38714), .DIN2(_34489), .Q(_39744) );
  nnd2s1 _39791_inst ( .DIN1(_30174), .DIN2(_39745), .Q(_39743) );
  nor2s1 _39792_inst ( .DIN1(_39746), .DIN2(_27500), .Q(
        ____3____________3_____) );
  nor2s1 _39793_inst ( .DIN1(_39747), .DIN2(_39748), .Q(_39746) );
  nnd2s1 _39794_inst ( .DIN1(_39749), .DIN2(_39750), .Q(_39748) );
  nor2s1 _39795_inst ( .DIN1(_39751), .DIN2(_39752), .Q(_39750) );
  nnd2s1 _39796_inst ( .DIN1(_39753), .DIN2(_39754), .Q(_39752) );
  hi1s1 _39797_inst ( .DIN(_39507), .Q(_39754) );
  nnd2s1 _39798_inst ( .DIN1(_39755), .DIN2(_39756), .Q(_39507) );
  nnd2s1 _39799_inst ( .DIN1(_39585), .DIN2(_39638), .Q(_39756) );
  nnd2s1 _39800_inst ( .DIN1(_39757), .DIN2(_39758), .Q(_39755) );
  or2s1 _39801_inst ( .DIN1(_39723), .DIN2(_39357), .Q(_39751) );
  nnd2s1 _39802_inst ( .DIN1(_39759), .DIN2(_39760), .Q(_39357) );
  nor2s1 _39803_inst ( .DIN1(_39761), .DIN2(_39762), .Q(_39760) );
  nnd2s1 _39804_inst ( .DIN1(_39763), .DIN2(_39764), .Q(_39762) );
  nnd2s1 _39805_inst ( .DIN1(_39545), .DIN2(_39710), .Q(_39764) );
  nnd2s1 _39806_inst ( .DIN1(_39554), .DIN2(_39765), .Q(_39763) );
  nnd2s1 _39807_inst ( .DIN1(_39766), .DIN2(_39767), .Q(_39761) );
  nnd2s1 _39808_inst ( .DIN1(_39768), .DIN2(_39769), .Q(_39767) );
  nnd2s1 _39809_inst ( .DIN1(_39770), .DIN2(_39666), .Q(_39769) );
  or2s1 _39810_inst ( .DIN1(_39771), .DIN2(_39441), .Q(_39766) );
  nor2s1 _39811_inst ( .DIN1(_39772), .DIN2(_39773), .Q(_39759) );
  nnd2s1 _39812_inst ( .DIN1(_39774), .DIN2(_39775), .Q(_39773) );
  hi1s1 _39813_inst ( .DIN(_39667), .Q(_39775) );
  nnd2s1 _39814_inst ( .DIN1(_39776), .DIN2(_39777), .Q(_39667) );
  nnd2s1 _39815_inst ( .DIN1(_39778), .DIN2(_39779), .Q(_39777) );
  nor2s1 _39816_inst ( .DIN1(_39780), .DIN2(_39372), .Q(_39778) );
  nnd2s1 _39817_inst ( .DIN1(_39533), .DIN2(_39781), .Q(_39772) );
  hi1s1 _39818_inst ( .DIN(_39506), .Q(_39781) );
  nnd2s1 _39819_inst ( .DIN1(_39782), .DIN2(_39728), .Q(_39506) );
  and2s1 _39820_inst ( .DIN1(_39783), .DIN2(_39784), .Q(_39533) );
  nor2s1 _39821_inst ( .DIN1(_39785), .DIN2(_39786), .Q(_39783) );
  nor2s1 _39822_inst ( .DIN1(_39390), .DIN2(_39787), .Q(_39786) );
  nnd2s1 _39823_inst ( .DIN1(_39640), .DIN2(_39788), .Q(_39723) );
  nnd2s1 _39824_inst ( .DIN1(_39789), .DIN2(_26838), .Q(_39788) );
  nnd2s1 _39825_inst ( .DIN1(_39790), .DIN2(_39791), .Q(_39640) );
  nnd2s1 _39826_inst ( .DIN1(_39792), .DIN2(_39793), .Q(_39791) );
  nnd2s1 _39827_inst ( .DIN1(_39794), .DIN2(_39795), .Q(_39792) );
  nor2s1 _39828_inst ( .DIN1(_39796), .DIN2(_39797), .Q(_39749) );
  nnd2s1 _39829_inst ( .DIN1(_39798), .DIN2(_39799), .Q(_39797) );
  hi1s1 _39830_inst ( .DIN(_39409), .Q(_39799) );
  nnd2s1 _39831_inst ( .DIN1(_39800), .DIN2(_39801), .Q(_39409) );
  nor2s1 _39832_inst ( .DIN1(_39802), .DIN2(_39803), .Q(_39801) );
  nor2s1 _39833_inst ( .DIN1(_39383), .DIN2(_39804), .Q(_39802) );
  nor2s1 _39834_inst ( .DIN1(_39805), .DIN2(_39427), .Q(_39800) );
  nnd2s1 _39835_inst ( .DIN1(_39806), .DIN2(_39690), .Q(_39427) );
  nnd2s1 _39836_inst ( .DIN1(_39807), .DIN2(_39768), .Q(_39690) );
  nor2s1 _39837_inst ( .DIN1(_39808), .DIN2(_39809), .Q(_39806) );
  nor2s1 _39838_inst ( .DIN1(_39810), .DIN2(_39811), .Q(_39809) );
  nnd2s1 _39839_inst ( .DIN1(_39812), .DIN2(_39813), .Q(_39811) );
  nnd2s1 _39840_inst ( .DIN1(_39814), .DIN2(_39815), .Q(_39810) );
  hi1s1 _39841_inst ( .DIN(_39816), .Q(_39808) );
  nnd2s1 _39842_inst ( .DIN1(_39817), .DIN2(_39818), .Q(_39747) );
  nor2s1 _39843_inst ( .DIN1(_39819), .DIN2(_39820), .Q(_39818) );
  nnd2s1 _39844_inst ( .DIN1(_39821), .DIN2(_39822), .Q(_39820) );
  nnd2s1 _39845_inst ( .DIN1(_39823), .DIN2(_39824), .Q(_39822) );
  nor2s1 _39846_inst ( .DIN1(_39430), .DIN2(_39825), .Q(_39823) );
  nnd2s1 _39847_inst ( .DIN1(_39826), .DIN2(_26838), .Q(_39821) );
  nnd2s1 _39848_inst ( .DIN1(_39827), .DIN2(_39828), .Q(_39826) );
  nor2s1 _39849_inst ( .DIN1(_39678), .DIN2(_39547), .Q(_39828) );
  and2s1 _39850_inst ( .DIN1(_39829), .DIN2(_39475), .Q(_39827) );
  nnd2s1 _39851_inst ( .DIN1(_39830), .DIN2(_39831), .Q(_39819) );
  nor2s1 _39852_inst ( .DIN1(_39832), .DIN2(_39833), .Q(_39817) );
  nnd2s1 _39853_inst ( .DIN1(_39691), .DIN2(_39834), .Q(_39833) );
  nnd2s1 _39854_inst ( .DIN1(_39677), .DIN2(_39768), .Q(_39834) );
  nnd2s1 _39855_inst ( .DIN1(_39578), .DIN2(_39638), .Q(_39691) );
  hi1s1 _39856_inst ( .DIN(_39835), .Q(_39578) );
  nnd2s1 _39857_inst ( .DIN1(_39836), .DIN2(_39837), .Q(
        ____3____________2_____) );
  nnd2s1 _39858_inst ( .DIN1(_39838), .DIN2(_39839), .Q(_39837) );
  xor2s1 _39859_inst ( .DIN1(_39840), .DIN2(_53389), .Q(_39839) );
  nor2s1 _39860_inst ( .DIN1(_28684), .DIN2(_39841), .Q(_39838) );
  nnd2s1 _39861_inst ( .DIN1(_39842), .DIN2(_39843), .Q(_39836) );
  nnd2s1 _39862_inst ( .DIN1(_39844), .DIN2(_39845), .Q(_39843) );
  nor2s1 _39863_inst ( .DIN1(_39846), .DIN2(_39847), .Q(_39845) );
  nnd2s1 _39864_inst ( .DIN1(_39848), .DIN2(_39411), .Q(_39847) );
  and2s1 _39865_inst ( .DIN1(_39849), .DIN2(_39850), .Q(_39411) );
  nor2s1 _39866_inst ( .DIN1(_39851), .DIN2(_39852), .Q(_39850) );
  nnd2s1 _39867_inst ( .DIN1(_39853), .DIN2(_39830), .Q(_39852) );
  nnd2s1 _39868_inst ( .DIN1(_39346), .DIN2(_39854), .Q(_39851) );
  nor2s1 _39869_inst ( .DIN1(_39855), .DIN2(_39856), .Q(_39849) );
  or2s1 _39870_inst ( .DIN1(_39857), .DIN2(_39498), .Q(_39856) );
  or2s1 _39871_inst ( .DIN1(_39452), .DIN2(_39858), .Q(_39498) );
  nor2s1 _39872_inst ( .DIN1(_39859), .DIN2(_39369), .Q(_39858) );
  nnd2s1 _39873_inst ( .DIN1(_39860), .DIN2(_39861), .Q(_39452) );
  nnd2s1 _39874_inst ( .DIN1(_39862), .DIN2(_39863), .Q(_39861) );
  nor2s1 _39875_inst ( .DIN1(_39380), .DIN2(_39864), .Q(_39863) );
  nor2s1 _39876_inst ( .DIN1(_39865), .DIN2(_39866), .Q(_39862) );
  nnd2s1 _39877_inst ( .DIN1(_39867), .DIN2(_39868), .Q(_39855) );
  or2s1 _39878_inst ( .DIN1(_39869), .DIN2(_39383), .Q(_39868) );
  nnd2s1 _39879_inst ( .DIN1(_39706), .DIN2(_39574), .Q(_39867) );
  nor2s1 _39880_inst ( .DIN1(_39358), .DIN2(_39805), .Q(_39848) );
  nnd2s1 _39881_inst ( .DIN1(_39870), .DIN2(_39871), .Q(_39805) );
  nnd2s1 _39882_inst ( .DIN1(_39623), .DIN2(_39765), .Q(_39871) );
  hi1s1 _39883_inst ( .DIN(_39872), .Q(_39623) );
  nnd2s1 _39884_inst ( .DIN1(_39873), .DIN2(_39874), .Q(_39358) );
  nor2s1 _39885_inst ( .DIN1(_39875), .DIN2(_39876), .Q(_39874) );
  nnd2s1 _39886_inst ( .DIN1(_39877), .DIN2(_39816), .Q(_39876) );
  nor2s1 _39887_inst ( .DIN1(_39878), .DIN2(_39380), .Q(_39875) );
  nor2s1 _39888_inst ( .DIN1(_39551), .DIN2(_39694), .Q(_39878) );
  nor2s1 _39889_inst ( .DIN1(_39879), .DIN2(_39497), .Q(_39873) );
  nnd2s1 _39890_inst ( .DIN1(_39880), .DIN2(_39881), .Q(_39497) );
  nnd2s1 _39891_inst ( .DIN1(_39765), .DIN2(_39882), .Q(_39881) );
  nnd2s1 _39892_inst ( .DIN1(_39883), .DIN2(_39557), .Q(_39882) );
  nnd2s1 _39893_inst ( .DIN1(_39884), .DIN2(_39789), .Q(_39880) );
  hi1s1 _39894_inst ( .DIN(_39614), .Q(_39789) );
  nor2s1 _39895_inst ( .DIN1(_39333), .DIN2(_39793), .Q(_39879) );
  nnd2s1 _39896_inst ( .DIN1(_39885), .DIN2(_39886), .Q(_39846) );
  nnd2s1 _39897_inst ( .DIN1(_39887), .DIN2(_26838), .Q(_39886) );
  nnd2s1 _39898_inst ( .DIN1(_39888), .DIN2(_39602), .Q(_39887) );
  nor2s1 _39899_inst ( .DIN1(_39381), .DIN2(_39610), .Q(_39888) );
  hi1s1 _39900_inst ( .DIN(_39391), .Q(_39610) );
  hi1s1 _39901_inst ( .DIN(_39437), .Q(_39381) );
  nor2s1 _39902_inst ( .DIN1(_39889), .DIN2(_39890), .Q(_39885) );
  nor2s1 _39903_inst ( .DIN1(_39891), .DIN2(_39892), .Q(_39844) );
  nnd2s1 _39904_inst ( .DIN1(_39893), .DIN2(_39894), .Q(_39892) );
  xor2s1 _39905_inst ( .DIN1(_37577), .DIN2(_39895), .Q(_39894) );
  nor2s1 _39906_inst ( .DIN1(_39896), .DIN2(_39897), .Q(_39895) );
  nor2s1 _39907_inst ( .DIN1(_39898), .DIN2(_39330), .Q(_39897) );
  nor2s1 _39908_inst ( .DIN1(_39635), .DIN2(_39899), .Q(_39898) );
  nor2s1 _39909_inst ( .DIN1(_39369), .DIN2(_39385), .Q(_39896) );
  nor2s1 _39910_inst ( .DIN1(_39796), .DIN2(_39900), .Q(_39893) );
  nnd2s1 _39911_inst ( .DIN1(_39901), .DIN2(_39902), .Q(_39796) );
  nor2s1 _39912_inst ( .DIN1(_39903), .DIN2(_39904), .Q(_39902) );
  nnd2s1 _39913_inst ( .DIN1(_39905), .DIN2(_39906), .Q(_39904) );
  nnd2s1 _39914_inst ( .DIN1(_39907), .DIN2(_39641), .Q(_39903) );
  nor2s1 _39915_inst ( .DIN1(_39908), .DIN2(_39909), .Q(_39901) );
  or2s1 _39916_inst ( .DIN1(_39910), .DIN2(_39449), .Q(_39909) );
  nnd2s1 _39917_inst ( .DIN1(_39911), .DIN2(_39912), .Q(_39449) );
  nnd2s1 _39918_inst ( .DIN1(_39566), .DIN2(_39706), .Q(_39912) );
  nor2s1 _39919_inst ( .DIN1(_39502), .DIN2(_39913), .Q(_39911) );
  nor2s1 _39920_inst ( .DIN1(_39914), .DIN2(_39915), .Q(_39913) );
  nnd2s1 _39921_inst ( .DIN1(_39814), .DIN2(_39916), .Q(_39915) );
  xnr2s1 _39922_inst ( .DIN1(_29049), .DIN2(_39917), .Q(_39908) );
  nnd2s1 _39923_inst ( .DIN1(_39918), .DIN2(_39919), .Q(_39917) );
  nor2s1 _39924_inst ( .DIN1(_39920), .DIN2(_39921), .Q(_39919) );
  nnd2s1 _39925_inst ( .DIN1(_39730), .DIN2(_39922), .Q(_39921) );
  nnd2s1 _39926_inst ( .DIN1(_39482), .DIN2(_39923), .Q(_39920) );
  nor2s1 _39927_inst ( .DIN1(_39711), .DIN2(_39924), .Q(_39918) );
  nnd2s1 _39928_inst ( .DIN1(_39925), .DIN2(_39926), .Q(_39924) );
  nnd2s1 _39929_inst ( .DIN1(_39927), .DIN2(_39928), .Q(_39926) );
  nnd2s1 _39930_inst ( .DIN1(_39929), .DIN2(_39930), .Q(_39711) );
  nnd2s1 _39931_inst ( .DIN1(_39931), .DIN2(_39932), .Q(_39930) );
  and2s1 _39932_inst ( .DIN1(_39933), .DIN2(_39934), .Q(_39931) );
  nnd2s1 _39933_inst ( .DIN1(_39935), .DIN2(_39936), .Q(_39891) );
  hi1s1 _39934_inst ( .DIN(_39493), .Q(_39936) );
  nnd2s1 _39935_inst ( .DIN1(_39937), .DIN2(_39938), .Q(_39493) );
  nnd2s1 _39936_inst ( .DIN1(_39939), .DIN2(_39940), .Q(_39938) );
  hi1s1 _39937_inst ( .DIN(_39941), .Q(_39940) );
  nnd2s1 _39938_inst ( .DIN1(_39575), .DIN2(_39710), .Q(_39937) );
  nor2s1 _39939_inst ( .DIN1(_39499), .DIN2(_39942), .Q(_39935) );
  nnd2s1 _39940_inst ( .DIN1(_39943), .DIN2(_39944), .Q(
        ____3____________1_____) );
  nor2s1 _39941_inst ( .DIN1(_39945), .DIN2(_39946), .Q(_39943) );
  nor2s1 _39942_inst ( .DIN1(_39947), .DIN2(_39948), .Q(_39946) );
  nnd2s1 _39943_inst ( .DIN1(_39949), .DIN2(_39950), .Q(_39948) );
  nor2s1 _39944_inst ( .DIN1(_39951), .DIN2(_39952), .Q(_39950) );
  nnd2s1 _39945_inst ( .DIN1(_39953), .DIN2(_39954), .Q(_39952) );
  nnd2s1 _39946_inst ( .DIN1(_39955), .DIN2(_39932), .Q(_39954) );
  nor2s1 _39947_inst ( .DIN1(_39956), .DIN2(_39957), .Q(_39955) );
  nor2s1 _39948_inst ( .DIN1(_39719), .DIN2(_39502), .Q(_39953) );
  and2s1 _39949_inst ( .DIN1(_39958), .DIN2(_39824), .Q(_39502) );
  nor2s1 _39950_inst ( .DIN1(_34359), .DIN2(_39485), .Q(_39958) );
  hi1s1 _39951_inst ( .DIN(_39922), .Q(_39719) );
  nnd2s1 _39952_inst ( .DIN1(_39959), .DIN2(_39960), .Q(_39922) );
  nor2s1 _39953_inst ( .DIN1(_39441), .DIN2(_39961), .Q(_39959) );
  nnd2s1 _39954_inst ( .DIN1(_39962), .DIN2(_39963), .Q(_39951) );
  nor2s1 _39955_inst ( .DIN1(_39339), .DIN2(_39964), .Q(_39963) );
  hi1s1 _39956_inst ( .DIN(_39965), .Q(_39964) );
  and2s1 _39957_inst ( .DIN1(_39966), .DIN2(_26838), .Q(_39339) );
  nnd2s1 _39958_inst ( .DIN1(_39967), .DIN2(_39968), .Q(_39966) );
  nor2s1 _39959_inst ( .DIN1(_39677), .DIN2(_39699), .Q(_39968) );
  nor2s1 _39960_inst ( .DIN1(_39969), .DIN2(_39970), .Q(_39967) );
  xor2s1 _39961_inst ( .DIN1(_31885), .DIN2(_39971), .Q(_39970) );
  nor2s1 _39962_inst ( .DIN1(_39972), .DIN2(_39973), .Q(_39971) );
  nnd2s1 _39963_inst ( .DIN1(_39633), .DIN2(_39556), .Q(_39973) );
  nnd2s1 _39964_inst ( .DIN1(_39391), .DIN2(_39859), .Q(_39972) );
  hi1s1 _39965_inst ( .DIN(_31307), .Q(_31885) );
  and2s1 _39966_inst ( .DIN1(_39860), .DIN2(_39877), .Q(_39962) );
  nnd2s1 _39967_inst ( .DIN1(_39974), .DIN2(_39975), .Q(_39860) );
  nor2s1 _39968_inst ( .DIN1(_39976), .DIN2(_39441), .Q(_39974) );
  nor2s1 _39969_inst ( .DIN1(_39977), .DIN2(_39978), .Q(_39949) );
  nnd2s1 _39970_inst ( .DIN1(_39979), .DIN2(_39980), .Q(_39978) );
  hi1s1 _39971_inst ( .DIN(_39981), .Q(_39980) );
  nor2s1 _39972_inst ( .DIN1(_39982), .DIN2(_39703), .Q(_39979) );
  nnd2s1 _39973_inst ( .DIN1(_39983), .DIN2(_39984), .Q(_39703) );
  nnd2s1 _39974_inst ( .DIN1(_39555), .DIN2(_39758), .Q(_39984) );
  nnd2s1 _39975_inst ( .DIN1(_39344), .DIN2(_26838), .Q(_39983) );
  nnd2s1 _39976_inst ( .DIN1(_39985), .DIN2(_39986), .Q(_39977) );
  nor2s1 _39977_inst ( .DIN1(_39987), .DIN2(_39988), .Q(_39985) );
  nor2s1 _39978_inst ( .DIN1(_39383), .DIN2(_39989), .Q(_39988) );
  nor2s1 _39979_inst ( .DIN1(_39380), .DIN2(_39829), .Q(_39987) );
  nor2s1 _39980_inst ( .DIN1(_39842), .DIN2(_39990), .Q(_39945) );
  xor2s1 _39981_inst ( .DIN1(_26466), .DIN2(_39840), .Q(_39990) );
  nnd2s1 _39982_inst ( .DIN1(_53438), .DIN2(_53390), .Q(_39840) );
  nnd2s1 _39983_inst ( .DIN1(_27325), .DIN2(_39991), .Q(
        ____3____________10_____) );
  nnd2s1 _39984_inst ( .DIN1(_39992), .DIN2(_39993), .Q(_39991) );
  nor2s1 _39985_inst ( .DIN1(_39994), .DIN2(_39995), .Q(_39993) );
  nnd2s1 _39986_inst ( .DIN1(_39996), .DIN2(_39986), .Q(_39995) );
  hi1s1 _39987_inst ( .DIN(_39351), .Q(_39986) );
  nnd2s1 _39988_inst ( .DIN1(_39997), .DIN2(_39998), .Q(_39351) );
  and2s1 _39989_inst ( .DIN1(_39831), .DIN2(_39482), .Q(_39998) );
  nnd2s1 _39990_inst ( .DIN1(_39999), .DIN2(_39768), .Q(_39482) );
  nnd2s1 _39991_inst ( .DIN1(_40000), .DIN2(_39934), .Q(_39831) );
  nor2s1 _39992_inst ( .DIN1(_40001), .DIN2(_39476), .Q(_40000) );
  nor2s1 _39993_inst ( .DIN1(_40002), .DIN2(_40003), .Q(_39997) );
  nor2s1 _39994_inst ( .DIN1(_39330), .DIN2(_40004), .Q(_40003) );
  nor2s1 _39995_inst ( .DIN1(_39383), .DIN2(_40005), .Q(_40002) );
  nor2s1 _39996_inst ( .DIN1(_39575), .DIN2(_40006), .Q(_40005) );
  hi1s1 _39997_inst ( .DIN(_40007), .Q(_39575) );
  nor2s1 _39998_inst ( .DIN1(_40008), .DIN2(_39832), .Q(_39996) );
  nor2s1 _39999_inst ( .DIN1(_39721), .DIN2(_39369), .Q(_39832) );
  nor2s1 _40000_inst ( .DIN1(_39383), .DIN2(_39331), .Q(_40008) );
  nnd2s1 _40001_inst ( .DIN1(_40009), .DIN2(_39830), .Q(_39994) );
  and2s1 _40002_inst ( .DIN1(_39816), .DIN2(_39403), .Q(_40009) );
  nor2s1 _40003_inst ( .DIN1(_40010), .DIN2(_40011), .Q(_39992) );
  nnd2s1 _40004_inst ( .DIN1(_40012), .DIN2(_40013), .Q(_40011) );
  hi1s1 _40005_inst ( .DIN(_39900), .Q(_40013) );
  nnd2s1 _40006_inst ( .DIN1(_40014), .DIN2(_40015), .Q(_39900) );
  nor2s1 _40007_inst ( .DIN1(_40016), .DIN2(_40017), .Q(_40015) );
  nor2s1 _40008_inst ( .DIN1(_39343), .DIN2(_39804), .Q(_40017) );
  hi1s1 _40009_inst ( .DIN(_39505), .Q(_40016) );
  nor2s1 _40010_inst ( .DIN1(_39429), .DIN2(_39803), .Q(_40014) );
  hi1s1 _40011_inst ( .DIN(_40018), .Q(_39803) );
  nor2s1 _40012_inst ( .DIN1(_39494), .DIN2(_39910), .Q(_40012) );
  nnd2s1 _40013_inst ( .DIN1(_39673), .DIN2(_40019), .Q(_39910) );
  nnd2s1 _40014_inst ( .DIN1(_39546), .DIN2(_40020), .Q(_40019) );
  hi1s1 _40015_inst ( .DIN(_39386), .Q(_39546) );
  nnd2s1 _40016_inst ( .DIN1(_40021), .DIN2(_39790), .Q(_39673) );
  nnd2s1 _40017_inst ( .DIN1(_40022), .DIN2(_40023), .Q(_39494) );
  nor2s1 _40018_inst ( .DIN1(_40024), .DIN2(_40025), .Q(_40023) );
  nnd2s1 _40019_inst ( .DIN1(_40026), .DIN2(_40027), .Q(_40025) );
  nor2s1 _40020_inst ( .DIN1(_40028), .DIN2(_40029), .Q(_40027) );
  nor2s1 _40021_inst ( .DIN1(_39383), .DIN2(_40030), .Q(_40029) );
  nor2s1 _40022_inst ( .DIN1(_39551), .DIN2(_39635), .Q(_40030) );
  nor2s1 _40023_inst ( .DIN1(_40031), .DIN2(_39485), .Q(_40028) );
  and2s1 _40024_inst ( .DIN1(_39407), .DIN2(_39770), .Q(_40031) );
  nor2s1 _40025_inst ( .DIN1(_40032), .DIN2(_39388), .Q(_40026) );
  nor2s1 _40026_inst ( .DIN1(_39476), .DIN2(_39602), .Q(_39388) );
  nnd2s1 _40027_inst ( .DIN1(_40033), .DIN2(_40034), .Q(_40024) );
  nor2s1 _40028_inst ( .DIN1(_40035), .DIN2(_39338), .Q(_40034) );
  hi1s1 _40029_inst ( .DIN(_39907), .Q(_39338) );
  nnd2s1 _40030_inst ( .DIN1(_40036), .DIN2(_40020), .Q(_39907) );
  hi1s1 _40031_inst ( .DIN(_39380), .Q(_40020) );
  nor2s1 _40032_inst ( .DIN1(_39889), .DIN2(_40037), .Q(_40033) );
  hi1s1 _40033_inst ( .DIN(_39729), .Q(_40037) );
  and2s1 _40034_inst ( .DIN1(_39939), .DIN2(_40038), .Q(_39889) );
  nor2s1 _40035_inst ( .DIN1(_39865), .DIN2(_39441), .Q(_39939) );
  nor2s1 _40036_inst ( .DIN1(_40039), .DIN2(_40040), .Q(_40022) );
  nnd2s1 _40037_inst ( .DIN1(_40041), .DIN2(_40042), .Q(_40040) );
  nor2s1 _40038_inst ( .DIN1(_40043), .DIN2(_39447), .Q(_40042) );
  nnd2s1 _40039_inst ( .DIN1(_40044), .DIN2(_40045), .Q(_39447) );
  xor2s1 _40040_inst ( .DIN1(_39890), .DIN2(_40046), .Q(_40045) );
  nor2s1 _40041_inst ( .DIN1(_40047), .DIN2(_40048), .Q(_40044) );
  nor2s1 _40042_inst ( .DIN1(_39588), .DIN2(_40049), .Q(_40048) );
  nnd2s1 _40043_inst ( .DIN1(_40050), .DIN2(_39638), .Q(_40049) );
  nor2s1 _40044_inst ( .DIN1(_40051), .DIN2(_40052), .Q(_40047) );
  nnd2s1 _40045_inst ( .DIN1(_40053), .DIN2(_39706), .Q(_40052) );
  nor2s1 _40046_inst ( .DIN1(_39685), .DIN2(_39982), .Q(_40041) );
  nnd2s1 _40047_inst ( .DIN1(_40054), .DIN2(_40055), .Q(_39982) );
  nor2s1 _40048_inst ( .DIN1(_39785), .DIN2(_40056), .Q(_40055) );
  hi1s1 _40049_inst ( .DIN(_39712), .Q(_40056) );
  nnd2s1 _40050_inst ( .DIN1(_40057), .DIN2(_39932), .Q(_39712) );
  hi1s1 _40051_inst ( .DIN(_39390), .Q(_39932) );
  nor2s1 _40052_inst ( .DIN1(_39956), .DIN2(_40058), .Q(_40057) );
  and2s1 _40053_inst ( .DIN1(_40059), .DIN2(_39638), .Q(_39785) );
  and2s1 _40054_inst ( .DIN1(_39923), .DIN2(_39853), .Q(_40054) );
  nnd2s1 _40055_inst ( .DIN1(_40060), .DIN2(_40061), .Q(_39923) );
  nor2s1 _40056_inst ( .DIN1(_39430), .DIN2(_40058), .Q(_40060) );
  nnd2s1 _40057_inst ( .DIN1(_40062), .DIN2(_40063), .Q(_39685) );
  or2s1 _40058_inst ( .DIN1(_39787), .DIN2(_39390), .Q(_40063) );
  nor2s1 _40059_inst ( .DIN1(_40064), .DIN2(_40065), .Q(_40062) );
  nor2s1 _40060_inst ( .DIN1(_39372), .DIN2(_39872), .Q(_40065) );
  nor2s1 _40061_inst ( .DIN1(_40066), .DIN2(_39633), .Q(_40064) );
  nnd2s1 _40062_inst ( .DIN1(_40067), .DIN2(_40068), .Q(_40039) );
  nor2s1 _40063_inst ( .DIN1(_39406), .DIN2(_39722), .Q(_40068) );
  nnd2s1 _40064_inst ( .DIN1(_40069), .DIN2(_40070), .Q(_39406) );
  nnd2s1 _40065_inst ( .DIN1(_40071), .DIN2(_40072), .Q(_40070) );
  nor2s1 _40066_inst ( .DIN1(_39380), .DIN2(_40073), .Q(_40072) );
  nnd2s1 _40067_inst ( .DIN1(_40074), .DIN2(_39813), .Q(_40069) );
  nor2s1 _40068_inst ( .DIN1(_39857), .DIN2(_39649), .Q(_40067) );
  nnd2s1 _40069_inst ( .DIN1(_40075), .DIN2(_40076), .Q(_39857) );
  nnd2s1 _40070_inst ( .DIN1(_40077), .DIN2(_40078), .Q(_40010) );
  hi1s1 _40071_inst ( .DIN(_39453), .Q(_40078) );
  nnd2s1 _40072_inst ( .DIN1(_40079), .DIN2(_40080), .Q(_39453) );
  nor2s1 _40073_inst ( .DIN1(_40081), .DIN2(_40082), .Q(_40080) );
  nnd2s1 _40074_inst ( .DIN1(_40083), .DIN2(_39929), .Q(_40082) );
  nnd2s1 _40075_inst ( .DIN1(_39344), .DIN2(_39758), .Q(_40083) );
  nnd2s1 _40076_inst ( .DIN1(_39672), .DIN2(_40084), .Q(_40081) );
  hi1s1 _40077_inst ( .DIN(_40085), .Q(_40084) );
  nnd2s1 _40078_inst ( .DIN1(_40086), .DIN2(_39927), .Q(_39672) );
  nor2s1 _40079_inst ( .DIN1(_39330), .DIN2(_40087), .Q(_40086) );
  nor2s1 _40080_inst ( .DIN1(_40088), .DIN2(_40089), .Q(_40079) );
  nnd2s1 _40081_inst ( .DIN1(_40090), .DIN2(_40091), .Q(_40089) );
  nnd2s1 _40082_inst ( .DIN1(_39678), .DIN2(_39638), .Q(_40091) );
  hi1s1 _40083_inst ( .DIN(_39859), .Q(_39678) );
  nnd2s1 _40084_inst ( .DIN1(_39603), .DIN2(_39790), .Q(_40090) );
  and2s1 _40085_inst ( .DIN1(_40092), .DIN2(_40093), .Q(_39603) );
  nor2s1 _40086_inst ( .DIN1(_40094), .DIN2(_40095), .Q(_40092) );
  nor2s1 _40087_inst ( .DIN1(_39614), .DIN2(_39390), .Q(_40088) );
  nor2s1 _40088_inst ( .DIN1(_39398), .DIN2(_40096), .Q(_40077) );
  nnd2s1 _40089_inst ( .DIN1(_40097), .DIN2(_40098), .Q(_39398) );
  nor2s1 _40090_inst ( .DIN1(_40099), .DIN2(_40100), .Q(_40098) );
  nnd2s1 _40091_inst ( .DIN1(_40101), .DIN2(_40102), .Q(_40100) );
  nnd2s1 _40092_inst ( .DIN1(_39566), .DIN2(_39710), .Q(_40102) );
  hi1s1 _40093_inst ( .DIN(_40103), .Q(_39566) );
  nnd2s1 _40094_inst ( .DIN1(_39345), .DIN2(_39758), .Q(_40101) );
  hi1s1 _40095_inst ( .DIN(_39989), .Q(_39345) );
  nnd2s1 _40096_inst ( .DIN1(_40104), .DIN2(_40105), .Q(_40099) );
  nnd2s1 _40097_inst ( .DIN1(_40106), .DIN2(_26838), .Q(_40104) );
  or2s1 _40098_inst ( .DIN1(_40107), .DIN2(_39709), .Q(_40106) );
  hi1s1 _40099_inst ( .DIN(_39431), .Q(_39709) );
  nor2s1 _40100_inst ( .DIN1(_40108), .DIN2(_40109), .Q(_40097) );
  nnd2s1 _40101_inst ( .DIN1(_40110), .DIN2(_39753), .Q(_40109) );
  and2s1 _40102_inst ( .DIN1(_40111), .DIN2(_40112), .Q(_39753) );
  nnd2s1 _40103_inst ( .DIN1(_39694), .DIN2(_26838), .Q(_40112) );
  hi1s1 _40104_inst ( .DIN(_39442), .Q(_39694) );
  or2s1 _40105_inst ( .DIN1(_39557), .DIN2(_39372), .Q(_40111) );
  hi1s1 _40106_inst ( .DIN(_39716), .Q(_40110) );
  nnd2s1 _40107_inst ( .DIN1(_40113), .DIN2(_40114), .Q(_39716) );
  nnd2s1 _40108_inst ( .DIN1(_39545), .DIN2(_39706), .Q(_40114) );
  hi1s1 _40109_inst ( .DIN(_39430), .Q(_39706) );
  nnd2s1 _40110_inst ( .DIN1(_40115), .DIN2(_39774), .Q(_40108) );
  nnd2s1 _40111_inst ( .DIN1(_40116), .DIN2(_40117), .Q(
        ____3____________0_____) );
  nnd2s1 _40112_inst ( .DIN1(_40118), .DIN2(_29658), .Q(_40117) );
  nor2s1 _40113_inst ( .DIN1(_27476), .DIN2(_36388), .Q(_29658) );
  nor2s1 _40114_inst ( .DIN1(_35370), .DIN2(_40119), .Q(_36388) );
  nor2s1 _40115_inst ( .DIN1(_26774), .DIN2(_26386), .Q(_40118) );
  nnd2s1 _40116_inst ( .DIN1(_27476), .DIN2(_40120), .Q(_40116) );
  nnd2s1 _40117_inst ( .DIN1(_40121), .DIN2(_40122), .Q(_40120) );
  nor2s1 _40118_inst ( .DIN1(_40123), .DIN2(_40124), .Q(_40122) );
  nnd2s1 _40119_inst ( .DIN1(_40125), .DIN2(_39728), .Q(_40124) );
  nnd2s1 _40120_inst ( .DIN1(_39622), .DIN2(_39765), .Q(_39728) );
  nnd2s1 _40121_inst ( .DIN1(_40126), .DIN2(_26838), .Q(_40125) );
  nnd2s1 _40122_inst ( .DIN1(_40127), .DIN2(_40128), .Q(_40126) );
  nor2s1 _40123_inst ( .DIN1(_40129), .DIN2(_40130), .Q(_40128) );
  nnd2s1 _40124_inst ( .DIN1(_40131), .DIN2(_40132), .Q(_40130) );
  nor2s1 _40125_inst ( .DIN1(_40133), .DIN2(_40134), .Q(_40132) );
  nnd2s1 _40126_inst ( .DIN1(_40103), .DIN2(_39407), .Q(_40134) );
  nnd2s1 _40127_inst ( .DIN1(_40135), .DIN2(_40050), .Q(_39407) );
  nor2s1 _40128_inst ( .DIN1(_40073), .DIN2(_39780), .Q(_40135) );
  nnd2s1 _40129_inst ( .DIN1(_40136), .DIN2(_40137), .Q(_40103) );
  nor2s1 _40130_inst ( .DIN1(_40138), .DIN2(_40139), .Q(_40136) );
  nor2s1 _40131_inst ( .DIN1(_40140), .DIN2(_40051), .Q(_40133) );
  nor2s1 _40132_inst ( .DIN1(_40053), .DIN2(_40141), .Q(_40140) );
  nor2s1 _40133_inst ( .DIN1(_40142), .DIN2(_40143), .Q(_40131) );
  nor2s1 _40134_inst ( .DIN1(_40144), .DIN2(_40145), .Q(_40143) );
  nor2s1 _40135_inst ( .DIN1(_40146), .DIN2(_40147), .Q(_40144) );
  nor2s1 _40136_inst ( .DIN1(_40148), .DIN2(_39587), .Q(_40146) );
  and2s1 _40137_inst ( .DIN1(_40149), .DIN2(_40150), .Q(_40148) );
  nor2s1 _40138_inst ( .DIN1(_40151), .DIN2(_40087), .Q(_40142) );
  nor2s1 _40139_inst ( .DIN1(_40152), .DIN2(_39927), .Q(_40151) );
  nor2s1 _40140_inst ( .DIN1(_40153), .DIN2(_39780), .Q(_40152) );
  nor2s1 _40141_inst ( .DIN1(_39814), .DIN2(_40154), .Q(_40153) );
  nnd2s1 _40142_inst ( .DIN1(_40155), .DIN2(_40156), .Q(_40129) );
  nor2s1 _40143_inst ( .DIN1(_40074), .DIN2(_40157), .Q(_40156) );
  nnd2s1 _40144_inst ( .DIN1(_40158), .DIN2(_39666), .Q(_40157) );
  nnd2s1 _40145_inst ( .DIN1(_40159), .DIN2(_40160), .Q(_39666) );
  nor2s1 _40146_inst ( .DIN1(_40161), .DIN2(_39865), .Q(_40160) );
  and2s1 _40147_inst ( .DIN1(_40162), .DIN2(_40163), .Q(_40074) );
  nor2s1 _40148_inst ( .DIN1(_40138), .DIN2(_39864), .Q(_40162) );
  nor2s1 _40149_inst ( .DIN1(_39545), .DIN2(_40164), .Q(_40155) );
  nnd2s1 _40150_inst ( .DIN1(_39442), .DIN2(_39391), .Q(_40164) );
  nnd2s1 _40151_inst ( .DIN1(_40165), .DIN2(_39815), .Q(_39391) );
  nor2s1 _40152_inst ( .DIN1(_40150), .DIN2(_40166), .Q(_40165) );
  nnd2s1 _40153_inst ( .DIN1(_40137), .DIN2(_40167), .Q(_39442) );
  and2s1 _40154_inst ( .DIN1(_40168), .DIN2(_40050), .Q(_39545) );
  nor2s1 _40155_inst ( .DIN1(_40169), .DIN2(_40170), .Q(_40127) );
  nnd2s1 _40156_inst ( .DIN1(_40171), .DIN2(_40172), .Q(_40170) );
  nor2s1 _40157_inst ( .DIN1(_40173), .DIN2(_40174), .Q(_40172) );
  nnd2s1 _40158_inst ( .DIN1(_40175), .DIN2(_40176), .Q(_40174) );
  nnd2s1 _40159_inst ( .DIN1(_40177), .DIN2(_26306), .Q(_40176) );
  xor2s1 _40160_inst ( .DIN1(_40178), .DIN2(_31462), .Q(_40173) );
  nnd2s1 _40161_inst ( .DIN1(_40179), .DIN2(_39869), .Q(_40178) );
  nor2s1 _40162_inst ( .DIN1(_39677), .DIN2(_39344), .Q(_39869) );
  hi1s1 _40163_inst ( .DIN(_39627), .Q(_39344) );
  nnd2s1 _40164_inst ( .DIN1(_40180), .DIN2(_40181), .Q(_39627) );
  hi1s1 _40165_inst ( .DIN(_39486), .Q(_39677) );
  nnd2s1 _40166_inst ( .DIN1(_40182), .DIN2(_40183), .Q(_39486) );
  nor2s1 _40167_inst ( .DIN1(_40001), .DIN2(_40184), .Q(_40182) );
  nor2s1 _40168_inst ( .DIN1(_39584), .DIN2(_39637), .Q(_40179) );
  nnd2s1 _40169_inst ( .DIN1(_39859), .DIN2(_39771), .Q(_39584) );
  nnd2s1 _40170_inst ( .DIN1(_40185), .DIN2(_40093), .Q(_39771) );
  nnd2s1 _40171_inst ( .DIN1(_40186), .DIN2(_40187), .Q(_39859) );
  nor2s1 _40172_inst ( .DIN1(_39699), .DIN2(_40107), .Q(_40171) );
  nnd2s1 _40173_inst ( .DIN1(_40188), .DIN2(_39835), .Q(_40107) );
  nnd2s1 _40174_inst ( .DIN1(_40189), .DIN2(_40167), .Q(_39835) );
  nor2s1 _40175_inst ( .DIN1(_39865), .DIN2(_40190), .Q(_40189) );
  nor2s1 _40176_inst ( .DIN1(_39554), .DIN2(_39334), .Q(_40188) );
  hi1s1 _40177_inst ( .DIN(_39477), .Q(_39334) );
  nnd2s1 _40178_inst ( .DIN1(_40167), .DIN2(_40163), .Q(_39477) );
  and2s1 _40179_inst ( .DIN1(_40191), .DIN2(_40163), .Q(_39554) );
  nor2s1 _40180_inst ( .DIN1(_40161), .DIN2(_40192), .Q(_40191) );
  nnd2s1 _40181_inst ( .DIN1(_39437), .DIN2(_39385), .Q(_39699) );
  nnd2s1 _40182_inst ( .DIN1(_40193), .DIN2(_40194), .Q(_39385) );
  hi1s1 _40183_inst ( .DIN(_39864), .Q(_40193) );
  nnd2s1 _40184_inst ( .DIN1(_40186), .DIN2(_40195), .Q(_39437) );
  nnd2s1 _40185_inst ( .DIN1(_40196), .DIN2(_40197), .Q(_40169) );
  nor2s1 _40186_inst ( .DIN1(_40198), .DIN2(_40199), .Q(_40197) );
  nnd2s1 _40187_inst ( .DIN1(_40200), .DIN2(_40201), .Q(_40199) );
  nnd2s1 _40188_inst ( .DIN1(_40202), .DIN2(_39625), .Q(_40201) );
  nnd2s1 _40189_inst ( .DIN1(_40203), .DIN2(_40204), .Q(_40202) );
  nor2s1 _40190_inst ( .DIN1(_39555), .DIN2(_40205), .Q(_40204) );
  hi1s1 _40191_inst ( .DIN(_39804), .Q(_39555) );
  nnd2s1 _40192_inst ( .DIN1(_40206), .DIN2(_40207), .Q(_39804) );
  nor2s1 _40193_inst ( .DIN1(_40208), .DIN2(_40209), .Q(_40206) );
  nor2s1 _40194_inst ( .DIN1(_40210), .DIN2(_40211), .Q(_40203) );
  nor2s1 _40195_inst ( .DIN1(_26356), .DIN2(_40212), .Q(_40211) );
  nnd2s1 _40196_inst ( .DIN1(_40050), .DIN2(_40213), .Q(_40200) );
  nor2s1 _40197_inst ( .DIN1(_40214), .DIN2(_40192), .Q(_40198) );
  nor2s1 _40198_inst ( .DIN1(_40215), .DIN2(_39572), .Q(_40214) );
  nor2s1 _40199_inst ( .DIN1(_40149), .DIN2(_39587), .Q(_40215) );
  nor2s1 _40200_inst ( .DIN1(_40216), .DIN2(_40217), .Q(_40196) );
  nor2s1 _40201_inst ( .DIN1(_40218), .DIN2(_40219), .Q(_40217) );
  nor2s1 _40202_inst ( .DIN1(_40220), .DIN2(_40221), .Q(_40218) );
  nor2s1 _40203_inst ( .DIN1(_40222), .DIN2(_40192), .Q(_40221) );
  nor2s1 _40204_inst ( .DIN1(_26359), .DIN2(_39588), .Q(_40220) );
  nor2s1 _40205_inst ( .DIN1(_40223), .DIN2(_40094), .Q(_40216) );
  nor2s1 _40206_inst ( .DIN1(_40224), .DIN2(_40225), .Q(_40223) );
  nor2s1 _40207_inst ( .DIN1(_40095), .DIN2(_40219), .Q(_40224) );
  nnd2s1 _40208_inst ( .DIN1(_39505), .DIN2(_39816), .Q(_40123) );
  nnd2s1 _40209_inst ( .DIN1(_39807), .DIN2(_40226), .Q(_39816) );
  hi1s1 _40210_inst ( .DIN(_39597), .Q(_39807) );
  nnd2s1 _40211_inst ( .DIN1(_40227), .DIN2(_40228), .Q(_39597) );
  nor2s1 _40212_inst ( .DIN1(_39976), .DIN2(_40073), .Q(_40227) );
  nnd2s1 _40213_inst ( .DIN1(_39622), .DIN2(_39758), .Q(_39505) );
  and2s1 _40214_inst ( .DIN1(_40229), .DIN2(_40093), .Q(_39622) );
  nor2s1 _40215_inst ( .DIN1(_40150), .DIN2(_39780), .Q(_40229) );
  nor2s1 _40216_inst ( .DIN1(_39981), .DIN2(_40230), .Q(_40121) );
  nnd2s1 _40217_inst ( .DIN1(_39644), .DIN2(_39451), .Q(_40230) );
  and2s1 _40218_inst ( .DIN1(_40231), .DIN2(_40232), .Q(_39451) );
  nor2s1 _40219_inst ( .DIN1(_40233), .DIN2(_40234), .Q(_40232) );
  nnd2s1 _40220_inst ( .DIN1(_40235), .DIN2(_40236), .Q(_40234) );
  hi1s1 _40221_inst ( .DIN(_39491), .Q(_40236) );
  nnd2s1 _40222_inst ( .DIN1(_40237), .DIN2(_40238), .Q(_39491) );
  nnd2s1 _40223_inst ( .DIN1(_40239), .DIN2(_39779), .Q(_40238) );
  hi1s1 _40224_inst ( .DIN(_40051), .Q(_39779) );
  nnd2s1 _40225_inst ( .DIN1(_40050), .DIN2(_40181), .Q(_40051) );
  nor2s1 _40226_inst ( .DIN1(_39383), .DIN2(_40145), .Q(_40239) );
  nnd2s1 _40227_inst ( .DIN1(_40240), .DIN2(_40147), .Q(_40237) );
  nor2s1 _40228_inst ( .DIN1(_40094), .DIN2(_40241), .Q(_40240) );
  nor2s1 _40229_inst ( .DIN1(_40032), .DIN2(_39327), .Q(_40235) );
  nnd2s1 _40230_inst ( .DIN1(_40242), .DIN2(_40115), .Q(_39327) );
  and2s1 _40231_inst ( .DIN1(_39925), .DIN2(_40243), .Q(_40115) );
  nnd2s1 _40232_inst ( .DIN1(_39680), .DIN2(_26838), .Q(_40243) );
  hi1s1 _40233_inst ( .DIN(_39626), .Q(_39680) );
  nnd2s1 _40234_inst ( .DIN1(_40159), .DIN2(_40244), .Q(_39626) );
  nor2s1 _40235_inst ( .DIN1(_40150), .DIN2(_39865), .Q(_40244) );
  and2s1 _40236_inst ( .DIN1(_40245), .DIN2(_40246), .Q(_39925) );
  nnd2s1 _40237_inst ( .DIN1(_40247), .DIN2(_40093), .Q(_40246) );
  and2s1 _40238_inst ( .DIN1(_40213), .DIN2(_39813), .Q(_40247) );
  hi1s1 _40239_inst ( .DIN(_39330), .Q(_39813) );
  nnd2s1 _40240_inst ( .DIN1(_39630), .DIN2(_26838), .Q(_39330) );
  hi1s1 _40241_inst ( .DIN(_40248), .Q(_39630) );
  nnd2s1 _40242_inst ( .DIN1(_39588), .DIN2(_40249), .Q(_40213) );
  nnd2s1 _40243_inst ( .DIN1(_40053), .DIN2(_40250), .Q(_40249) );
  hi1s1 _40244_inst ( .DIN(_39927), .Q(_39588) );
  nnd2s1 _40245_inst ( .DIN1(_39585), .DIN2(_40251), .Q(_40245) );
  and2s1 _40246_inst ( .DIN1(_40252), .DIN2(_40253), .Q(_39585) );
  nor2s1 _40247_inst ( .DIN1(_40161), .DIN2(_39976), .Q(_40253) );
  and2s1 _40248_inst ( .DIN1(_40254), .DIN2(_40255), .Q(_40252) );
  nor2s1 _40249_inst ( .DIN1(_40256), .DIN2(_40257), .Q(_40242) );
  nor2s1 _40250_inst ( .DIN1(_39343), .DIN2(_39872), .Q(_40257) );
  nnd2s1 _40251_inst ( .DIN1(_40258), .DIN2(_40228), .Q(_39872) );
  nor2s1 _40252_inst ( .DIN1(_39383), .DIN2(_39386), .Q(_40256) );
  nnd2s1 _40253_inst ( .DIN1(_40259), .DIN2(_40137), .Q(_39386) );
  xor2s1 _40254_inst ( .DIN1(_29450), .DIN2(_40168), .Q(_40259) );
  nor2s1 _40255_inst ( .DIN1(_40192), .DIN2(_40073), .Q(_40168) );
  nor2s1 _40256_inst ( .DIN1(_39737), .DIN2(_39787), .Q(_40032) );
  nnd2s1 _40257_inst ( .DIN1(_40260), .DIN2(_40261), .Q(_39787) );
  nor2s1 _40258_inst ( .DIN1(_40262), .DIN2(_34359), .Q(_40261) );
  nor2s1 _40259_inst ( .DIN1(_39956), .DIN2(_40208), .Q(_40260) );
  nnd2s1 _40260_inst ( .DIN1(_40263), .DIN2(_40264), .Q(_40233) );
  nnd2s1 _40261_inst ( .DIN1(_39899), .DIN2(_26838), .Q(_40264) );
  hi1s1 _40262_inst ( .DIN(_39633), .Q(_39899) );
  nnd2s1 _40263_inst ( .DIN1(_40265), .DIN2(_40266), .Q(_39633) );
  nor2s1 _40264_inst ( .DIN1(_40073), .DIN2(_39865), .Q(_40265) );
  nor2s1 _40265_inst ( .DIN1(_40267), .DIN2(_40268), .Q(_40263) );
  nor2s1 _40266_inst ( .DIN1(_40066), .DIN2(_39331), .Q(_40268) );
  nnd2s1 _40267_inst ( .DIN1(_40269), .DIN2(_40270), .Q(_39331) );
  and2s1 _40268_inst ( .DIN1(_39695), .DIN2(_39551), .Q(_40267) );
  nor2s1 _40269_inst ( .DIN1(_39957), .DIN2(_39976), .Q(_39551) );
  nor2s1 _40270_inst ( .DIN1(_40271), .DIN2(_40272), .Q(_40231) );
  nnd2s1 _40271_inst ( .DIN1(_40273), .DIN2(_40274), .Q(_40272) );
  xor2s1 _40272_inst ( .DIN1(_40275), .DIN2(_32005), .Q(_40274) );
  nnd2s1 _40273_inst ( .DIN1(_40276), .DIN2(_39784), .Q(_40275) );
  and2s1 _40274_inst ( .DIN1(_40105), .DIN2(_39854), .Q(_39784) );
  nnd2s1 _40275_inst ( .DIN1(_40059), .DIN2(_40251), .Q(_39854) );
  and2s1 _40276_inst ( .DIN1(_40277), .DIN2(_40270), .Q(_40059) );
  nor2s1 _40277_inst ( .DIN1(_40150), .DIN2(_40001), .Q(_40277) );
  nnd2s1 _40278_inst ( .DIN1(_40278), .DIN2(_40147), .Q(_40105) );
  nor2s1 _40279_inst ( .DIN1(_40145), .DIN2(_39485), .Q(_40278) );
  hi1s1 _40280_inst ( .DIN(_39352), .Q(_40276) );
  nnd2s1 _40281_inst ( .DIN1(_40279), .DIN2(_39504), .Q(_39352) );
  nnd2s1 _40282_inst ( .DIN1(_40280), .DIN2(_39790), .Q(_39504) );
  xor2s1 _40283_inst ( .DIN1(_40177), .DIN2(_29450), .Q(_40280) );
  and2s1 _40284_inst ( .DIN1(_40281), .DIN2(_40163), .Q(_40177) );
  nor2s1 _40285_inst ( .DIN1(_40150), .DIN2(_40192), .Q(_40281) );
  and2s1 _40286_inst ( .DIN1(_40076), .DIN2(_39870), .Q(_40279) );
  nnd2s1 _40287_inst ( .DIN1(_40282), .DIN2(_40061), .Q(_39870) );
  nor2s1 _40288_inst ( .DIN1(_40241), .DIN2(_40058), .Q(_40282) );
  nnd2s1 _40289_inst ( .DIN1(_39758), .DIN2(_40210), .Q(_40076) );
  and2s1 _40290_inst ( .DIN1(_40283), .DIN2(_40284), .Q(_40210) );
  nor2s1 _40291_inst ( .DIN1(_39976), .DIN2(_39864), .Q(_40284) );
  nor2s1 _40292_inst ( .DIN1(_40190), .DIN2(_39780), .Q(_40283) );
  nor2s1 _40293_inst ( .DIN1(_39649), .DIN2(_40043), .Q(_40273) );
  nnd2s1 _40294_inst ( .DIN1(_40285), .DIN2(_40286), .Q(_40043) );
  nnd2s1 _40295_inst ( .DIN1(_40287), .DIN2(_39927), .Q(_40286) );
  nor2s1 _40296_inst ( .DIN1(_40138), .DIN2(_40161), .Q(_39927) );
  nor2s1 _40297_inst ( .DIN1(_39383), .DIN2(_39587), .Q(_40287) );
  nnd2s1 _40298_inst ( .DIN1(_40288), .DIN2(_40141), .Q(_40285) );
  nor2s1 _40299_inst ( .DIN1(_39476), .DIN2(_40289), .Q(_40288) );
  nnd2s1 _40300_inst ( .DIN1(_39346), .DIN2(_40290), .Q(_39649) );
  or2s1 _40301_inst ( .DIN1(_40158), .DIN2(_39390), .Q(_40290) );
  nnd2s1 _40302_inst ( .DIN1(_40291), .DIN2(_40181), .Q(_40158) );
  nor2s1 _40303_inst ( .DIN1(_39780), .DIN2(_39587), .Q(_40291) );
  hi1s1 _40304_inst ( .DIN(_40163), .Q(_39587) );
  nnd2s1 _40305_inst ( .DIN1(_40292), .DIN2(_40141), .Q(_39346) );
  hi1s1 _40306_inst ( .DIN(_39780), .Q(_40141) );
  nor2s1 _40307_inst ( .DIN1(_39333), .DIN2(_40289), .Q(_40292) );
  hi1s1 _40308_inst ( .DIN(_40147), .Q(_40289) );
  nnd2s1 _40309_inst ( .DIN1(_40293), .DIN2(_39905), .Q(_40271) );
  and2s1 _40310_inst ( .DIN1(_40294), .DIN2(_40295), .Q(_39905) );
  nnd2s1 _40311_inst ( .DIN1(_39638), .DIN2(_39637), .Q(_40295) );
  nnd2s1 _40312_inst ( .DIN1(_40296), .DIN2(_40297), .Q(_39637) );
  nnd2s1 _40313_inst ( .DIN1(_40298), .DIN2(_40137), .Q(_40297) );
  nor2s1 _40314_inst ( .DIN1(_40145), .DIN2(_40073), .Q(_40298) );
  nnd2s1 _40315_inst ( .DIN1(_40050), .DIN2(_40167), .Q(_40296) );
  nor2s1 _40316_inst ( .DIN1(_39780), .DIN2(_40161), .Q(_40167) );
  nor2s1 _40317_inst ( .DIN1(_40299), .DIN2(_40300), .Q(_40294) );
  nor2s1 _40318_inst ( .DIN1(_39737), .DIN2(_40301), .Q(_40300) );
  nnd2s1 _40319_inst ( .DIN1(_39975), .DIN2(_39815), .Q(_40301) );
  nor2s1 _40320_inst ( .DIN1(_40302), .DIN2(_40303), .Q(_40299) );
  nnd2s1 _40321_inst ( .DIN1(_39573), .DIN2(_26838), .Q(_40303) );
  hi1s1 _40322_inst ( .DIN(_39572), .Q(_40302) );
  nor2s1 _40323_inst ( .DIN1(_39724), .DIN2(_39942), .Q(_40293) );
  nnd2s1 _40324_inst ( .DIN1(_40304), .DIN2(_40305), .Q(_39942) );
  nnd2s1 _40325_inst ( .DIN1(_39547), .DIN2(_39710), .Q(_40305) );
  nor2s1 _40326_inst ( .DIN1(_39941), .DIN2(_40209), .Q(_39547) );
  nor2s1 _40327_inst ( .DIN1(_40306), .DIN2(_40307), .Q(_40304) );
  nor2s1 _40328_inst ( .DIN1(_39343), .DIN2(_39475), .Q(_40307) );
  nnd2s1 _40329_inst ( .DIN1(_40308), .DIN2(_39812), .Q(_39475) );
  hi1s1 _40330_inst ( .DIN(_39961), .Q(_39812) );
  nor2s1 _40331_inst ( .DIN1(_39865), .DIN2(_40095), .Q(_40308) );
  hi1s1 _40332_inst ( .DIN(_40181), .Q(_40095) );
  nor2s1 _40333_inst ( .DIN1(_39383), .DIN2(_40309), .Q(_40306) );
  nor2s1 _40334_inst ( .DIN1(_40006), .DIN2(_40310), .Q(_40309) );
  nnd2s1 _40335_inst ( .DIN1(_39556), .DIN2(_39989), .Q(_40310) );
  nnd2s1 _40336_inst ( .DIN1(_40311), .DIN2(_40195), .Q(_39989) );
  nor2s1 _40337_inst ( .DIN1(_40166), .DIN2(_40073), .Q(_40311) );
  nnd2s1 _40338_inst ( .DIN1(_40312), .DIN2(_39815), .Q(_39556) );
  nor2s1 _40339_inst ( .DIN1(_40161), .DIN2(_40166), .Q(_40312) );
  nnd2s1 _40340_inst ( .DIN1(_39598), .DIN2(_39636), .Q(_40006) );
  nnd2s1 _40341_inst ( .DIN1(_39814), .DIN2(_40194), .Q(_39636) );
  nnd2s1 _40342_inst ( .DIN1(_40313), .DIN2(_40314), .Q(_39598) );
  nor2s1 _40343_inst ( .DIN1(_40001), .DIN2(_40315), .Q(_40313) );
  nnd2s1 _40344_inst ( .DIN1(_40316), .DIN2(_40317), .Q(_39724) );
  nor2s1 _40345_inst ( .DIN1(_40318), .DIN2(_40319), .Q(_40317) );
  nnd2s1 _40346_inst ( .DIN1(_40320), .DIN2(_40321), .Q(_40319) );
  nnd2s1 _40347_inst ( .DIN1(_39382), .DIN2(_39695), .Q(_40321) );
  hi1s1 _40348_inst ( .DIN(_39829), .Q(_39382) );
  nnd2s1 _40349_inst ( .DIN1(_40322), .DIN2(_40323), .Q(_39829) );
  nor2s1 _40350_inst ( .DIN1(_39956), .DIN2(_40324), .Q(_40323) );
  nor2s1 _40351_inst ( .DIN1(_40208), .DIN2(_39825), .Q(_40322) );
  nnd2s1 _40352_inst ( .DIN1(_39635), .DIN2(_26838), .Q(_40320) );
  nnd2s1 _40353_inst ( .DIN1(_39965), .DIN2(_39404), .Q(_40318) );
  nnd2s1 _40354_inst ( .DIN1(_40036), .DIN2(_39695), .Q(_39404) );
  nor2s1 _40355_inst ( .DIN1(_39976), .DIN2(_40325), .Q(_40036) );
  nnd2s1 _40356_inst ( .DIN1(_40326), .DIN2(_39537), .Q(_39965) );
  nnd2s1 _40357_inst ( .DIN1(_39557), .DIN2(_39602), .Q(_40326) );
  nnd2s1 _40358_inst ( .DIN1(_40180), .DIN2(_40250), .Q(_39602) );
  nor2s1 _40359_inst ( .DIN1(_40166), .DIN2(_40001), .Q(_40180) );
  nnd2s1 _40360_inst ( .DIN1(_40327), .DIN2(_40328), .Q(_39557) );
  nor2s1 _40361_inst ( .DIN1(_40329), .DIN2(_40330), .Q(_40316) );
  nnd2s1 _40362_inst ( .DIN1(_39798), .DIN2(_40331), .Q(_40330) );
  hi1s1 _40363_inst ( .DIN(_40096), .Q(_40331) );
  nnd2s1 _40364_inst ( .DIN1(_40332), .DIN2(_40333), .Q(_40096) );
  nnd2s1 _40365_inst ( .DIN1(_40334), .DIN2(_39824), .Q(_40333) );
  nor2s1 _40366_inst ( .DIN1(_34359), .DIN2(_39735), .Q(_40334) );
  nor2s1 _40367_inst ( .DIN1(_40335), .DIN2(_39401), .Q(_40332) );
  and2s1 _40368_inst ( .DIN1(_40071), .DIN2(_40336), .Q(_39401) );
  nor2s1 _40369_inst ( .DIN1(_39476), .DIN2(_40149), .Q(_40336) );
  nor2s1 _40370_inst ( .DIN1(_39780), .DIN2(_40087), .Q(_40071) );
  nnd2s1 _40371_inst ( .DIN1(_40337), .DIN2(_53440), .Q(_39780) );
  hi1s1 _40372_inst ( .DIN(_39641), .Q(_40335) );
  nnd2s1 _40373_inst ( .DIN1(_40053), .DIN2(_40338), .Q(_39641) );
  nnd2s1 _40374_inst ( .DIN1(_40339), .DIN2(_40340), .Q(_40338) );
  nnd2s1 _40375_inst ( .DIN1(_40341), .DIN2(_40050), .Q(_40340) );
  nor2s1 _40376_inst ( .DIN1(_40222), .DIN2(_39390), .Q(_40341) );
  nnd2s1 _40377_inst ( .DIN1(_39928), .DIN2(_39814), .Q(_40339) );
  and2s1 _40378_inst ( .DIN1(_40342), .DIN2(_40343), .Q(_39798) );
  nor2s1 _40379_inst ( .DIN1(_40035), .DIN2(_40344), .Q(_40343) );
  nor2s1 _40380_inst ( .DIN1(_39957), .DIN2(_40345), .Q(_40344) );
  nnd2s1 _40381_inst ( .DIN1(_39884), .DIN2(_39815), .Q(_40345) );
  and2s1 _40382_inst ( .DIN1(_40205), .DIN2(_39758), .Q(_40035) );
  hi1s1 _40383_inst ( .DIN(_39372), .Q(_39758) );
  and2s1 _40384_inst ( .DIN1(_40159), .DIN2(_40346), .Q(_40205) );
  nor2s1 _40385_inst ( .DIN1(_39956), .DIN2(_40139), .Q(_40346) );
  nor2s1 _40386_inst ( .DIN1(_40190), .DIN2(_40192), .Q(_40159) );
  nor2s1 _40387_inst ( .DIN1(_40347), .DIN2(_39499), .Q(_40342) );
  nnd2s1 _40388_inst ( .DIN1(_40348), .DIN2(_40349), .Q(_39499) );
  nnd2s1 _40389_inst ( .DIN1(_39999), .DIN2(_40226), .Q(_40349) );
  nor2s1 _40390_inst ( .DIN1(_40325), .DIN2(_40001), .Q(_39999) );
  nnd2s1 _40391_inst ( .DIN1(_40350), .DIN2(_34370), .Q(_40325) );
  hi1s1 _40392_inst ( .DIN(_34359), .Q(_34370) );
  nor2s1 _40393_inst ( .DIN1(_40145), .DIN2(_40161), .Q(_40350) );
  or2s1 _40394_inst ( .DIN1(_40066), .DIN2(_40004), .Q(_40348) );
  nnd2s1 _40395_inst ( .DIN1(_39960), .DIN2(_40270), .Q(_40004) );
  nor2s1 _40396_inst ( .DIN1(_39383), .DIN2(_40007), .Q(_40347) );
  nnd2s1 _40397_inst ( .DIN1(_40194), .DIN2(_40154), .Q(_40007) );
  xor2s1 _40398_inst ( .DIN1(_31269), .DIN2(_40351), .Q(_40329) );
  and2s1 _40399_inst ( .DIN1(_39782), .DIN2(_39853), .Q(_40351) );
  nnd2s1 _40400_inst ( .DIN1(_40352), .DIN2(_40353), .Q(_39853) );
  xnr2s1 _40401_inst ( .DIN1(_40354), .DIN2(_31975), .Q(_40353) );
  nnd2s1 _40402_inst ( .DIN1(_40266), .DIN2(_39815), .Q(_40354) );
  hi1s1 _40403_inst ( .DIN(_40355), .Q(_40266) );
  nor2s1 _40404_inst ( .DIN1(_39383), .DIN2(_40150), .Q(_40352) );
  nnd2s1 _40405_inst ( .DIN1(_40021), .DIN2(_39736), .Q(_39782) );
  and2s1 _40406_inst ( .DIN1(_40258), .DIN2(_40270), .Q(_40021) );
  hi1s1 _40407_inst ( .DIN(_39866), .Q(_40270) );
  nor2s1 _40408_inst ( .DIN1(_39865), .DIN2(_40149), .Q(_40258) );
  and2s1 _40409_inst ( .DIN1(_40356), .DIN2(_40357), .Q(_39644) );
  nor2s1 _40410_inst ( .DIN1(_40358), .DIN2(_40359), .Q(_40357) );
  nnd2s1 _40411_inst ( .DIN1(_40360), .DIN2(_39730), .Q(_40359) );
  nnd2s1 _40412_inst ( .DIN1(_40361), .DIN2(_39638), .Q(_39730) );
  nnd2s1 _40413_inst ( .DIN1(_39757), .DIN2(_39765), .Q(_40360) );
  hi1s1 _40414_inst ( .DIN(_39343), .Q(_39765) );
  nnd2s1 _40415_inst ( .DIN1(_39625), .DIN2(_39537), .Q(_39343) );
  hi1s1 _40416_inst ( .DIN(_39883), .Q(_39757) );
  nnd2s1 _40417_inst ( .DIN1(_40362), .DIN2(_40363), .Q(_39883) );
  nor2s1 _40418_inst ( .DIN1(_40138), .DIN2(_40073), .Q(_40362) );
  nnd2s1 _40419_inst ( .DIN1(_40364), .DIN2(_39403), .Q(_40358) );
  nnd2s1 _40420_inst ( .DIN1(_40361), .DIN2(_40251), .Q(_39403) );
  and2s1 _40421_inst ( .DIN1(_40365), .DIN2(_40137), .Q(_40361) );
  hi1s1 _40422_inst ( .DIN(_40087), .Q(_40137) );
  nor2s1 _40423_inst ( .DIN1(_39864), .DIN2(_40192), .Q(_40365) );
  and2s1 _40424_inst ( .DIN1(_40113), .DIN2(_39877), .Q(_40364) );
  nnd2s1 _40425_inst ( .DIN1(_39537), .DIN2(_40366), .Q(_39877) );
  nnd2s1 _40426_inst ( .DIN1(_39373), .DIN2(_39368), .Q(_40366) );
  nnd2s1 _40427_inst ( .DIN1(_40367), .DIN2(_40328), .Q(_39368) );
  nor2s1 _40428_inst ( .DIN1(_40166), .DIN2(_40149), .Q(_40367) );
  nnd2s1 _40429_inst ( .DIN1(_40368), .DIN2(_39814), .Q(_39373) );
  nor2s1 _40430_inst ( .DIN1(_40001), .DIN2(_40355), .Q(_40368) );
  nnd2s1 _40431_inst ( .DIN1(_39934), .DIN2(_40369), .Q(_40113) );
  nnd2s1 _40432_inst ( .DIN1(_40370), .DIN2(_40371), .Q(_40369) );
  or2s1 _40433_inst ( .DIN1(_39333), .DIN2(_40001), .Q(_40371) );
  nnd2s1 _40434_inst ( .DIN1(_40372), .DIN2(_53442), .Q(_40001) );
  nor2s1 _40435_inst ( .DIN1(_53436), .DIN2(_53443), .Q(_40372) );
  nnd2s1 _40436_inst ( .DIN1(_39884), .DIN2(_39933), .Q(_40370) );
  hi1s1 _40437_inst ( .DIN(_39737), .Q(_39884) );
  nor2s1 _40438_inst ( .DIN1(_39866), .DIN2(_40161), .Q(_39934) );
  nnd2s1 _40439_inst ( .DIN1(_40373), .DIN2(_53392), .Q(_40161) );
  nor2s1 _40440_inst ( .DIN1(_40374), .DIN2(_40375), .Q(_40356) );
  nnd2s1 _40441_inst ( .DIN1(_40018), .DIN2(_40075), .Q(_40375) );
  and2s1 _40442_inst ( .DIN1(_40376), .DIN2(_40377), .Q(_40075) );
  nnd2s1 _40443_inst ( .DIN1(_40378), .DIN2(_40147), .Q(_40377) );
  xor2s1 _40444_inst ( .DIN1(_30186), .DIN2(_40379), .Q(_40147) );
  nor2s1 _40445_inst ( .DIN1(_40190), .DIN2(_40380), .Q(_40379) );
  nnd2s1 _40446_inst ( .DIN1(_39814), .DIN2(_39933), .Q(_40380) );
  nor2s1 _40447_inst ( .DIN1(_40094), .DIN2(_39430), .Q(_40378) );
  or2s1 _40448_inst ( .DIN1(_40175), .DIN2(_39380), .Q(_40376) );
  xnr2s1 _40449_inst ( .DIN1(_34338), .DIN2(_40381), .Q(_40175) );
  nor2s1 _40450_inst ( .DIN1(_40382), .DIN2(_40383), .Q(_40381) );
  nnd2s1 _40451_inst ( .DIN1(_40384), .DIN2(_39815), .Q(_40383) );
  hi1s1 _40452_inst ( .DIN(_39956), .Q(_39815) );
  nnd2s1 _40453_inst ( .DIN1(_40154), .DIN2(_39916), .Q(_40382) );
  hi1s1 _40454_inst ( .DIN(_40073), .Q(_40154) );
  xor2s1 _40455_inst ( .DIN1(_29994), .DIN2(_40385), .Q(_40018) );
  nor2s1 _40456_inst ( .DIN1(_40386), .DIN2(_39670), .Q(_40385) );
  nor2s1 _40457_inst ( .DIN1(_39770), .DIN2(_39735), .Q(_39670) );
  nnd2s1 _40458_inst ( .DIN1(_40387), .DIN2(_40388), .Q(_39770) );
  nor2s1 _40459_inst ( .DIN1(_34359), .DIN2(_39865), .Q(_40388) );
  nor2s1 _40460_inst ( .DIN1(_40324), .DIN2(_40208), .Q(_40387) );
  nor2s1 _40461_inst ( .DIN1(_39369), .DIN2(_40389), .Q(_40386) );
  nnd2s1 _40462_inst ( .DIN1(_40038), .DIN2(_40195), .Q(_40389) );
  hi1s1 _40463_inst ( .DIN(_39957), .Q(_40038) );
  nnd2s1 _40464_inst ( .DIN1(_40181), .DIN2(_40228), .Q(_39957) );
  and2s1 _40465_inst ( .DIN1(_40207), .DIN2(_26238), .Q(_40228) );
  nnd2s1 _40466_inst ( .DIN1(_40390), .DIN2(_40391), .Q(_29994) );
  nor2s1 _40467_inst ( .DIN1(_40392), .DIN2(_40393), .Q(_40391) );
  nnd2s1 _40468_inst ( .DIN1(_40394), .DIN2(_40395), .Q(_40393) );
  nor2s1 _40469_inst ( .DIN1(_40396), .DIN2(_40397), .Q(_40392) );
  nor2s1 _40470_inst ( .DIN1(_40398), .DIN2(_40399), .Q(_40390) );
  nnd2s1 _40471_inst ( .DIN1(_40400), .DIN2(_39774), .Q(_40374) );
  and2s1 _40472_inst ( .DIN1(_40401), .DIN2(_40402), .Q(_39774) );
  nnd2s1 _40473_inst ( .DIN1(_40403), .DIN2(_39960), .Q(_40402) );
  nor2s1 _40474_inst ( .DIN1(_39976), .DIN2(_40139), .Q(_39960) );
  nor2s1 _40475_inst ( .DIN1(_39961), .DIN2(_39369), .Q(_40403) );
  nnd2s1 _40476_inst ( .DIN1(_40185), .DIN2(_39928), .Q(_40401) );
  hi1s1 _40477_inst ( .DIN(_39914), .Q(_39928) );
  nnd2s1 _40478_inst ( .DIN1(_40163), .DIN2(_39638), .Q(_39914) );
  nor2s1 _40479_inst ( .DIN1(_40190), .DIN2(_40404), .Q(_40163) );
  nor2s1 _40480_inst ( .DIN1(_40145), .DIN2(_40150), .Q(_40185) );
  hi1s1 _40481_inst ( .DIN(_39916), .Q(_40145) );
  nor2s1 _40482_inst ( .DIN1(_26238), .DIN2(_40262), .Q(_39916) );
  hi1s1 _40483_inst ( .DIN(_39355), .Q(_40400) );
  nnd2s1 _40484_inst ( .DIN1(_40405), .DIN2(_39906), .Q(_39355) );
  and2s1 _40485_inst ( .DIN1(_40406), .DIN2(_40407), .Q(_39906) );
  nor2s1 _40486_inst ( .DIN1(_40408), .DIN2(_40409), .Q(_40407) );
  nnd2s1 _40487_inst ( .DIN1(_40410), .DIN2(_40411), .Q(_40409) );
  nnd2s1 _40488_inst ( .DIN1(_40412), .DIN2(_40413), .Q(_40411) );
  hi1s1 _40489_inst ( .DIN(_40212), .Q(_40413) );
  nnd2s1 _40490_inst ( .DIN1(_40414), .DIN2(_40093), .Q(_40212) );
  nor2s1 _40491_inst ( .DIN1(_26228), .DIN2(_40208), .Q(_40414) );
  nor2s1 _40492_inst ( .DIN1(_26356), .DIN2(_39372), .Q(_40412) );
  nnd2s1 _40493_inst ( .DIN1(_39619), .DIN2(_39537), .Q(_39372) );
  hi1s1 _40494_inst ( .DIN(_39625), .Q(_39619) );
  nnd2s1 _40495_inst ( .DIN1(_40415), .DIN2(_27651), .Q(_39625) );
  nnd2s1 _40496_inst ( .DIN1(_40416), .DIN2(_39824), .Q(_40410) );
  and2s1 _40497_inst ( .DIN1(_40417), .DIN2(_40254), .Q(_39824) );
  nor2s1 _40498_inst ( .DIN1(_40241), .DIN2(_39825), .Q(_40416) );
  nor2s1 _40499_inst ( .DIN1(_39369), .DIN2(_40418), .Q(_40408) );
  nnd2s1 _40500_inst ( .DIN1(_39975), .DIN2(_39933), .Q(_40418) );
  hi1s1 _40501_inst ( .DIN(_39976), .Q(_39933) );
  hi1s1 _40502_inst ( .DIN(_40058), .Q(_39975) );
  nnd2s1 _40503_inst ( .DIN1(_40419), .DIN2(_40255), .Q(_40058) );
  nor2s1 _40504_inst ( .DIN1(_40262), .DIN2(_40208), .Q(_40419) );
  nnd2s1 _40505_inst ( .DIN1(_40250), .DIN2(_53440), .Q(_40208) );
  nor2s1 _40506_inst ( .DIN1(_39722), .DIN2(_40420), .Q(_40406) );
  nnd2s1 _40507_inst ( .DIN1(_40421), .DIN2(_40422), .Q(_40420) );
  nnd2s1 _40508_inst ( .DIN1(_40423), .DIN2(_39537), .Q(_40422) );
  nnd2s1 _40509_inst ( .DIN1(_39374), .DIN2(_39431), .Q(_40423) );
  nnd2s1 _40510_inst ( .DIN1(_40424), .DIN2(_40050), .Q(_39431) );
  and2s1 _40511_inst ( .DIN1(_40328), .DIN2(_40384), .Q(_40050) );
  and2s1 _40512_inst ( .DIN1(_40425), .DIN2(_26288), .Q(_40328) );
  nor2s1 _40513_inst ( .DIN1(_40139), .DIN2(_40192), .Q(_40424) );
  nnd2s1 _40514_inst ( .DIN1(_40426), .DIN2(_40093), .Q(_39374) );
  hi1s1 _40515_inst ( .DIN(_40219), .Q(_40093) );
  nnd2s1 _40516_inst ( .DIN1(_40384), .DIN2(_40187), .Q(_40219) );
  nor2s1 _40517_inst ( .DIN1(_40138), .DIN2(_40222), .Q(_40426) );
  hi1s1 _40518_inst ( .DIN(_40250), .Q(_40222) );
  nor2s1 _40519_inst ( .DIN1(_40184), .DIN2(_26437), .Q(_40250) );
  hi1s1 _40520_inst ( .DIN(_39478), .Q(_40421) );
  xor2s1 _40521_inst ( .DIN1(_40427), .DIN2(_27956), .Q(_39478) );
  hi1s1 _40522_inst ( .DIN(_37195), .Q(_27956) );
  nnd2s1 _40523_inst ( .DIN1(_40428), .DIN2(_40269), .Q(_40427) );
  nor2s1 _40524_inst ( .DIN1(_39956), .DIN2(_40149), .Q(_40269) );
  nor2s1 _40525_inst ( .DIN1(_39961), .DIN2(_40066), .Q(_40428) );
  nnd2s1 _40526_inst ( .DIN1(_40248), .DIN2(_39537), .Q(_40066) );
  nnd2s1 _40527_inst ( .DIN1(_40429), .DIN2(______[6]), .Q(_40248) );
  nor2s1 _40528_inst ( .DIN1(______[15]), .DIN2(______[14]), .Q(_40429) );
  nnd2s1 _40529_inst ( .DIN1(_40430), .DIN2(_40431), .Q(_39961) );
  nor2s1 _40530_inst ( .DIN1(_26238), .DIN2(_34359), .Q(_40430) );
  nnd2s1 _40531_inst ( .DIN1(_40432), .DIN2(_40433), .Q(_39722) );
  nnd2s1 _40532_inst ( .DIN1(_40225), .DIN2(_40434), .Q(_40433) );
  nor2s1 _40533_inst ( .DIN1(_40094), .DIN2(_39441), .Q(_40434) );
  nor2s1 _40534_inst ( .DIN1(_40149), .DIN2(_40087), .Q(_40225) );
  nnd2s1 _40535_inst ( .DIN1(_40435), .DIN2(_39572), .Q(_40432) );
  nor2s1 _40536_inst ( .DIN1(_40087), .DIN2(_40150), .Q(_39572) );
  nnd2s1 _40537_inst ( .DIN1(_40061), .DIN2(_40384), .Q(_40087) );
  hi1s1 _40538_inst ( .DIN(_40190), .Q(_40384) );
  nnd2s1 _40539_inst ( .DIN1(_26587), .DIN2(_26286), .Q(_40190) );
  hi1s1 _40540_inst ( .DIN(_40209), .Q(_40061) );
  nnd2s1 _40541_inst ( .DIN1(_40436), .DIN2(_53436), .Q(_40209) );
  nor2s1 _40542_inst ( .DIN1(_53442), .DIN2(_26288), .Q(_40436) );
  nor2s1 _40543_inst ( .DIN1(_40192), .DIN2(_39390), .Q(_40435) );
  hi1s1 _40544_inst ( .DIN(_40053), .Q(_40192) );
  nor2s1 _40545_inst ( .DIN1(_40324), .DIN2(_53440), .Q(_40053) );
  nor2s1 _40546_inst ( .DIN1(_39696), .DIN2(_40437), .Q(_40405) );
  nor2s1 _40547_inst ( .DIN1(_39941), .DIN2(_40438), .Q(_40437) );
  nnd2s1 _40548_inst ( .DIN1(_40251), .DIN2(_40195), .Q(_40438) );
  hi1s1 _40549_inst ( .DIN(_39865), .Q(_40195) );
  hi1s1 _40550_inst ( .DIN(_39369), .Q(_40251) );
  nnd2s1 _40551_inst ( .DIN1(_39579), .DIN2(_39537), .Q(_39369) );
  nnd2s1 _40552_inst ( .DIN1(_40439), .DIN2(_40181), .Q(_39941) );
  nor2s1 _40553_inst ( .DIN1(_40184), .DIN2(_53392), .Q(_40181) );
  nnd2s1 _40554_inst ( .DIN1(_53435), .DIN2(_26211), .Q(_40184) );
  nor2s1 _40555_inst ( .DIN1(_34359), .DIN2(_40138), .Q(_40439) );
  hi1s1 _40556_inst ( .DIN(_39830), .Q(_39696) );
  nnd2s1 _40557_inst ( .DIN1(_40440), .DIN2(_40417), .Q(_39830) );
  nor2s1 _40558_inst ( .DIN1(_39864), .DIN2(_39865), .Q(_40417) );
  nnd2s1 _40559_inst ( .DIN1(_40314), .DIN2(_53392), .Q(_39864) );
  nor2s1 _40560_inst ( .DIN1(_39436), .DIN2(_39866), .Q(_40440) );
  nnd2s1 _40561_inst ( .DIN1(_40207), .DIN2(_53440), .Q(_39866) );
  and2s1 _40562_inst ( .DIN1(_40255), .DIN2(_40431), .Q(_40207) );
  hi1s1 _40563_inst ( .DIN(_39825), .Q(_40255) );
  nnd2s1 _40564_inst ( .DIN1(_53439), .DIN2(_26286), .Q(_39825) );
  nnd2s1 _40565_inst ( .DIN1(_40441), .DIN2(_40442), .Q(_39981) );
  nor2s1 _40566_inst ( .DIN1(_40085), .DIN2(_40443), .Q(_40442) );
  nor2s1 _40567_inst ( .DIN1(_39383), .DIN2(_39614), .Q(_40443) );
  nnd2s1 _40568_inst ( .DIN1(_39794), .DIN2(_40194), .Q(_39614) );
  nor2s1 _40569_inst ( .DIN1(_40444), .DIN2(_40166), .Q(_40194) );
  nor2s1 _40570_inst ( .DIN1(_39793), .DIN2(_40445), .Q(_40085) );
  nor2s1 _40571_inst ( .DIN1(_39736), .DIN2(_39790), .Q(_40445) );
  nnd2s1 _40572_inst ( .DIN1(_40446), .DIN2(_40373), .Q(_39793) );
  nor2s1 _40573_inst ( .DIN1(_26211), .DIN2(_26686), .Q(_40373) );
  nor2s1 _40574_inst ( .DIN1(_40315), .DIN2(_39956), .Q(_40446) );
  nnd2s1 _40575_inst ( .DIN1(_40447), .DIN2(_53436), .Q(_39956) );
  nor2s1 _40576_inst ( .DIN1(_53442), .DIN2(_53443), .Q(_40447) );
  and2s1 _40577_inst ( .DIN1(_39776), .DIN2(_39350), .Q(_40441) );
  and2s1 _40578_inst ( .DIN1(_40448), .DIN2(_40449), .Q(_39350) );
  nor2s1 _40579_inst ( .DIN1(_40450), .DIN2(_40451), .Q(_40449) );
  nnd2s1 _40580_inst ( .DIN1(_40452), .DIN2(_39729), .Q(_40451) );
  nnd2s1 _40581_inst ( .DIN1(_39574), .DIN2(_39710), .Q(_39729) );
  hi1s1 _40582_inst ( .DIN(_40241), .Q(_39710) );
  nnd2s1 _40583_inst ( .DIN1(_39567), .DIN2(_39537), .Q(_40241) );
  hi1s1 _40584_inst ( .DIN(_40453), .Q(_39574) );
  nnd2s1 _40585_inst ( .DIN1(_40454), .DIN2(_39790), .Q(_40452) );
  hi1s1 _40586_inst ( .DIN(_39476), .Q(_39790) );
  nnd2s1 _40587_inst ( .DIN1(_39604), .DIN2(_39537), .Q(_39476) );
  hi1s1 _40588_inst ( .DIN(_39601), .Q(_39604) );
  nor2s1 _40589_inst ( .DIN1(_40453), .DIN2(_39430), .Q(_40450) );
  nnd2s1 _40590_inst ( .DIN1(_39568), .DIN2(_39537), .Q(_39430) );
  hi1s1 _40591_inst ( .DIN(_39567), .Q(_39568) );
  nnd2s1 _40592_inst ( .DIN1(_40455), .DIN2(______[15]), .Q(_39567) );
  nor2s1 _40593_inst ( .DIN1(______[6]), .DIN2(_27651), .Q(_40455) );
  nnd2s1 _40594_inst ( .DIN1(_40456), .DIN2(_39794), .Q(_40453) );
  hi1s1 _40595_inst ( .DIN(_40139), .Q(_39794) );
  nor2s1 _40596_inst ( .DIN1(_40166), .DIN2(_39865), .Q(_40456) );
  nnd2s1 _40597_inst ( .DIN1(_40457), .DIN2(_53442), .Q(_39865) );
  nor2s1 _40598_inst ( .DIN1(_53436), .DIN2(_26288), .Q(_40457) );
  nor2s1 _40599_inst ( .DIN1(_39704), .DIN2(_40458), .Q(_40448) );
  or2s1 _40600_inst ( .DIN1(_39429), .DIN2(_39479), .Q(_40458) );
  nnd2s1 _40601_inst ( .DIN1(_39929), .DIN2(_40459), .Q(_39479) );
  nnd2s1 _40602_inst ( .DIN1(_40460), .DIN2(_39638), .Q(_40459) );
  hi1s1 _40603_inst ( .DIN(_39441), .Q(_39638) );
  nnd2s1 _40604_inst ( .DIN1(_39580), .DIN2(_39537), .Q(_39441) );
  hi1s1 _40605_inst ( .DIN(_39579), .Q(_39580) );
  nnd2s1 _40606_inst ( .DIN1(_40461), .DIN2(______[15]), .Q(_39579) );
  nor2s1 _40607_inst ( .DIN1(______[14]), .DIN2(_28646), .Q(_40461) );
  nnd2s1 _40608_inst ( .DIN1(_40462), .DIN2(_40186), .Q(_39929) );
  hi1s1 _40609_inst ( .DIN(_40463), .Q(_40186) );
  nor2s1 _40610_inst ( .DIN1(_39380), .DIN2(_40404), .Q(_40462) );
  nnd2s1 _40611_inst ( .DIN1(_39549), .DIN2(_39537), .Q(_39380) );
  hi1s1 _40612_inst ( .DIN(_40464), .Q(_39549) );
  nnd2s1 _40613_inst ( .DIN1(_39713), .DIN2(_40465), .Q(_39429) );
  nnd2s1 _40614_inst ( .DIN1(_40454), .DIN2(_39736), .Q(_40465) );
  hi1s1 _40615_inst ( .DIN(_39333), .Q(_39736) );
  nnd2s1 _40616_inst ( .DIN1(_39601), .DIN2(_39537), .Q(_39333) );
  nnd2s1 _40617_inst ( .DIN1(_40466), .DIN2(______[15]), .Q(_39601) );
  nor2s1 _40618_inst ( .DIN1(______[6]), .DIN2(______[14]), .Q(_40466) );
  nor2s1 _40619_inst ( .DIN1(_40467), .DIN2(_40139), .Q(_40454) );
  nnd2s1 _40620_inst ( .DIN1(_40468), .DIN2(_53392), .Q(_40139) );
  nnd2s1 _40621_inst ( .DIN1(_39768), .DIN2(_40469), .Q(_39713) );
  hi1s1 _40622_inst ( .DIN(_39485), .Q(_39768) );
  nnd2s1 _40623_inst ( .DIN1(_39595), .DIN2(_39537), .Q(_39485) );
  hi1s1 _40624_inst ( .DIN(_39594), .Q(_39595) );
  nnd2s1 _40625_inst ( .DIN1(_40470), .DIN2(_40471), .Q(_39704) );
  nnd2s1 _40626_inst ( .DIN1(_40472), .DIN2(_39695), .Q(_40471) );
  hi1s1 _40627_inst ( .DIN(_39436), .Q(_39695) );
  nnd2s1 _40628_inst ( .DIN1(_39537), .DIN2(_40464), .Q(_39436) );
  nnd2s1 _40629_inst ( .DIN1(_40473), .DIN2(______[15]), .Q(_40464) );
  nor2s1 _40630_inst ( .DIN1(_28646), .DIN2(_27651), .Q(_40473) );
  nor2s1 _40631_inst ( .DIN1(_40404), .DIN2(_40463), .Q(_40472) );
  nnd2s1 _40632_inst ( .DIN1(_40183), .DIN2(_40468), .Q(_40463) );
  hi1s1 _40633_inst ( .DIN(_40315), .Q(_40183) );
  nnd2s1 _40634_inst ( .DIN1(_40226), .DIN2(_40469), .Q(_40470) );
  and2s1 _40635_inst ( .DIN1(_40327), .DIN2(_40187), .Q(_40469) );
  hi1s1 _40636_inst ( .DIN(_40444), .Q(_40187) );
  nor2s1 _40637_inst ( .DIN1(_40315), .DIN2(_40474), .Q(_40327) );
  nnd2s1 _40638_inst ( .DIN1(_40475), .DIN2(_40476), .Q(_40315) );
  nor2s1 _40639_inst ( .DIN1(_26437), .DIN2(_40094), .Q(_40475) );
  hi1s1 _40640_inst ( .DIN(_39573), .Q(_40094) );
  nor2s1 _40641_inst ( .DIN1(_40262), .DIN2(_53440), .Q(_39573) );
  nnd2s1 _40642_inst ( .DIN1(_26356), .DIN2(_26228), .Q(_40262) );
  hi1s1 _40643_inst ( .DIN(_39735), .Q(_40226) );
  nnd2s1 _40644_inst ( .DIN1(_39594), .DIN2(_39537), .Q(_39735) );
  nnd2s1 _40645_inst ( .DIN1(_40477), .DIN2(______[14]), .Q(_39594) );
  nor2s1 _40646_inst ( .DIN1(______[15]), .DIN2(_28646), .Q(_40477) );
  nor2s1 _40647_inst ( .DIN1(_39890), .DIN2(_40478), .Q(_39776) );
  nor2s1 _40648_inst ( .DIN1(_39390), .DIN2(_39392), .Q(_40478) );
  nnd2s1 _40649_inst ( .DIN1(_39612), .DIN2(_39537), .Q(_39390) );
  hi1s1 _40650_inst ( .DIN(_39611), .Q(_39612) );
  nor2s1 _40651_inst ( .DIN1(_39392), .DIN2(_39737), .Q(_39890) );
  nnd2s1 _40652_inst ( .DIN1(_39611), .DIN2(_39537), .Q(_39737) );
  nnd2s1 _40653_inst ( .DIN1(_40415), .DIN2(______[14]), .Q(_39611) );
  nor2s1 _40654_inst ( .DIN1(______[6]), .DIN2(______[15]), .Q(_40415) );
  nnd2s1 _40655_inst ( .DIN1(_40479), .DIN2(_39814), .Q(_39392) );
  hi1s1 _40656_inst ( .DIN(_40149), .Q(_39814) );
  nnd2s1 _40657_inst ( .DIN1(_40314), .DIN2(_26437), .Q(_40149) );
  hi1s1 _40658_inst ( .DIN(_40474), .Q(_40314) );
  nnd2s1 _40659_inst ( .DIN1(_26686), .DIN2(_26211), .Q(_40474) );
  nor2s1 _40660_inst ( .DIN1(_40444), .DIN2(_40355), .Q(_40479) );
  nnd2s1 _40661_inst ( .DIN1(_40476), .DIN2(_40254), .Q(_40355) );
  nor2s1 _40662_inst ( .DIN1(_40324), .DIN2(_26238), .Q(_40254) );
  nnd2s1 _40663_inst ( .DIN1(_53437), .DIN2(_26228), .Q(_40324) );
  nor2s1 _40664_inst ( .DIN1(_53439), .DIN2(_26286), .Q(_40476) );
  nnd2s1 _40665_inst ( .DIN1(_40480), .DIN2(_53436), .Q(_40444) );
  nor2s1 _40666_inst ( .DIN1(_53443), .DIN2(_26466), .Q(_40480) );
  hi1s1 _40667_inst ( .DIN(_27453), .Q(_27476) );
  nnd2s1 _40668_inst ( .DIN1(_29560), .DIN2(_38162), .Q(_27453) );
  hi1s1 _40669_inst ( .DIN(_29555), .Q(_29560) );
  nnd2s1 _40670_inst ( .DIN1(_27247), .DIN2(_33489), .Q(_29555) );
  hi1s1 _40671_inst ( .DIN(_31026), .Q(_27247) );
  nnd2s1 _40672_inst ( .DIN1(_40481), .DIN2(_35369), .Q(_31026) );
  nor2s1 _40673_inst ( .DIN1(_38165), .DIN2(_40482), .Q(_40481) );
  nnd2s1 _40674_inst ( .DIN1(_40483), .DIN2(_40484), .Q(
        ____2____________9_____) );
  nnd2s1 _40675_inst ( .DIN1(_40485), .DIN2(_53408), .Q(_40484) );
  nor2s1 _40676_inst ( .DIN1(_40486), .DIN2(_28684), .Q(_40485) );
  nnd2s1 _40677_inst ( .DIN1(_35940), .DIN2(_40487), .Q(_40483) );
  nnd2s1 _40678_inst ( .DIN1(_40488), .DIN2(_40489), .Q(_40487) );
  nor2s1 _40679_inst ( .DIN1(_40490), .DIN2(_40491), .Q(_40489) );
  nnd2s1 _40680_inst ( .DIN1(_40492), .DIN2(_40493), .Q(_40491) );
  nnd2s1 _40681_inst ( .DIN1(_40494), .DIN2(_40495), .Q(_40493) );
  nor2s1 _40682_inst ( .DIN1(_40496), .DIN2(_40497), .Q(_40492) );
  nor2s1 _40683_inst ( .DIN1(_40498), .DIN2(_40499), .Q(_40497) );
  nnd2s1 _40684_inst ( .DIN1(_40500), .DIN2(_40501), .Q(_40490) );
  hi1s1 _40685_inst ( .DIN(_40502), .Q(_40501) );
  nor2s1 _40686_inst ( .DIN1(_40503), .DIN2(_40504), .Q(_40500) );
  nor2s1 _40687_inst ( .DIN1(_40505), .DIN2(_40506), .Q(_40488) );
  or2s1 _40688_inst ( .DIN1(_40507), .DIN2(_40508), .Q(_40506) );
  nnd2s1 _40689_inst ( .DIN1(_40509), .DIN2(_40510), .Q(_40505) );
  nor2s1 _40690_inst ( .DIN1(_40511), .DIN2(_40512), .Q(_40509) );
  nnd2s1 _40691_inst ( .DIN1(_40513), .DIN2(_40514), .Q(
        ____2____________8_____) );
  nnd2s1 _40692_inst ( .DIN1(_40515), .DIN2(_40516), .Q(_40514) );
  nor2s1 _40693_inst ( .DIN1(_40517), .DIN2(_27066), .Q(_40515) );
  xor2s1 _40694_inst ( .DIN1(_40518), .DIN2(_53411), .Q(_40517) );
  nnd2s1 _40695_inst ( .DIN1(_40519), .DIN2(_40520), .Q(_40513) );
  nnd2s1 _40696_inst ( .DIN1(_40521), .DIN2(_40522), .Q(_40520) );
  nor2s1 _40697_inst ( .DIN1(_40523), .DIN2(_40524), .Q(_40522) );
  nnd2s1 _40698_inst ( .DIN1(_40525), .DIN2(_40526), .Q(_40524) );
  nor2s1 _40699_inst ( .DIN1(_40527), .DIN2(_40528), .Q(_40526) );
  nor2s1 _40700_inst ( .DIN1(_40529), .DIN2(_40499), .Q(_40528) );
  nor2s1 _40701_inst ( .DIN1(_40530), .DIN2(_40531), .Q(_40525) );
  nor2s1 _40702_inst ( .DIN1(_40532), .DIN2(_40533), .Q(_40530) );
  nnd2s1 _40703_inst ( .DIN1(_40534), .DIN2(_40535), .Q(_40523) );
  nor2s1 _40704_inst ( .DIN1(_40536), .DIN2(_40537), .Q(_40535) );
  nor2s1 _40705_inst ( .DIN1(_40538), .DIN2(_40498), .Q(_40537) );
  nor2s1 _40706_inst ( .DIN1(_40494), .DIN2(_40539), .Q(_40538) );
  hi1s1 _40707_inst ( .DIN(_40540), .Q(_40536) );
  nor2s1 _40708_inst ( .DIN1(_40541), .DIN2(_40542), .Q(_40534) );
  nor2s1 _40709_inst ( .DIN1(_40543), .DIN2(_40544), .Q(_40542) );
  and2s1 _40710_inst ( .DIN1(_40545), .DIN2(_40546), .Q(_40541) );
  nor2s1 _40711_inst ( .DIN1(_40547), .DIN2(_40548), .Q(_40521) );
  nnd2s1 _40712_inst ( .DIN1(_40549), .DIN2(_40550), .Q(_40548) );
  nor2s1 _40713_inst ( .DIN1(_40551), .DIN2(_40552), .Q(_40549) );
  nnd2s1 _40714_inst ( .DIN1(_40553), .DIN2(_40554), .Q(_40547) );
  nor2s1 _40715_inst ( .DIN1(_40555), .DIN2(_40556), .Q(_40554) );
  nor2s1 _40716_inst ( .DIN1(_40557), .DIN2(_40558), .Q(_40553) );
  nnd2s1 _40717_inst ( .DIN1(_40559), .DIN2(_40560), .Q(
        ____2____________7_____) );
  nor2s1 _40718_inst ( .DIN1(_40561), .DIN2(_40562), .Q(_40559) );
  nor2s1 _40719_inst ( .DIN1(_40563), .DIN2(_40564), .Q(_40562) );
  nnd2s1 _40720_inst ( .DIN1(_40565), .DIN2(_40566), .Q(_40564) );
  nor2s1 _40721_inst ( .DIN1(_40567), .DIN2(_40568), .Q(_40566) );
  nnd2s1 _40722_inst ( .DIN1(_40569), .DIN2(_40570), .Q(_40568) );
  nor2s1 _40723_inst ( .DIN1(_40571), .DIN2(_40572), .Q(_40570) );
  nor2s1 _40724_inst ( .DIN1(_40573), .DIN2(_40574), .Q(_40572) );
  nor2s1 _40725_inst ( .DIN1(_40575), .DIN2(_40576), .Q(_40571) );
  nor2s1 _40726_inst ( .DIN1(_40577), .DIN2(_40578), .Q(_40569) );
  nor2s1 _40727_inst ( .DIN1(_40579), .DIN2(_40580), .Q(_40578) );
  nor2s1 _40728_inst ( .DIN1(_26842), .DIN2(_40582), .Q(_40577) );
  nnd2s1 _40729_inst ( .DIN1(_40583), .DIN2(_40584), .Q(_40567) );
  nor2s1 _40730_inst ( .DIN1(_40585), .DIN2(_40586), .Q(_40584) );
  and2s1 _40731_inst ( .DIN1(_40587), .DIN2(_40588), .Q(_40583) );
  nor2s1 _40732_inst ( .DIN1(_40589), .DIN2(_40590), .Q(_40565) );
  nnd2s1 _40733_inst ( .DIN1(_40591), .DIN2(_40592), .Q(_40590) );
  nor2s1 _40734_inst ( .DIN1(_40593), .DIN2(_40594), .Q(_40592) );
  nor2s1 _40735_inst ( .DIN1(_40595), .DIN2(_40596), .Q(_40591) );
  nnd2s1 _40736_inst ( .DIN1(_40597), .DIN2(_40598), .Q(_40589) );
  nor2s1 _40737_inst ( .DIN1(_40512), .DIN2(_40599), .Q(_40598) );
  nnd2s1 _40738_inst ( .DIN1(_40600), .DIN2(_40601), .Q(_40512) );
  nor2s1 _40739_inst ( .DIN1(_40602), .DIN2(_40603), .Q(_40601) );
  nnd2s1 _40740_inst ( .DIN1(_40604), .DIN2(_40605), .Q(_40603) );
  hi1s1 _40741_inst ( .DIN(_40606), .Q(_40605) );
  nnd2s1 _40742_inst ( .DIN1(_40607), .DIN2(_40608), .Q(_40604) );
  nor2s1 _40743_inst ( .DIN1(_40609), .DIN2(_40610), .Q(_40600) );
  nor2s1 _40744_inst ( .DIN1(_40558), .DIN2(_40611), .Q(_40597) );
  nnd2s1 _40745_inst ( .DIN1(_40612), .DIN2(_40613), .Q(_40558) );
  nor2s1 _40746_inst ( .DIN1(_40614), .DIN2(_40615), .Q(_40613) );
  nnd2s1 _40747_inst ( .DIN1(_40616), .DIN2(_40617), .Q(_40615) );
  nnd2s1 _40748_inst ( .DIN1(_40618), .DIN2(_40619), .Q(_40614) );
  nor2s1 _40749_inst ( .DIN1(_40620), .DIN2(_40621), .Q(_40612) );
  or2s1 _40750_inst ( .DIN1(_40622), .DIN2(_40623), .Q(_40621) );
  nor2s1 _40751_inst ( .DIN1(_40519), .DIN2(_40624), .Q(_40561) );
  nor2s1 _40752_inst ( .DIN1(_26988), .DIN2(_40625), .Q(_40624) );
  nnd2s1 _40753_inst ( .DIN1(_40626), .DIN2(_40518), .Q(_40625) );
  nnd2s1 _40754_inst ( .DIN1(_26208), .DIN2(_26443), .Q(_40626) );
  nnd2s1 _40755_inst ( .DIN1(_40627), .DIN2(_40628), .Q(
        ____2____________6_____) );
  nnd2s1 _40756_inst ( .DIN1(_40629), .DIN2(_40516), .Q(_40628) );
  nor2s1 _40757_inst ( .DIN1(_40630), .DIN2(_27448), .Q(_40629) );
  xor2s1 _40758_inst ( .DIN1(_40518), .DIN2(_53400), .Q(_40630) );
  nnd2s1 _40759_inst ( .DIN1(_40519), .DIN2(_40631), .Q(_40627) );
  nnd2s1 _40760_inst ( .DIN1(_40632), .DIN2(_40633), .Q(_40631) );
  nor2s1 _40761_inst ( .DIN1(_40634), .DIN2(_40635), .Q(_40633) );
  nnd2s1 _40762_inst ( .DIN1(_40636), .DIN2(_40637), .Q(_40635) );
  nnd2s1 _40763_inst ( .DIN1(_40638), .DIN2(_40639), .Q(_40637) );
  nor2s1 _40764_inst ( .DIN1(_40640), .DIN2(_40641), .Q(_40636) );
  nor2s1 _40765_inst ( .DIN1(_40642), .DIN2(_40532), .Q(_40641) );
  nor2s1 _40766_inst ( .DIN1(_40498), .DIN2(_40643), .Q(_40640) );
  nnd2s1 _40767_inst ( .DIN1(_40644), .DIN2(_40645), .Q(_40634) );
  nor2s1 _40768_inst ( .DIN1(_40646), .DIN2(_40647), .Q(_40645) );
  nor2s1 _40769_inst ( .DIN1(_40648), .DIN2(_40649), .Q(_40647) );
  nor2s1 _40770_inst ( .DIN1(_40650), .DIN2(_40651), .Q(_40644) );
  nor2s1 _40771_inst ( .DIN1(_40652), .DIN2(_40653), .Q(_40651) );
  nor2s1 _40772_inst ( .DIN1(_40654), .DIN2(_40655), .Q(_40650) );
  nor2s1 _40773_inst ( .DIN1(_40656), .DIN2(_40657), .Q(_40632) );
  nnd2s1 _40774_inst ( .DIN1(_40658), .DIN2(_40659), .Q(_40657) );
  nor2s1 _40775_inst ( .DIN1(_40660), .DIN2(_40661), .Q(_40658) );
  nnd2s1 _40776_inst ( .DIN1(_40662), .DIN2(_40663), .Q(_40656) );
  hi1s1 _40777_inst ( .DIN(_40611), .Q(_40663) );
  nnd2s1 _40778_inst ( .DIN1(_40664), .DIN2(_40665), .Q(_40611) );
  nor2s1 _40779_inst ( .DIN1(_40666), .DIN2(_40667), .Q(_40665) );
  nnd2s1 _40780_inst ( .DIN1(_40668), .DIN2(_40669), .Q(_40667) );
  nnd2s1 _40781_inst ( .DIN1(_40670), .DIN2(_40671), .Q(_40666) );
  nor2s1 _40782_inst ( .DIN1(_40502), .DIN2(_40672), .Q(_40670) );
  nor2s1 _40783_inst ( .DIN1(_40673), .DIN2(_40674), .Q(_40664) );
  or2s1 _40784_inst ( .DIN1(_40675), .DIN2(_40676), .Q(_40674) );
  nnd2s1 _40785_inst ( .DIN1(_40677), .DIN2(_40678), .Q(_40673) );
  hi1s1 _40786_inst ( .DIN(_40679), .Q(_40678) );
  and2s1 _40787_inst ( .DIN1(_40680), .DIN2(_40681), .Q(_40677) );
  nor2s1 _40788_inst ( .DIN1(_40682), .DIN2(_40683), .Q(_40662) );
  xor2s1 _40789_inst ( .DIN1(_40684), .DIN2(_40046), .Q(_40683) );
  hi1s1 _40790_inst ( .DIN(_31768), .Q(_40046) );
  nnd2s1 _40791_inst ( .DIN1(_40685), .DIN2(_40686), .Q(_40684) );
  nnd2s1 _40792_inst ( .DIN1(_40687), .DIN2(_29686), .Q(
        ____2____________5_____) );
  nnd2s1 _40793_inst ( .DIN1(_29689), .DIN2(_31291), .Q(_29686) );
  nor2s1 _40794_inst ( .DIN1(_40688), .DIN2(_40689), .Q(_40687) );
  nor2s1 _40795_inst ( .DIN1(_29689), .DIN2(_40690), .Q(_40689) );
  nnd2s1 _40796_inst ( .DIN1(_40691), .DIN2(_40692), .Q(_40690) );
  nor2s1 _40797_inst ( .DIN1(_40693), .DIN2(_40694), .Q(_40692) );
  nnd2s1 _40798_inst ( .DIN1(_40695), .DIN2(_40696), .Q(_40694) );
  nor2s1 _40799_inst ( .DIN1(_40697), .DIN2(_40698), .Q(_40696) );
  nor2s1 _40800_inst ( .DIN1(_40699), .DIN2(_40700), .Q(_40697) );
  nor2s1 _40801_inst ( .DIN1(_40701), .DIN2(_40702), .Q(_40695) );
  hi1s1 _40802_inst ( .DIN(_40703), .Q(_40702) );
  xor2s1 _40803_inst ( .DIN1(_40704), .DIN2(_36757), .Q(_40701) );
  nnd2s1 _40804_inst ( .DIN1(_40705), .DIN2(_40706), .Q(_40693) );
  nor2s1 _40805_inst ( .DIN1(_40707), .DIN2(_40708), .Q(_40706) );
  hi1s1 _40806_inst ( .DIN(_40709), .Q(_40708) );
  nor2s1 _40807_inst ( .DIN1(_40710), .DIN2(_40711), .Q(_40705) );
  nor2s1 _40808_inst ( .DIN1(_40498), .DIN2(_40574), .Q(_40711) );
  nor2s1 _40809_inst ( .DIN1(_40712), .DIN2(_40713), .Q(_40691) );
  nnd2s1 _40810_inst ( .DIN1(_40714), .DIN2(_40715), .Q(_40713) );
  hi1s1 _40811_inst ( .DIN(_40716), .Q(_40715) );
  nor2s1 _40812_inst ( .DIN1(_40717), .DIN2(_40718), .Q(_40714) );
  nnd2s1 _40813_inst ( .DIN1(_40719), .DIN2(_40720), .Q(_40712) );
  nor2s1 _40814_inst ( .DIN1(_40721), .DIN2(_40722), .Q(_40720) );
  nor2s1 _40815_inst ( .DIN1(_40723), .DIN2(_40724), .Q(_40719) );
  nor2s1 _40816_inst ( .DIN1(_27154), .DIN2(_40725), .Q(_40688) );
  nor2s1 _40817_inst ( .DIN1(_40726), .DIN2(_40727), .Q(_40725) );
  nnd2s1 _40818_inst ( .DIN1(_40728), .DIN2(_40729), .Q(_40727) );
  nnd2s1 _40819_inst ( .DIN1(_31292), .DIN2(_26564), .Q(_40729) );
  nor2s1 _40820_inst ( .DIN1(_26440), .DIN2(_26239), .Q(_31292) );
  nnd2s1 _40821_inst ( .DIN1(_53393), .DIN2(_26440), .Q(_40728) );
  nor2s1 _40822_inst ( .DIN1(_53394), .DIN2(_53395), .Q(_40726) );
  hi1s1 _40823_inst ( .DIN(_29689), .Q(_27154) );
  nnd2s1 _40824_inst ( .DIN1(_40730), .DIN2(_40731), .Q(_29689) );
  nor2s1 _40825_inst ( .DIN1(_27161), .DIN2(_40732), .Q(_40730) );
  hi1s1 _40826_inst ( .DIN(_31291), .Q(_27161) );
  nnd2s1 _40827_inst ( .DIN1(_40733), .DIN2(_40734), .Q(
        ____2____________4_____) );
  nnd2s1 _40828_inst ( .DIN1(_29390), .DIN2(_40735), .Q(_40734) );
  xor2s1 _40829_inst ( .DIN1(_52850), .DIN2(_53396), .Q(_40735) );
  nor2s1 _40830_inst ( .DIN1(_28250), .DIN2(_38919), .Q(_29390) );
  nnd2s1 _40831_inst ( .DIN1(_28250), .DIN2(_40736), .Q(_40733) );
  nnd2s1 _40832_inst ( .DIN1(_40737), .DIN2(_40738), .Q(_40736) );
  nor2s1 _40833_inst ( .DIN1(_40739), .DIN2(_40740), .Q(_40738) );
  nnd2s1 _40834_inst ( .DIN1(_40741), .DIN2(_40742), .Q(_40740) );
  nor2s1 _40835_inst ( .DIN1(_40743), .DIN2(_40744), .Q(_40742) );
  nor2s1 _40836_inst ( .DIN1(_40745), .DIN2(_40700), .Q(_40744) );
  nor2s1 _40837_inst ( .DIN1(_40602), .DIN2(_40746), .Q(_40741) );
  nor2s1 _40838_inst ( .DIN1(_40498), .DIN2(_40747), .Q(_40746) );
  nor2s1 _40839_inst ( .DIN1(_40544), .DIN2(_40748), .Q(_40602) );
  nnd2s1 _40840_inst ( .DIN1(_40749), .DIN2(_40750), .Q(_40739) );
  nor2s1 _40841_inst ( .DIN1(_40751), .DIN2(_40752), .Q(_40750) );
  hi1s1 _40842_inst ( .DIN(_40671), .Q(_40752) );
  nnd2s1 _40843_inst ( .DIN1(_40753), .DIN2(_40754), .Q(_40671) );
  nnd2s1 _40844_inst ( .DIN1(_40755), .DIN2(_40756), .Q(_40753) );
  nor2s1 _40845_inst ( .DIN1(_40757), .DIN2(_40646), .Q(_40749) );
  nor2s1 _40846_inst ( .DIN1(_40758), .DIN2(_40759), .Q(_40737) );
  nnd2s1 _40847_inst ( .DIN1(_40760), .DIN2(_40761), .Q(_40759) );
  nor2s1 _40848_inst ( .DIN1(_40594), .DIN2(_40762), .Q(_40761) );
  nnd2s1 _40849_inst ( .DIN1(_40763), .DIN2(_40764), .Q(_40594) );
  or2s1 _40850_inst ( .DIN1(_40765), .DIN2(_40573), .Q(_40764) );
  nor2s1 _40851_inst ( .DIN1(_40766), .DIN2(_40767), .Q(_40763) );
  nor2s1 _40852_inst ( .DIN1(_26842), .DIN2(_40768), .Q(_40767) );
  nor2s1 _40853_inst ( .DIN1(_40769), .DIN2(_40770), .Q(_40768) );
  nor2s1 _40854_inst ( .DIN1(_40771), .DIN2(_40772), .Q(_40760) );
  hi1s1 _40855_inst ( .DIN(_40773), .Q(_40771) );
  nnd2s1 _40856_inst ( .DIN1(_40774), .DIN2(_40775), .Q(_40758) );
  nor2s1 _40857_inst ( .DIN1(_40511), .DIN2(_40776), .Q(_40775) );
  nor2s1 _40858_inst ( .DIN1(_40777), .DIN2(_40778), .Q(_40776) );
  nor2s1 _40859_inst ( .DIN1(_40654), .DIN2(_40582), .Q(_40511) );
  nor2s1 _40860_inst ( .DIN1(_40779), .DIN2(_40623), .Q(_40774) );
  nnd2s1 _40861_inst ( .DIN1(_40780), .DIN2(_40781), .Q(_40623) );
  nnd2s1 _40862_inst ( .DIN1(_40782), .DIN2(_40783), .Q(_40781) );
  nor2s1 _40863_inst ( .DIN1(_40784), .DIN2(_40710), .Q(_40780) );
  hi1s1 _40864_inst ( .DIN(_28241), .Q(_28250) );
  nnd2s1 _40865_inst ( .DIN1(_40785), .DIN2(_40786), .Q(_28241) );
  nor2s1 _40866_inst ( .DIN1(_40732), .DIN2(_37418), .Q(_40785) );
  nnd2s1 _40867_inst ( .DIN1(_40787), .DIN2(_28026), .Q(
        ____2____________3_____) );
  nnd2s1 _40868_inst ( .DIN1(_40786), .DIN2(_28016), .Q(_28026) );
  nor2s1 _40869_inst ( .DIN1(_40788), .DIN2(_40789), .Q(_40787) );
  nor2s1 _40870_inst ( .DIN1(_28016), .DIN2(_40790), .Q(_40789) );
  nnd2s1 _40871_inst ( .DIN1(_40791), .DIN2(_40792), .Q(_40790) );
  nor2s1 _40872_inst ( .DIN1(_40793), .DIN2(_40794), .Q(_40792) );
  nnd2s1 _40873_inst ( .DIN1(_40795), .DIN2(_40510), .Q(_40794) );
  and2s1 _40874_inst ( .DIN1(_40796), .DIN2(_40797), .Q(_40510) );
  nor2s1 _40875_inst ( .DIN1(_40798), .DIN2(_40799), .Q(_40797) );
  nnd2s1 _40876_inst ( .DIN1(_40680), .DIN2(_40800), .Q(_40799) );
  nnd2s1 _40877_inst ( .DIN1(_40801), .DIN2(_40686), .Q(_40680) );
  nor2s1 _40878_inst ( .DIN1(_40802), .DIN2(_40529), .Q(_40798) );
  nor2s1 _40879_inst ( .DIN1(_40782), .DIN2(_40803), .Q(_40802) );
  nor2s1 _40880_inst ( .DIN1(_40804), .DIN2(_40805), .Q(_40796) );
  and2s1 _40881_inst ( .DIN1(_40608), .DIN2(_40806), .Q(_40804) );
  nor2s1 _40882_inst ( .DIN1(_40807), .DIN2(_40808), .Q(_40795) );
  hi1s1 _40883_inst ( .DIN(_40809), .Q(_40808) );
  nor2s1 _40884_inst ( .DIN1(_40649), .DIN2(_40810), .Q(_40807) );
  nnd2s1 _40885_inst ( .DIN1(_40811), .DIN2(_40812), .Q(_40793) );
  nor2s1 _40886_inst ( .DIN1(_40813), .DIN2(_40814), .Q(_40812) );
  hi1s1 _40887_inst ( .DIN(_40815), .Q(_40813) );
  nor2s1 _40888_inst ( .DIN1(_40816), .DIN2(_40817), .Q(_40811) );
  nor2s1 _40889_inst ( .DIN1(_40818), .DIN2(_40819), .Q(_40817) );
  nor2s1 _40890_inst ( .DIN1(_40820), .DIN2(_40529), .Q(_40816) );
  nor2s1 _40891_inst ( .DIN1(_40769), .DIN2(_40821), .Q(_40820) );
  hi1s1 _40892_inst ( .DIN(_40499), .Q(_40769) );
  nor2s1 _40893_inst ( .DIN1(_40822), .DIN2(_40823), .Q(_40791) );
  nnd2s1 _40894_inst ( .DIN1(_40824), .DIN2(_40825), .Q(_40823) );
  hi1s1 _40895_inst ( .DIN(_40826), .Q(_40825) );
  nor2s1 _40896_inst ( .DIN1(_40827), .DIN2(_40762), .Q(_40824) );
  nnd2s1 _40897_inst ( .DIN1(_40828), .DIN2(_40829), .Q(_40762) );
  nor2s1 _40898_inst ( .DIN1(_40830), .DIN2(_40831), .Q(_40829) );
  nnd2s1 _40899_inst ( .DIN1(_40832), .DIN2(_40833), .Q(_40831) );
  nnd2s1 _40900_inst ( .DIN1(_40834), .DIN2(_40835), .Q(_40833) );
  nnd2s1 _40901_inst ( .DIN1(_40836), .DIN2(_40837), .Q(_40830) );
  nor2s1 _40902_inst ( .DIN1(_40838), .DIN2(_40527), .Q(_40836) );
  nor2s1 _40903_inst ( .DIN1(_40818), .DIN2(_40839), .Q(_40527) );
  nor2s1 _40904_inst ( .DIN1(_40840), .DIN2(_40841), .Q(_40828) );
  nnd2s1 _40905_inst ( .DIN1(_40842), .DIN2(_40843), .Q(_40841) );
  hi1s1 _40906_inst ( .DIN(_40724), .Q(_40843) );
  nnd2s1 _40907_inst ( .DIN1(_40844), .DIN2(_40845), .Q(_40724) );
  nnd2s1 _40908_inst ( .DIN1(_40539), .DIN2(_40495), .Q(_40845) );
  hi1s1 _40909_inst ( .DIN(_40643), .Q(_40539) );
  nor2s1 _40910_inst ( .DIN1(_40846), .DIN2(_40847), .Q(_40844) );
  nor2s1 _40911_inst ( .DIN1(_26842), .DIN2(_40848), .Q(_40847) );
  nor2s1 _40912_inst ( .DIN1(_40849), .DIN2(_40850), .Q(_40846) );
  nnd2s1 _40913_inst ( .DIN1(_40851), .DIN2(_40852), .Q(_40840) );
  nor2s1 _40914_inst ( .DIN1(_40622), .DIN2(_40593), .Q(_40851) );
  nnd2s1 _40915_inst ( .DIN1(_40853), .DIN2(_40854), .Q(_40593) );
  nnd2s1 _40916_inst ( .DIN1(_40855), .DIN2(_40856), .Q(_40854) );
  nor2s1 _40917_inst ( .DIN1(_34893), .DIN2(_40857), .Q(_40855) );
  nnd2s1 _40918_inst ( .DIN1(_40858), .DIN2(_40859), .Q(_40822) );
  nor2s1 _40919_inst ( .DIN1(_40860), .DIN2(_40861), .Q(_40859) );
  nor2s1 _40920_inst ( .DIN1(_40596), .DIN2(_40862), .Q(_40858) );
  nor2s1 _40921_inst ( .DIN1(_28024), .DIN2(_40863), .Q(_40788) );
  nor2s1 _40922_inst ( .DIN1(_27291), .DIN2(_26356), .Q(_40863) );
  hi1s1 _40923_inst ( .DIN(_28016), .Q(_28024) );
  nnd2s1 _40924_inst ( .DIN1(_40864), .DIN2(_40786), .Q(_28016) );
  and2s1 _40925_inst ( .DIN1(_40865), .DIN2(_40866), .Q(_40786) );
  nor2s1 _40926_inst ( .DIN1(_37417), .DIN2(_40867), .Q(_40865) );
  nor2s1 _40927_inst ( .DIN1(_40732), .DIN2(_40868), .Q(_40864) );
  nor2s1 _40928_inst ( .DIN1(_40869), .DIN2(_27235), .Q(
        ____2____________2_____) );
  nor2s1 _40929_inst ( .DIN1(_40870), .DIN2(_40871), .Q(_40869) );
  nnd2s1 _40930_inst ( .DIN1(_40872), .DIN2(_40873), .Q(_40871) );
  nor2s1 _40931_inst ( .DIN1(_40874), .DIN2(_40875), .Q(_40873) );
  or2s1 _40932_inst ( .DIN1(_40660), .DIN2(_40531), .Q(_40875) );
  nnd2s1 _40933_inst ( .DIN1(_40703), .DIN2(_40876), .Q(_40531) );
  xor2s1 _40934_inst ( .DIN1(_31569), .DIN2(_40877), .Q(_40703) );
  nor2s1 _40935_inst ( .DIN1(_40878), .DIN2(_40672), .Q(_40877) );
  nor2s1 _40936_inst ( .DIN1(_40879), .DIN2(_40498), .Q(_40672) );
  nnd2s1 _40937_inst ( .DIN1(_40880), .DIN2(_40881), .Q(_40660) );
  nor2s1 _40938_inst ( .DIN1(_40882), .DIN2(_40883), .Q(_40881) );
  nnd2s1 _40939_inst ( .DIN1(_40884), .DIN2(_40885), .Q(_40883) );
  nnd2s1 _40940_inst ( .DIN1(_40886), .DIN2(_40887), .Q(_40885) );
  nnd2s1 _40941_inst ( .DIN1(_40888), .DIN2(_40889), .Q(_40884) );
  nor2s1 _40942_inst ( .DIN1(_40722), .DIN2(_40862), .Q(_40880) );
  nnd2s1 _40943_inst ( .DIN1(_40890), .DIN2(_40891), .Q(_40862) );
  xor2s1 _40944_inst ( .DIN1(_29579), .DIN2(_40892), .Q(_40891) );
  nnd2s1 _40945_inst ( .DIN1(_40893), .DIN2(_40894), .Q(_40892) );
  nor2s1 _40946_inst ( .DIN1(_40895), .DIN2(_40896), .Q(_40893) );
  nor2s1 _40947_inst ( .DIN1(_40897), .DIN2(_40898), .Q(_40890) );
  nnd2s1 _40948_inst ( .DIN1(_40899), .DIN2(_40900), .Q(_40722) );
  nnd2s1 _40949_inst ( .DIN1(_40901), .DIN2(_40902), .Q(_40900) );
  nor2s1 _40950_inst ( .DIN1(_40654), .DIN2(_40903), .Q(_40901) );
  nor2s1 _40951_inst ( .DIN1(_40904), .DIN2(_40905), .Q(_40872) );
  nnd2s1 _40952_inst ( .DIN1(_40906), .DIN2(_40907), .Q(_40870) );
  nor2s1 _40953_inst ( .DIN1(_40908), .DIN2(_40909), .Q(_40907) );
  nnd2s1 _40954_inst ( .DIN1(_40910), .DIN2(_40911), .Q(_40909) );
  nnd2s1 _40955_inst ( .DIN1(_40782), .DIN2(_40495), .Q(_40911) );
  hi1s1 _40956_inst ( .DIN(_40912), .Q(_40782) );
  nor2s1 _40957_inst ( .DIN1(_40745), .DIN2(_40913), .Q(_40908) );
  nor2s1 _40958_inst ( .DIN1(_40914), .DIN2(_40915), .Q(_40906) );
  nnd2s1 _40959_inst ( .DIN1(_40916), .DIN2(_40917), .Q(_40915) );
  hi1s1 _40960_inst ( .DIN(_40918), .Q(_40917) );
  nnd2s1 _40961_inst ( .DIN1(_40919), .DIN2(_40920), .Q(
        ____2____________1_____) );
  nnd2s1 _40962_inst ( .DIN1(_40921), .DIN2(_35502), .Q(_40920) );
  nnd2s1 _40963_inst ( .DIN1(_40922), .DIN2(_35501), .Q(_40921) );
  xor2s1 _40964_inst ( .DIN1(_40923), .DIN2(_40924), .Q(_40922) );
  and2s1 _40965_inst ( .DIN1(_26218), .DIN2(_52847), .Q(_40924) );
  xor2s1 _40966_inst ( .DIN1(_26469), .DIN2(_53156), .Q(_40923) );
  nnd2s1 _40967_inst ( .DIN1(_40925), .DIN2(_27895), .Q(_40919) );
  nor2s1 _40968_inst ( .DIN1(_40926), .DIN2(_40927), .Q(_40925) );
  nnd2s1 _40969_inst ( .DIN1(_40928), .DIN2(_40929), .Q(_40927) );
  nor2s1 _40970_inst ( .DIN1(_40930), .DIN2(_40931), .Q(_40929) );
  nnd2s1 _40971_inst ( .DIN1(_40899), .DIN2(_40932), .Q(_40931) );
  hi1s1 _40972_inst ( .DIN(_40933), .Q(_40899) );
  or2s1 _40973_inst ( .DIN1(_40557), .DIN2(_40609), .Q(_40930) );
  nnd2s1 _40974_inst ( .DIN1(_40934), .DIN2(_40935), .Q(_40609) );
  nnd2s1 _40975_inst ( .DIN1(_40936), .DIN2(_40937), .Q(_40935) );
  nnd2s1 _40976_inst ( .DIN1(_40889), .DIN2(_40938), .Q(_40934) );
  or2s1 _40977_inst ( .DIN1(_40939), .DIN2(_40940), .Q(_40557) );
  or2s1 _40978_inst ( .DIN1(_40504), .DIN2(_40941), .Q(_40939) );
  nor2s1 _40979_inst ( .DIN1(_40942), .DIN2(_40896), .Q(_40941) );
  nor2s1 _40980_inst ( .DIN1(_40943), .DIN2(_40944), .Q(_40928) );
  or2s1 _40981_inst ( .DIN1(_40945), .DIN2(_40874), .Q(_40944) );
  nnd2s1 _40982_inst ( .DIN1(_40946), .DIN2(_40947), .Q(_40874) );
  nor2s1 _40983_inst ( .DIN1(_40948), .DIN2(_40949), .Q(_40947) );
  nnd2s1 _40984_inst ( .DIN1(_40950), .DIN2(_40587), .Q(_40949) );
  nor2s1 _40985_inst ( .DIN1(_40814), .DIN2(_40710), .Q(_40950) );
  nor2s1 _40986_inst ( .DIN1(_40951), .DIN2(_26842), .Q(_40710) );
  nnd2s1 _40987_inst ( .DIN1(_40952), .DIN2(_40953), .Q(_40948) );
  nor2s1 _40988_inst ( .DIN1(_40954), .DIN2(_40585), .Q(_40953) );
  hi1s1 _40989_inst ( .DIN(_40955), .Q(_40954) );
  nor2s1 _40990_inst ( .DIN1(_40956), .DIN2(_40957), .Q(_40952) );
  nor2s1 _40991_inst ( .DIN1(_40958), .DIN2(_40959), .Q(_40946) );
  nnd2s1 _40992_inst ( .DIN1(_40960), .DIN2(_40773), .Q(_40959) );
  nor2s1 _40993_inst ( .DIN1(_40961), .DIN2(_40551), .Q(_40773) );
  nnd2s1 _40994_inst ( .DIN1(_40962), .DIN2(_40963), .Q(_40551) );
  nor2s1 _40995_inst ( .DIN1(_40707), .DIN2(_40964), .Q(_40963) );
  nor2s1 _40996_inst ( .DIN1(_40965), .DIN2(_40966), .Q(_40964) );
  and2s1 _40997_inst ( .DIN1(_40967), .DIN2(_40754), .Q(_40707) );
  nor2s1 _40998_inst ( .DIN1(_40968), .DIN2(_40969), .Q(_40962) );
  nor2s1 _40999_inst ( .DIN1(_40579), .DIN2(_40970), .Q(_40968) );
  nor2s1 _41000_inst ( .DIN1(_40971), .DIN2(_40972), .Q(_40579) );
  or2s1 _41001_inst ( .DIN1(_40502), .DIN2(_40973), .Q(_40961) );
  nor2s1 _41002_inst ( .DIN1(_40777), .DIN2(_40974), .Q(_40973) );
  nor2s1 _41003_inst ( .DIN1(_40529), .DIN2(_40975), .Q(_40502) );
  nor2s1 _41004_inst ( .DIN1(_40976), .DIN2(_40599), .Q(_40960) );
  nnd2s1 _41005_inst ( .DIN1(_40977), .DIN2(_40978), .Q(_40958) );
  nor2s1 _41006_inst ( .DIN1(_40766), .DIN2(_40979), .Q(_40978) );
  nor2s1 _41007_inst ( .DIN1(_40850), .DIN2(_40756), .Q(_40979) );
  hi1s1 _41008_inst ( .DIN(_40980), .Q(_40766) );
  nor2s1 _41009_inst ( .DIN1(_40981), .DIN2(_40982), .Q(_40977) );
  nnd2s1 _41010_inst ( .DIN1(_40983), .DIN2(_40984), .Q(_40926) );
  nor2s1 _41011_inst ( .DIN1(_40985), .DIN2(_40986), .Q(_40984) );
  nnd2s1 _41012_inst ( .DIN1(_40987), .DIN2(_40988), .Q(_40986) );
  nnd2s1 _41013_inst ( .DIN1(_40989), .DIN2(_40990), .Q(_40988) );
  xor2s1 _41014_inst ( .DIN1(_40991), .DIN2(_40992), .Q(_40990) );
  nor2s1 _41015_inst ( .DIN1(_40993), .DIN2(_40994), .Q(_40992) );
  nnd2s1 _41016_inst ( .DIN1(_40995), .DIN2(_40937), .Q(_40987) );
  nnd2s1 _41017_inst ( .DIN1(_40617), .DIN2(_40709), .Q(_40985) );
  nor2s1 _41018_inst ( .DIN1(_40996), .DIN2(_40997), .Q(_40983) );
  nnd2s1 _41019_inst ( .DIN1(_40998), .DIN2(_40999), .Q(_40997) );
  nnd2s1 _41020_inst ( .DIN1(_41000), .DIN2(_41001), .Q(_40999) );
  nnd2s1 _41021_inst ( .DIN1(_40801), .DIN2(_41002), .Q(_40998) );
  nnd2s1 _41022_inst ( .DIN1(_41003), .DIN2(_41004), .Q(
        ____2____________13_____) );
  nnd2s1 _41023_inst ( .DIN1(_41005), .DIN2(_35938), .Q(_41004) );
  xor2s1 _41024_inst ( .DIN1(_53406), .DIN2(_53408), .Q(_41005) );
  nnd2s1 _41025_inst ( .DIN1(_35940), .DIN2(_41006), .Q(_41003) );
  nnd2s1 _41026_inst ( .DIN1(_41007), .DIN2(_41008), .Q(_41006) );
  nor2s1 _41027_inst ( .DIN1(_41009), .DIN2(_41010), .Q(_41008) );
  nnd2s1 _41028_inst ( .DIN1(_41011), .DIN2(_41012), .Q(_41010) );
  nor2s1 _41029_inst ( .DIN1(_41013), .DIN2(_40969), .Q(_41012) );
  nor2s1 _41030_inst ( .DIN1(_40498), .DIN2(_41014), .Q(_40969) );
  nor2s1 _41031_inst ( .DIN1(_40573), .DIN2(_40879), .Q(_41013) );
  nor2s1 _41032_inst ( .DIN1(_41015), .DIN2(_41016), .Q(_41011) );
  nor2s1 _41033_inst ( .DIN1(_26842), .DIN2(_40643), .Q(_41015) );
  nnd2s1 _41034_inst ( .DIN1(_41017), .DIN2(_41018), .Q(_41009) );
  nor2s1 _41035_inst ( .DIN1(_41019), .DIN2(_40757), .Q(_41018) );
  hi1s1 _41036_inst ( .DIN(_40669), .Q(_41019) );
  nnd2s1 _41037_inst ( .DIN1(_40967), .DIN2(_40546), .Q(_40669) );
  nor2s1 _41038_inst ( .DIN1(_41020), .DIN2(_40981), .Q(_41017) );
  nor2s1 _41039_inst ( .DIN1(_40896), .DIN2(_41021), .Q(_40981) );
  nor2s1 _41040_inst ( .DIN1(_41022), .DIN2(_41023), .Q(_41007) );
  nnd2s1 _41041_inst ( .DIN1(_41024), .DIN2(_41025), .Q(_41023) );
  xor2s1 _41042_inst ( .DIN1(_41026), .DIN2(_32548), .Q(_41025) );
  nor2s1 _41043_inst ( .DIN1(_40661), .DIN2(_40716), .Q(_41024) );
  nnd2s1 _41044_inst ( .DIN1(_41027), .DIN2(_41028), .Q(_40716) );
  nor2s1 _41045_inst ( .DIN1(_41029), .DIN2(_41030), .Q(_41028) );
  nnd2s1 _41046_inst ( .DIN1(_41031), .DIN2(_41032), .Q(_41030) );
  or2s1 _41047_inst ( .DIN1(_40819), .DIN2(_40818), .Q(_41031) );
  hi1s1 _41048_inst ( .DIN(_41033), .Q(_40818) );
  nnd2s1 _41049_inst ( .DIN1(_41034), .DIN2(_41035), .Q(_41029) );
  hi1s1 _41050_inst ( .DIN(_41036), .Q(_41035) );
  nor2s1 _41051_inst ( .DIN1(_40751), .DIN2(_40957), .Q(_41034) );
  and2s1 _41052_inst ( .DIN1(_41037), .DIN2(_40608), .Q(_40957) );
  nor2s1 _41053_inst ( .DIN1(_41038), .DIN2(_41039), .Q(_41027) );
  nnd2s1 _41054_inst ( .DIN1(_41040), .DIN2(_41041), .Q(_41039) );
  hi1s1 _41055_inst ( .DIN(_41042), .Q(_41041) );
  xor2s1 _41056_inst ( .DIN1(_41043), .DIN2(_41044), .Q(_41040) );
  nor2s1 _41057_inst ( .DIN1(_41045), .DIN2(_41046), .Q(_41044) );
  or2s1 _41058_inst ( .DIN1(_40552), .DIN2(_41047), .Q(_41046) );
  nnd2s1 _41059_inst ( .DIN1(_41048), .DIN2(_41049), .Q(_40552) );
  or2s1 _41060_inst ( .DIN1(_40756), .DIN2(_26842), .Q(_41049) );
  nor2s1 _41061_inst ( .DIN1(_41050), .DIN2(_40814), .Q(_41048) );
  and2s1 _41062_inst ( .DIN1(_41051), .DIN2(_40972), .Q(_40814) );
  nnd2s1 _41063_inst ( .DIN1(_41052), .DIN2(_40852), .Q(_41038) );
  and2s1 _41064_inst ( .DIN1(_41053), .DIN2(_41054), .Q(_40852) );
  nnd2s1 _41065_inst ( .DIN1(_41055), .DIN2(_41056), .Q(_41054) );
  nor2s1 _41066_inst ( .DIN1(_41057), .DIN2(_41058), .Q(_41053) );
  nor2s1 _41067_inst ( .DIN1(_26842), .DIN2(_40533), .Q(_41058) );
  nor2s1 _41068_inst ( .DIN1(_41059), .DIN2(_40653), .Q(_41057) );
  nor2s1 _41069_inst ( .DIN1(_41060), .DIN2(_41061), .Q(_41052) );
  nor2s1 _41070_inst ( .DIN1(_41062), .DIN2(_41063), .Q(_41060) );
  nnd2s1 _41071_inst ( .DIN1(_41064), .DIN2(_41065), .Q(_40661) );
  nor2s1 _41072_inst ( .DIN1(_40496), .DIN2(_41066), .Q(_41065) );
  nor2s1 _41073_inst ( .DIN1(_40529), .DIN2(_40951), .Q(_41066) );
  and2s1 _41074_inst ( .DIN1(_41067), .DIN2(_41068), .Q(_40496) );
  nor2s1 _41075_inst ( .DIN1(_41069), .DIN2(_41070), .Q(_41064) );
  xor2s1 _41076_inst ( .DIN1(_41071), .DIN2(_41072), .Q(_41070) );
  nnd2s1 _41077_inst ( .DIN1(_41073), .DIN2(_40686), .Q(_41071) );
  nor2s1 _41078_inst ( .DIN1(_40649), .DIN2(_40839), .Q(_41069) );
  nnd2s1 _41079_inst ( .DIN1(_41074), .DIN2(_41075), .Q(_41022) );
  nor2s1 _41080_inst ( .DIN1(_41076), .DIN2(_40556), .Q(_41075) );
  nnd2s1 _41081_inst ( .DIN1(_41077), .DIN2(_41078), .Q(_40556) );
  nnd2s1 _41082_inst ( .DIN1(_40995), .DIN2(_41079), .Q(_41078) );
  hi1s1 _41083_inst ( .DIN(_41080), .Q(_40995) );
  nnd2s1 _41084_inst ( .DIN1(_41081), .DIN2(_40888), .Q(_41077) );
  nor2s1 _41085_inst ( .DIN1(_41082), .DIN2(_40933), .Q(_41074) );
  nnd2s1 _41086_inst ( .DIN1(_41083), .DIN2(_41084), .Q(_40933) );
  nor2s1 _41087_inst ( .DIN1(_41085), .DIN2(_40606), .Q(_41084) );
  nor2s1 _41088_inst ( .DIN1(_41086), .DIN2(_41087), .Q(_41083) );
  nor2s1 _41089_inst ( .DIN1(_26842), .DIN2(_41088), .Q(_41086) );
  nor2s1 _41090_inst ( .DIN1(_41089), .DIN2(_41090), .Q(_41088) );
  nnd2s1 _41091_inst ( .DIN1(_41091), .DIN2(_36504), .Q(
        ____2____________12_____) );
  nnd2s1 _41092_inst ( .DIN1(_40486), .DIN2(_36511), .Q(_36504) );
  hi1s1 _41093_inst ( .DIN(_35938), .Q(_40486) );
  nnd2s1 _41094_inst ( .DIN1(_30043), .DIN2(_38283), .Q(_35938) );
  hi1s1 _41095_inst ( .DIN(_28071), .Q(_30043) );
  nor2s1 _41096_inst ( .DIN1(_41092), .DIN2(_41093), .Q(_41091) );
  nor2s1 _41097_inst ( .DIN1(_36511), .DIN2(_41094), .Q(_41093) );
  nnd2s1 _41098_inst ( .DIN1(_41095), .DIN2(_41096), .Q(_41094) );
  nor2s1 _41099_inst ( .DIN1(_41097), .DIN2(_41098), .Q(_41096) );
  nnd2s1 _41100_inst ( .DIN1(_41099), .DIN2(_41100), .Q(_41098) );
  nnd2s1 _41101_inst ( .DIN1(_41089), .DIN2(_40608), .Q(_41100) );
  hi1s1 _41102_inst ( .DIN(_40544), .Q(_41089) );
  nnd2s1 _41103_inst ( .DIN1(_41101), .DIN2(_33822), .Q(_40544) );
  nor2s1 _41104_inst ( .DIN1(_41102), .DIN2(_39027), .Q(_41101) );
  nor2s1 _41105_inst ( .DIN1(_41103), .DIN2(_41104), .Q(_41099) );
  nor2s1 _41106_inst ( .DIN1(_41105), .DIN2(_40896), .Q(_41104) );
  nor2s1 _41107_inst ( .DIN1(_41081), .DIN2(_40889), .Q(_41105) );
  nor2s1 _41108_inst ( .DIN1(_40965), .DIN2(_41106), .Q(_41103) );
  nnd2s1 _41109_inst ( .DIN1(_41107), .DIN2(_41108), .Q(_41097) );
  nor2s1 _41110_inst ( .DIN1(_41109), .DIN2(_40743), .Q(_41108) );
  and2s1 _41111_inst ( .DIN1(_41073), .DIN2(_40639), .Q(_40743) );
  nor2s1 _41112_inst ( .DIN1(_41110), .DIN2(_41111), .Q(_41107) );
  nor2s1 _41113_inst ( .DIN1(_40498), .DIN2(_40951), .Q(_41111) );
  nor2s1 _41114_inst ( .DIN1(_41112), .DIN2(_41113), .Q(_41095) );
  nnd2s1 _41115_inst ( .DIN1(_41114), .DIN2(_40842), .Q(_41113) );
  and2s1 _41116_inst ( .DIN1(_41115), .DIN2(_41116), .Q(_40842) );
  xor2s1 _41117_inst ( .DIN1(_33214), .DIN2(_41117), .Q(_41116) );
  nor2s1 _41118_inst ( .DIN1(_41118), .DIN2(_41119), .Q(_41117) );
  hi1s1 _41119_inst ( .DIN(_41120), .Q(_41118) );
  nor2s1 _41120_inst ( .DIN1(_41020), .DIN2(_41121), .Q(_41115) );
  hi1s1 _41121_inst ( .DIN(_40617), .Q(_41020) );
  nnd2s1 _41122_inst ( .DIN1(_41122), .DIN2(_40902), .Q(_40617) );
  nor2s1 _41123_inst ( .DIN1(_26842), .DIN2(_40903), .Q(_41122) );
  nor2s1 _41124_inst ( .DIN1(_41061), .DIN2(_40717), .Q(_41114) );
  nnd2s1 _41125_inst ( .DIN1(_41123), .DIN2(_41124), .Q(_40717) );
  nor2s1 _41126_inst ( .DIN1(_41125), .DIN2(_41126), .Q(_41124) );
  nnd2s1 _41127_inst ( .DIN1(_40980), .DIN2(_40588), .Q(_41126) );
  nnd2s1 _41128_inst ( .DIN1(_41127), .DIN2(_41068), .Q(_40980) );
  nor2s1 _41129_inst ( .DIN1(_26842), .DIN2(_34890), .Q(_41127) );
  nor2s1 _41130_inst ( .DIN1(_40903), .DIN2(_41128), .Q(_41125) );
  nnd2s1 _41131_inst ( .DIN1(_41129), .DIN2(_40495), .Q(_41128) );
  nor2s1 _41132_inst ( .DIN1(_40805), .DIN2(_41130), .Q(_41123) );
  nor2s1 _41133_inst ( .DIN1(_41131), .DIN2(_40839), .Q(_41130) );
  nor2s1 _41134_inst ( .DIN1(_40965), .DIN2(_40655), .Q(_40805) );
  nnd2s1 _41135_inst ( .DIN1(_41132), .DIN2(_41133), .Q(_41061) );
  nor2s1 _41136_inst ( .DIN1(_41134), .DIN2(_41135), .Q(_41133) );
  nnd2s1 _41137_inst ( .DIN1(_40616), .DIN2(_41136), .Q(_41135) );
  nnd2s1 _41138_inst ( .DIN1(_41137), .DIN2(_40754), .Q(_40616) );
  hi1s1 _41139_inst ( .DIN(_41138), .Q(_41137) );
  nor2s1 _41140_inst ( .DIN1(_40974), .DIN2(_40532), .Q(_41134) );
  nor2s1 _41141_inst ( .DIN1(_41139), .DIN2(_41140), .Q(_41132) );
  nor2s1 _41142_inst ( .DIN1(_40573), .DIN2(_40975), .Q(_41140) );
  nor2s1 _41143_inst ( .DIN1(_40654), .DIN2(_40755), .Q(_41139) );
  nnd2s1 _41144_inst ( .DIN1(_41141), .DIN2(_40659), .Q(_41112) );
  and2s1 _41145_inst ( .DIN1(_41142), .DIN2(_41143), .Q(_40659) );
  nor2s1 _41146_inst ( .DIN1(_41144), .DIN2(_41145), .Q(_41143) );
  nnd2s1 _41147_inst ( .DIN1(_41146), .DIN2(_41147), .Q(_41145) );
  nor2s1 _41148_inst ( .DIN1(_41148), .DIN2(_41149), .Q(_41147) );
  nor2s1 _41149_inst ( .DIN1(_40649), .DIN2(_41150), .Q(_41148) );
  nor2s1 _41150_inst ( .DIN1(_40508), .DIN2(_40620), .Q(_41146) );
  nnd2s1 _41151_inst ( .DIN1(_40800), .DIN2(_40910), .Q(_40620) );
  nnd2s1 _41152_inst ( .DIN1(_40803), .DIN2(_40783), .Q(_40910) );
  nnd2s1 _41153_inst ( .DIN1(_41151), .DIN2(_41152), .Q(_40800) );
  nor2s1 _41154_inst ( .DIN1(_41153), .DIN2(_40649), .Q(_41151) );
  nnd2s1 _41155_inst ( .DIN1(_41154), .DIN2(_41155), .Q(_40508) );
  nnd2s1 _41156_inst ( .DIN1(_40835), .DIN2(_40938), .Q(_41155) );
  hi1s1 _41157_inst ( .DIN(_40942), .Q(_40835) );
  xor2s1 _41158_inst ( .DIN1(_37577), .DIN2(_41156), .Q(_41154) );
  nnd2s1 _41159_inst ( .DIN1(_40993), .DIN2(_41033), .Q(_41156) );
  nnd2s1 _41160_inst ( .DIN1(_41157), .DIN2(_41158), .Q(_41144) );
  nor2s1 _41161_inst ( .DIN1(_40784), .DIN2(_41159), .Q(_41158) );
  nor2s1 _41162_inst ( .DIN1(_41160), .DIN2(_40896), .Q(_41159) );
  and2s1 _41163_inst ( .DIN1(_41161), .DIN2(_41033), .Q(_40784) );
  nor2s1 _41164_inst ( .DIN1(_41162), .DIN2(_41163), .Q(_41157) );
  nor2s1 _41165_inst ( .DIN1(_40654), .DIN2(_41080), .Q(_41163) );
  nor2s1 _41166_inst ( .DIN1(_41164), .DIN2(_40532), .Q(_41162) );
  nor2s1 _41167_inst ( .DIN1(_41165), .DIN2(_41166), .Q(_41142) );
  nnd2s1 _41168_inst ( .DIN1(_41167), .DIN2(_40932), .Q(_41166) );
  and2s1 _41169_inst ( .DIN1(_41168), .DIN2(_41169), .Q(_40932) );
  nor2s1 _41170_inst ( .DIN1(_40503), .DIN2(_41170), .Q(_41169) );
  hi1s1 _41171_inst ( .DIN(_41171), .Q(_40503) );
  nor2s1 _41172_inst ( .DIN1(_41172), .DIN2(_41173), .Q(_41168) );
  nor2s1 _41173_inst ( .DIN1(_40778), .DIN2(_40532), .Q(_41173) );
  nor2s1 _41174_inst ( .DIN1(_41174), .DIN2(_40498), .Q(_41172) );
  nor2s1 _41175_inst ( .DIN1(_41175), .DIN2(_41176), .Q(_41174) );
  nor2s1 _41176_inst ( .DIN1(_41045), .DIN2(_41082), .Q(_41167) );
  nnd2s1 _41177_inst ( .DIN1(_41177), .DIN2(_41178), .Q(_41082) );
  nnd2s1 _41178_inst ( .DIN1(_41179), .DIN2(_40608), .Q(_41178) );
  hi1s1 _41179_inst ( .DIN(_40543), .Q(_40608) );
  or2s1 _41180_inst ( .DIN1(_40574), .DIN2(_40573), .Q(_41177) );
  nnd2s1 _41181_inst ( .DIN1(_41180), .DIN2(_41181), .Q(_41045) );
  nor2s1 _41182_inst ( .DIN1(_40586), .DIN2(_41182), .Q(_41181) );
  nor2s1 _41183_inst ( .DIN1(_40498), .DIN2(_40912), .Q(_41182) );
  nor2s1 _41184_inst ( .DIN1(_40610), .DIN2(_40596), .Q(_41180) );
  nnd2s1 _41185_inst ( .DIN1(_41183), .DIN2(_41184), .Q(_40596) );
  or2s1 _41186_inst ( .DIN1(_40966), .DIN2(_40654), .Q(_41184) );
  nnd2s1 _41187_inst ( .DIN1(_41185), .DIN2(_40971), .Q(_41183) );
  nnd2s1 _41188_inst ( .DIN1(_41186), .DIN2(_41187), .Q(_41165) );
  nor2s1 _41189_inst ( .DIN1(_41188), .DIN2(_41189), .Q(_41187) );
  and2s1 _41190_inst ( .DIN1(_40550), .DIN2(_41190), .Q(_41186) );
  and2s1 _41191_inst ( .DIN1(_41191), .DIN2(_40704), .Q(_40550) );
  nnd2s1 _41192_inst ( .DIN1(_41192), .DIN2(_40938), .Q(_40704) );
  nor2s1 _41193_inst ( .DIN1(_41193), .DIN2(_41194), .Q(_41191) );
  nor2s1 _41194_inst ( .DIN1(_41059), .DIN2(_40896), .Q(_41194) );
  nor2s1 _41195_inst ( .DIN1(_40498), .DIN2(_41195), .Q(_41193) );
  nor2s1 _41196_inst ( .DIN1(_40860), .DIN2(_41087), .Q(_41141) );
  nnd2s1 _41197_inst ( .DIN1(_41196), .DIN2(_41197), .Q(_41087) );
  nor2s1 _41198_inst ( .DIN1(_41198), .DIN2(_41199), .Q(_41197) );
  nnd2s1 _41199_inst ( .DIN1(_41200), .DIN2(_40619), .Q(_41199) );
  nnd2s1 _41200_inst ( .DIN1(_40546), .DIN2(_40545), .Q(_41200) );
  nnd2s1 _41201_inst ( .DIN1(_41201), .DIN2(_41202), .Q(_40545) );
  nnd2s1 _41202_inst ( .DIN1(_41203), .DIN2(_41204), .Q(_41202) );
  nor2s1 _41203_inst ( .DIN1(_36337), .DIN2(_38990), .Q(_41204) );
  nor2s1 _41204_inst ( .DIN1(_34762), .DIN2(_34193), .Q(_41203) );
  nnd2s1 _41205_inst ( .DIN1(_41068), .DIN2(_27653), .Q(_41201) );
  nor2s1 _41206_inst ( .DIN1(_26842), .DIN2(_40499), .Q(_41198) );
  nor2s1 _41207_inst ( .DIN1(_40595), .DIN2(_41205), .Q(_41196) );
  or2s1 _41208_inst ( .DIN1(_41206), .DIN2(_40622), .Q(_41205) );
  nnd2s1 _41209_inst ( .DIN1(_41207), .DIN2(_41208), .Q(_40622) );
  or2s1 _41210_inst ( .DIN1(_41209), .DIN2(_40529), .Q(_41208) );
  nnd2s1 _41211_inst ( .DIN1(_41210), .DIN2(_40546), .Q(_41207) );
  nnd2s1 _41212_inst ( .DIN1(_41211), .DIN2(_41212), .Q(_40595) );
  nnd2s1 _41213_inst ( .DIN1(_40494), .DIN2(_40754), .Q(_41212) );
  hi1s1 _41214_inst ( .DIN(_40747), .Q(_40494) );
  and2s1 _41215_inst ( .DIN1(_41213), .DIN2(_41214), .Q(_41211) );
  nor2s1 _41216_inst ( .DIN1(_35940), .DIN2(_41215), .Q(_41092) );
  nor2s1 _41217_inst ( .DIN1(_41216), .DIN2(_26771), .Q(_41215) );
  xor2s1 _41218_inst ( .DIN1(_35939), .DIN2(_53398), .Q(_41216) );
  nnd2s1 _41219_inst ( .DIN1(_53408), .DIN2(_53406), .Q(_35939) );
  hi1s1 _41220_inst ( .DIN(_36511), .Q(_35940) );
  nnd2s1 _41221_inst ( .DIN1(_41217), .DIN2(_37955), .Q(_36511) );
  nor2s1 _41222_inst ( .DIN1(_36976), .DIN2(_36492), .Q(_37955) );
  hi1s1 _41223_inst ( .DIN(_38283), .Q(_36976) );
  nor2s1 _41224_inst ( .DIN1(_38072), .DIN2(_28071), .Q(_41217) );
  nnd2s1 _41225_inst ( .DIN1(_41218), .DIN2(_41219), .Q(_28071) );
  and2s1 _41226_inst ( .DIN1(_41220), .DIN2(_38284), .Q(_41219) );
  and2s1 _41227_inst ( .DIN1(_36021), .DIN2(_41221), .Q(_41218) );
  nnd2s1 _41228_inst ( .DIN1(_41222), .DIN2(_40560), .Q(
        ____2____________11_____) );
  nor2s1 _41229_inst ( .DIN1(_41223), .DIN2(_41224), .Q(_41222) );
  nor2s1 _41230_inst ( .DIN1(_40563), .DIN2(_41225), .Q(_41224) );
  xor2s1 _41231_inst ( .DIN1(_41226), .DIN2(_29579), .Q(_41225) );
  nnd2s1 _41232_inst ( .DIN1(_41227), .DIN2(_41228), .Q(_41226) );
  nor2s1 _41233_inst ( .DIN1(_41229), .DIN2(_41230), .Q(_41228) );
  nnd2s1 _41234_inst ( .DIN1(_41231), .DIN2(_41232), .Q(_41230) );
  and2s1 _41235_inst ( .DIN1(_41136), .DIN2(_41233), .Q(_41232) );
  nnd2s1 _41236_inst ( .DIN1(_41234), .DIN2(_40989), .Q(_41136) );
  nor2s1 _41237_inst ( .DIN1(_40895), .DIN2(_41235), .Q(_41234) );
  nor2s1 _41238_inst ( .DIN1(_41119), .DIN2(_41236), .Q(_41231) );
  nor2s1 _41239_inst ( .DIN1(_40879), .DIN2(_40529), .Q(_41119) );
  nnd2s1 _41240_inst ( .DIN1(_41237), .DIN2(_41238), .Q(_41229) );
  nor2s1 _41241_inst ( .DIN1(_41036), .DIN2(_40838), .Q(_41238) );
  and2s1 _41242_inst ( .DIN1(_41239), .DIN2(_40989), .Q(_40838) );
  nor2s1 _41243_inst ( .DIN1(_33520), .DIN2(_41240), .Q(_41239) );
  nor2s1 _41244_inst ( .DIN1(_40777), .DIN2(_41164), .Q(_41036) );
  and2s1 _41245_inst ( .DIN1(_40668), .DIN2(_41241), .Q(_41237) );
  nnd2s1 _41246_inst ( .DIN1(_41037), .DIN2(_41242), .Q(_40668) );
  nor2s1 _41247_inst ( .DIN1(_41243), .DIN2(_41244), .Q(_41227) );
  nnd2s1 _41248_inst ( .DIN1(_41245), .DIN2(_41246), .Q(_41244) );
  xor2s1 _41249_inst ( .DIN1(_32716), .DIN2(_41247), .Q(_41246) );
  nor2s1 _41250_inst ( .DIN1(_40904), .DIN2(_40943), .Q(_41247) );
  nnd2s1 _41251_inst ( .DIN1(_41248), .DIN2(_41249), .Q(_40943) );
  or2s1 _41252_inst ( .DIN1(_40576), .DIN2(_40575), .Q(_41249) );
  or2s1 _41253_inst ( .DIN1(_40655), .DIN2(_40654), .Q(_41248) );
  nnd2s1 _41254_inst ( .DIN1(_40618), .DIN2(_41250), .Q(_40904) );
  nnd2s1 _41255_inst ( .DIN1(_41251), .DIN2(_41252), .Q(_41250) );
  nor2s1 _41256_inst ( .DIN1(_40699), .DIN2(_34893), .Q(_41252) );
  nor2s1 _41257_inst ( .DIN1(_41253), .DIN2(_41254), .Q(_41251) );
  nnd2s1 _41258_inst ( .DIN1(_41179), .DIN2(_41255), .Q(_40618) );
  xnr2s1 _41259_inst ( .DIN1(_29049), .DIN2(_40806), .Q(_41179) );
  nor2s1 _41260_inst ( .DIN1(_41256), .DIN2(_41257), .Q(_41245) );
  nnd2s1 _41261_inst ( .DIN1(_41258), .DIN2(_41259), .Q(_41243) );
  nor2s1 _41262_inst ( .DIN1(_41260), .DIN2(_41261), .Q(_41259) );
  nor2s1 _41263_inst ( .DIN1(_40573), .DIN2(_40765), .Q(_41261) );
  nor2s1 _41264_inst ( .DIN1(_40529), .DIN2(_40574), .Q(_41260) );
  nor2s1 _41265_inst ( .DIN1(_40507), .DIN2(_41262), .Q(_41258) );
  nnd2s1 _41266_inst ( .DIN1(_41263), .DIN2(_41264), .Q(_40507) );
  nor2s1 _41267_inst ( .DIN1(_41265), .DIN2(_41266), .Q(_41264) );
  nnd2s1 _41268_inst ( .DIN1(_41267), .DIN2(_40837), .Q(_41266) );
  nnd2s1 _41269_inst ( .DIN1(_41176), .DIN2(_40783), .Q(_40837) );
  nor2s1 _41270_inst ( .DIN1(_41268), .DIN2(_41269), .Q(_41267) );
  nor2s1 _41271_inst ( .DIN1(_40777), .DIN2(_41138), .Q(_41269) );
  and2s1 _41272_inst ( .DIN1(_41033), .DIN2(_40994), .Q(_41268) );
  nnd2s1 _41273_inst ( .DIN1(_40649), .DIN2(_41131), .Q(_41033) );
  nnd2s1 _41274_inst ( .DIN1(_41270), .DIN2(_41120), .Q(_41265) );
  nnd2s1 _41275_inst ( .DIN1(_41001), .DIN2(_41271), .Q(_41120) );
  hi1s1 _41276_inst ( .DIN(_40642), .Q(_41001) );
  nor2s1 _41277_inst ( .DIN1(_40585), .DIN2(_41272), .Q(_41270) );
  hi1s1 _41278_inst ( .DIN(_41214), .Q(_41272) );
  and2s1 _41279_inst ( .DIN1(_40546), .DIN2(_41273), .Q(_40585) );
  nor2s1 _41280_inst ( .DIN1(_41274), .DIN2(_41275), .Q(_41263) );
  nnd2s1 _41281_inst ( .DIN1(_41276), .DIN2(_41277), .Q(_41275) );
  hi1s1 _41282_inst ( .DIN(_41278), .Q(_41277) );
  nor2s1 _41283_inst ( .DIN1(_41016), .DIN2(_40679), .Q(_41276) );
  nnd2s1 _41284_inst ( .DIN1(_41279), .DIN2(_41280), .Q(_40679) );
  nor2s1 _41285_inst ( .DIN1(_41281), .DIN2(_41282), .Q(_41280) );
  hi1s1 _41286_inst ( .DIN(_41283), .Q(_41281) );
  nor2s1 _41287_inst ( .DIN1(_41284), .DIN2(_40982), .Q(_41279) );
  nor2s1 _41288_inst ( .DIN1(_40529), .DIN2(_41014), .Q(_41284) );
  nnd2s1 _41289_inst ( .DIN1(_41285), .DIN2(_41286), .Q(_41016) );
  nor2s1 _41290_inst ( .DIN1(_41109), .DIN2(_41287), .Q(_41286) );
  nor2s1 _41291_inst ( .DIN1(_40575), .DIN2(_41288), .Q(_41287) );
  nor2s1 _41292_inst ( .DIN1(_40940), .DIN2(_40882), .Q(_41285) );
  nnd2s1 _41293_inst ( .DIN1(_41289), .DIN2(_41290), .Q(_40882) );
  nnd2s1 _41294_inst ( .DIN1(_41291), .DIN2(_40971), .Q(_41290) );
  nnd2s1 _41295_inst ( .DIN1(_41292), .DIN2(_41293), .Q(_40940) );
  nnd2s1 _41296_inst ( .DIN1(_40685), .DIN2(_41002), .Q(_41293) );
  hi1s1 _41297_inst ( .DIN(_41294), .Q(_40685) );
  nnd2s1 _41298_inst ( .DIN1(_40972), .DIN2(_41291), .Q(_41292) );
  hi1s1 _41299_inst ( .DIN(_40849), .Q(_41291) );
  nnd2s1 _41300_inst ( .DIN1(_41295), .DIN2(_40809), .Q(_41274) );
  nor2s1 _41301_inst ( .DIN1(_41296), .DIN2(_40721), .Q(_40809) );
  nnd2s1 _41302_inst ( .DIN1(_41297), .DIN2(_41298), .Q(_40721) );
  nor2s1 _41303_inst ( .DIN1(_41299), .DIN2(_41300), .Q(_41298) );
  nor2s1 _41304_inst ( .DIN1(_41301), .DIN2(_40778), .Q(_41300) );
  nor2s1 _41305_inst ( .DIN1(_41302), .DIN2(_41303), .Q(_41297) );
  nor2s1 _41306_inst ( .DIN1(_40965), .DIN2(_41080), .Q(_41303) );
  hi1s1 _41307_inst ( .DIN(_40937), .Q(_40965) );
  nor2s1 _41308_inst ( .DIN1(_40573), .DIN2(_41304), .Q(_41302) );
  or2s1 _41309_inst ( .DIN1(_41170), .DIN2(_41305), .Q(_41296) );
  nor2s1 _41310_inst ( .DIN1(_26842), .DIN2(_40652), .Q(_41305) );
  nor2s1 _41311_inst ( .DIN1(_40700), .DIN2(_26842), .Q(_41170) );
  nnd2s1 _41312_inst ( .DIN1(_41306), .DIN2(_41307), .Q(_40700) );
  nor2s1 _41313_inst ( .DIN1(_41308), .DIN2(_40996), .Q(_41295) );
  nnd2s1 _41314_inst ( .DIN1(_41309), .DIN2(_41310), .Q(_40996) );
  or2s1 _41315_inst ( .DIN1(_41160), .DIN2(_41062), .Q(_41310) );
  nnd2s1 _41316_inst ( .DIN1(_40770), .DIN2(_40754), .Q(_41309) );
  hi1s1 _41317_inst ( .DIN(_41311), .Q(_40770) );
  nor2s1 _41318_inst ( .DIN1(_41312), .DIN2(_41313), .Q(_41308) );
  nor2s1 _41319_inst ( .DIN1(_40519), .DIN2(_41314), .Q(_41223) );
  nor2s1 _41320_inst ( .DIN1(_27365), .DIN2(_26208), .Q(_41314) );
  nnd2s1 _41321_inst ( .DIN1(_41315), .DIN2(_40560), .Q(
        ____2____________10_____) );
  nnd2s1 _41322_inst ( .DIN1(_41316), .DIN2(_40563), .Q(_40560) );
  nor2s1 _41323_inst ( .DIN1(_41317), .DIN2(_41318), .Q(_41315) );
  nor2s1 _41324_inst ( .DIN1(_40563), .DIN2(_41319), .Q(_41318) );
  nnd2s1 _41325_inst ( .DIN1(_41320), .DIN2(_41321), .Q(_41319) );
  nor2s1 _41326_inst ( .DIN1(_41322), .DIN2(_41323), .Q(_41321) );
  nnd2s1 _41327_inst ( .DIN1(_41324), .DIN2(_41325), .Q(_41323) );
  nor2s1 _41328_inst ( .DIN1(_41326), .DIN2(_41282), .Q(_41325) );
  nor2s1 _41329_inst ( .DIN1(_41301), .DIN2(_40974), .Q(_41282) );
  hi1s1 _41330_inst ( .DIN(_41271), .Q(_41301) );
  nor2s1 _41331_inst ( .DIN1(_41327), .DIN2(_41328), .Q(_41326) );
  nnd2s1 _41332_inst ( .DIN1(_41329), .DIN2(_40937), .Q(_41328) );
  nnd2s1 _41333_inst ( .DIN1(_41330), .DIN2(_40654), .Q(_40937) );
  nor2s1 _41334_inst ( .DIN1(_41331), .DIN2(_40898), .Q(_41324) );
  nor2s1 _41335_inst ( .DIN1(_40543), .DIN2(_39537), .Q(_40898) );
  nor2s1 _41336_inst ( .DIN1(_40777), .DIN2(_40533), .Q(_41331) );
  nnd2s1 _41337_inst ( .DIN1(_41332), .DIN2(_41333), .Q(_41322) );
  nor2s1 _41338_inst ( .DIN1(_41334), .DIN2(_41335), .Q(_41333) );
  nnd2s1 _41339_inst ( .DIN1(_40876), .DIN2(_41171), .Q(_41335) );
  nnd2s1 _41340_inst ( .DIN1(_41336), .DIN2(_41337), .Q(_41171) );
  nor2s1 _41341_inst ( .DIN1(_41338), .DIN2(_41339), .Q(_41337) );
  nnd2s1 _41342_inst ( .DIN1(_40686), .DIN2(_41340), .Q(_41339) );
  hi1s1 _41343_inst ( .DIN(_40699), .Q(_40686) );
  nor2s1 _41344_inst ( .DIN1(_41341), .DIN2(_40518), .Q(_41336) );
  nnd2s1 _41345_inst ( .DIN1(_40607), .DIN2(_41255), .Q(_40876) );
  hi1s1 _41346_inst ( .DIN(_41342), .Q(_41334) );
  nor2s1 _41347_inst ( .DIN1(_40586), .DIN2(_41343), .Q(_41332) );
  nor2s1 _41348_inst ( .DIN1(_40654), .DIN2(_41311), .Q(_41343) );
  hi1s1 _41349_inst ( .DIN(_41344), .Q(_40586) );
  nor2s1 _41350_inst ( .DIN1(_41345), .DIN2(_41346), .Q(_41320) );
  nnd2s1 _41351_inst ( .DIN1(_41347), .DIN2(_41348), .Q(_41346) );
  nor2s1 _41352_inst ( .DIN1(_40718), .DIN2(_40772), .Q(_41348) );
  nnd2s1 _41353_inst ( .DIN1(_41349), .DIN2(_41350), .Q(_40772) );
  nor2s1 _41354_inst ( .DIN1(_41351), .DIN2(_41352), .Q(_41350) );
  nnd2s1 _41355_inst ( .DIN1(_41353), .DIN2(_40619), .Q(_41352) );
  nnd2s1 _41356_inst ( .DIN1(_41354), .DIN2(_41355), .Q(_40619) );
  nor2s1 _41357_inst ( .DIN1(_34893), .DIN2(_41253), .Q(_41355) );
  nor2s1 _41358_inst ( .DIN1(_41254), .DIN2(_40745), .Q(_41354) );
  nnd2s1 _41359_inst ( .DIN1(_41079), .DIN2(_41356), .Q(_41353) );
  nnd2s1 _41360_inst ( .DIN1(_40655), .DIN2(_41080), .Q(_41356) );
  nnd2s1 _41361_inst ( .DIN1(_41357), .DIN2(_41358), .Q(_41080) );
  nor2s1 _41362_inst ( .DIN1(_41338), .DIN2(_41359), .Q(_41357) );
  nnd2s1 _41363_inst ( .DIN1(_40709), .DIN2(_41214), .Q(_41351) );
  nnd2s1 _41364_inst ( .DIN1(_41360), .DIN2(_41361), .Q(_41214) );
  nnd2s1 _41365_inst ( .DIN1(_41242), .DIN2(_40806), .Q(_40709) );
  nor2s1 _41366_inst ( .DIN1(_41153), .DIN2(_40903), .Q(_40806) );
  nor2s1 _41367_inst ( .DIN1(_41362), .DIN2(_41363), .Q(_41349) );
  nnd2s1 _41368_inst ( .DIN1(_41364), .DIN2(_41365), .Q(_41363) );
  hi1s1 _41369_inst ( .DIN(_41366), .Q(_41365) );
  xor2s1 _41370_inst ( .DIN1(_41367), .DIN2(_41368), .Q(_41364) );
  nor2s1 _41371_inst ( .DIN1(_41369), .DIN2(_41370), .Q(_41368) );
  nnd2s1 _41372_inst ( .DIN1(_41371), .DIN2(_41372), .Q(_41370) );
  nor2s1 _41373_inst ( .DIN1(_40675), .DIN2(_41373), .Q(_41372) );
  nor2s1 _41374_inst ( .DIN1(_41042), .DIN2(_40827), .Q(_41371) );
  nnd2s1 _41375_inst ( .DIN1(_41374), .DIN2(_41375), .Q(_40827) );
  nor2s1 _41376_inst ( .DIN1(_41376), .DIN2(_41377), .Q(_41375) );
  nnd2s1 _41377_inst ( .DIN1(_41233), .DIN2(_41032), .Q(_41377) );
  or2s1 _41378_inst ( .DIN1(_41195), .DIN2(_40529), .Q(_41032) );
  nnd2s1 _41379_inst ( .DIN1(_41378), .DIN2(_41379), .Q(_41376) );
  hi1s1 _41380_inst ( .DIN(_41050), .Q(_41379) );
  nor2s1 _41381_inst ( .DIN1(_40653), .DIN2(_41160), .Q(_41050) );
  nnd2s1 _41382_inst ( .DIN1(_41380), .DIN2(_41381), .Q(_41160) );
  nor2s1 _41383_inst ( .DIN1(_40606), .DIN2(_40504), .Q(_41378) );
  nor2s1 _41384_inst ( .DIN1(_41164), .DIN2(_26842), .Q(_40504) );
  nnd2s1 _41385_inst ( .DIN1(_41382), .DIN2(_41381), .Q(_41164) );
  hi1s1 _41386_inst ( .DIN(_41383), .Q(_41381) );
  nor2s1 _41387_inst ( .DIN1(_41384), .DIN2(_41385), .Q(_40606) );
  nor2s1 _41388_inst ( .DIN1(_41386), .DIN2(_41387), .Q(_41374) );
  nnd2s1 _41389_inst ( .DIN1(_41388), .DIN2(_41389), .Q(_41387) );
  hi1s1 _41390_inst ( .DIN(_40676), .Q(_41389) );
  xor2s1 _41391_inst ( .DIN1(_40723), .DIN2(_31658), .Q(_41388) );
  nnd2s1 _41392_inst ( .DIN1(_41390), .DIN2(_41391), .Q(_40723) );
  hi1s1 _41393_inst ( .DIN(_41189), .Q(_41391) );
  nor2s1 _41394_inst ( .DIN1(_41392), .DIN2(_41393), .Q(_41390) );
  nor2s1 _41395_inst ( .DIN1(_40699), .DIN2(_41288), .Q(_41393) );
  nor2s1 _41396_inst ( .DIN1(_40745), .DIN2(_41294), .Q(_41392) );
  nnd2s1 _41397_inst ( .DIN1(_41394), .DIN2(_41395), .Q(_41294) );
  nor2s1 _41398_inst ( .DIN1(_53414), .DIN2(_41396), .Q(_41394) );
  nnd2s1 _41399_inst ( .DIN1(_41397), .DIN2(_41398), .Q(_41386) );
  hi1s1 _41400_inst ( .DIN(_40610), .Q(_41398) );
  nnd2s1 _41401_inst ( .DIN1(_41399), .DIN2(_41400), .Q(_40610) );
  nnd2s1 _41402_inst ( .DIN1(_41401), .DIN2(_41402), .Q(_41400) );
  nor2s1 _41403_inst ( .DIN1(_27630), .DIN2(_40777), .Q(_41401) );
  nor2s1 _41404_inst ( .DIN1(_41403), .DIN2(_41404), .Q(_41397) );
  nor2s1 _41405_inst ( .DIN1(_41063), .DIN2(_40653), .Q(_41404) );
  nor2s1 _41406_inst ( .DIN1(_41405), .DIN2(_40649), .Q(_41403) );
  nnd2s1 _41407_inst ( .DIN1(_41406), .DIN2(_41407), .Q(_41042) );
  nnd2s1 _41408_inst ( .DIN1(_40936), .DIN2(_40886), .Q(_41407) );
  hi1s1 _41409_inst ( .DIN(_41106), .Q(_40936) );
  nnd2s1 _41410_inst ( .DIN1(_40801), .DIN2(_40639), .Q(_41406) );
  hi1s1 _41411_inst ( .DIN(_40913), .Q(_40801) );
  nnd2s1 _41412_inst ( .DIN1(_41408), .DIN2(_41409), .Q(_41369) );
  nor2s1 _41413_inst ( .DIN1(_41410), .DIN2(_41411), .Q(_41409) );
  or2s1 _41414_inst ( .DIN1(_40878), .DIN2(_41109), .Q(_41411) );
  hi1s1 _41415_inst ( .DIN(_40587), .Q(_41109) );
  nnd2s1 _41416_inst ( .DIN1(_41412), .DIN2(_41413), .Q(_40587) );
  nor2s1 _41417_inst ( .DIN1(_40529), .DIN2(_41414), .Q(_41413) );
  nor2s1 _41418_inst ( .DIN1(_39133), .DIN2(_41415), .Q(_41412) );
  nor2s1 _41419_inst ( .DIN1(_40576), .DIN2(_40745), .Q(_40878) );
  nor2s1 _41420_inst ( .DIN1(_40648), .DIN2(_41131), .Q(_41410) );
  and2s1 _41421_inst ( .DIN1(_40810), .DIN2(_40819), .Q(_40648) );
  nor2s1 _41422_inst ( .DIN1(_41416), .DIN2(_40982), .Q(_41408) );
  xor2s1 _41423_inst ( .DIN1(_41417), .DIN2(_32716), .Q(_40982) );
  nnd2s1 _41424_inst ( .DIN1(_41418), .DIN2(_41419), .Q(_41417) );
  nnd2s1 _41425_inst ( .DIN1(_41067), .DIN2(_41420), .Q(_41419) );
  nor2s1 _41426_inst ( .DIN1(_41330), .DIN2(_34890), .Q(_41067) );
  nor2s1 _41427_inst ( .DIN1(_41421), .DIN2(_41422), .Q(_41418) );
  nor2s1 _41428_inst ( .DIN1(_40895), .DIN2(_41423), .Q(_41422) );
  nnd2s1 _41429_inst ( .DIN1(_41129), .DIN2(_41056), .Q(_41423) );
  nor2s1 _41430_inst ( .DIN1(_41424), .DIN2(_41425), .Q(_41421) );
  or2s1 _41431_inst ( .DIN1(_33139), .DIN2(_41102), .Q(_41425) );
  nnd2s1 _41432_inst ( .DIN1(_41426), .DIN2(_41427), .Q(_41362) );
  nnd2s1 _41433_inst ( .DIN1(_40834), .DIN2(_41428), .Q(_41426) );
  nnd2s1 _41434_inst ( .DIN1(_41429), .DIN2(_41430), .Q(_40718) );
  nor2s1 _41435_inst ( .DIN1(_41431), .DIN2(_41432), .Q(_41430) );
  nnd2s1 _41436_inst ( .DIN1(_41433), .DIN2(_41283), .Q(_41432) );
  nnd2s1 _41437_inst ( .DIN1(_41434), .DIN2(_41435), .Q(_41283) );
  nor2s1 _41438_inst ( .DIN1(_40543), .DIN2(_41436), .Q(_41434) );
  nnd2s1 _41439_inst ( .DIN1(_41437), .DIN2(_40989), .Q(_41433) );
  nor2s1 _41440_inst ( .DIN1(_41256), .DIN2(_41438), .Q(_41429) );
  nnd2s1 _41441_inst ( .DIN1(_41190), .DIN2(_40681), .Q(_41438) );
  hi1s1 _41442_inst ( .DIN(_41439), .Q(_40681) );
  nor2s1 _41443_inst ( .DIN1(_40599), .DIN2(_41440), .Q(_41190) );
  and2s1 _41444_inst ( .DIN1(_41273), .DIN2(_41271), .Q(_41440) );
  nnd2s1 _41445_inst ( .DIN1(_40955), .DIN2(_41441), .Q(_41256) );
  nnd2s1 _41446_inst ( .DIN1(_41161), .DIN2(_40989), .Q(_40955) );
  hi1s1 _41447_inst ( .DIN(_40649), .Q(_40989) );
  nor2s1 _41448_inst ( .DIN1(_40826), .DIN2(_41257), .Q(_41347) );
  nnd2s1 _41449_inst ( .DIN1(_41442), .DIN2(_41443), .Q(_41257) );
  nor2s1 _41450_inst ( .DIN1(_41444), .DIN2(_41445), .Q(_41443) );
  nnd2s1 _41451_inst ( .DIN1(_41446), .DIN2(_40540), .Q(_41445) );
  nnd2s1 _41452_inst ( .DIN1(_41447), .DIN2(_40886), .Q(_40540) );
  hi1s1 _41453_inst ( .DIN(_40654), .Q(_40886) );
  nor2s1 _41454_inst ( .DIN1(_34890), .DIN2(_41448), .Q(_41447) );
  nnd2s1 _41455_inst ( .DIN1(_41079), .DIN2(_41449), .Q(_41446) );
  nnd2s1 _41456_inst ( .DIN1(_40755), .DIN2(_40966), .Q(_41449) );
  nnd2s1 _41457_inst ( .DIN1(_41450), .DIN2(_41451), .Q(_40966) );
  nor2s1 _41458_inst ( .DIN1(_41452), .DIN2(_34211), .Q(_41450) );
  nor2s1 _41459_inst ( .DIN1(_41453), .DIN2(_40498), .Q(_41444) );
  and2s1 _41460_inst ( .DIN1(_40499), .DIN2(_40951), .Q(_41453) );
  nnd2s1 _41461_inst ( .DIN1(_41454), .DIN2(_41455), .Q(_40951) );
  nor2s1 _41462_inst ( .DIN1(_36336), .DIN2(_39027), .Q(_41454) );
  nnd2s1 _41463_inst ( .DIN1(_41456), .DIN2(_33945), .Q(_40499) );
  nor2s1 _41464_inst ( .DIN1(_41102), .DIN2(_39026), .Q(_41456) );
  nor2s1 _41465_inst ( .DIN1(_41457), .DIN2(_41458), .Q(_41442) );
  nnd2s1 _41466_inst ( .DIN1(_41459), .DIN2(_41460), .Q(_41458) );
  nnd2s1 _41467_inst ( .DIN1(_41000), .DIN2(_40967), .Q(_41460) );
  nor2s1 _41468_inst ( .DIN1(_41461), .DIN2(_41452), .Q(_40967) );
  nnd2s1 _41469_inst ( .DIN1(_41185), .DIN2(_40972), .Q(_41459) );
  hi1s1 _41470_inst ( .DIN(_40850), .Q(_40972) );
  hi1s1 _41471_inst ( .DIN(_40970), .Q(_41185) );
  nnd2s1 _41472_inst ( .DIN1(_41462), .DIN2(_41455), .Q(_40970) );
  nor2s1 _41473_inst ( .DIN1(_27630), .DIN2(_36308), .Q(_41462) );
  nor2s1 _41474_inst ( .DIN1(_26842), .DIN2(_40747), .Q(_41457) );
  nnd2s1 _41475_inst ( .DIN1(_41463), .DIN2(_41464), .Q(_40826) );
  nor2s1 _41476_inst ( .DIN1(_41465), .DIN2(_41466), .Q(_41463) );
  hi1s1 _41477_inst ( .DIN(_41467), .Q(_41466) );
  nnd2s1 _41478_inst ( .DIN1(_41468), .DIN2(_41469), .Q(_41345) );
  nor2s1 _41479_inst ( .DIN1(_41470), .DIN2(_41149), .Q(_41469) );
  nor2s1 _41480_inst ( .DIN1(_40498), .DIN2(_40765), .Q(_41149) );
  nor2s1 _41481_inst ( .DIN1(_41062), .DIN2(_40942), .Q(_41470) );
  nor2s1 _41482_inst ( .DIN1(_41471), .DIN2(_41206), .Q(_41468) );
  nor2s1 _41483_inst ( .DIN1(_39969), .DIN2(_41313), .Q(_41471) );
  nor2s1 _41484_inst ( .DIN1(_40519), .DIN2(_41472), .Q(_41317) );
  xor2s1 _41485_inst ( .DIN1(_53418), .DIN2(_53420), .Q(_41472) );
  nnd2s1 _41486_inst ( .DIN1(_41473), .DIN2(_41474), .Q(
        ____2____________0_____) );
  nnd2s1 _41487_inst ( .DIN1(_28010), .DIN2(_41475), .Q(_41474) );
  nnd2s1 _41488_inst ( .DIN1(_41476), .DIN2(_41477), .Q(_41475) );
  nor2s1 _41489_inst ( .DIN1(_41478), .DIN2(_41479), .Q(_41477) );
  nnd2s1 _41490_inst ( .DIN1(_41480), .DIN2(_41481), .Q(_41479) );
  nor2s1 _41491_inst ( .DIN1(_41482), .DIN2(_41483), .Q(_41481) );
  nor2s1 _41492_inst ( .DIN1(_41461), .DIN2(_41484), .Q(_41483) );
  nnd2s1 _41493_inst ( .DIN1(_27653), .DIN2(_41271), .Q(_41484) );
  nnd2s1 _41494_inst ( .DIN1(_40532), .DIN2(_40777), .Q(_41271) );
  nor2s1 _41495_inst ( .DIN1(_41485), .DIN2(_41486), .Q(_41482) );
  nnd2s1 _41496_inst ( .DIN1(_41487), .DIN2(_41255), .Q(_41486) );
  hi1s1 _41497_inst ( .DIN(_41436), .Q(_41487) );
  nor2s1 _41498_inst ( .DIN1(_41488), .DIN2(_41489), .Q(_41480) );
  nor2s1 _41499_inst ( .DIN1(_40748), .DIN2(_41490), .Q(_41489) );
  nor2s1 _41500_inst ( .DIN1(_41491), .DIN2(_26793), .Q(_41488) );
  nor2s1 _41501_inst ( .DIN1(_41492), .DIN2(_41493), .Q(_41491) );
  nnd2s1 _41502_inst ( .DIN1(_41494), .DIN2(_41495), .Q(_41493) );
  nnd2s1 _41503_inst ( .DIN1(_39031), .DIN2(_41496), .Q(_41495) );
  nnd2s1 _41504_inst ( .DIN1(_41461), .DIN2(_41497), .Q(_41496) );
  nnd2s1 _41505_inst ( .DIN1(_41498), .DIN2(_33275), .Q(_41497) );
  nnd2s1 _41506_inst ( .DIN1(_41420), .DIN2(_39193), .Q(_41494) );
  nnd2s1 _41507_inst ( .DIN1(_40912), .DIN2(_41209), .Q(_41492) );
  nnd2s1 _41508_inst ( .DIN1(_41499), .DIN2(_33946), .Q(_41209) );
  nor2s1 _41509_inst ( .DIN1(_34890), .DIN2(_41485), .Q(_41499) );
  nnd2s1 _41510_inst ( .DIN1(_41500), .DIN2(_41501), .Q(_40912) );
  nor2s1 _41511_inst ( .DIN1(_41253), .DIN2(_39257), .Q(_41501) );
  nnd2s1 _41512_inst ( .DIN1(_41502), .DIN2(_41503), .Q(_41478) );
  nor2s1 _41513_inst ( .DIN1(_41504), .DIN2(_41465), .Q(_41503) );
  nor2s1 _41514_inst ( .DIN1(_40756), .DIN2(_40857), .Q(_41465) );
  nnd2s1 _41515_inst ( .DIN1(_41402), .DIN2(_34960), .Q(_40756) );
  hi1s1 _41516_inst ( .DIN(_41399), .Q(_41504) );
  nnd2s1 _41517_inst ( .DIN1(_41505), .DIN2(_41506), .Q(_41399) );
  nor2s1 _41518_inst ( .DIN1(_41452), .DIN2(_41102), .Q(_41506) );
  nor2s1 _41519_inst ( .DIN1(_40857), .DIN2(_41507), .Q(_41505) );
  nor2s1 _41520_inst ( .DIN1(_41508), .DIN2(_40646), .Q(_41502) );
  nor2s1 _41521_inst ( .DIN1(_40532), .DIN2(_41138), .Q(_40646) );
  nnd2s1 _41522_inst ( .DIN1(_41509), .DIN2(_41510), .Q(_41138) );
  nor2s1 _41523_inst ( .DIN1(_39301), .DIN2(_34204), .Q(_41509) );
  hi1s1 _41524_inst ( .DIN(_41233), .Q(_41508) );
  nnd2s1 _41525_inst ( .DIN1(_40888), .DIN2(_41192), .Q(_41233) );
  hi1s1 _41526_inst ( .DIN(_41021), .Q(_41192) );
  nnd2s1 _41527_inst ( .DIN1(_41511), .DIN2(_41455), .Q(_41021) );
  nor2s1 _41528_inst ( .DIN1(_41512), .DIN2(_41513), .Q(_41476) );
  nnd2s1 _41529_inst ( .DIN1(_41514), .DIN2(_41515), .Q(_41513) );
  nor2s1 _41530_inst ( .DIN1(_40905), .DIN2(_40945), .Q(_41515) );
  nnd2s1 _41531_inst ( .DIN1(_41516), .DIN2(_41517), .Q(_40945) );
  nor2s1 _41532_inst ( .DIN1(_41518), .DIN2(_41519), .Q(_41517) );
  nnd2s1 _41533_inst ( .DIN1(_41464), .DIN2(_41520), .Q(_41519) );
  hi1s1 _41534_inst ( .DIN(_41236), .Q(_41520) );
  nor2s1 _41535_inst ( .DIN1(_40580), .DIN2(_40857), .Q(_41236) );
  nnd2s1 _41536_inst ( .DIN1(_41361), .DIN2(_40495), .Q(_41464) );
  and2s1 _41537_inst ( .DIN1(_41521), .DIN2(_34531), .Q(_41361) );
  nor2s1 _41538_inst ( .DIN1(_41522), .DIN2(_33931), .Q(_41521) );
  nnd2s1 _41539_inst ( .DIN1(_41342), .DIN2(_40815), .Q(_41518) );
  nnd2s1 _41540_inst ( .DIN1(_41523), .DIN2(_40856), .Q(_40815) );
  nor2s1 _41541_inst ( .DIN1(_40529), .DIN2(_39032), .Q(_41523) );
  nnd2s1 _41542_inst ( .DIN1(_41524), .DIN2(_41525), .Q(_41342) );
  nor2s1 _41543_inst ( .DIN1(_40699), .DIN2(_34638), .Q(_41525) );
  nor2s1 _41544_inst ( .DIN1(_41254), .DIN2(_33825), .Q(_41524) );
  nor2s1 _41545_inst ( .DIN1(_41526), .DIN2(_41527), .Q(_41516) );
  nnd2s1 _41546_inst ( .DIN1(_41528), .DIN2(_41441), .Q(_41527) );
  nnd2s1 _41547_inst ( .DIN1(_40803), .DIN2(_41360), .Q(_41441) );
  and2s1 _41548_inst ( .DIN1(_41529), .DIN2(_41530), .Q(_40803) );
  or2s1 _41549_inst ( .DIN1(_40879), .DIN2(_40573), .Q(_41528) );
  nnd2s1 _41550_inst ( .DIN1(_41531), .DIN2(_41532), .Q(_40879) );
  nor2s1 _41551_inst ( .DIN1(_37778), .DIN2(_34638), .Q(_41532) );
  nor2s1 _41552_inst ( .DIN1(_33520), .DIN2(_41253), .Q(_41531) );
  xor2s1 _41553_inst ( .DIN1(_27840), .DIN2(_41533), .Q(_41526) );
  nor2s1 _41554_inst ( .DIN1(_41121), .DIN2(_40751), .Q(_41533) );
  and2s1 _41555_inst ( .DIN1(_41242), .DIN2(_40607), .Q(_40751) );
  nor2s1 _41556_inst ( .DIN1(_41235), .DIN2(_41327), .Q(_40607) );
  and2s1 _41557_inst ( .DIN1(_41051), .DIN2(_40971), .Q(_41121) );
  and2s1 _41558_inst ( .DIN1(_41534), .DIN2(_34765), .Q(_41051) );
  nor2s1 _41559_inst ( .DIN1(_41522), .DIN2(_34204), .Q(_41534) );
  nnd2s1 _41560_inst ( .DIN1(_41535), .DIN2(_41536), .Q(_40905) );
  nnd2s1 _41561_inst ( .DIN1(_41056), .DIN2(_40994), .Q(_41536) );
  nnd2s1 _41562_inst ( .DIN1(_41537), .DIN2(_41150), .Q(_40994) );
  hi1s1 _41563_inst ( .DIN(_41055), .Q(_41150) );
  nor2s1 _41564_inst ( .DIN1(_41359), .DIN2(_41538), .Q(_41055) );
  and2s1 _41565_inst ( .DIN1(_40839), .DIN2(_40819), .Q(_41537) );
  nnd2s1 _41566_inst ( .DIN1(_41539), .DIN2(_41380), .Q(_40819) );
  nor2s1 _41567_inst ( .DIN1(_41341), .DIN2(_41540), .Q(_41539) );
  nnd2s1 _41568_inst ( .DIN1(_41541), .DIN2(_41358), .Q(_40839) );
  nor2s1 _41569_inst ( .DIN1(_41540), .DIN2(_41542), .Q(_41541) );
  nor2s1 _41570_inst ( .DIN1(_41543), .DIN2(_41544), .Q(_41535) );
  nor2s1 _41571_inst ( .DIN1(_40942), .DIN2(_40653), .Q(_41544) );
  nnd2s1 _41572_inst ( .DIN1(_41545), .DIN2(_41546), .Q(_40942) );
  nor2s1 _41573_inst ( .DIN1(_41547), .DIN2(_41338), .Q(_41546) );
  nor2s1 _41574_inst ( .DIN1(_41396), .DIN2(_41548), .Q(_41545) );
  hi1s1 _41575_inst ( .DIN(_41358), .Q(_41548) );
  nor2s1 _41576_inst ( .DIN1(_41330), .DIN2(_40655), .Q(_41543) );
  nnd2s1 _41577_inst ( .DIN1(_41549), .DIN2(_41380), .Q(_40655) );
  nor2s1 _41578_inst ( .DIN1(_41026), .DIN2(_41550), .Q(_41514) );
  xor2s1 _41579_inst ( .DIN1(_31222), .DIN2(_41551), .Q(_41550) );
  nnd2s1 _41580_inst ( .DIN1(_41552), .DIN2(_41553), .Q(_41551) );
  nnd2s1 _41581_inst ( .DIN1(_41000), .DIN2(_41554), .Q(_41553) );
  nnd2s1 _41582_inst ( .DIN1(_41555), .DIN2(_41556), .Q(_41554) );
  nor2s1 _41583_inst ( .DIN1(_41210), .DIN2(_41557), .Q(_41556) );
  hi1s1 _41584_inst ( .DIN(_40974), .Q(_41557) );
  nnd2s1 _41585_inst ( .DIN1(_41558), .DIN2(_41559), .Q(_40974) );
  nor2s1 _41586_inst ( .DIN1(_38990), .DIN2(_34211), .Q(_41559) );
  nor2s1 _41587_inst ( .DIN1(_36336), .DIN2(_34762), .Q(_41558) );
  and2s1 _41588_inst ( .DIN1(_41560), .DIN2(_41511), .Q(_41210) );
  nor2s1 _41589_inst ( .DIN1(_36308), .DIN2(_41452), .Q(_41511) );
  nor2s1 _41590_inst ( .DIN1(_38990), .DIN2(_34193), .Q(_41560) );
  hi1s1 _41591_inst ( .DIN(_33945), .Q(_34193) );
  nor2s1 _41592_inst ( .DIN1(_41561), .DIN2(_41562), .Q(_41555) );
  nor2s1 _41593_inst ( .DIN1(_41448), .DIN2(_39133), .Q(_41562) );
  nor2s1 _41594_inst ( .DIN1(_41563), .DIN2(_34762), .Q(_41561) );
  nor2s1 _41595_inst ( .DIN1(_41564), .DIN2(_41420), .Q(_41563) );
  nor2s1 _41596_inst ( .DIN1(_41102), .DIN2(_33139), .Q(_41564) );
  nor2s1 _41597_inst ( .DIN1(_41565), .DIN2(_41566), .Q(_41552) );
  nor2s1 _41598_inst ( .DIN1(_41567), .DIN2(_40850), .Q(_41566) );
  nor2s1 _41599_inst ( .DIN1(_41568), .DIN2(_41569), .Q(_41567) );
  nor2s1 _41600_inst ( .DIN1(_41448), .DIN2(_39027), .Q(_41569) );
  nor2s1 _41601_inst ( .DIN1(_41415), .DIN2(_41570), .Q(_41568) );
  nnd2s1 _41602_inst ( .DIN1(_34017), .DIN2(_39255), .Q(_41570) );
  nor2s1 _41603_inst ( .DIN1(_41571), .DIN2(_40654), .Q(_41565) );
  nor2s1 _41604_inst ( .DIN1(_41572), .DIN2(_41573), .Q(_41571) );
  nor2s1 _41605_inst ( .DIN1(_34890), .DIN2(_41574), .Q(_41572) );
  nnd2s1 _41606_inst ( .DIN1(_41575), .DIN2(_41576), .Q(_41026) );
  nnd2s1 _41607_inst ( .DIN1(_41161), .DIN2(_41056), .Q(_41576) );
  and2s1 _41608_inst ( .DIN1(_41577), .DIN2(_41455), .Q(_41161) );
  hi1s1 _41609_inst ( .DIN(_41384), .Q(_41455) );
  nnd2s1 _41610_inst ( .DIN1(_33946), .DIN2(_38132), .Q(_41384) );
  hi1s1 _41611_inst ( .DIN(_38990), .Q(_38132) );
  hi1s1 _41612_inst ( .DIN(_41110), .Q(_41575) );
  nor2s1 _41613_inst ( .DIN1(_40576), .DIN2(_40699), .Q(_41110) );
  nnd2s1 _41614_inst ( .DIN1(_41529), .DIN2(_33930), .Q(_40576) );
  nor2s1 _41615_inst ( .DIN1(_41522), .DIN2(_34638), .Q(_41529) );
  nnd2s1 _41616_inst ( .DIN1(_41578), .DIN2(_41579), .Q(_41512) );
  nor2s1 _41617_inst ( .DIN1(_41580), .DIN2(_41431), .Q(_41579) );
  nor2s1 _41618_inst ( .DIN1(_40573), .DIN2(_41014), .Q(_41431) );
  nnd2s1 _41619_inst ( .DIN1(_41581), .DIN2(_34960), .Q(_41014) );
  nor2s1 _41620_inst ( .DIN1(_33139), .DIN2(_41485), .Q(_41581) );
  nor2s1 _41621_inst ( .DIN1(_40529), .DIN2(_40747), .Q(_41580) );
  nnd2s1 _41622_inst ( .DIN1(_41582), .DIN2(_41583), .Q(_40747) );
  nor2s1 _41623_inst ( .DIN1(_36337), .DIN2(_39026), .Q(_41583) );
  nor2s1 _41624_inst ( .DIN1(_41278), .DIN2(_40555), .Q(_41578) );
  nnd2s1 _41625_inst ( .DIN1(_41584), .DIN2(_41585), .Q(_40555) );
  nor2s1 _41626_inst ( .DIN1(_41586), .DIN2(_41587), .Q(_41585) );
  nnd2s1 _41627_inst ( .DIN1(_41588), .DIN2(_41589), .Q(_41587) );
  nnd2s1 _41628_inst ( .DIN1(_41090), .DIN2(_41079), .Q(_41589) );
  hi1s1 _41629_inst ( .DIN(_40582), .Q(_41090) );
  nnd2s1 _41630_inst ( .DIN1(_41590), .DIN2(_41451), .Q(_40582) );
  nor2s1 _41631_inst ( .DIN1(_33139), .DIN2(_34762), .Q(_41590) );
  nor2s1 _41632_inst ( .DIN1(_41591), .DIN2(_41592), .Q(_41588) );
  nor2s1 _41633_inst ( .DIN1(_26842), .DIN2(_40755), .Q(_41592) );
  nnd2s1 _41634_inst ( .DIN1(_41593), .DIN2(_33822), .Q(_40755) );
  hi1s1 _41635_inst ( .DIN(_34190), .Q(_33822) );
  nor2s1 _41636_inst ( .DIN1(_40857), .DIN2(_40849), .Q(_41591) );
  nnd2s1 _41637_inst ( .DIN1(_41594), .DIN2(_41595), .Q(_40849) );
  nor2s1 _41638_inst ( .DIN1(_26208), .DIN2(_41547), .Q(_41595) );
  nor2s1 _41639_inst ( .DIN1(_41596), .DIN2(_41597), .Q(_41594) );
  nnd2s1 _41640_inst ( .DIN1(_41598), .DIN2(_41599), .Q(_41586) );
  nor2s1 _41641_inst ( .DIN1(_41085), .DIN2(_40956), .Q(_41599) );
  and2s1 _41642_inst ( .DIN1(_41360), .DIN2(_40821), .Q(_40956) );
  nnd2s1 _41643_inst ( .DIN1(_40574), .DIN2(_40765), .Q(_40821) );
  nnd2s1 _41644_inst ( .DIN1(_41600), .DIN2(_40894), .Q(_40765) );
  nor2s1 _41645_inst ( .DIN1(_33825), .DIN2(_34638), .Q(_41600) );
  nnd2s1 _41646_inst ( .DIN1(_41601), .DIN2(_34642), .Q(_40574) );
  nor2s1 _41647_inst ( .DIN1(_34205), .DIN2(_41522), .Q(_41601) );
  or2s1 _41648_inst ( .DIN1(_33520), .DIN2(_27596), .Q(_41522) );
  hi1s1 _41649_inst ( .DIN(_40498), .Q(_41360) );
  hi1s1 _41650_inst ( .DIN(_40853), .Q(_41085) );
  nnd2s1 _41651_inst ( .DIN1(_41573), .DIN2(_41079), .Q(_40853) );
  and2s1 _41652_inst ( .DIN1(_41582), .DIN2(_41577), .Q(_41573) );
  nor2s1 _41653_inst ( .DIN1(_39027), .DIN2(_36337), .Q(_41577) );
  nor2s1 _41654_inst ( .DIN1(_38465), .DIN2(_41507), .Q(_41582) );
  hi1s1 _41655_inst ( .DIN(_33946), .Q(_41507) );
  nor2s1 _41656_inst ( .DIN1(_41602), .DIN2(_41603), .Q(_33946) );
  nor2s1 _41657_inst ( .DIN1(_40757), .DIN2(_41604), .Q(_41598) );
  hi1s1 _41658_inst ( .DIN(_41289), .Q(_41604) );
  nnd2s1 _41659_inst ( .DIN1(_41605), .DIN2(_41606), .Q(_41289) );
  nor2s1 _41660_inst ( .DIN1(_41341), .DIN2(_41607), .Q(_41606) );
  nnd2s1 _41661_inst ( .DIN1(_41608), .DIN2(_41340), .Q(_41607) );
  hi1s1 _41662_inst ( .DIN(_41609), .Q(_41340) );
  nor2s1 _41663_inst ( .DIN1(_40518), .DIN2(_40745), .Q(_41605) );
  and2s1 _41664_inst ( .DIN1(_41000), .DIN2(_41273), .Q(_40757) );
  and2s1 _41665_inst ( .DIN1(_39193), .DIN2(_41610), .Q(_41273) );
  hi1s1 _41666_inst ( .DIN(_40532), .Q(_41000) );
  nnd2s1 _41667_inst ( .DIN1(_41611), .DIN2(_40754), .Q(_40532) );
  xor2s1 _41668_inst ( .DIN1(_31569), .DIN2(_41612), .Q(_41611) );
  nor2s1 _41669_inst ( .DIN1(_41613), .DIN2(_41614), .Q(_41584) );
  nnd2s1 _41670_inst ( .DIN1(_41615), .DIN2(_41616), .Q(_41614) );
  hi1s1 _41671_inst ( .DIN(_40914), .Q(_41616) );
  nnd2s1 _41672_inst ( .DIN1(_41617), .DIN2(_41618), .Q(_40914) );
  nor2s1 _41673_inst ( .DIN1(_41299), .DIN2(_40698), .Q(_41618) );
  nor2s1 _41674_inst ( .DIN1(_40777), .DIN2(_40642), .Q(_40698) );
  nnd2s1 _41675_inst ( .DIN1(_41306), .DIN2(_41619), .Q(_40642) );
  and2s1 _41676_inst ( .DIN1(_41073), .DIN2(_40754), .Q(_41299) );
  nor2s1 _41677_inst ( .DIN1(_41542), .DIN2(_41383), .Q(_41073) );
  hi1s1 _41678_inst ( .DIN(_41306), .Q(_41542) );
  nor2s1 _41679_inst ( .DIN1(_41076), .DIN2(_41620), .Q(_41617) );
  xor2s1 _41680_inst ( .DIN1(_28613), .DIN2(_41621), .Q(_41620) );
  nnd2s1 _41681_inst ( .DIN1(_41241), .DIN2(_41622), .Q(_41621) );
  nnd2s1 _41682_inst ( .DIN1(_40638), .DIN2(_41002), .Q(_41622) );
  hi1s1 _41683_inst ( .DIN(_41288), .Q(_40638) );
  nnd2s1 _41684_inst ( .DIN1(_41623), .DIN2(_41358), .Q(_41288) );
  nor2s1 _41685_inst ( .DIN1(_41624), .DIN2(_41603), .Q(_41358) );
  nor2s1 _41686_inst ( .DIN1(_41540), .DIN2(_41359), .Q(_41623) );
  nnd2s1 _41687_inst ( .DIN1(_41625), .DIN2(_53401), .Q(_41359) );
  nnd2s1 _41688_inst ( .DIN1(_40993), .DIN2(_41056), .Q(_41241) );
  hi1s1 _41689_inst ( .DIN(_41405), .Q(_40993) );
  nnd2s1 _41690_inst ( .DIN1(_41380), .DIN2(_41307), .Q(_41405) );
  nnd2s1 _41691_inst ( .DIN1(_41626), .DIN2(_41427), .Q(_41076) );
  nnd2s1 _41692_inst ( .DIN1(_41175), .DIN2(_40495), .Q(_41427) );
  hi1s1 _41693_inst ( .DIN(_41304), .Q(_41175) );
  nnd2s1 _41694_inst ( .DIN1(_41627), .DIN2(_41395), .Q(_41304) );
  nor2s1 _41695_inst ( .DIN1(_53407), .DIN2(_41609), .Q(_41627) );
  or2s1 _41696_inst ( .DIN1(_40778), .DIN2(_40777), .Q(_41626) );
  nnd2s1 _41697_inst ( .DIN1(_41628), .DIN2(_41629), .Q(_40778) );
  nor2s1 _41698_inst ( .DIN1(_26208), .DIN2(_41630), .Q(_41629) );
  nor2s1 _41699_inst ( .DIN1(_41596), .DIN2(_41383), .Q(_41628) );
  nnd2s1 _41700_inst ( .DIN1(_41631), .DIN2(_41608), .Q(_41383) );
  nor2s1 _41701_inst ( .DIN1(_41632), .DIN2(_41633), .Q(_41631) );
  nor2s1 _41702_inst ( .DIN1(_41262), .DIN2(_41047), .Q(_41615) );
  nnd2s1 _41703_inst ( .DIN1(_41634), .DIN2(_41635), .Q(_41047) );
  nor2s1 _41704_inst ( .DIN1(_41636), .DIN2(_41637), .Q(_41635) );
  or2s1 _41705_inst ( .DIN1(_40860), .DIN2(_41188), .Q(_41637) );
  or2s1 _41706_inst ( .DIN1(_41416), .DIN2(_40779), .Q(_41188) );
  nor2s1 _41707_inst ( .DIN1(_40850), .DIN2(_40580), .Q(_40779) );
  nnd2s1 _41708_inst ( .DIN1(_41638), .DIN2(_40902), .Q(_40580) );
  nnd2s1 _41709_inst ( .DIN1(_41639), .DIN2(_41640), .Q(_41416) );
  nnd2s1 _41710_inst ( .DIN1(_41641), .DIN2(_41451), .Q(_41640) );
  nor2s1 _41711_inst ( .DIN1(_40529), .DIN2(_41436), .Q(_41641) );
  nnd2s1 _41712_inst ( .DIN1(_33934), .DIN2(_27653), .Q(_41436) );
  hi1s1 _41713_inst ( .DIN(_34191), .Q(_33934) );
  nnd2s1 _41714_inst ( .DIN1(_39383), .DIN2(_41242), .Q(_41639) );
  hi1s1 _41715_inst ( .DIN(_40748), .Q(_41242) );
  nnd2s1 _41716_inst ( .DIN1(_41642), .DIN2(_41329), .Q(_39537) );
  hi1s1 _41717_inst ( .DIN(_41643), .Q(_41329) );
  nnd2s1 _41718_inst ( .DIN1(_41644), .DIN2(_41645), .Q(_40860) );
  nnd2s1 _41719_inst ( .DIN1(_41646), .DIN2(_40856), .Q(_41645) );
  nor2s1 _41720_inst ( .DIN1(_34893), .DIN2(_40850), .Q(_41646) );
  nnd2s1 _41721_inst ( .DIN1(_40754), .DIN2(_41647), .Q(_40850) );
  nnd2s1 _41722_inst ( .DIN1(_41648), .DIN2(______[8]), .Q(_41647) );
  nor2s1 _41723_inst ( .DIN1(______[26]), .DIN2(______[15]), .Q(_41648) );
  nnd2s1 _41724_inst ( .DIN1(_41649), .DIN2(_39031), .Q(_41644) );
  hi1s1 _41725_inst ( .DIN(_39133), .Q(_39031) );
  nor2s1 _41726_inst ( .DIN1(_41448), .DIN2(_40777), .Q(_41649) );
  hi1s1 _41727_inst ( .DIN(_40546), .Q(_40777) );
  nnd2s1 _41728_inst ( .DIN1(_40832), .DIN2(_41650), .Q(_41636) );
  nnd2s1 _41729_inst ( .DIN1(_40897), .DIN2(_39969), .Q(_41650) );
  hi1s1 _41730_inst ( .DIN(_41313), .Q(_40897) );
  nnd2s1 _41731_inst ( .DIN1(_41500), .DIN2(_41651), .Q(_41313) );
  nor2s1 _41732_inst ( .DIN1(_39032), .DIN2(_41652), .Q(_41651) );
  nnd2s1 _41733_inst ( .DIN1(_33821), .DIN2(_40754), .Q(_41652) );
  hi1s1 _41734_inst ( .DIN(_40682), .Q(_40832) );
  xor2s1 _41735_inst ( .DIN1(_34235), .DIN2(_41653), .Q(_40682) );
  nor2s1 _41736_inst ( .DIN1(_41424), .DIN2(_41574), .Q(_41653) );
  nor2s1 _41737_inst ( .DIN1(_40676), .DIN2(_41654), .Q(_41634) );
  nnd2s1 _41738_inst ( .DIN1(_41655), .DIN2(_40916), .Q(_41654) );
  and2s1 _41739_inst ( .DIN1(_41656), .DIN2(_41657), .Q(_40916) );
  nnd2s1 _41740_inst ( .DIN1(_41428), .DIN2(_40754), .Q(_41657) );
  hi1s1 _41741_inst ( .DIN(_40652), .Q(_41428) );
  nnd2s1 _41742_inst ( .DIN1(_41625), .DIN2(_41395), .Q(_40652) );
  nor2s1 _41743_inst ( .DIN1(_53407), .DIN2(_41658), .Q(_41625) );
  nnd2s1 _41744_inst ( .DIN1(_41176), .DIN2(_40495), .Q(_41656) );
  and2s1 _41745_inst ( .DIN1(_41659), .DIN2(_41660), .Q(_41176) );
  nor2s1 _41746_inst ( .DIN1(_53414), .DIN2(_26208), .Q(_41660) );
  nor2s1 _41747_inst ( .DIN1(_41596), .DIN2(_41661), .Q(_41659) );
  hi1s1 _41748_inst ( .DIN(_40976), .Q(_41655) );
  nnd2s1 _41749_inst ( .DIN1(_41467), .DIN2(_41662), .Q(_40976) );
  or2s1 _41750_inst ( .DIN1(_40810), .DIN2(_41131), .Q(_41662) );
  nnd2s1 _41751_inst ( .DIN1(_41663), .DIN2(_34765), .Q(_40810) );
  nor2s1 _41752_inst ( .DIN1(_41643), .DIN2(_34204), .Q(_41663) );
  nnd2s1 _41753_inst ( .DIN1(_41593), .DIN2(_41664), .Q(_41467) );
  nor2s1 _41754_inst ( .DIN1(_26842), .DIN2(_34211), .Q(_41664) );
  nor2s1 _41755_inst ( .DIN1(_39026), .DIN2(_41485), .Q(_41593) );
  hi1s1 _41756_inst ( .DIN(_41435), .Q(_41485) );
  nor2s1 _41757_inst ( .DIN1(_36336), .DIN2(_38466), .Q(_41435) );
  nnd2s1 _41758_inst ( .DIN1(_41665), .DIN2(_41666), .Q(_40676) );
  nnd2s1 _41759_inst ( .DIN1(_41667), .DIN2(_41668), .Q(_41666) );
  nor2s1 _41760_inst ( .DIN1(_33139), .DIN2(_41669), .Q(_41668) );
  nnd2s1 _41761_inst ( .DIN1(_40971), .DIN2(_41670), .Q(_41669) );
  hi1s1 _41762_inst ( .DIN(_40857), .Q(_40971) );
  nor2s1 _41763_inst ( .DIN1(_38465), .DIN2(_39133), .Q(_41667) );
  nnd2s1 _41764_inst ( .DIN1(_41437), .DIN2(_41056), .Q(_41665) );
  hi1s1 _41765_inst ( .DIN(_41131), .Q(_41056) );
  and2s1 _41766_inst ( .DIN1(_41500), .DIN2(_41638), .Q(_41437) );
  nor2s1 _41767_inst ( .DIN1(_34205), .DIN2(_34893), .Q(_41638) );
  nor2s1 _41768_inst ( .DIN1(_33518), .DIN2(_34913), .Q(_41500) );
  nnd2s1 _41769_inst ( .DIN1(_41671), .DIN2(_41672), .Q(_41262) );
  nor2s1 _41770_inst ( .DIN1(_40675), .DIN2(_41673), .Q(_41672) );
  nnd2s1 _41771_inst ( .DIN1(_41674), .DIN2(_41675), .Q(_41673) );
  nnd2s1 _41772_inst ( .DIN1(_40834), .DIN2(_40889), .Q(_41675) );
  hi1s1 _41773_inst ( .DIN(_41063), .Q(_40889) );
  nnd2s1 _41774_inst ( .DIN1(_41676), .DIN2(_41530), .Q(_41063) );
  nor2s1 _41775_inst ( .DIN1(_39032), .DIN2(_41254), .Q(_41676) );
  hi1s1 _41776_inst ( .DIN(_41206), .Q(_41674) );
  nnd2s1 _41777_inst ( .DIN1(_41677), .DIN2(_41678), .Q(_41206) );
  nnd2s1 _41778_inst ( .DIN1(_41679), .DIN2(_41498), .Q(_41678) );
  nor2s1 _41779_inst ( .DIN1(_41680), .DIN2(_33139), .Q(_41679) );
  nor2s1 _41780_inst ( .DIN1(_41681), .DIN2(_41682), .Q(_41680) );
  nor2s1 _41781_inst ( .DIN1(_27630), .DIN2(_40649), .Q(_41682) );
  nnd2s1 _41782_inst ( .DIN1(_41683), .DIN2(_41684), .Q(_40649) );
  hi1s1 _41783_inst ( .DIN(_27653), .Q(_27630) );
  nor2s1 _41784_inst ( .DIN1(_41452), .DIN2(_40857), .Q(_41681) );
  or2s1 _41785_inst ( .DIN1(_41490), .DIN2(_40543), .Q(_41677) );
  nnd2s1 _41786_inst ( .DIN1(_41685), .DIN2(_41451), .Q(_41490) );
  nor2s1 _41787_inst ( .DIN1(_41414), .DIN2(_34890), .Q(_41685) );
  nnd2s1 _41788_inst ( .DIN1(_41686), .DIN2(_41687), .Q(_40675) );
  nnd2s1 _41789_inst ( .DIN1(_41688), .DIN2(_41402), .Q(_41687) );
  hi1s1 _41790_inst ( .DIN(_41461), .Q(_41402) );
  nnd2s1 _41791_inst ( .DIN1(_41689), .DIN2(_33275), .Q(_41461) );
  nor2s1 _41792_inst ( .DIN1(_38466), .DIN2(_36308), .Q(_41689) );
  nor2s1 _41793_inst ( .DIN1(_40529), .DIN2(_39133), .Q(_41688) );
  nnd2s1 _41794_inst ( .DIN1(_41690), .DIN2(_41691), .Q(_39133) );
  nor2s1 _41795_inst ( .DIN1(_41692), .DIN2(_41693), .Q(_41686) );
  nor2s1 _41796_inst ( .DIN1(_41385), .DIN2(_41694), .Q(_41693) );
  nnd2s1 _41797_inst ( .DIN1(_34017), .DIN2(_41695), .Q(_41694) );
  nnd2s1 _41798_inst ( .DIN1(_41696), .DIN2(_40546), .Q(_41385) );
  nor2s1 _41799_inst ( .DIN1(_36308), .DIN2(_34890), .Q(_41696) );
  nor2s1 _41800_inst ( .DIN1(_41697), .DIN2(_41698), .Q(_41692) );
  nnd2s1 _41801_inst ( .DIN1(_41530), .DIN2(_40639), .Q(_41698) );
  hi1s1 _41802_inst ( .DIN(_40745), .Q(_40639) );
  nnd2s1 _41803_inst ( .DIN1(_34766), .DIN2(_40902), .Q(_41697) );
  nor2s1 _41804_inst ( .DIN1(_40599), .DIN2(_41699), .Q(_41671) );
  or2s1 _41805_inst ( .DIN1(_41189), .DIN2(_41373), .Q(_41699) );
  nnd2s1 _41806_inst ( .DIN1(_40588), .DIN2(_41700), .Q(_41373) );
  nnd2s1 _41807_inst ( .DIN1(_41701), .DIN2(_41152), .Q(_41700) );
  nor2s1 _41808_inst ( .DIN1(_34204), .DIN2(_34638), .Q(_41152) );
  nor2s1 _41809_inst ( .DIN1(_41131), .DIN2(_41153), .Q(_41701) );
  nnd2s1 _41810_inst ( .DIN1(_41702), .DIN2(_40856), .Q(_40588) );
  nor2s1 _41811_inst ( .DIN1(_41153), .DIN2(_33931), .Q(_40856) );
  nnd2s1 _41812_inst ( .DIN1(_41703), .DIN2(_41704), .Q(_33931) );
  hi1s1 _41813_inst ( .DIN(_41510), .Q(_41153) );
  nor2s1 _41814_inst ( .DIN1(_34913), .DIN2(_33520), .Q(_41510) );
  nor2s1 _41815_inst ( .DIN1(_40498), .DIN2(_39032), .Q(_41702) );
  nnd2s1 _41816_inst ( .DIN1(_41705), .DIN2(_41706), .Q(_41189) );
  nnd2s1 _41817_inst ( .DIN1(_41707), .DIN2(_34960), .Q(_41706) );
  hi1s1 _41818_inst ( .DIN(_39027), .Q(_34960) );
  nnd2s1 _41819_inst ( .DIN1(_41708), .DIN2(_41690), .Q(_39027) );
  nor2s1 _41820_inst ( .DIN1(_41448), .DIN2(_40857), .Q(_41707) );
  hi1s1 _41821_inst ( .DIN(_41068), .Q(_41448) );
  nor2s1 _41822_inst ( .DIN1(_41414), .DIN2(_41102), .Q(_41068) );
  nnd2s1 _41823_inst ( .DIN1(_41670), .DIN2(_41695), .Q(_41102) );
  hi1s1 _41824_inst ( .DIN(_38466), .Q(_41695) );
  hi1s1 _41825_inst ( .DIN(_36337), .Q(_41670) );
  nnd2s1 _41826_inst ( .DIN1(_41709), .DIN2(_53406), .Q(_36337) );
  nor2s1 _41827_inst ( .DIN1(_53407), .DIN2(_26283), .Q(_41709) );
  hi1s1 _41828_inst ( .DIN(_33275), .Q(_41414) );
  nor2s1 _41829_inst ( .DIN1(_41602), .DIN2(_41633), .Q(_33275) );
  nnd2s1 _41830_inst ( .DIN1(_39193), .DIN2(_41710), .Q(_41705) );
  nnd2s1 _41831_inst ( .DIN1(_41711), .DIN2(_41712), .Q(_41710) );
  nnd2s1 _41832_inst ( .DIN1(_41713), .DIN2(_40834), .Q(_41712) );
  hi1s1 _41833_inst ( .DIN(_40896), .Q(_40834) );
  nor2s1 _41834_inst ( .DIN1(_41415), .DIN2(_34190), .Q(_41713) );
  nnd2s1 _41835_inst ( .DIN1(_41714), .DIN2(_41715), .Q(_34190) );
  hi1s1 _41836_inst ( .DIN(_41498), .Q(_41415) );
  nnd2s1 _41837_inst ( .DIN1(_41420), .DIN2(_40495), .Q(_41711) );
  hi1s1 _41838_inst ( .DIN(_40529), .Q(_40495) );
  hi1s1 _41839_inst ( .DIN(_41574), .Q(_41420) );
  nnd2s1 _41840_inst ( .DIN1(_41451), .DIN2(_33945), .Q(_41574) );
  nor2s1 _41841_inst ( .DIN1(_41633), .DIN2(_41716), .Q(_33945) );
  nor2s1 _41842_inst ( .DIN1(_38465), .DIN2(_36308), .Q(_41451) );
  hi1s1 _41843_inst ( .DIN(_39026), .Q(_39193) );
  nnd2s1 _41844_inst ( .DIN1(_41708), .DIN2(_41717), .Q(_39026) );
  nnd2s1 _41845_inst ( .DIN1(_41718), .DIN2(_41719), .Q(_40599) );
  nnd2s1 _41846_inst ( .DIN1(_41720), .DIN2(_41721), .Q(_41719) );
  nor2s1 _41847_inst ( .DIN1(_38990), .DIN2(_36336), .Q(_41721) );
  nor2s1 _41848_inst ( .DIN1(_34191), .DIN2(_41424), .Q(_41720) );
  nnd2s1 _41849_inst ( .DIN1(_34891), .DIN2(_40546), .Q(_41424) );
  nor2s1 _41850_inst ( .DIN1(_41612), .DIN2(_26842), .Q(_40546) );
  nnd2s1 _41851_inst ( .DIN1(_41722), .DIN2(______[15]), .Q(_41612) );
  hi1s1 _41852_inst ( .DIN(_34762), .Q(_34891) );
  nnd2s1 _41853_inst ( .DIN1(_41691), .DIN2(_41723), .Q(_34762) );
  nnd2s1 _41854_inst ( .DIN1(_41724), .DIN2(_40894), .Q(_41718) );
  nor2s1 _41855_inst ( .DIN1(_27596), .DIN2(_41725), .Q(_40894) );
  nor2s1 _41856_inst ( .DIN1(_40895), .DIN2(_40653), .Q(_41724) );
  nnd2s1 _41857_inst ( .DIN1(_34531), .DIN2(_33821), .Q(_40895) );
  hi1s1 _41858_inst ( .DIN(_39301), .Q(_34531) );
  nnd2s1 _41859_inst ( .DIN1(_41726), .DIN2(_41727), .Q(_41613) );
  hi1s1 _41860_inst ( .DIN(_40861), .Q(_41727) );
  nnd2s1 _41861_inst ( .DIN1(_41728), .DIN2(_41729), .Q(_40861) );
  nnd2s1 _41862_inst ( .DIN1(_41079), .DIN2(_40887), .Q(_41729) );
  nnd2s1 _41863_inst ( .DIN1(_41311), .DIN2(_41106), .Q(_40887) );
  nnd2s1 _41864_inst ( .DIN1(_41730), .DIN2(_41530), .Q(_41106) );
  hi1s1 _41865_inst ( .DIN(_33825), .Q(_41530) );
  nnd2s1 _41866_inst ( .DIN1(_41731), .DIN2(_53409), .Q(_33825) );
  xor2s1 _41867_inst ( .DIN1(_34338), .DIN2(_41732), .Q(_41730) );
  nor2s1 _41868_inst ( .DIN1(_39301), .DIN2(_41254), .Q(_41732) );
  nnd2s1 _41869_inst ( .DIN1(_41733), .DIN2(_41734), .Q(_39301) );
  nnd2s1 _41870_inst ( .DIN1(_41642), .DIN2(_41129), .Q(_41311) );
  nor2s1 _41871_inst ( .DIN1(_34205), .DIN2(_34638), .Q(_41642) );
  hi1s1 _41872_inst ( .DIN(_34766), .Q(_34638) );
  xor2s1 _41873_inst ( .DIN1(_41735), .DIN2(_30912), .Q(_34766) );
  nnd2s1 _41874_inst ( .DIN1(_41690), .DIN2(_41736), .Q(_41735) );
  hi1s1 _41875_inst ( .DIN(_33821), .Q(_34205) );
  nor2s1 _41876_inst ( .DIN1(_41632), .DIN2(_41603), .Q(_33821) );
  or2s1 _41877_inst ( .DIN1(_40498), .DIN2(_40975), .Q(_41728) );
  nnd2s1 _41878_inst ( .DIN1(_39255), .DIN2(_41610), .Q(_40975) );
  and2s1 _41879_inst ( .DIN1(_41737), .DIN2(_36310), .Q(_41610) );
  xor2s1 _41880_inst ( .DIN1(_32362), .DIN2(_41738), .Q(_41737) );
  nor2s1 _41881_inst ( .DIN1(_34211), .DIN2(_38466), .Q(_41738) );
  nnd2s1 _41882_inst ( .DIN1(_41739), .DIN2(_53405), .Q(_38466) );
  hi1s1 _41883_inst ( .DIN(_33932), .Q(_34211) );
  xor2s1 _41884_inst ( .DIN1(_41740), .DIN2(_29168), .Q(_33932) );
  hi1s1 _41885_inst ( .DIN(_32657), .Q(_29168) );
  nnd2s1 _41886_inst ( .DIN1(_41731), .DIN2(_26578), .Q(_41740) );
  nor2s1 _41887_inst ( .DIN1(_41602), .DIN2(_53411), .Q(_41731) );
  or2s1 _41888_inst ( .DIN1(_53410), .DIN2(_53412), .Q(_41602) );
  hi1s1 _41889_inst ( .DIN(_41452), .Q(_39255) );
  nnd2s1 _41890_inst ( .DIN1(_41733), .DIN2(_41708), .Q(_41452) );
  nor2s1 _41891_inst ( .DIN1(_26443), .DIN2(_26274), .Q(_41708) );
  nor2s1 _41892_inst ( .DIN1(_41741), .DIN2(_41366), .Q(_41726) );
  xnr2s1 _41893_inst ( .DIN1(_41742), .DIN2(_31975), .Q(_41366) );
  nnd2s1 _41894_inst ( .DIN1(_41037), .DIN2(_41255), .Q(_41742) );
  nnd2s1 _41895_inst ( .DIN1(_40748), .DIN2(_40543), .Q(_41255) );
  nnd2s1 _41896_inst ( .DIN1(_41743), .DIN2(_41684), .Q(_40543) );
  nnd2s1 _41897_inst ( .DIN1(_40754), .DIN2(_41744), .Q(_40748) );
  nnd2s1 _41898_inst ( .DIN1(_41745), .DIN2(______[26]), .Q(_41744) );
  nor2s1 _41899_inst ( .DIN1(______[8]), .DIN2(______[15]), .Q(_41745) );
  and2s1 _41900_inst ( .DIN1(_41746), .DIN2(_41498), .Q(_41037) );
  nor2s1 _41901_inst ( .DIN1(_38465), .DIN2(_36336), .Q(_41498) );
  nnd2s1 _41902_inst ( .DIN1(_41747), .DIN2(_53407), .Q(_36336) );
  nnd2s1 _41903_inst ( .DIN1(_41748), .DIN2(_53402), .Q(_38465) );
  nor2s1 _41904_inst ( .DIN1(_53405), .DIN2(_26218), .Q(_41748) );
  nor2s1 _41905_inst ( .DIN1(_34890), .DIN2(_34191), .Q(_41746) );
  nnd2s1 _41906_inst ( .DIN1(_41749), .DIN2(_41703), .Q(_34191) );
  nnd2s1 _41907_inst ( .DIN1(_41734), .DIN2(_41690), .Q(_34890) );
  and2s1 _41908_inst ( .DIN1(_53408), .DIN2(_53403), .Q(_41690) );
  nor2s1 _41909_inst ( .DIN1(_40575), .DIN2(_40913), .Q(_41741) );
  nnd2s1 _41910_inst ( .DIN1(_41750), .DIN2(_40902), .Q(_40913) );
  nor2s1 _41911_inst ( .DIN1(_34204), .DIN2(_39257), .Q(_41750) );
  hi1s1 _41912_inst ( .DIN(_41002), .Q(_40575) );
  nnd2s1 _41913_inst ( .DIN1(_40745), .DIN2(_40699), .Q(_41002) );
  nnd2s1 _41914_inst ( .DIN1(_41751), .DIN2(______[26]), .Q(_40699) );
  nnd2s1 _41915_inst ( .DIN1(_40754), .DIN2(_41752), .Q(_40745) );
  nnd2s1 _41916_inst ( .DIN1(_41743), .DIN2(______[15]), .Q(_41752) );
  nor2s1 _41917_inst ( .DIN1(______[8]), .DIN2(_27365), .Q(_41743) );
  nnd2s1 _41918_inst ( .DIN1(_41753), .DIN2(_41754), .Q(_41278) );
  nor2s1 _41919_inst ( .DIN1(_41755), .DIN2(_41756), .Q(_41754) );
  nnd2s1 _41920_inst ( .DIN1(_41344), .DIN2(_41213), .Q(_41756) );
  nnd2s1 _41921_inst ( .DIN1(_41757), .DIN2(_41758), .Q(_41213) );
  hi1s1 _41922_inst ( .DIN(_41327), .Q(_41758) );
  nnd2s1 _41923_inst ( .DIN1(_34642), .DIN2(_33930), .Q(_41327) );
  hi1s1 _41924_inst ( .DIN(_34204), .Q(_33930) );
  nnd2s1 _41925_inst ( .DIN1(_41714), .DIN2(_41704), .Q(_34204) );
  hi1s1 _41926_inst ( .DIN(_41632), .Q(_41704) );
  nnd2s1 _41927_inst ( .DIN1(_53412), .DIN2(_53410), .Q(_41632) );
  hi1s1 _41928_inst ( .DIN(_34893), .Q(_34642) );
  nnd2s1 _41929_inst ( .DIN1(_41734), .DIN2(_41717), .Q(_34893) );
  nor2s1 _41930_inst ( .DIN1(_53401), .DIN2(_53414), .Q(_41734) );
  nor2s1 _41931_inst ( .DIN1(_41643), .DIN2(_40654), .Q(_41757) );
  nnd2s1 _41932_inst ( .DIN1(_40754), .DIN2(_41759), .Q(_40654) );
  nnd2s1 _41933_inst ( .DIN1(_41760), .DIN2(______[15]), .Q(_41759) );
  nnd2s1 _41934_inst ( .DIN1(_38133), .DIN2(_36530), .Q(_41643) );
  hi1s1 _41935_inst ( .DIN(_37778), .Q(_36530) );
  hi1s1 _41936_inst ( .DIN(_41725), .Q(_38133) );
  nnd2s1 _41937_inst ( .DIN1(_41761), .DIN2(_41762), .Q(_41344) );
  nor2s1 _41938_inst ( .DIN1(_40498), .DIN2(_41235), .Q(_41761) );
  hi1s1 _41939_inst ( .DIN(_41129), .Q(_41235) );
  xor2s1 _41940_inst ( .DIN1(_41763), .DIN2(_27093), .Q(_41129) );
  nnd2s1 _41941_inst ( .DIN1(_38314), .DIN2(_27585), .Q(_41763) );
  hi1s1 _41942_inst ( .DIN(_27596), .Q(_27585) );
  nnd2s1 _41943_inst ( .DIN1(_41764), .DIN2(_53406), .Q(_27596) );
  nor2s1 _41944_inst ( .DIN1(_26208), .DIN2(_26283), .Q(_41764) );
  hi1s1 _41945_inst ( .DIN(_33518), .Q(_38314) );
  nnd2s1 _41946_inst ( .DIN1(_41765), .DIN2(_53404), .Q(_33518) );
  nor2s1 _41947_inst ( .DIN1(_53402), .DIN2(_26240), .Q(_41765) );
  nor2s1 _41948_inst ( .DIN1(_41254), .DIN2(_41766), .Q(_41755) );
  nnd2s1 _41949_inst ( .DIN1(_41762), .DIN2(_41079), .Q(_41766) );
  hi1s1 _41950_inst ( .DIN(_41330), .Q(_41079) );
  nnd2s1 _41951_inst ( .DIN1(_41751), .DIN2(_26809), .Q(_41330) );
  and2s1 _41952_inst ( .DIN1(_41767), .DIN2(______[15]), .Q(_41751) );
  nor2s1 _41953_inst ( .DIN1(______[8]), .DIN2(_26842), .Q(_41767) );
  hi1s1 _41954_inst ( .DIN(_40903), .Q(_41762) );
  nnd2s1 _41955_inst ( .DIN1(_34894), .DIN2(_33824), .Q(_40903) );
  hi1s1 _41956_inst ( .DIN(_41253), .Q(_33824) );
  hi1s1 _41957_inst ( .DIN(_39032), .Q(_34894) );
  nnd2s1 _41958_inst ( .DIN1(_41717), .DIN2(_41691), .Q(_39032) );
  hi1s1 _41959_inst ( .DIN(_41630), .Q(_41691) );
  hi1s1 _41960_inst ( .DIN(_40902), .Q(_41254) );
  nor2s1 _41961_inst ( .DIN1(_34913), .DIN2(_41725), .Q(_40902) );
  nnd2s1 _41962_inst ( .DIN1(_41768), .DIN2(_53402), .Q(_41725) );
  nor2s1 _41963_inst ( .DIN1(_26240), .DIN2(_26218), .Q(_41768) );
  nnd2s1 _41964_inst ( .DIN1(_41747), .DIN2(_26208), .Q(_34913) );
  nor2s1 _41965_inst ( .DIN1(_53400), .DIN2(_53406), .Q(_41747) );
  nor2s1 _41966_inst ( .DIN1(_40918), .DIN2(_41439), .Q(_41753) );
  nnd2s1 _41967_inst ( .DIN1(_41769), .DIN2(_41770), .Q(_41439) );
  nnd2s1 _41968_inst ( .DIN1(_41771), .DIN2(_41772), .Q(_41770) );
  nor2s1 _41969_inst ( .DIN1(_40857), .DIN2(_41773), .Q(_41772) );
  nnd2s1 _41970_inst ( .DIN1(_36310), .DIN2(_27653), .Q(_41773) );
  nor2s1 _41971_inst ( .DIN1(_41658), .DIN2(_53401), .Q(_27653) );
  hi1s1 _41972_inst ( .DIN(_36308), .Q(_36310) );
  nnd2s1 _41973_inst ( .DIN1(_41774), .DIN2(_53400), .Q(_36308) );
  nor2s1 _41974_inst ( .DIN1(_53406), .DIN2(_26208), .Q(_41774) );
  nnd2s1 _41975_inst ( .DIN1(_41722), .DIN2(_41684), .Q(_40857) );
  nor2s1 _41976_inst ( .DIN1(______[26]), .DIN2(_27066), .Q(_41722) );
  nor2s1 _41977_inst ( .DIN1(_38990), .DIN2(_33139), .Q(_41771) );
  hi1s1 _41978_inst ( .DIN(_34017), .Q(_33139) );
  nor2s1 _41979_inst ( .DIN1(_41624), .DIN2(_41633), .Q(_34017) );
  nnd2s1 _41980_inst ( .DIN1(_53411), .DIN2(_26578), .Q(_41633) );
  hi1s1 _41981_inst ( .DIN(_41749), .Q(_41624) );
  nnd2s1 _41982_inst ( .DIN1(_41739), .DIN2(_26240), .Q(_38990) );
  nor2s1 _41983_inst ( .DIN1(_53402), .DIN2(_53404), .Q(_41739) );
  nnd2s1 _41984_inst ( .DIN1(_41775), .DIN2(_41776), .Q(_41769) );
  hi1s1 _41985_inst ( .DIN(_41240), .Q(_41776) );
  nnd2s1 _41986_inst ( .DIN1(_41777), .DIN2(_34765), .Q(_41240) );
  hi1s1 _41987_inst ( .DIN(_39257), .Q(_34765) );
  nnd2s1 _41988_inst ( .DIN1(_41736), .DIN2(_41717), .Q(_39257) );
  nor2s1 _41989_inst ( .DIN1(_53403), .DIN2(_53408), .Q(_41717) );
  hi1s1 _41990_inst ( .DIN(_41547), .Q(_41736) );
  nor2s1 _41991_inst ( .DIN1(_37778), .DIN2(_41253), .Q(_41777) );
  nnd2s1 _41992_inst ( .DIN1(_41703), .DIN2(_41715), .Q(_41253) );
  hi1s1 _41993_inst ( .DIN(_41716), .Q(_41715) );
  nor2s1 _41994_inst ( .DIN1(_26578), .DIN2(_53411), .Q(_41703) );
  nnd2s1 _41995_inst ( .DIN1(_41778), .DIN2(_53400), .Q(_37778) );
  nor2s1 _41996_inst ( .DIN1(_53406), .DIN2(_53407), .Q(_41778) );
  nor2s1 _41997_inst ( .DIN1(_33520), .DIN2(_41131), .Q(_41775) );
  nnd2s1 _41998_inst ( .DIN1(_40754), .DIN2(_41779), .Q(_41131) );
  nnd2s1 _41999_inst ( .DIN1(_41780), .DIN2(______[26]), .Q(_41779) );
  nor2s1 _42000_inst ( .DIN1(______[15]), .DIN2(_27066), .Q(_41780) );
  nnd2s1 _42001_inst ( .DIN1(_41781), .DIN2(_53402), .Q(_33520) );
  nor2s1 _42002_inst ( .DIN1(_53404), .DIN2(_53405), .Q(_41781) );
  nnd2s1 _42003_inst ( .DIN1(_41782), .DIN2(_41783), .Q(_40918) );
  or2s1 _42004_inst ( .DIN1(_41059), .DIN2(_41062), .Q(_41783) );
  hi1s1 _42005_inst ( .DIN(_40938), .Q(_41062) );
  nnd2s1 _42006_inst ( .DIN1(_40653), .DIN2(_40896), .Q(_40938) );
  nnd2s1 _42007_inst ( .DIN1(_41784), .DIN2(_40754), .Q(_40896) );
  hi1s1 _42008_inst ( .DIN(_40888), .Q(_40653) );
  xor2s1 _42009_inst ( .DIN1(_32753), .DIN2(_41785), .Q(_40888) );
  nor2s1 _42010_inst ( .DIN1(_41784), .DIN2(_26842), .Q(_41785) );
  and2s1 _42011_inst ( .DIN1(_41683), .DIN2(______[15]), .Q(_41784) );
  nor2s1 _42012_inst ( .DIN1(_27066), .DIN2(_27365), .Q(_41683) );
  nnd2s1 _42013_inst ( .DIN1(_41549), .DIN2(_41306), .Q(_41059) );
  nor2s1 _42014_inst ( .DIN1(_40518), .DIN2(_41658), .Q(_41306) );
  nnd2s1 _42015_inst ( .DIN1(_53401), .DIN2(_53407), .Q(_40518) );
  nor2s1 _42016_inst ( .DIN1(_41338), .DIN2(_41341), .Q(_41549) );
  nor2s1 _42017_inst ( .DIN1(_41786), .DIN2(_41787), .Q(_41782) );
  nor2s1 _42018_inst ( .DIN1(_40573), .DIN2(_41195), .Q(_41787) );
  nnd2s1 _42019_inst ( .DIN1(_41380), .DIN2(_41619), .Q(_41195) );
  hi1s1 _42020_inst ( .DIN(_41597), .Q(_41619) );
  nnd2s1 _42021_inst ( .DIN1(_41788), .DIN2(_41789), .Q(_41597) );
  nor2s1 _42022_inst ( .DIN1(_41396), .DIN2(_41630), .Q(_41380) );
  nnd2s1 _42023_inst ( .DIN1(_53414), .DIN2(_26443), .Q(_41630) );
  hi1s1 _42024_inst ( .DIN(_40783), .Q(_40573) );
  nnd2s1 _42025_inst ( .DIN1(_40529), .DIN2(_40498), .Q(_40783) );
  nnd2s1 _42026_inst ( .DIN1(_40754), .DIN2(_41790), .Q(_40498) );
  nnd2s1 _42027_inst ( .DIN1(_41760), .DIN2(_39248), .Q(_41790) );
  hi1s1 _42028_inst ( .DIN(______[15]), .Q(_39248) );
  nnd2s1 _42029_inst ( .DIN1(_41760), .DIN2(_41684), .Q(_40529) );
  nor2s1 _42030_inst ( .DIN1(______[15]), .DIN2(_26842), .Q(_41684) );
  nor2s1 _42031_inst ( .DIN1(______[8]), .DIN2(______[26]), .Q(_41760) );
  nor2s1 _42032_inst ( .DIN1(_26842), .DIN2(_41791), .Q(_41786) );
  nor2s1 _42033_inst ( .DIN1(_41081), .DIN2(_41792), .Q(_41791) );
  nnd2s1 _42034_inst ( .DIN1(_40533), .DIN2(_40643), .Q(_41792) );
  nnd2s1 _42035_inst ( .DIN1(_41793), .DIN2(_41395), .Q(_40643) );
  nor2s1 _42036_inst ( .DIN1(_26208), .DIN2(_41658), .Q(_41793) );
  nnd2s1 _42037_inst ( .DIN1(_41723), .DIN2(_26274), .Q(_41658) );
  nnd2s1 _42038_inst ( .DIN1(_41794), .DIN2(_41395), .Q(_40533) );
  hi1s1 _42039_inst ( .DIN(_41661), .Q(_41395) );
  nnd2s1 _42040_inst ( .DIN1(_41795), .DIN2(_41789), .Q(_41661) );
  hi1s1 _42041_inst ( .DIN(_41540), .Q(_41789) );
  nnd2s1 _42042_inst ( .DIN1(_41796), .DIN2(_41797), .Q(_41540) );
  nor2s1 _42043_inst ( .DIN1(_53405), .DIN2(_41798), .Q(_41797) );
  nnd2s1 _42044_inst ( .DIN1(_26696), .DIN2(_26283), .Q(_41798) );
  nor2s1 _42045_inst ( .DIN1(_26615), .DIN2(_26218), .Q(_41796) );
  nor2s1 _42046_inst ( .DIN1(_26443), .DIN2(_41341), .Q(_41795) );
  nnd2s1 _42047_inst ( .DIN1(_41749), .DIN2(_41714), .Q(_41341) );
  nor2s1 _42048_inst ( .DIN1(_53409), .DIN2(_53411), .Q(_41714) );
  nor2s1 _42049_inst ( .DIN1(_26707), .DIN2(_53412), .Q(_41749) );
  nor2s1 _42050_inst ( .DIN1(_26208), .DIN2(_41609), .Q(_41794) );
  nnd2s1 _42051_inst ( .DIN1(_53414), .DIN2(_41723), .Q(_41609) );
  nor2s1 _42052_inst ( .DIN1(_26515), .DIN2(_53408), .Q(_41723) );
  hi1s1 _42053_inst ( .DIN(_40848), .Q(_41081) );
  nnd2s1 _42054_inst ( .DIN1(_41382), .DIN2(_41307), .Q(_40848) );
  hi1s1 _42055_inst ( .DIN(_41538), .Q(_41307) );
  nnd2s1 _42056_inst ( .DIN1(_41788), .DIN2(_41608), .Q(_41538) );
  hi1s1 _42057_inst ( .DIN(_41338), .Q(_41608) );
  nnd2s1 _42058_inst ( .DIN1(_41799), .DIN2(_41800), .Q(_41338) );
  nor2s1 _42059_inst ( .DIN1(_26615), .DIN2(_41801), .Q(_41800) );
  nnd2s1 _42060_inst ( .DIN1(_26218), .DIN2(_26283), .Q(_41801) );
  nor2s1 _42061_inst ( .DIN1(_26240), .DIN2(_26696), .Q(_41799) );
  nor2s1 _42062_inst ( .DIN1(_41603), .DIN2(_41716), .Q(_41788) );
  nnd2s1 _42063_inst ( .DIN1(_53412), .DIN2(_26707), .Q(_41716) );
  nnd2s1 _42064_inst ( .DIN1(_53409), .DIN2(_53411), .Q(_41603) );
  nor2s1 _42065_inst ( .DIN1(_41547), .DIN2(_41396), .Q(_41382) );
  nnd2s1 _42066_inst ( .DIN1(_41733), .DIN2(_26208), .Q(_41396) );
  hi1s1 _42067_inst ( .DIN(_41596), .Q(_41733) );
  nnd2s1 _42068_inst ( .DIN1(_53408), .DIN2(_26515), .Q(_41596) );
  nnd2s1 _42069_inst ( .DIN1(_53401), .DIN2(_26274), .Q(_41547) );
  hi1s1 _42070_inst ( .DIN(_27749), .Q(_28010) );
  nnd2s1 _42071_inst ( .DIN1(_41802), .DIN2(_28253), .Q(_27749) );
  hi1s1 _42072_inst ( .DIN(_31037), .Q(_28253) );
  nnd2s1 _42073_inst ( .DIN1(_34214), .DIN2(_35994), .Q(_31037) );
  nor2s1 _42074_inst ( .DIN1(_35342), .DIN2(_35511), .Q(_41802) );
  nnd2s1 _42075_inst ( .DIN1(_28178), .DIN2(_26362), .Q(_41473) );
  nnd2s1 _42076_inst ( .DIN1(_41803), .DIN2(_41804), .Q(
        ____1____________9_____) );
  nnd2s1 _42077_inst ( .DIN1(_41805), .DIN2(_41806), .Q(_41804) );
  xor2s1 _42078_inst ( .DIN1(_53445), .DIN2(_53456), .Q(_41805) );
  nnd2s1 _42079_inst ( .DIN1(_41807), .DIN2(_41808), .Q(_41803) );
  nnd2s1 _42080_inst ( .DIN1(_41809), .DIN2(_41810), .Q(_41808) );
  nor2s1 _42081_inst ( .DIN1(_41811), .DIN2(_41812), .Q(_41810) );
  nnd2s1 _42082_inst ( .DIN1(_41813), .DIN2(_41814), .Q(_41812) );
  nor2s1 _42083_inst ( .DIN1(_41815), .DIN2(_41816), .Q(_41814) );
  xor2s1 _42084_inst ( .DIN1(_32330), .DIN2(_41817), .Q(_41816) );
  and2s1 _42085_inst ( .DIN1(_41818), .DIN2(_41819), .Q(_41817) );
  nor2s1 _42086_inst ( .DIN1(_41820), .DIN2(_41821), .Q(_41813) );
  nnd2s1 _42087_inst ( .DIN1(_41822), .DIN2(_41823), .Q(_41811) );
  nor2s1 _42088_inst ( .DIN1(_41824), .DIN2(_41825), .Q(_41823) );
  nnd2s1 _42089_inst ( .DIN1(_41826), .DIN2(_41827), .Q(_41825) );
  nor2s1 _42090_inst ( .DIN1(_41828), .DIN2(_41829), .Q(_41822) );
  and2s1 _42091_inst ( .DIN1(_41830), .DIN2(_41831), .Q(_41829) );
  hi1s1 _42092_inst ( .DIN(_41832), .Q(_41828) );
  nor2s1 _42093_inst ( .DIN1(_41833), .DIN2(_41834), .Q(_41809) );
  nnd2s1 _42094_inst ( .DIN1(_41835), .DIN2(_41836), .Q(_41834) );
  nor2s1 _42095_inst ( .DIN1(_41837), .DIN2(_41838), .Q(_41836) );
  nor2s1 _42096_inst ( .DIN1(_41839), .DIN2(_41840), .Q(_41835) );
  nnd2s1 _42097_inst ( .DIN1(_41841), .DIN2(_41842), .Q(_41833) );
  nor2s1 _42098_inst ( .DIN1(_41843), .DIN2(_41844), .Q(_41842) );
  or2s1 _42099_inst ( .DIN1(_41845), .DIN2(_41846), .Q(_41844) );
  nor2s1 _42100_inst ( .DIN1(_41847), .DIN2(_41848), .Q(_41841) );
  nnd2s1 _42101_inst ( .DIN1(_41849), .DIN2(_41850), .Q(
        ____1____________8_____) );
  nnd2s1 _42102_inst ( .DIN1(_41851), .DIN2(_41852), .Q(_41850) );
  nnd2s1 _42103_inst ( .DIN1(_41853), .DIN2(______[18]), .Q(_41851) );
  nor2s1 _42104_inst ( .DIN1(_41854), .DIN2(_41855), .Q(_41853) );
  nor2s1 _42105_inst ( .DIN1(_26212), .DIN2(_41856), .Q(_41855) );
  nor2s1 _42106_inst ( .DIN1(_53422), .DIN2(_41857), .Q(_41854) );
  nor2s1 _42107_inst ( .DIN1(_26285), .DIN2(_26212), .Q(_41857) );
  nor2s1 _42108_inst ( .DIN1(_41858), .DIN2(_41859), .Q(_41849) );
  nor2s1 _42109_inst ( .DIN1(_41860), .DIN2(_41861), .Q(_41859) );
  nnd2s1 _42110_inst ( .DIN1(_41862), .DIN2(_41863), .Q(_41861) );
  nor2s1 _42111_inst ( .DIN1(_41864), .DIN2(_41865), .Q(_41863) );
  nnd2s1 _42112_inst ( .DIN1(_41866), .DIN2(_41867), .Q(_41865) );
  or2s1 _42113_inst ( .DIN1(_41868), .DIN2(_41869), .Q(_41864) );
  nor2s1 _42114_inst ( .DIN1(_41870), .DIN2(_41871), .Q(_41862) );
  nnd2s1 _42115_inst ( .DIN1(_41872), .DIN2(_41873), .Q(_41871) );
  xor2s1 _42116_inst ( .DIN1(_34151), .DIN2(_41874), .Q(_41872) );
  nor2s1 _42117_inst ( .DIN1(_41875), .DIN2(_41876), .Q(_41874) );
  nnd2s1 _42118_inst ( .DIN1(_41877), .DIN2(_41878), .Q(_41876) );
  nor2s1 _42119_inst ( .DIN1(_41879), .DIN2(_41880), .Q(_41877) );
  nnd2s1 _42120_inst ( .DIN1(_41881), .DIN2(_41882), .Q(_41875) );
  nor2s1 _42121_inst ( .DIN1(_41883), .DIN2(_41884), .Q(_41881) );
  hi1s1 _42122_inst ( .DIN(_41885), .Q(_41883) );
  nnd2s1 _42123_inst ( .DIN1(_41886), .DIN2(_41887), .Q(_41870) );
  hi1s1 _42124_inst ( .DIN(_41888), .Q(_41886) );
  nnd2s1 _42125_inst ( .DIN1(_41889), .DIN2(_41890), .Q(_41860) );
  nor2s1 _42126_inst ( .DIN1(_41891), .DIN2(_41892), .Q(_41890) );
  nnd2s1 _42127_inst ( .DIN1(_41893), .DIN2(_41894), .Q(_41892) );
  nnd2s1 _42128_inst ( .DIN1(_41895), .DIN2(_41896), .Q(_41894) );
  nnd2s1 _42129_inst ( .DIN1(_41897), .DIN2(_41898), .Q(_41891) );
  nnd2s1 _42130_inst ( .DIN1(_41899), .DIN2(_41900), .Q(_41898) );
  nor2s1 _42131_inst ( .DIN1(_41901), .DIN2(_41902), .Q(_41897) );
  nor2s1 _42132_inst ( .DIN1(_41903), .DIN2(_41904), .Q(_41902) );
  xor2s1 _42133_inst ( .DIN1(_32657), .DIN2(_41905), .Q(_41904) );
  nor2s1 _42134_inst ( .DIN1(_41906), .DIN2(_41907), .Q(_41905) );
  nnd2s1 _42135_inst ( .DIN1(_41908), .DIN2(_41909), .Q(_41907) );
  nnd2s1 _42136_inst ( .DIN1(_41910), .DIN2(_41911), .Q(_32657) );
  nor2s1 _42137_inst ( .DIN1(_41912), .DIN2(_41913), .Q(_41911) );
  nor2s1 _42138_inst ( .DIN1(_41914), .DIN2(_41915), .Q(_41910) );
  nor2s1 _42139_inst ( .DIN1(_41916), .DIN2(_41917), .Q(_41889) );
  or2s1 _42140_inst ( .DIN1(_41918), .DIN2(_41919), .Q(_41917) );
  nnd2s1 _42141_inst ( .DIN1(_41920), .DIN2(_41921), .Q(_41916) );
  nnd2s1 _42142_inst ( .DIN1(_41922), .DIN2(_41923), .Q(
        ____1____________7_____) );
  nor2s1 _42143_inst ( .DIN1(_41924), .DIN2(_41925), .Q(_41922) );
  nor2s1 _42144_inst ( .DIN1(_41852), .DIN2(_41926), .Q(_41925) );
  nnd2s1 _42145_inst ( .DIN1(_41927), .DIN2(_41928), .Q(_41926) );
  nor2s1 _42146_inst ( .DIN1(_41929), .DIN2(_41930), .Q(_41928) );
  nnd2s1 _42147_inst ( .DIN1(_41931), .DIN2(_41932), .Q(_41930) );
  nor2s1 _42148_inst ( .DIN1(_41933), .DIN2(_41934), .Q(_41931) );
  nor2s1 _42149_inst ( .DIN1(_41935), .DIN2(_41936), .Q(_41933) );
  nnd2s1 _42150_inst ( .DIN1(_41937), .DIN2(_41938), .Q(_41929) );
  nor2s1 _42151_inst ( .DIN1(_41939), .DIN2(_41940), .Q(_41938) );
  nor2s1 _42152_inst ( .DIN1(_41941), .DIN2(_41942), .Q(_41937) );
  nor2s1 _42153_inst ( .DIN1(_41943), .DIN2(_41944), .Q(_41942) );
  nor2s1 _42154_inst ( .DIN1(_41945), .DIN2(_41946), .Q(_41943) );
  hi1s1 _42155_inst ( .DIN(_41878), .Q(_41941) );
  nor2s1 _42156_inst ( .DIN1(_41947), .DIN2(_41948), .Q(_41927) );
  nnd2s1 _42157_inst ( .DIN1(_41949), .DIN2(_41950), .Q(_41948) );
  nor2s1 _42158_inst ( .DIN1(_41951), .DIN2(_41952), .Q(_41949) );
  nnd2s1 _42159_inst ( .DIN1(_41953), .DIN2(_41954), .Q(_41947) );
  hi1s1 _42160_inst ( .DIN(_41955), .Q(_41954) );
  nor2s1 _42161_inst ( .DIN1(_41956), .DIN2(_41957), .Q(_41953) );
  xor2s1 _42162_inst ( .DIN1(_36757), .DIN2(_41958), .Q(_41957) );
  nor2s1 _42163_inst ( .DIN1(_41959), .DIN2(_41960), .Q(_41958) );
  or2s1 _42164_inst ( .DIN1(_41961), .DIN2(_41962), .Q(_41960) );
  or2s1 _42165_inst ( .DIN1(_41963), .DIN2(_41821), .Q(_41959) );
  nnd2s1 _42166_inst ( .DIN1(_41964), .DIN2(_41965), .Q(_41821) );
  nor2s1 _42167_inst ( .DIN1(_41966), .DIN2(_41967), .Q(_41965) );
  nnd2s1 _42168_inst ( .DIN1(_41968), .DIN2(_41969), .Q(_41967) );
  nnd2s1 _42169_inst ( .DIN1(_41970), .DIN2(_39969), .Q(_41968) );
  or2s1 _42170_inst ( .DIN1(_41879), .DIN2(_41971), .Q(_41966) );
  nor2s1 _42171_inst ( .DIN1(_41972), .DIN2(_41973), .Q(_41964) );
  nnd2s1 _42172_inst ( .DIN1(_41974), .DIN2(_41975), .Q(_41973) );
  hi1s1 _42173_inst ( .DIN(_41976), .Q(_41974) );
  nor2s1 _42174_inst ( .DIN1(_41977), .DIN2(_41978), .Q(_41924) );
  nor2s1 _42175_inst ( .DIN1(_41979), .DIN2(_28684), .Q(_41978) );
  xor2s1 _42176_inst ( .DIN1(_41856), .DIN2(_41980), .Q(_41979) );
  xor2s1 _42177_inst ( .DIN1(_53424), .DIN2(_53425), .Q(_41980) );
  nnd2s1 _42178_inst ( .DIN1(_53424), .DIN2(_53422), .Q(_41856) );
  nnd2s1 _42179_inst ( .DIN1(_41981), .DIN2(_41982), .Q(
        ____1____________6_____) );
  nnd2s1 _42180_inst ( .DIN1(_41983), .DIN2(_41984), .Q(_41982) );
  xor2s1 _42181_inst ( .DIN1(_53413), .DIN2(_26345), .Q(_41983) );
  nnd2s1 _42182_inst ( .DIN1(_28056), .DIN2(_41985), .Q(_41981) );
  nnd2s1 _42183_inst ( .DIN1(_41986), .DIN2(_41987), .Q(_41985) );
  nor2s1 _42184_inst ( .DIN1(_41988), .DIN2(_41989), .Q(_41987) );
  nnd2s1 _42185_inst ( .DIN1(_41990), .DIN2(_41991), .Q(_41989) );
  and2s1 _42186_inst ( .DIN1(_41992), .DIN2(_41993), .Q(_41991) );
  nor2s1 _42187_inst ( .DIN1(_41994), .DIN2(_41995), .Q(_41990) );
  nor2s1 _42188_inst ( .DIN1(_41996), .DIN2(_41997), .Q(_41995) );
  nnd2s1 _42189_inst ( .DIN1(_37193), .DIN2(_28597), .Q(_41997) );
  nnd2s1 _42190_inst ( .DIN1(_41998), .DIN2(_41999), .Q(_41988) );
  nor2s1 _42191_inst ( .DIN1(_42000), .DIN2(_42001), .Q(_41999) );
  or2s1 _42192_inst ( .DIN1(_41971), .DIN2(_42002), .Q(_42001) );
  and2s1 _42193_inst ( .DIN1(_42003), .DIN2(_42004), .Q(_41998) );
  nor2s1 _42194_inst ( .DIN1(_42005), .DIN2(_42006), .Q(_41986) );
  nnd2s1 _42195_inst ( .DIN1(_42007), .DIN2(_42008), .Q(_42006) );
  nor2s1 _42196_inst ( .DIN1(_41955), .DIN2(_42009), .Q(_42008) );
  nnd2s1 _42197_inst ( .DIN1(_42010), .DIN2(_42011), .Q(_41955) );
  nnd2s1 _42198_inst ( .DIN1(_41819), .DIN2(_42012), .Q(_42010) );
  nor2s1 _42199_inst ( .DIN1(_42013), .DIN2(_42014), .Q(_42007) );
  nnd2s1 _42200_inst ( .DIN1(_42015), .DIN2(_42016), .Q(_42005) );
  nor2s1 _42201_inst ( .DIN1(_42017), .DIN2(_42018), .Q(_42016) );
  nnd2s1 _42202_inst ( .DIN1(_42019), .DIN2(_42020), .Q(_42018) );
  nnd2s1 _42203_inst ( .DIN1(_42021), .DIN2(_42022), .Q(_42020) );
  nnd2s1 _42204_inst ( .DIN1(_42023), .DIN2(_42024), .Q(_42022) );
  nnd2s1 _42205_inst ( .DIN1(_42025), .DIN2(_42026), .Q(_42019) );
  nor2s1 _42206_inst ( .DIN1(_41846), .DIN2(_41888), .Q(_42015) );
  nnd2s1 _42207_inst ( .DIN1(_42027), .DIN2(_42028), .Q(_41846) );
  nor2s1 _42208_inst ( .DIN1(_42029), .DIN2(_42030), .Q(_42027) );
  nor2s1 _42209_inst ( .DIN1(_35930), .DIN2(_42031), .Q(_42029) );
  nnd2s1 _42210_inst ( .DIN1(_42032), .DIN2(_42021), .Q(_42031) );
  nnd2s1 _42211_inst ( .DIN1(_42033), .DIN2(_41923), .Q(
        ____1____________5_____) );
  nor2s1 _42212_inst ( .DIN1(_42034), .DIN2(_42035), .Q(_42033) );
  nor2s1 _42213_inst ( .DIN1(_41852), .DIN2(_42036), .Q(_42035) );
  nnd2s1 _42214_inst ( .DIN1(_42037), .DIN2(_42038), .Q(_42036) );
  nor2s1 _42215_inst ( .DIN1(_42039), .DIN2(_42040), .Q(_42038) );
  nnd2s1 _42216_inst ( .DIN1(_42041), .DIN2(_42042), .Q(_42040) );
  nor2s1 _42217_inst ( .DIN1(_42043), .DIN2(_42044), .Q(_42042) );
  nnd2s1 _42218_inst ( .DIN1(_42045), .DIN2(_42046), .Q(_42044) );
  nor2s1 _42219_inst ( .DIN1(_42047), .DIN2(_42048), .Q(_42041) );
  nor2s1 _42220_inst ( .DIN1(_42049), .DIN2(_42050), .Q(_42048) );
  nor2s1 _42221_inst ( .DIN1(_42051), .DIN2(_42052), .Q(_42047) );
  nor2s1 _42222_inst ( .DIN1(_42053), .DIN2(_42054), .Q(_42051) );
  nnd2s1 _42223_inst ( .DIN1(_42055), .DIN2(_42056), .Q(_42039) );
  nor2s1 _42224_inst ( .DIN1(_42057), .DIN2(_42058), .Q(_42056) );
  nnd2s1 _42225_inst ( .DIN1(_42059), .DIN2(_42060), .Q(_42058) );
  hi1s1 _42226_inst ( .DIN(_42061), .Q(_42059) );
  hi1s1 _42227_inst ( .DIN(_42062), .Q(_42057) );
  nor2s1 _42228_inst ( .DIN1(_42063), .DIN2(_42064), .Q(_42055) );
  nor2s1 _42229_inst ( .DIN1(_42065), .DIN2(_42066), .Q(_42037) );
  nnd2s1 _42230_inst ( .DIN1(_42067), .DIN2(_42068), .Q(_42066) );
  nor2s1 _42231_inst ( .DIN1(_42069), .DIN2(_42070), .Q(_42068) );
  nnd2s1 _42232_inst ( .DIN1(_42071), .DIN2(_42072), .Q(_42070) );
  hi1s1 _42233_inst ( .DIN(_42073), .Q(_42071) );
  nor2s1 _42234_inst ( .DIN1(_42074), .DIN2(_42075), .Q(_42067) );
  hi1s1 _42235_inst ( .DIN(_42076), .Q(_42074) );
  nnd2s1 _42236_inst ( .DIN1(_42077), .DIN2(_42078), .Q(_42065) );
  nor2s1 _42237_inst ( .DIN1(_41845), .DIN2(_42079), .Q(_42078) );
  nnd2s1 _42238_inst ( .DIN1(_42080), .DIN2(_42081), .Q(_42079) );
  xor2s1 _42239_inst ( .DIN1(_30367), .DIN2(_42082), .Q(_42081) );
  nor2s1 _42240_inst ( .DIN1(_42083), .DIN2(_42084), .Q(_42082) );
  hi1s1 _42241_inst ( .DIN(_42085), .Q(_42080) );
  nnd2s1 _42242_inst ( .DIN1(_42086), .DIN2(_42087), .Q(_41845) );
  nor2s1 _42243_inst ( .DIN1(_41901), .DIN2(_42088), .Q(_42087) );
  nnd2s1 _42244_inst ( .DIN1(_42089), .DIN2(_42090), .Q(_42088) );
  nor2s1 _42245_inst ( .DIN1(_42091), .DIN2(_42092), .Q(_42086) );
  nor2s1 _42246_inst ( .DIN1(_41903), .DIN2(_42093), .Q(_42092) );
  nor2s1 _42247_inst ( .DIN1(_42094), .DIN2(_42095), .Q(_42091) );
  nor2s1 _42248_inst ( .DIN1(_41952), .DIN2(_42096), .Q(_42077) );
  nnd2s1 _42249_inst ( .DIN1(_42097), .DIN2(_42098), .Q(_41952) );
  nor2s1 _42250_inst ( .DIN1(_42099), .DIN2(_42100), .Q(_42098) );
  nnd2s1 _42251_inst ( .DIN1(_42101), .DIN2(_42102), .Q(_42100) );
  nor2s1 _42252_inst ( .DIN1(_42103), .DIN2(_42017), .Q(_42101) );
  nor2s1 _42253_inst ( .DIN1(_42104), .DIN2(_42105), .Q(_42017) );
  nor2s1 _42254_inst ( .DIN1(_41903), .DIN2(_42106), .Q(_42103) );
  nnd2s1 _42255_inst ( .DIN1(_42107), .DIN2(_42108), .Q(_42099) );
  and2s1 _42256_inst ( .DIN1(_42109), .DIN2(_42110), .Q(_42108) );
  nor2s1 _42257_inst ( .DIN1(_42111), .DIN2(_42112), .Q(_42107) );
  and2s1 _42258_inst ( .DIN1(_42113), .DIN2(_42114), .Q(_42112) );
  nor2s1 _42259_inst ( .DIN1(_41935), .DIN2(_42115), .Q(_42111) );
  nor2s1 _42260_inst ( .DIN1(_42116), .DIN2(_42117), .Q(_42097) );
  nnd2s1 _42261_inst ( .DIN1(_42118), .DIN2(_42119), .Q(_42117) );
  nor2s1 _42262_inst ( .DIN1(_42120), .DIN2(_42121), .Q(_42118) );
  nnd2s1 _42263_inst ( .DIN1(_42122), .DIN2(_42123), .Q(_42116) );
  nor2s1 _42264_inst ( .DIN1(_42124), .DIN2(_42125), .Q(_42123) );
  hi1s1 _42265_inst ( .DIN(_42126), .Q(_42124) );
  nor2s1 _42266_inst ( .DIN1(_41848), .DIN2(_41839), .Q(_42122) );
  nor2s1 _42267_inst ( .DIN1(_41977), .DIN2(_42127), .Q(_42034) );
  nor2s1 _42268_inst ( .DIN1(_27774), .DIN2(_26699), .Q(_42127) );
  nnd2s1 _42269_inst ( .DIN1(_42128), .DIN2(_39944), .Q(
        ____1____________4_____) );
  nnd2s1 _42270_inst ( .DIN1(_42129), .DIN2(_42130), .Q(_39944) );
  nor2s1 _42271_inst ( .DIN1(_39842), .DIN2(_42131), .Q(_42129) );
  nor2s1 _42272_inst ( .DIN1(_42132), .DIN2(_42133), .Q(_42128) );
  nor2s1 _42273_inst ( .DIN1(_39947), .DIN2(_42134), .Q(_42133) );
  nnd2s1 _42274_inst ( .DIN1(_42135), .DIN2(_42136), .Q(_42134) );
  nor2s1 _42275_inst ( .DIN1(_42137), .DIN2(_42138), .Q(_42136) );
  nnd2s1 _42276_inst ( .DIN1(_42139), .DIN2(_42140), .Q(_42138) );
  nor2s1 _42277_inst ( .DIN1(_42141), .DIN2(_42142), .Q(_42140) );
  nnd2s1 _42278_inst ( .DIN1(_42143), .DIN2(_42144), .Q(_42142) );
  or2s1 _42279_inst ( .DIN1(_42050), .DIN2(_41935), .Q(_42144) );
  nnd2s1 _42280_inst ( .DIN1(_42145), .DIN2(_41818), .Q(_42143) );
  and2s1 _42281_inst ( .DIN1(_42146), .DIN2(_41896), .Q(_42141) );
  nor2s1 _42282_inst ( .DIN1(_42147), .DIN2(_42148), .Q(_42139) );
  nnd2s1 _42283_inst ( .DIN1(_42149), .DIN2(_42150), .Q(_42148) );
  nnd2s1 _42284_inst ( .DIN1(_42151), .DIN2(_42152), .Q(_42150) );
  or2s1 _42285_inst ( .DIN1(_42024), .DIN2(_42153), .Q(_42149) );
  nor2s1 _42286_inst ( .DIN1(_41312), .DIN2(_42045), .Q(_42147) );
  nnd2s1 _42287_inst ( .DIN1(_42154), .DIN2(_42155), .Q(_42137) );
  nor2s1 _42288_inst ( .DIN1(_42156), .DIN2(_42157), .Q(_42155) );
  nnd2s1 _42289_inst ( .DIN1(_42158), .DIN2(_42109), .Q(_42157) );
  hi1s1 _42290_inst ( .DIN(_41882), .Q(_42156) );
  nnd2s1 _42291_inst ( .DIN1(_42159), .DIN2(_42160), .Q(_41882) );
  nor2s1 _42292_inst ( .DIN1(_37199), .DIN2(_42161), .Q(_42159) );
  nor2s1 _42293_inst ( .DIN1(_42162), .DIN2(_42163), .Q(_42154) );
  nnd2s1 _42294_inst ( .DIN1(_42164), .DIN2(_41832), .Q(_42163) );
  nor2s1 _42295_inst ( .DIN1(_42165), .DIN2(_42166), .Q(_42135) );
  nnd2s1 _42296_inst ( .DIN1(_42167), .DIN2(_42168), .Q(_42166) );
  nor2s1 _42297_inst ( .DIN1(_42169), .DIN2(_42170), .Q(_42168) );
  nnd2s1 _42298_inst ( .DIN1(_42171), .DIN2(_42076), .Q(_42170) );
  nor2s1 _42299_inst ( .DIN1(_42172), .DIN2(_42173), .Q(_42076) );
  nnd2s1 _42300_inst ( .DIN1(_42174), .DIN2(_42175), .Q(_42172) );
  hi1s1 _42301_inst ( .DIN(_42176), .Q(_42175) );
  nor2s1 _42302_inst ( .DIN1(_42177), .DIN2(_42178), .Q(_42167) );
  nnd2s1 _42303_inst ( .DIN1(_42179), .DIN2(_42180), .Q(_42178) );
  hi1s1 _42304_inst ( .DIN(_42181), .Q(_42180) );
  nnd2s1 _42305_inst ( .DIN1(_42182), .DIN2(_42183), .Q(_42165) );
  nor2s1 _42306_inst ( .DIN1(_41962), .DIN2(_42184), .Q(_42183) );
  nnd2s1 _42307_inst ( .DIN1(_42185), .DIN2(_42186), .Q(_42184) );
  nnd2s1 _42308_inst ( .DIN1(_42187), .DIN2(_42188), .Q(_41962) );
  or2s1 _42309_inst ( .DIN1(_42189), .DIN2(_42190), .Q(_42188) );
  xor2s1 _42310_inst ( .DIN1(_29599), .DIN2(_42191), .Q(_42187) );
  nnd2s1 _42311_inst ( .DIN1(_42192), .DIN2(_42160), .Q(_42191) );
  nor2s1 _42312_inst ( .DIN1(_42069), .DIN2(_42193), .Q(_42182) );
  or2s1 _42313_inst ( .DIN1(_42194), .DIN2(_42195), .Q(_42193) );
  nnd2s1 _42314_inst ( .DIN1(_42196), .DIN2(_42197), .Q(_42069) );
  nor2s1 _42315_inst ( .DIN1(_42198), .DIN2(_42199), .Q(_42196) );
  nor2s1 _42316_inst ( .DIN1(_42083), .DIN2(_42200), .Q(_42199) );
  hi1s1 _42317_inst ( .DIN(_42201), .Q(_42198) );
  nor2s1 _42318_inst ( .DIN1(_39842), .DIN2(_42202), .Q(_42132) );
  nor2s1 _42319_inst ( .DIN1(_42203), .DIN2(_27291), .Q(_42202) );
  xor2s1 _42320_inst ( .DIN1(_26369), .DIN2(_53478), .Q(_42203) );
  nnd2s1 _42321_inst ( .DIN1(_42204), .DIN2(_42205), .Q(
        ____1____________3_____) );
  nnd2s1 _42322_inst ( .DIN1(_40516), .DIN2(_42206), .Q(_42205) );
  xor2s1 _42323_inst ( .DIN1(_26274), .DIN2(_42207), .Q(_42206) );
  nor2s1 _42324_inst ( .DIN1(_40519), .DIN2(_41316), .Q(_40516) );
  and2s1 _42325_inst ( .DIN1(_42208), .DIN2(_34090), .Q(_41316) );
  hi1s1 _42326_inst ( .DIN(_36024), .Q(_34090) );
  nnd2s1 _42327_inst ( .DIN1(_42209), .DIN2(_38284), .Q(_36024) );
  nor2s1 _42328_inst ( .DIN1(_36977), .DIN2(_35997), .Q(_42208) );
  nnd2s1 _42329_inst ( .DIN1(_40519), .DIN2(_42210), .Q(_42204) );
  nnd2s1 _42330_inst ( .DIN1(_42211), .DIN2(_42212), .Q(_42210) );
  nor2s1 _42331_inst ( .DIN1(_42213), .DIN2(_42214), .Q(_42212) );
  nnd2s1 _42332_inst ( .DIN1(_42215), .DIN2(_42216), .Q(_42214) );
  nor2s1 _42333_inst ( .DIN1(_42217), .DIN2(_42218), .Q(_42216) );
  nor2s1 _42334_inst ( .DIN1(_42219), .DIN2(_41944), .Q(_42218) );
  nor2s1 _42335_inst ( .DIN1(_39969), .DIN2(_42045), .Q(_42217) );
  nor2s1 _42336_inst ( .DIN1(_41972), .DIN2(_42220), .Q(_42215) );
  nnd2s1 _42337_inst ( .DIN1(_42221), .DIN2(_42222), .Q(_41972) );
  and2s1 _42338_inst ( .DIN1(_42158), .DIN2(_42223), .Q(_42222) );
  or2s1 _42339_inst ( .DIN1(_42224), .DIN2(_42225), .Q(_42158) );
  nor2s1 _42340_inst ( .DIN1(_42226), .DIN2(_42227), .Q(_42221) );
  nor2s1 _42341_inst ( .DIN1(_42228), .DIN2(_42229), .Q(_42226) );
  nnd2s1 _42342_inst ( .DIN1(_42230), .DIN2(_42231), .Q(_42229) );
  nnd2s1 _42343_inst ( .DIN1(_42232), .DIN2(_42233), .Q(_42213) );
  nor2s1 _42344_inst ( .DIN1(_41940), .DIN2(_42234), .Q(_42233) );
  hi1s1 _42345_inst ( .DIN(_42235), .Q(_41940) );
  nor2s1 _42346_inst ( .DIN1(_41880), .DIN2(_42162), .Q(_42232) );
  hi1s1 _42347_inst ( .DIN(_42236), .Q(_41880) );
  nor2s1 _42348_inst ( .DIN1(_42237), .DIN2(_42238), .Q(_42211) );
  nnd2s1 _42349_inst ( .DIN1(_42239), .DIN2(_42240), .Q(_42238) );
  nor2s1 _42350_inst ( .DIN1(_42241), .DIN2(_42242), .Q(_42239) );
  nnd2s1 _42351_inst ( .DIN1(_42243), .DIN2(_42244), .Q(_42237) );
  nor2s1 _42352_inst ( .DIN1(_41843), .DIN2(_42120), .Q(_42244) );
  nnd2s1 _42353_inst ( .DIN1(_42245), .DIN2(_42246), .Q(_42120) );
  nor2s1 _42354_inst ( .DIN1(_42247), .DIN2(_42248), .Q(_42245) );
  nor2s1 _42355_inst ( .DIN1(_42249), .DIN2(_42250), .Q(_42248) );
  nor2s1 _42356_inst ( .DIN1(_42094), .DIN2(_42251), .Q(_42247) );
  hi1s1 _42357_inst ( .DIN(_41900), .Q(_42094) );
  nnd2s1 _42358_inst ( .DIN1(_42252), .DIN2(_42253), .Q(_41843) );
  nnd2s1 _42359_inst ( .DIN1(_42254), .DIN2(_42032), .Q(_42253) );
  nor2s1 _42360_inst ( .DIN1(_42255), .DIN2(_42083), .Q(_42254) );
  and2s1 _42361_inst ( .DIN1(_42256), .DIN2(_42164), .Q(_42252) );
  nnd2s1 _42362_inst ( .DIN1(_42257), .DIN2(_42258), .Q(_42164) );
  nor2s1 _42363_inst ( .DIN1(_42075), .DIN2(_42177), .Q(_42243) );
  nnd2s1 _42364_inst ( .DIN1(_42259), .DIN2(_42260), .Q(_42075) );
  nor2s1 _42365_inst ( .DIN1(_42261), .DIN2(_42262), .Q(_42260) );
  nnd2s1 _42366_inst ( .DIN1(_42263), .DIN2(_41826), .Q(_42262) );
  nnd2s1 _42367_inst ( .DIN1(_42026), .DIN2(_42264), .Q(_41826) );
  nnd2s1 _42368_inst ( .DIN1(_42265), .DIN2(_42021), .Q(_42263) );
  nor2s1 _42369_inst ( .DIN1(_42266), .DIN2(_42267), .Q(_42259) );
  nor2s1 _42370_inst ( .DIN1(_42225), .DIN2(_42268), .Q(_42266) );
  hi1s1 _42371_inst ( .DIN(_40563), .Q(_40519) );
  nnd2s1 _42372_inst ( .DIN1(_42269), .DIN2(_28182), .Q(_40563) );
  hi1s1 _42373_inst ( .DIN(_28146), .Q(_28182) );
  nnd2s1 _42374_inst ( .DIN1(_42209), .DIN2(_42270), .Q(_28146) );
  nor2s1 _42375_inst ( .DIN1(_36019), .DIN2(_38282), .Q(_42269) );
  nnd2s1 _42376_inst ( .DIN1(_42271), .DIN2(_38261), .Q(_38282) );
  nor2s1 _42377_inst ( .DIN1(_36492), .DIN2(_38031), .Q(_42271) );
  hi1s1 _42378_inst ( .DIN(_36022), .Q(_36492) );
  hi1s1 _42379_inst ( .DIN(_41221), .Q(_36019) );
  nnd2s1 _42380_inst ( .DIN1(_42272), .DIN2(_41923), .Q(
        ____1____________2_____) );
  nor2s1 _42381_inst ( .DIN1(_42273), .DIN2(_42274), .Q(_42272) );
  nor2s1 _42382_inst ( .DIN1(_41852), .DIN2(_42275), .Q(_42274) );
  nnd2s1 _42383_inst ( .DIN1(_42276), .DIN2(_42277), .Q(_42275) );
  nor2s1 _42384_inst ( .DIN1(_42278), .DIN2(_42279), .Q(_42277) );
  nnd2s1 _42385_inst ( .DIN1(_42280), .DIN2(_42281), .Q(_42279) );
  nor2s1 _42386_inst ( .DIN1(_41869), .DIN2(_42282), .Q(_42281) );
  nnd2s1 _42387_inst ( .DIN1(_42197), .DIN2(_42283), .Q(_42282) );
  nnd2s1 _42388_inst ( .DIN1(_42284), .DIN2(_41896), .Q(_42283) );
  nnd2s1 _42389_inst ( .DIN1(_42152), .DIN2(_42285), .Q(_42197) );
  nnd2s1 _42390_inst ( .DIN1(_42286), .DIN2(_42287), .Q(_41869) );
  nor2s1 _42391_inst ( .DIN1(_42288), .DIN2(_42289), .Q(_42287) );
  nnd2s1 _42392_inst ( .DIN1(_42046), .DIN2(_42235), .Q(_42289) );
  nnd2s1 _42393_inst ( .DIN1(_42290), .DIN2(_35101), .Q(_42235) );
  nnd2s1 _42394_inst ( .DIN1(_42291), .DIN2(_42292), .Q(_42046) );
  nor2s1 _42395_inst ( .DIN1(_37199), .DIN2(_42293), .Q(_42291) );
  hi1s1 _42396_inst ( .DIN(_42294), .Q(_42288) );
  nor2s1 _42397_inst ( .DIN1(_42295), .DIN2(_42296), .Q(_42286) );
  nor2s1 _42398_inst ( .DIN1(_41903), .DIN2(_42297), .Q(_42296) );
  nor2s1 _42399_inst ( .DIN1(_42298), .DIN2(_42225), .Q(_42295) );
  nor2s1 _42400_inst ( .DIN1(_41868), .DIN2(_42299), .Q(_42280) );
  nnd2s1 _42401_inst ( .DIN1(_42300), .DIN2(_42301), .Q(_41868) );
  nnd2s1 _42402_inst ( .DIN1(_42302), .DIN2(_42151), .Q(_42301) );
  nor2s1 _42403_inst ( .DIN1(_42303), .DIN2(_42304), .Q(_42300) );
  and2s1 _42404_inst ( .DIN1(_42305), .DIN2(_41896), .Q(_42304) );
  nnd2s1 _42405_inst ( .DIN1(_42306), .DIN2(_42307), .Q(_42278) );
  nor2s1 _42406_inst ( .DIN1(_42162), .DIN2(_42308), .Q(_42307) );
  nnd2s1 _42407_inst ( .DIN1(_42309), .DIN2(_42310), .Q(_42308) );
  and2s1 _42408_inst ( .DIN1(_42311), .DIN2(_26837), .Q(_42162) );
  nor2s1 _42409_inst ( .DIN1(_42313), .DIN2(_42314), .Q(_42306) );
  nor2s1 _42410_inst ( .DIN1(_42249), .DIN2(_42189), .Q(_42314) );
  and2s1 _42411_inst ( .DIN1(_42292), .DIN2(_42315), .Q(_42313) );
  nor2s1 _42412_inst ( .DIN1(_42316), .DIN2(_42317), .Q(_42276) );
  nnd2s1 _42413_inst ( .DIN1(_42318), .DIN2(_42319), .Q(_42317) );
  nor2s1 _42414_inst ( .DIN1(_42320), .DIN2(_42321), .Q(_42319) );
  nnd2s1 _42415_inst ( .DIN1(_42322), .DIN2(_42323), .Q(_42321) );
  hi1s1 _42416_inst ( .DIN(_42241), .Q(_42323) );
  nnd2s1 _42417_inst ( .DIN1(_42324), .DIN2(_42325), .Q(_42241) );
  nor2s1 _42418_inst ( .DIN1(_42326), .DIN2(_42327), .Q(_42325) );
  nnd2s1 _42419_inst ( .DIN1(_42328), .DIN2(_42062), .Q(_42327) );
  nnd2s1 _42420_inst ( .DIN1(_42329), .DIN2(_42231), .Q(_42328) );
  nor2s1 _42421_inst ( .DIN1(_37318), .DIN2(_42330), .Q(_42329) );
  nor2s1 _42422_inst ( .DIN1(_42052), .DIN2(_42331), .Q(_42326) );
  nor2s1 _42423_inst ( .DIN1(_41848), .DIN2(_41919), .Q(_42324) );
  nnd2s1 _42424_inst ( .DIN1(_42332), .DIN2(_42333), .Q(_41919) );
  nnd2s1 _42425_inst ( .DIN1(_41819), .DIN2(_41818), .Q(_42333) );
  or2s1 _42426_inst ( .DIN1(_42105), .DIN2(_41935), .Q(_42332) );
  nnd2s1 _42427_inst ( .DIN1(_42334), .DIN2(_42335), .Q(_41848) );
  nnd2s1 _42428_inst ( .DIN1(_42336), .DIN2(_42337), .Q(_42335) );
  nor2s1 _42429_inst ( .DIN1(_35533), .DIN2(_42104), .Q(_42337) );
  nor2s1 _42430_inst ( .DIN1(_36066), .DIN2(_42338), .Q(_42336) );
  xor2s1 _42431_inst ( .DIN1(_41367), .DIN2(_42339), .Q(_42334) );
  nnd2s1 _42432_inst ( .DIN1(_42340), .DIN2(_42341), .Q(_42339) );
  nor2s1 _42433_inst ( .DIN1(_42342), .DIN2(_36207), .Q(_42340) );
  hi1s1 _42434_inst ( .DIN(_42343), .Q(_42320) );
  nor2s1 _42435_inst ( .DIN1(_42344), .DIN2(_42345), .Q(_42318) );
  hi1s1 _42436_inst ( .DIN(_42346), .Q(_42345) );
  nnd2s1 _42437_inst ( .DIN1(_42347), .DIN2(_42348), .Q(_42316) );
  nor2s1 _42438_inst ( .DIN1(_42349), .DIN2(_42350), .Q(_42348) );
  or2s1 _42439_inst ( .DIN1(_42013), .DIN2(_41951), .Q(_42350) );
  nnd2s1 _42440_inst ( .DIN1(_42351), .DIN2(_42352), .Q(_41951) );
  nnd2s1 _42441_inst ( .DIN1(_42026), .DIN2(_26837), .Q(_42352) );
  nor2s1 _42442_inst ( .DIN1(_42353), .DIN2(_36455), .Q(_42026) );
  nnd2s1 _42443_inst ( .DIN1(_42053), .DIN2(_41896), .Q(_42351) );
  hi1s1 _42444_inst ( .DIN(_42354), .Q(_42053) );
  nnd2s1 _42445_inst ( .DIN1(_42355), .DIN2(_42356), .Q(_42013) );
  nor2s1 _42446_inst ( .DIN1(_42357), .DIN2(_42358), .Q(_42356) );
  nnd2s1 _42447_inst ( .DIN1(_42359), .DIN2(_26816), .Q(_42358) );
  nor2s1 _42448_inst ( .DIN1(_42361), .DIN2(_42362), .Q(_42359) );
  nor2s1 _42449_inst ( .DIN1(_42363), .DIN2(_41909), .Q(_42362) );
  nnd2s1 _42450_inst ( .DIN1(_42364), .DIN2(_42365), .Q(_42357) );
  nor2s1 _42451_inst ( .DIN1(_42366), .DIN2(_42367), .Q(_42365) );
  hi1s1 _42452_inst ( .DIN(_42368), .Q(_42366) );
  nor2s1 _42453_inst ( .DIN1(_42234), .DIN2(_41824), .Q(_42364) );
  hi1s1 _42454_inst ( .DIN(_42369), .Q(_41824) );
  and2s1 _42455_inst ( .DIN1(_42370), .DIN2(_42371), .Q(_42234) );
  nor2s1 _42456_inst ( .DIN1(_42372), .DIN2(_42373), .Q(_42355) );
  nnd2s1 _42457_inst ( .DIN1(_42374), .DIN2(_42375), .Q(_42373) );
  nor2s1 _42458_inst ( .DIN1(_42096), .DIN2(_42194), .Q(_42374) );
  nnd2s1 _42459_inst ( .DIN1(_42376), .DIN2(_42377), .Q(_42194) );
  nor2s1 _42460_inst ( .DIN1(_42378), .DIN2(_41879), .Q(_42377) );
  nor2s1 _42461_inst ( .DIN1(_42379), .DIN2(_41903), .Q(_41879) );
  and2s1 _42462_inst ( .DIN1(_42380), .DIN2(_42381), .Q(_42376) );
  nnd2s1 _42463_inst ( .DIN1(_42382), .DIN2(_42383), .Q(_42096) );
  nor2s1 _42464_inst ( .DIN1(_41884), .DIN2(_42384), .Q(_42383) );
  nor2s1 _42465_inst ( .DIN1(_41944), .DIN2(_42385), .Q(_42384) );
  and2s1 _42466_inst ( .DIN1(_42386), .DIN2(_35101), .Q(_41884) );
  nor2s1 _42467_inst ( .DIN1(_42387), .DIN2(_42388), .Q(_42386) );
  nor2s1 _42468_inst ( .DIN1(_41847), .DIN2(_42389), .Q(_42382) );
  nnd2s1 _42469_inst ( .DIN1(_42390), .DIN2(_42391), .Q(_41847) );
  hi1s1 _42470_inst ( .DIN(_42392), .Q(_42390) );
  nnd2s1 _42471_inst ( .DIN1(_42393), .DIN2(_42394), .Q(_42372) );
  nor2s1 _42472_inst ( .DIN1(_42395), .DIN2(_41918), .Q(_42394) );
  nnd2s1 _42473_inst ( .DIN1(_42396), .DIN2(_42223), .Q(_41918) );
  nnd2s1 _42474_inst ( .DIN1(_42397), .DIN2(_36063), .Q(_42223) );
  nor2s1 _42475_inst ( .DIN1(_42083), .DIN2(_42330), .Q(_42397) );
  nor2s1 _42476_inst ( .DIN1(_41961), .DIN2(_42398), .Q(_42393) );
  nnd2s1 _42477_inst ( .DIN1(_42399), .DIN2(_42400), .Q(_41961) );
  nnd2s1 _42478_inst ( .DIN1(_42401), .DIN2(_42402), .Q(_42400) );
  nor2s1 _42479_inst ( .DIN1(_42403), .DIN2(_42169), .Q(_42347) );
  nnd2s1 _42480_inst ( .DIN1(_42404), .DIN2(_42405), .Q(_42169) );
  or2s1 _42481_inst ( .DIN1(_42406), .DIN2(_42407), .Q(_42405) );
  nnd2s1 _42482_inst ( .DIN1(_42160), .DIN2(_42408), .Q(_42404) );
  nor2s1 _42483_inst ( .DIN1(_41977), .DIN2(_42409), .Q(_42273) );
  nor2s1 _42484_inst ( .DIN1(_27448), .DIN2(_26285), .Q(_42409) );
  nnd2s1 _42485_inst ( .DIN1(_42410), .DIN2(_41923), .Q(
        ____1____________1_____) );
  nor2s1 _42486_inst ( .DIN1(_42411), .DIN2(_42412), .Q(_42410) );
  nor2s1 _42487_inst ( .DIN1(_41852), .DIN2(_42413), .Q(_42412) );
  nnd2s1 _42488_inst ( .DIN1(_42414), .DIN2(_42415), .Q(_42413) );
  nor2s1 _42489_inst ( .DIN1(_42416), .DIN2(_42417), .Q(_42415) );
  nnd2s1 _42490_inst ( .DIN1(_42418), .DIN2(_42419), .Q(_42417) );
  nor2s1 _42491_inst ( .DIN1(_42420), .DIN2(_42421), .Q(_42419) );
  nnd2s1 _42492_inst ( .DIN1(_42391), .DIN2(_41878), .Q(_42421) );
  nnd2s1 _42493_inst ( .DIN1(_42025), .DIN2(_42311), .Q(_41878) );
  nnd2s1 _42494_inst ( .DIN1(_42422), .DIN2(_42264), .Q(_42391) );
  hi1s1 _42495_inst ( .DIN(_42423), .Q(_42422) );
  nor2s1 _42496_inst ( .DIN1(_42379), .DIN2(_42225), .Q(_42420) );
  nor2s1 _42497_inst ( .DIN1(_42424), .DIN2(_42425), .Q(_42418) );
  nor2s1 _42498_inst ( .DIN1(_42426), .DIN2(_42052), .Q(_42425) );
  nor2s1 _42499_inst ( .DIN1(_42427), .DIN2(_42284), .Q(_42426) );
  nor2s1 _42500_inst ( .DIN1(_41935), .DIN2(_42105), .Q(_42424) );
  nnd2s1 _42501_inst ( .DIN1(_42428), .DIN2(_42429), .Q(_42416) );
  nor2s1 _42502_inst ( .DIN1(_42430), .DIN2(_42431), .Q(_42429) );
  nnd2s1 _42503_inst ( .DIN1(_41993), .DIN2(_42368), .Q(_42431) );
  nnd2s1 _42504_inst ( .DIN1(_42432), .DIN2(_42230), .Q(_41993) );
  nor2s1 _42505_inst ( .DIN1(_42104), .DIN2(_42330), .Q(_42432) );
  hi1s1 _42506_inst ( .DIN(_42433), .Q(_42430) );
  and2s1 _42507_inst ( .DIN1(_42434), .DIN2(_42045), .Q(_42428) );
  nor2s1 _42508_inst ( .DIN1(_42435), .DIN2(_42436), .Q(_42414) );
  nnd2s1 _42509_inst ( .DIN1(_42437), .DIN2(_42438), .Q(_42436) );
  nor2s1 _42510_inst ( .DIN1(_42181), .DIN2(_42439), .Q(_42438) );
  nnd2s1 _42511_inst ( .DIN1(_42440), .DIN2(_42119), .Q(_42439) );
  and2s1 _42512_inst ( .DIN1(_42441), .DIN2(_42442), .Q(_42119) );
  nnd2s1 _42513_inst ( .DIN1(_42443), .DIN2(_42032), .Q(_42442) );
  nor2s1 _42514_inst ( .DIN1(_42255), .DIN2(_42052), .Q(_42443) );
  nnd2s1 _42515_inst ( .DIN1(_42371), .DIN2(_42444), .Q(_42441) );
  hi1s1 _42516_inst ( .DIN(_42267), .Q(_42440) );
  nnd2s1 _42517_inst ( .DIN1(_42445), .DIN2(_42446), .Q(_42267) );
  nor2s1 _42518_inst ( .DIN1(_42447), .DIN2(_42448), .Q(_42446) );
  nnd2s1 _42519_inst ( .DIN1(_41885), .DIN2(_41992), .Q(_42448) );
  nnd2s1 _42520_inst ( .DIN1(_42449), .DIN2(_42450), .Q(_41885) );
  nor2s1 _42521_inst ( .DIN1(_42407), .DIN2(_35930), .Q(_42449) );
  hi1s1 _42522_inst ( .DIN(_42451), .Q(_42447) );
  nor2s1 _42523_inst ( .DIN1(_42452), .DIN2(_42453), .Q(_42445) );
  nnd2s1 _42524_inst ( .DIN1(_42454), .DIN2(_42310), .Q(_42453) );
  nor2s1 _42525_inst ( .DIN1(_42049), .DIN2(_41936), .Q(_42452) );
  nnd2s1 _42526_inst ( .DIN1(_42455), .DIN2(_42456), .Q(_42181) );
  nor2s1 _42527_inst ( .DIN1(_41901), .DIN2(_42457), .Q(_42456) );
  nor2s1 _42528_inst ( .DIN1(_42052), .DIN2(_42084), .Q(_42457) );
  hi1s1 _42529_inst ( .DIN(_42309), .Q(_41901) );
  nor2s1 _42530_inst ( .DIN1(_42458), .DIN2(_42403), .Q(_42455) );
  nnd2s1 _42531_inst ( .DIN1(_42459), .DIN2(_42460), .Q(_42403) );
  nnd2s1 _42532_inst ( .DIN1(_42461), .DIN2(_42401), .Q(_42460) );
  or2s1 _42533_inst ( .DIN1(_42462), .DIN2(_42093), .Q(_42459) );
  and2s1 _42534_inst ( .DIN1(_42463), .DIN2(_42302), .Q(_42458) );
  nor2s1 _42535_inst ( .DIN1(_42242), .DIN2(_42464), .Q(_42437) );
  nnd2s1 _42536_inst ( .DIN1(_42465), .DIN2(_42466), .Q(_42242) );
  nor2s1 _42537_inst ( .DIN1(_42467), .DIN2(_42468), .Q(_42466) );
  nnd2s1 _42538_inst ( .DIN1(_42469), .DIN2(_42470), .Q(_42468) );
  nnd2s1 _42539_inst ( .DIN1(_42231), .DIN2(_42471), .Q(_42469) );
  nnd2s1 _42540_inst ( .DIN1(_42472), .DIN2(_42380), .Q(_42467) );
  nor2s1 _42541_inst ( .DIN1(_42473), .DIN2(_42474), .Q(_42465) );
  nnd2s1 _42542_inst ( .DIN1(_42475), .DIN2(_42375), .Q(_42474) );
  and2s1 _42543_inst ( .DIN1(_42201), .DIN2(_42476), .Q(_42375) );
  nnd2s1 _42544_inst ( .DIN1(_42477), .DIN2(_42292), .Q(_42476) );
  nor2s1 _42545_inst ( .DIN1(_42353), .DIN2(_36202), .Q(_42477) );
  nnd2s1 _42546_inst ( .DIN1(_42478), .DIN2(_42479), .Q(_42201) );
  nor2s1 _42547_inst ( .DIN1(_42083), .DIN2(_37318), .Q(_42478) );
  nnd2s1 _42548_inst ( .DIN1(_41921), .DIN2(_42480), .Q(_42473) );
  nor2s1 _42549_inst ( .DIN1(_42481), .DIN2(_42482), .Q(_41921) );
  and2s1 _42550_inst ( .DIN1(_42054), .DIN2(_41896), .Q(_42482) );
  nnd2s1 _42551_inst ( .DIN1(_42483), .DIN2(_42484), .Q(_42435) );
  nor2s1 _42552_inst ( .DIN1(_41976), .DIN2(_42485), .Q(_42484) );
  nnd2s1 _42553_inst ( .DIN1(_42486), .DIN2(_42487), .Q(_42485) );
  nnd2s1 _42554_inst ( .DIN1(_42401), .DIN2(_42488), .Q(_42487) );
  nnd2s1 _42555_inst ( .DIN1(_42489), .DIN2(_42251), .Q(_42488) );
  nnd2s1 _42556_inst ( .DIN1(_42490), .DIN2(_41818), .Q(_42486) );
  nnd2s1 _42557_inst ( .DIN1(_42491), .DIN2(_42492), .Q(_41976) );
  nnd2s1 _42558_inst ( .DIN1(_41906), .DIN2(_26837), .Q(_42492) );
  nor2s1 _42559_inst ( .DIN1(_41994), .DIN2(_42493), .Q(_42491) );
  hi1s1 _42560_inst ( .DIN(_42494), .Q(_42493) );
  and2s1 _42561_inst ( .DIN1(_42495), .DIN2(_42401), .Q(_41994) );
  nor2s1 _42562_inst ( .DIN1(_42496), .DIN2(_41837), .Q(_42483) );
  nnd2s1 _42563_inst ( .DIN1(_42497), .DIN2(_42498), .Q(_41837) );
  nor2s1 _42564_inst ( .DIN1(_42499), .DIN2(_42500), .Q(_42498) );
  nnd2s1 _42565_inst ( .DIN1(_42501), .DIN2(_42109), .Q(_42500) );
  or2s1 _42566_inst ( .DIN1(_42502), .DIN2(_41903), .Q(_42109) );
  nnd2s1 _42567_inst ( .DIN1(_42503), .DIN2(_26837), .Q(_42501) );
  nnd2s1 _42568_inst ( .DIN1(_41909), .DIN2(_42189), .Q(_42503) );
  and2s1 _42569_inst ( .DIN1(_41896), .DIN2(_42504), .Q(_42499) );
  nor2s1 _42570_inst ( .DIN1(_42505), .DIN2(_42176), .Q(_42497) );
  nnd2s1 _42571_inst ( .DIN1(_42506), .DIN2(_42507), .Q(_42176) );
  nnd2s1 _42572_inst ( .DIN1(_42508), .DIN2(_26837), .Q(_42507) );
  nor2s1 _42573_inst ( .DIN1(_42509), .DIN2(_42052), .Q(_42505) );
  nor2s1 _42574_inst ( .DIN1(_53421), .DIN2(_41977), .Q(_42411) );
  nor2s1 _42575_inst ( .DIN1(_42510), .DIN2(_27593), .Q(
        ____1____________11_____) );
  nnd2s1 _42576_inst ( .DIN1(_42511), .DIN2(_35721), .Q(_27593) );
  nor2s1 _42577_inst ( .DIN1(_35301), .DIN2(_39319), .Q(_42511) );
  nor2s1 _42578_inst ( .DIN1(_42512), .DIN2(_42513), .Q(_42510) );
  nnd2s1 _42579_inst ( .DIN1(_42514), .DIN2(_42515), .Q(_42513) );
  nor2s1 _42580_inst ( .DIN1(_42516), .DIN2(_42517), .Q(_42515) );
  nnd2s1 _42581_inst ( .DIN1(_41950), .DIN2(_41867), .Q(_42517) );
  and2s1 _42582_inst ( .DIN1(_42518), .DIN2(_42519), .Q(_41867) );
  nor2s1 _42583_inst ( .DIN1(_42520), .DIN2(_42521), .Q(_42519) );
  nnd2s1 _42584_inst ( .DIN1(_42522), .DIN2(_42523), .Q(_42521) );
  nnd2s1 _42585_inst ( .DIN1(_41970), .DIN2(_41312), .Q(_42523) );
  nnd2s1 _42586_inst ( .DIN1(_42461), .DIN2(_41900), .Q(_42522) );
  nnd2s1 _42587_inst ( .DIN1(_41832), .DIN2(_41992), .Q(_42520) );
  nnd2s1 _42588_inst ( .DIN1(_42524), .DIN2(_42160), .Q(_41992) );
  nor2s1 _42589_inst ( .DIN1(_36201), .DIN2(_42161), .Q(_42524) );
  nnd2s1 _42590_inst ( .DIN1(_42402), .DIN2(_41900), .Q(_41832) );
  nor2s1 _42591_inst ( .DIN1(_42395), .DIN2(_42525), .Q(_42518) );
  nnd2s1 _42592_inst ( .DIN1(_42480), .DIN2(_41932), .Q(_42525) );
  nnd2s1 _42593_inst ( .DIN1(_42265), .DIN2(_42231), .Q(_41932) );
  nnd2s1 _42594_inst ( .DIN1(_42192), .DIN2(_26837), .Q(_42480) );
  nnd2s1 _42595_inst ( .DIN1(_42526), .DIN2(_41975), .Q(_42395) );
  nnd2s1 _42596_inst ( .DIN1(_42527), .DIN2(_26837), .Q(_41975) );
  hi1s1 _42597_inst ( .DIN(_42084), .Q(_42527) );
  nnd2s1 _42598_inst ( .DIN1(_42528), .DIN2(_42264), .Q(_42526) );
  nor2s1 _42599_inst ( .DIN1(_42529), .DIN2(_42299), .Q(_41950) );
  nnd2s1 _42600_inst ( .DIN1(_42090), .DIN2(_42530), .Q(_42299) );
  nnd2s1 _42601_inst ( .DIN1(_42290), .DIN2(_42531), .Q(_42530) );
  hi1s1 _42602_inst ( .DIN(_37199), .Q(_42531) );
  or2s1 _42603_inst ( .DIN1(_42367), .DIN2(_42532), .Q(_42529) );
  nor2s1 _42604_inst ( .DIN1(_42533), .DIN2(_41909), .Q(_42532) );
  hi1s1 _42605_inst ( .DIN(_42534), .Q(_41909) );
  and2s1 _42606_inst ( .DIN1(_42292), .DIN2(_42535), .Q(_42367) );
  nnd2s1 _42607_inst ( .DIN1(_42536), .DIN2(_42537), .Q(_42535) );
  nnd2s1 _42608_inst ( .DIN1(_42538), .DIN2(_42539), .Q(_42516) );
  hi1s1 _42609_inst ( .DIN(_41838), .Q(_42539) );
  nnd2s1 _42610_inst ( .DIN1(_42540), .DIN2(_42102), .Q(_41838) );
  nnd2s1 _42611_inst ( .DIN1(_42463), .DIN2(_42541), .Q(_42102) );
  nor2s1 _42612_inst ( .DIN1(_42542), .DIN2(_42543), .Q(_42540) );
  nor2s1 _42613_inst ( .DIN1(_42330), .DIN2(_42544), .Q(_42543) );
  nnd2s1 _42614_inst ( .DIN1(_37334), .DIN2(_42021), .Q(_42544) );
  nor2s1 _42615_inst ( .DIN1(_42545), .DIN2(_42546), .Q(_42542) );
  nnd2s1 _42616_inst ( .DIN1(_37193), .DIN2(_42547), .Q(_42546) );
  nor2s1 _42617_inst ( .DIN1(_42303), .DIN2(_42548), .Q(_42538) );
  xor2s1 _42618_inst ( .DIN1(_42549), .DIN2(_27418), .Q(_42548) );
  hi1s1 _42619_inst ( .DIN(_32753), .Q(_27418) );
  nnd2s1 _42620_inst ( .DIN1(_42302), .DIN2(_42550), .Q(_42549) );
  nor2s1 _42621_inst ( .DIN1(_42551), .DIN2(_42104), .Q(_42303) );
  hi1s1 _42622_inst ( .DIN(_42552), .Q(_42551) );
  nor2s1 _42623_inst ( .DIN1(_42553), .DIN2(_42554), .Q(_42514) );
  nnd2s1 _42624_inst ( .DIN1(_42555), .DIN2(_42171), .Q(_42554) );
  and2s1 _42625_inst ( .DIN1(_42294), .DIN2(_42556), .Q(_42171) );
  nnd2s1 _42626_inst ( .DIN1(_42152), .DIN2(_41946), .Q(_42556) );
  nnd2s1 _42627_inst ( .DIN1(_41831), .DIN2(_42114), .Q(_42294) );
  nnd2s1 _42628_inst ( .DIN1(_42557), .DIN2(_42072), .Q(_42553) );
  and2s1 _42629_inst ( .DIN1(_42434), .DIN2(_42558), .Q(_42072) );
  nnd2s1 _42630_inst ( .DIN1(_42292), .DIN2(_41895), .Q(_42558) );
  nnd2s1 _42631_inst ( .DIN1(_42559), .DIN2(_35101), .Q(_42434) );
  hi1s1 _42632_inst ( .DIN(_35930), .Q(_35101) );
  nor2s1 _42633_inst ( .DIN1(_42161), .DIN2(_42407), .Q(_42559) );
  nnd2s1 _42634_inst ( .DIN1(_42560), .DIN2(_42561), .Q(_42512) );
  nor2s1 _42635_inst ( .DIN1(_42562), .DIN2(_42563), .Q(_42561) );
  nnd2s1 _42636_inst ( .DIN1(_42564), .DIN2(_42565), .Q(_42563) );
  nnd2s1 _42637_inst ( .DIN1(_42315), .DIN2(_42258), .Q(_42565) );
  or2s1 _42638_inst ( .DIN1(_42502), .DIN2(_42363), .Q(_42564) );
  nnd2s1 _42639_inst ( .DIN1(_42566), .DIN2(_42506), .Q(_42562) );
  nnd2s1 _42640_inst ( .DIN1(_41945), .DIN2(_26837), .Q(_42506) );
  hi1s1 _42641_inst ( .DIN(_42298), .Q(_41945) );
  nnd2s1 _42642_inst ( .DIN1(_42567), .DIN2(_42568), .Q(_42298) );
  nor2s1 _42643_inst ( .DIN1(_41971), .DIN2(_42378), .Q(_42566) );
  and2s1 _42644_inst ( .DIN1(_42569), .DIN2(_42570), .Q(_42378) );
  nor2s1 _42645_inst ( .DIN1(_39040), .DIN2(_42407), .Q(_42569) );
  nor2s1 _42646_inst ( .DIN1(_42571), .DIN2(_42104), .Q(_41971) );
  nor2s1 _42647_inst ( .DIN1(_42572), .DIN2(_42573), .Q(_42560) );
  nnd2s1 _42648_inst ( .DIN1(_42574), .DIN2(_42575), .Q(_42573) );
  nnd2s1 _42649_inst ( .DIN1(_42114), .DIN2(_42113), .Q(_42575) );
  nnd2s1 _42650_inst ( .DIN1(_41906), .DIN2(_41896), .Q(_42574) );
  nnd2s1 _42651_inst ( .DIN1(_42576), .DIN2(_42577), .Q(_42572) );
  nnd2s1 _42652_inst ( .DIN1(_42152), .DIN2(_42578), .Q(_42577) );
  nnd2s1 _42653_inst ( .DIN1(_42219), .DIN2(_42379), .Q(_42578) );
  nnd2s1 _42654_inst ( .DIN1(_42292), .DIN2(_42508), .Q(_42576) );
  hi1s1 _42655_inst ( .DIN(_42297), .Q(_42508) );
  nnd2s1 _42656_inst ( .DIN1(_42579), .DIN2(_42580), .Q(
        ____1____________10_____) );
  nnd2s1 _42657_inst ( .DIN1(_42581), .DIN2(_41852), .Q(_42580) );
  xor2s1 _42658_inst ( .DIN1(_26298), .DIN2(_53414), .Q(_42581) );
  nor2s1 _42659_inst ( .DIN1(_41858), .DIN2(_42582), .Q(_42579) );
  nor2s1 _42660_inst ( .DIN1(_42583), .DIN2(_42584), .Q(_42582) );
  nnd2s1 _42661_inst ( .DIN1(_42585), .DIN2(_42586), .Q(_42584) );
  nor2s1 _42662_inst ( .DIN1(_42587), .DIN2(_42588), .Q(_42586) );
  nnd2s1 _42663_inst ( .DIN1(_41866), .DIN2(_42589), .Q(_42588) );
  and2s1 _42664_inst ( .DIN1(_42590), .DIN2(_42591), .Q(_41866) );
  nor2s1 _42665_inst ( .DIN1(_42592), .DIN2(_42593), .Q(_42591) );
  nnd2s1 _42666_inst ( .DIN1(_42494), .DIN2(_42369), .Q(_42593) );
  nnd2s1 _42667_inst ( .DIN1(_42444), .DIN2(_26837), .Q(_42369) );
  nnd2s1 _42668_inst ( .DIN1(_42312), .DIN2(_42594), .Q(_42494) );
  nnd2s1 _42669_inst ( .DIN1(_42385), .DIN2(_42024), .Q(_42594) );
  nnd2s1 _42670_inst ( .DIN1(_42595), .DIN2(_42596), .Q(_42024) );
  nor2s1 _42671_inst ( .DIN1(_42597), .DIN2(_42598), .Q(_42595) );
  nnd2s1 _42672_inst ( .DIN1(_42599), .DIN2(_42600), .Q(_42385) );
  nnd2s1 _42673_inst ( .DIN1(_42399), .DIN2(_42003), .Q(_42592) );
  nnd2s1 _42674_inst ( .DIN1(_42601), .DIN2(_26837), .Q(_42003) );
  nnd2s1 _42675_inst ( .DIN1(_42093), .DIN2(_42189), .Q(_42601) );
  nnd2s1 _42676_inst ( .DIN1(_42602), .DIN2(_42603), .Q(_42189) );
  nnd2s1 _42677_inst ( .DIN1(_42292), .DIN2(_42504), .Q(_42399) );
  nor2s1 _42678_inst ( .DIN1(_41852), .DIN2(_42604), .Q(_42590) );
  nnd2s1 _42679_inst ( .DIN1(_42185), .DIN2(_42246), .Q(_42604) );
  and2s1 _42680_inst ( .DIN1(_42605), .DIN2(_42606), .Q(_42185) );
  nnd2s1 _42681_inst ( .DIN1(_42607), .DIN2(_42371), .Q(_42606) );
  nor2s1 _42682_inst ( .DIN1(_42000), .DIN2(_42608), .Q(_42605) );
  nor2s1 _42683_inst ( .DIN1(_42609), .DIN2(_42423), .Q(_42608) );
  nnd2s1 _42684_inst ( .DIN1(_42610), .DIN2(_42611), .Q(_42587) );
  nnd2s1 _42685_inst ( .DIN1(_42534), .DIN2(_42264), .Q(_42610) );
  nor2s1 _42686_inst ( .DIN1(_42612), .DIN2(_42613), .Q(_42534) );
  nor2s1 _42687_inst ( .DIN1(_42614), .DIN2(_42615), .Q(_42585) );
  nnd2s1 _42688_inst ( .DIN1(_42555), .DIN2(_42322), .Q(_42615) );
  and2s1 _42689_inst ( .DIN1(_42616), .DIN2(_42179), .Q(_42322) );
  and2s1 _42690_inst ( .DIN1(_42617), .DIN2(_42618), .Q(_42179) );
  nnd2s1 _42691_inst ( .DIN1(_42495), .DIN2(_42371), .Q(_42618) );
  nnd2s1 _42692_inst ( .DIN1(_42265), .DIN2(_26837), .Q(_42617) );
  hi1s1 _42693_inst ( .DIN(_42023), .Q(_42265) );
  nor2s1 _42694_inst ( .DIN1(_41970), .DIN2(_42619), .Q(_42616) );
  nor2s1 _42695_inst ( .DIN1(_42533), .DIN2(_42502), .Q(_42619) );
  nnd2s1 _42696_inst ( .DIN1(_42568), .DIN2(_42603), .Q(_42502) );
  hi1s1 _42697_inst ( .DIN(_42045), .Q(_41970) );
  nnd2s1 _42698_inst ( .DIN1(_42620), .DIN2(_42621), .Q(_42045) );
  nor2s1 _42699_inst ( .DIN1(_41903), .DIN2(_36202), .Q(_42620) );
  and2s1 _42700_inst ( .DIN1(_42622), .DIN2(_42623), .Q(_42555) );
  nor2s1 _42701_inst ( .DIN1(_42624), .DIN2(_42625), .Q(_42623) );
  nnd2s1 _42702_inst ( .DIN1(_42626), .DIN2(_42627), .Q(_42624) );
  nnd2s1 _42703_inst ( .DIN1(_42160), .DIN2(_42628), .Q(_42627) );
  nnd2s1 _42704_inst ( .DIN1(_42629), .DIN2(_42630), .Q(_42628) );
  and2s1 _42705_inst ( .DIN1(_42631), .DIN2(_42632), .Q(_42626) );
  nor2s1 _42706_inst ( .DIN1(_42633), .DIN2(_42634), .Q(_42622) );
  nnd2s1 _42707_inst ( .DIN1(_42635), .DIN2(_42343), .Q(_42634) );
  nor2s1 _42708_inst ( .DIN1(_42227), .DIN2(_42636), .Q(_42343) );
  and2s1 _42709_inst ( .DIN1(_42257), .DIN2(_41896), .Q(_42636) );
  nnd2s1 _42710_inst ( .DIN1(_42637), .DIN2(_42638), .Q(_42227) );
  nnd2s1 _42711_inst ( .DIN1(_42639), .DIN2(_37012), .Q(_42638) );
  nor2s1 _42712_inst ( .DIN1(_42462), .DIN2(_42640), .Q(_42639) );
  nnd2s1 _42713_inst ( .DIN1(_42641), .DIN2(_42479), .Q(_42637) );
  nor2s1 _42714_inst ( .DIN1(_36065), .DIN2(_42387), .Q(_42641) );
  xor2s1 _42715_inst ( .DIN1(_42642), .DIN2(_28195), .Q(_42635) );
  hi1s1 _42716_inst ( .DIN(_41043), .Q(_28195) );
  nnd2s1 _42717_inst ( .DIN1(_42643), .DIN2(_42644), .Q(_42642) );
  nor2s1 _42718_inst ( .DIN1(_42645), .DIN2(_42646), .Q(_42644) );
  nnd2s1 _42719_inst ( .DIN1(_42110), .DIN2(_42433), .Q(_42646) );
  nnd2s1 _42720_inst ( .DIN1(_42370), .DIN2(_26837), .Q(_42433) );
  nnd2s1 _42721_inst ( .DIN1(_42004), .DIN2(_41827), .Q(_42645) );
  nnd2s1 _42722_inst ( .DIN1(_42264), .DIN2(_42311), .Q(_41827) );
  and2s1 _42723_inst ( .DIN1(_42647), .DIN2(_28595), .Q(_42311) );
  hi1s1 _42724_inst ( .DIN(_35688), .Q(_28595) );
  nor2s1 _42725_inst ( .DIN1(_36201), .DIN2(_37923), .Q(_42647) );
  nnd2s1 _42726_inst ( .DIN1(_42648), .DIN2(_36208), .Q(_42004) );
  hi1s1 _42727_inst ( .DIN(_42649), .Q(_36208) );
  nor2s1 _42728_inst ( .DIN1(_42650), .DIN2(_42388), .Q(_42648) );
  nor2s1 _42729_inst ( .DIN1(_42651), .DIN2(_42652), .Q(_42643) );
  nnd2s1 _42730_inst ( .DIN1(_42360), .DIN2(_42381), .Q(_42652) );
  xnr2s1 _42731_inst ( .DIN1(_42454), .DIN2(_27840), .Q(_42381) );
  xor2s1 _42732_inst ( .DIN1(_27338), .DIN2(_42653), .Q(_42360) );
  nor2s1 _42733_inst ( .DIN1(_42650), .DIN2(_42224), .Q(_42653) );
  nnd2s1 _42734_inst ( .DIN1(_42475), .DIN2(_41887), .Q(_42633) );
  and2s1 _42735_inst ( .DIN1(_42654), .DIN2(_42655), .Q(_41887) );
  nor2s1 _42736_inst ( .DIN1(_42656), .DIN2(_42657), .Q(_42655) );
  nor2s1 _42737_inst ( .DIN1(_42052), .DIN2(_42200), .Q(_42657) );
  hi1s1 _42738_inst ( .DIN(_42310), .Q(_42656) );
  nnd2s1 _42739_inst ( .DIN1(_42302), .DIN2(_26842), .Q(_42310) );
  nor2s1 _42740_inst ( .DIN1(_42658), .DIN2(_41963), .Q(_42654) );
  nnd2s1 _42741_inst ( .DIN1(_42659), .DIN2(_42660), .Q(_41963) );
  nnd2s1 _42742_inst ( .DIN1(_42408), .DIN2(_41818), .Q(_42660) );
  nnd2s1 _42743_inst ( .DIN1(_42462), .DIN2(_42661), .Q(_41818) );
  and2s1 _42744_inst ( .DIN1(_42662), .DIN2(_42663), .Q(_42475) );
  nnd2s1 _42745_inst ( .DIN1(_42664), .DIN2(_42665), .Q(_42663) );
  nor2s1 _42746_inst ( .DIN1(_37034), .DIN2(_42407), .Q(_42664) );
  or2s1 _42747_inst ( .DIN1(_42177), .DIN2(_42014), .Q(_42614) );
  nnd2s1 _42748_inst ( .DIN1(_42666), .DIN2(_42667), .Q(_42014) );
  nor2s1 _42749_inst ( .DIN1(_42668), .DIN2(_42669), .Q(_42667) );
  nor2s1 _42750_inst ( .DIN1(_42083), .DIN2(_42297), .Q(_42669) );
  nnd2s1 _42751_inst ( .DIN1(_42670), .DIN2(_42671), .Q(_42297) );
  nor2s1 _42752_inst ( .DIN1(_42598), .DIN2(_42672), .Q(_42670) );
  nor2s1 _42753_inst ( .DIN1(_42673), .DIN2(_41944), .Q(_42668) );
  nor2s1 _42754_inst ( .DIN1(_41946), .DIN2(_42285), .Q(_42673) );
  hi1s1 _42755_inst ( .DIN(_42219), .Q(_42285) );
  hi1s1 _42756_inst ( .DIN(_42674), .Q(_41946) );
  nor2s1 _42757_inst ( .DIN1(_42173), .DIN2(_42195), .Q(_42666) );
  nnd2s1 _42758_inst ( .DIN1(_42675), .DIN2(_42676), .Q(_42173) );
  hi1s1 _42759_inst ( .DIN(_42677), .Q(_42675) );
  nnd2s1 _42760_inst ( .DIN1(_42678), .DIN2(_42679), .Q(_42177) );
  nor2s1 _42761_inst ( .DIN1(_42680), .DIN2(_42681), .Q(_42679) );
  or2s1 _42762_inst ( .DIN1(_42121), .DIN2(_41888), .Q(_42681) );
  nnd2s1 _42763_inst ( .DIN1(_42682), .DIN2(_42683), .Q(_41888) );
  nor2s1 _42764_inst ( .DIN1(_42684), .DIN2(_42685), .Q(_42683) );
  nor2s1 _42765_inst ( .DIN1(_39313), .DIN2(_42686), .Q(_42685) );
  or2s1 _42766_inst ( .DIN1(_42687), .DIN2(_42533), .Q(_42686) );
  nor2s1 _42767_inst ( .DIN1(_42228), .DIN2(_42688), .Q(_42684) );
  nnd2s1 _42768_inst ( .DIN1(_36060), .DIN2(_42292), .Q(_42688) );
  nor2s1 _42769_inst ( .DIN1(_42689), .DIN2(_42690), .Q(_42682) );
  nor2s1 _42770_inst ( .DIN1(_42049), .DIN2(_42115), .Q(_42690) );
  nor2s1 _42771_inst ( .DIN1(_42407), .DIN2(_42691), .Q(_42689) );
  nnd2s1 _42772_inst ( .DIN1(_37334), .DIN2(_42692), .Q(_42691) );
  nnd2s1 _42773_inst ( .DIN1(_42693), .DIN2(_41873), .Q(_42121) );
  and2s1 _42774_inst ( .DIN1(_42694), .DIN2(_42695), .Q(_41873) );
  nnd2s1 _42775_inst ( .DIN1(_42696), .DIN2(_42570), .Q(_42695) );
  nor2s1 _42776_inst ( .DIN1(_37211), .DIN2(_37670), .Q(_42570) );
  nor2s1 _42777_inst ( .DIN1(_39040), .DIN2(_42153), .Q(_42696) );
  nnd2s1 _42778_inst ( .DIN1(_42697), .DIN2(_42698), .Q(_42694) );
  nor2s1 _42779_inst ( .DIN1(_35686), .DIN2(_37323), .Q(_42697) );
  nor2s1 _42780_inst ( .DIN1(_42699), .DIN2(_42700), .Q(_42693) );
  nor2s1 _42781_inst ( .DIN1(_42342), .DIN2(_42701), .Q(_42699) );
  nnd2s1 _42782_inst ( .DIN1(_42702), .DIN2(_42703), .Q(_42680) );
  nor2s1 _42783_inst ( .DIN1(_42704), .DIN2(_42705), .Q(_42678) );
  nnd2s1 _42784_inst ( .DIN1(_42706), .DIN2(_42557), .Q(_42705) );
  and2s1 _42785_inst ( .DIN1(_42707), .DIN2(_42708), .Q(_42557) );
  nor2s1 _42786_inst ( .DIN1(_42361), .DIN2(_42709), .Q(_42708) );
  nnd2s1 _42787_inst ( .DIN1(_42089), .DIN2(_42368), .Q(_42709) );
  nnd2s1 _42788_inst ( .DIN1(_42710), .DIN2(_41830), .Q(_42089) );
  hi1s1 _42789_inst ( .DIN(_41969), .Q(_42361) );
  nnd2s1 _42790_inst ( .DIN1(_42711), .DIN2(_42712), .Q(_41969) );
  nor2s1 _42791_inst ( .DIN1(_37810), .DIN2(_42533), .Q(_42712) );
  nor2s1 _42792_inst ( .DIN1(_35270), .DIN2(_39042), .Q(_42711) );
  nor2s1 _42793_inst ( .DIN1(_42030), .DIN2(_42713), .Q(_42707) );
  nor2s1 _42794_inst ( .DIN1(_42387), .DIN2(_42714), .Q(_42713) );
  nor2s1 _42795_inst ( .DIN1(_41903), .DIN2(_42354), .Q(_42030) );
  nnd2s1 _42796_inst ( .DIN1(_42715), .DIN2(_37467), .Q(_42354) );
  nor2s1 _42797_inst ( .DIN1(_35104), .DIN2(_35686), .Q(_42715) );
  hi1s1 _42798_inst ( .DIN(_42349), .Q(_42706) );
  nnd2s1 _42799_inst ( .DIN1(_42716), .DIN2(_42717), .Q(_42349) );
  nor2s1 _42800_inst ( .DIN1(_42064), .DIN2(_42718), .Q(_42717) );
  hi1s1 _42801_inst ( .DIN(_42719), .Q(_42718) );
  nor2s1 _42802_inst ( .DIN1(_42043), .DIN2(_42720), .Q(_42716) );
  nor2s1 _42803_inst ( .DIN1(_42049), .DIN2(_42571), .Q(_42720) );
  and2s1 _42804_inst ( .DIN1(_42721), .DIN2(_42698), .Q(_42043) );
  hi1s1 _42805_inst ( .DIN(_41996), .Q(_42698) );
  nnd2s1 _42806_inst ( .DIN1(_36694), .DIN2(_42312), .Q(_41996) );
  nor2s1 _42807_inst ( .DIN1(_36065), .DIN2(_39311), .Q(_42721) );
  xor2s1 _42808_inst ( .DIN1(_33214), .DIN2(_42722), .Q(_42704) );
  nnd2s1 _42809_inst ( .DIN1(_42723), .DIN2(_42724), .Q(_42722) );
  nnd2s1 _42810_inst ( .DIN1(_41896), .DIN2(_42725), .Q(_42724) );
  nnd2s1 _42811_inst ( .DIN1(_42528), .DIN2(_42025), .Q(_42723) );
  hi1s1 _42812_inst ( .DIN(_42726), .Q(_42528) );
  nnd2s1 _42813_inst ( .DIN1(_42727), .DIN2(_42728), .Q(_42583) );
  nor2s1 _42814_inst ( .DIN1(_42729), .DIN2(_42730), .Q(_42728) );
  nnd2s1 _42815_inst ( .DIN1(_42731), .DIN2(_42309), .Q(_42730) );
  nnd2s1 _42816_inst ( .DIN1(_42732), .DIN2(_41830), .Q(_42309) );
  nnd2s1 _42817_inst ( .DIN1(_42256), .DIN2(_42062), .Q(_42729) );
  nnd2s1 _42818_inst ( .DIN1(_42733), .DIN2(_42114), .Q(_42062) );
  nnd2s1 _42819_inst ( .DIN1(_42734), .DIN2(_42032), .Q(_42256) );
  nor2s1 _42820_inst ( .DIN1(_42661), .DIN2(_37199), .Q(_42734) );
  nor2s1 _42821_inst ( .DIN1(_42735), .DIN2(_42736), .Q(_42727) );
  nnd2s1 _42822_inst ( .DIN1(_42737), .DIN2(_42738), .Q(_42736) );
  or2s1 _42823_inst ( .DIN1(_42250), .DIN2(_42190), .Q(_42738) );
  nnd2s1 _42824_inst ( .DIN1(_42152), .DIN2(_42550), .Q(_42737) );
  nnd2s1 _42825_inst ( .DIN1(_42739), .DIN2(_42740), .Q(_42735) );
  nnd2s1 _42826_inst ( .DIN1(_41830), .DIN2(_42113), .Q(_42740) );
  nnd2s1 _42827_inst ( .DIN1(_42250), .DIN2(_42741), .Q(_42113) );
  nnd2s1 _42828_inst ( .DIN1(_41906), .DIN2(_42292), .Q(_42739) );
  and2s1 _42829_inst ( .DIN1(_42600), .DIN2(_42742), .Q(_41906) );
  hi1s1 _42830_inst ( .DIN(_41923), .Q(_41858) );
  nnd2s1 _42831_inst ( .DIN1(_42743), .DIN2(_42744), .Q(_41923) );
  nor2s1 _42832_inst ( .DIN1(_41977), .DIN2(_42745), .Q(_42744) );
  nnd2s1 _42833_inst ( .DIN1(_29742), .DIN2(_27446), .Q(_42745) );
  hi1s1 _42834_inst ( .DIN(_41852), .Q(_41977) );
  nnd2s1 _42835_inst ( .DIN1(_42746), .DIN2(_42747), .Q(_41852) );
  nor2s1 _42836_inst ( .DIN1(_29288), .DIN2(_32810), .Q(_42747) );
  nor2s1 _42837_inst ( .DIN1(_27317), .DIN2(_42748), .Q(_42746) );
  nnd2s1 _42838_inst ( .DIN1(_42749), .DIN2(_27446), .Q(_27317) );
  nor2s1 _42839_inst ( .DIN1(_42750), .DIN2(_27310), .Q(_42749) );
  nor2s1 _42840_inst ( .DIN1(_27433), .DIN2(_31404), .Q(_42743) );
  nnd2s1 _42841_inst ( .DIN1(_42751), .DIN2(_42752), .Q(_27433) );
  nor2s1 _42842_inst ( .DIN1(_29288), .DIN2(_42753), .Q(_42752) );
  nor2s1 _42843_inst ( .DIN1(_29433), .DIN2(_32810), .Q(_42751) );
  nnd2s1 _42844_inst ( .DIN1(_42754), .DIN2(_42755), .Q(
        ____1____________0_____) );
  nnd2s1 _42845_inst ( .DIN1(_42756), .DIN2(_29082), .Q(_42755) );
  xor2s1 _42846_inst ( .DIN1(_33835), .DIN2(_53426), .Q(_42756) );
  nnd2s1 _42847_inst ( .DIN1(_53428), .DIN2(_53427), .Q(_33835) );
  nnd2s1 _42848_inst ( .DIN1(_29083), .DIN2(_42757), .Q(_42754) );
  nnd2s1 _42849_inst ( .DIN1(_42758), .DIN2(_42759), .Q(_42757) );
  nor2s1 _42850_inst ( .DIN1(_42760), .DIN2(_42761), .Q(_42759) );
  nnd2s1 _42851_inst ( .DIN1(_42762), .DIN2(_42763), .Q(_42761) );
  nnd2s1 _42852_inst ( .DIN1(_42012), .DIN2(_42764), .Q(_42763) );
  nnd2s1 _42853_inst ( .DIN1(_42765), .DIN2(_42766), .Q(_42764) );
  nnd2s1 _42854_inst ( .DIN1(_37012), .DIN2(_42767), .Q(_42766) );
  nnd2s1 _42855_inst ( .DIN1(_42490), .DIN2(_53131), .Q(_42765) );
  nnd2s1 _42856_inst ( .DIN1(_42401), .DIN2(_42768), .Q(_42762) );
  nnd2s1 _42857_inst ( .DIN1(_42769), .DIN2(_42770), .Q(_42768) );
  nor2s1 _42858_inst ( .DIN1(_42771), .DIN2(_42444), .Q(_42770) );
  and2s1 _42859_inst ( .DIN1(_42742), .DIN2(_42603), .Q(_42444) );
  nor2s1 _42860_inst ( .DIN1(_42772), .DIN2(_42773), .Q(_42769) );
  nor2s1 _42861_inst ( .DIN1(_35270), .DIN2(_42774), .Q(_42773) );
  nor2s1 _42862_inst ( .DIN1(_42338), .DIN2(_42775), .Q(_42772) );
  nnd2s1 _42863_inst ( .DIN1(_37033), .DIN2(_35433), .Q(_42775) );
  hi1s1 _42864_inst ( .DIN(_35103), .Q(_37033) );
  nnd2s1 _42865_inst ( .DIN1(_42776), .DIN2(_42777), .Q(_42760) );
  nnd2s1 _42866_inst ( .DIN1(_42733), .DIN2(_41830), .Q(_42777) );
  nor2s1 _42867_inst ( .DIN1(_42330), .DIN2(_36065), .Q(_42733) );
  nor2s1 _42868_inst ( .DIN1(_42064), .DIN2(_42778), .Q(_42776) );
  nor2s1 _42869_inst ( .DIN1(_42779), .DIN2(_42780), .Q(_42778) );
  nnd2s1 _42870_inst ( .DIN1(_36199), .DIN2(_42264), .Q(_42780) );
  and2s1 _42871_inst ( .DIN1(_42781), .DIN2(_42230), .Q(_42064) );
  nor2s1 _42872_inst ( .DIN1(_41903), .DIN2(_42330), .Q(_42781) );
  nor2s1 _42873_inst ( .DIN1(_42782), .DIN2(_42783), .Q(_42758) );
  nnd2s1 _42874_inst ( .DIN1(_42784), .DIN2(_42346), .Q(_42783) );
  nor2s1 _42875_inst ( .DIN1(_42658), .DIN2(_42785), .Q(_42346) );
  and2s1 _42876_inst ( .DIN1(_42786), .DIN2(_42787), .Q(_42785) );
  nnd2s1 _42877_inst ( .DIN1(_42115), .DIN2(_42788), .Q(_42787) );
  nnd2s1 _42878_inst ( .DIN1(_42789), .DIN2(_37193), .Q(_42788) );
  hi1s1 _42879_inst ( .DIN(_37323), .Q(_37193) );
  nnd2s1 _42880_inst ( .DIN1(_42479), .DIN2(_37012), .Q(_42115) );
  hi1s1 _42881_inst ( .DIN(_36949), .Q(_37012) );
  nnd2s1 _42882_inst ( .DIN1(_42790), .DIN2(_42791), .Q(_36949) );
  xor2s1 _42883_inst ( .DIN1(_32716), .DIN2(_42792), .Q(_42658) );
  and2s1 _42884_inst ( .DIN1(_37189), .DIN2(_42290), .Q(_42792) );
  nor2s1 _42885_inst ( .DIN1(_42161), .DIN2(_41903), .Q(_42290) );
  xor2s1 _42886_inst ( .DIN1(_42793), .DIN2(_30912), .Q(_42784) );
  hi1s1 _42887_inst ( .DIN(_30360), .Q(_30912) );
  nnd2s1 _42888_inst ( .DIN1(_42794), .DIN2(_42795), .Q(_30360) );
  nor2s1 _42889_inst ( .DIN1(_42796), .DIN2(_42797), .Q(_42795) );
  nor2s1 _42890_inst ( .DIN1(_42798), .DIN2(_42799), .Q(_42794) );
  nnd2s1 _42891_inst ( .DIN1(_42800), .DIN2(_42801), .Q(_42793) );
  nor2s1 _42892_inst ( .DIN1(_42802), .DIN2(_42803), .Q(_42801) );
  nnd2s1 _42893_inst ( .DIN1(_42396), .DIN2(_42804), .Q(_42803) );
  hi1s1 _42894_inst ( .DIN(_41820), .Q(_42804) );
  nnd2s1 _42895_inst ( .DIN1(_42805), .DIN2(_42806), .Q(_41820) );
  nor2s1 _42896_inst ( .DIN1(_42125), .DIN2(_42807), .Q(_42806) );
  nnd2s1 _42897_inst ( .DIN1(_42731), .DIN2(_42470), .Q(_42807) );
  or2s1 _42898_inst ( .DIN1(_42200), .DIN2(_41903), .Q(_42470) );
  nnd2s1 _42899_inst ( .DIN1(_42808), .DIN2(_37467), .Q(_42200) );
  nor2s1 _42900_inst ( .DIN1(_35686), .DIN2(_36065), .Q(_42808) );
  nnd2s1 _42901_inst ( .DIN1(_42192), .DIN2(_42012), .Q(_42731) );
  and2s1 _42902_inst ( .DIN1(_42809), .DIN2(_37189), .Q(_42192) );
  nor2s1 _42903_inst ( .DIN1(_37670), .DIN2(_39314), .Q(_42809) );
  nnd2s1 _42904_inst ( .DIN1(_42810), .DIN2(_42811), .Q(_42125) );
  and2s1 _42905_inst ( .DIN1(_42368), .DIN2(_42380), .Q(_42811) );
  nnd2s1 _42906_inst ( .DIN1(_42812), .DIN2(_42665), .Q(_42380) );
  nor2s1 _42907_inst ( .DIN1(_37995), .DIN2(_39312), .Q(_42665) );
  nor2s1 _42908_inst ( .DIN1(_42153), .DIN2(_37034), .Q(_42812) );
  nnd2s1 _42909_inst ( .DIN1(_42813), .DIN2(_42814), .Q(_42368) );
  nor2s1 _42910_inst ( .DIN1(_36065), .DIN2(_42338), .Q(_42814) );
  nor2s1 _42911_inst ( .DIN1(_42407), .DIN2(_39042), .Q(_42813) );
  nor2s1 _42912_inst ( .DIN1(_42815), .DIN2(_42816), .Q(_42810) );
  nor2s1 _42913_inst ( .DIN1(_42609), .DIN2(_42726), .Q(_42816) );
  nnd2s1 _42914_inst ( .DIN1(_42567), .DIN2(_42742), .Q(_42726) );
  nor2s1 _42915_inst ( .DIN1(_42817), .DIN2(_42597), .Q(_42742) );
  nor2s1 _42916_inst ( .DIN1(_42025), .DIN2(_42264), .Q(_42609) );
  hi1s1 _42917_inst ( .DIN(_42363), .Q(_42264) );
  nor2s1 _42918_inst ( .DIN1(_42649), .DIN2(_42818), .Q(_42815) );
  nnd2s1 _42919_inst ( .DIN1(_42152), .DIN2(_42819), .Q(_42818) );
  nor2s1 _42920_inst ( .DIN1(_41956), .DIN2(_42625), .Q(_42805) );
  nnd2s1 _42921_inst ( .DIN1(_42820), .DIN2(_42821), .Q(_42625) );
  hi1s1 _42922_inst ( .DIN(_42220), .Q(_42821) );
  nnd2s1 _42923_inst ( .DIN1(_42822), .DIN2(_42823), .Q(_42220) );
  nnd2s1 _42924_inst ( .DIN1(_41896), .DIN2(_42305), .Q(_42823) );
  nnd2s1 _42925_inst ( .DIN1(_42824), .DIN2(_42825), .Q(_42305) );
  or2s1 _42926_inst ( .DIN1(_36202), .DIN2(_42353), .Q(_42825) );
  nnd2s1 _42927_inst ( .DIN1(_38017), .DIN2(_37673), .Q(_42353) );
  nnd2s1 _42928_inst ( .DIN1(_42032), .DIN2(_37194), .Q(_42824) );
  hi1s1 _42929_inst ( .DIN(_42161), .Q(_42032) );
  nnd2s1 _42930_inst ( .DIN1(_42284), .DIN2(_42312), .Q(_42822) );
  hi1s1 _42931_inst ( .DIN(_41908), .Q(_42284) );
  nnd2s1 _42932_inst ( .DIN1(_42826), .DIN2(_36203), .Q(_41908) );
  nor2s1 _42933_inst ( .DIN1(_42338), .DIN2(_39042), .Q(_42826) );
  and2s1 _42934_inst ( .DIN1(_42451), .DIN2(_42827), .Q(_42820) );
  or2s1 _42935_inst ( .DIN1(_42105), .DIN2(_42049), .Q(_42827) );
  nor2s1 _42936_inst ( .DIN1(_42547), .DIN2(_42786), .Q(_42049) );
  hi1s1 _42937_inst ( .DIN(_42104), .Q(_42547) );
  nnd2s1 _42938_inst ( .DIN1(_42828), .DIN2(_36063), .Q(_42105) );
  nor2s1 _42939_inst ( .DIN1(_35533), .DIN2(_42338), .Q(_42828) );
  nnd2s1 _42940_inst ( .DIN1(_42829), .DIN2(_36063), .Q(_42451) );
  nor2s1 _42941_inst ( .DIN1(_42330), .DIN2(_42052), .Q(_42829) );
  nnd2s1 _42942_inst ( .DIN1(_42830), .DIN2(_42831), .Q(_41956) );
  nor2s1 _42943_inst ( .DIN1(_42832), .DIN2(_42833), .Q(_42831) );
  nnd2s1 _42944_inst ( .DIN1(_42834), .DIN2(_42454), .Q(_42833) );
  nnd2s1 _42945_inst ( .DIN1(_42835), .DIN2(_42450), .Q(_42454) );
  nor2s1 _42946_inst ( .DIN1(_37923), .DIN2(_39040), .Q(_42450) );
  nor2s1 _42947_inst ( .DIN1(_42153), .DIN2(_35930), .Q(_42835) );
  nnd2s1 _42948_inst ( .DIN1(_42836), .DIN2(_36063), .Q(_42834) );
  nor2s1 _42949_inst ( .DIN1(_42533), .DIN2(_42774), .Q(_42836) );
  nor2s1 _42950_inst ( .DIN1(_42837), .DIN2(_42838), .Q(_42832) );
  nnd2s1 _42951_inst ( .DIN1(_37334), .DIN2(_42258), .Q(_42838) );
  nor2s1 _42952_inst ( .DIN1(_42496), .DIN2(_42839), .Q(_42830) );
  nnd2s1 _42953_inst ( .DIN1(_42611), .DIN2(_42840), .Q(_42839) );
  nnd2s1 _42954_inst ( .DIN1(_42370), .DIN2(_42401), .Q(_42840) );
  nor2s1 _42955_inst ( .DIN1(_35930), .DIN2(_42293), .Q(_42370) );
  nnd2s1 _42956_inst ( .DIN1(_42151), .DIN2(_42312), .Q(_42611) );
  hi1s1 _42957_inst ( .DIN(_42268), .Q(_42151) );
  nnd2s1 _42958_inst ( .DIN1(_42841), .DIN2(_42567), .Q(_42268) );
  nor2s1 _42959_inst ( .DIN1(_42842), .DIN2(_42817), .Q(_42841) );
  nnd2s1 _42960_inst ( .DIN1(_42843), .DIN2(_42844), .Q(_42496) );
  nnd2s1 _42961_inst ( .DIN1(_26842), .DIN2(_42152), .Q(_42844) );
  hi1s1 _42962_inst ( .DIN(_40754), .Q(_40581) );
  nnd2s1 _42963_inst ( .DIN1(_42845), .DIN2(_42846), .Q(_40754) );
  nor2s1 _42964_inst ( .DIN1(_37211), .DIN2(_37995), .Q(_42845) );
  nor2s1 _42965_inst ( .DIN1(_42847), .DIN2(_42848), .Q(_42843) );
  nor2s1 _42966_inst ( .DIN1(_42161), .DIN2(_42849), .Q(_42848) );
  nnd2s1 _42967_inst ( .DIN1(_42012), .DIN2(_37197), .Q(_42849) );
  nor2s1 _42968_inst ( .DIN1(_35930), .DIN2(_42850), .Q(_42847) );
  nnd2s1 _42969_inst ( .DIN1(_42819), .DIN2(_42401), .Q(_42850) );
  nor2s1 _42970_inst ( .DIN1(_42700), .DIN2(_42851), .Q(_42396) );
  and2s1 _42971_inst ( .DIN1(_42152), .DIN2(_42463), .Q(_42851) );
  nor2s1 _42972_inst ( .DIN1(_42852), .DIN2(_42853), .Q(_42463) );
  hi1s1 _42973_inst ( .DIN(_42225), .Q(_42152) );
  nnd2s1 _42974_inst ( .DIN1(_42854), .DIN2(_42855), .Q(_42700) );
  nnd2s1 _42975_inst ( .DIN1(_42856), .DIN2(_42857), .Q(_42855) );
  nor2s1 _42976_inst ( .DIN1(_41935), .DIN2(_35930), .Q(_42856) );
  nnd2s1 _42977_inst ( .DIN1(_42858), .DIN2(_42231), .Q(_42854) );
  nor2s1 _42978_inst ( .DIN1(_36066), .DIN2(_42859), .Q(_42858) );
  nnd2s1 _42979_inst ( .DIN1(_42860), .DIN2(_42028), .Q(_42802) );
  and2s1 _42980_inst ( .DIN1(_42861), .DIN2(_42862), .Q(_42028) );
  nor2s1 _42981_inst ( .DIN1(_42863), .DIN2(_42864), .Q(_42862) );
  nnd2s1 _42982_inst ( .DIN1(_42865), .DIN2(_42472), .Q(_42864) );
  nnd2s1 _42983_inst ( .DIN1(_42408), .DIN2(_42012), .Q(_42472) );
  and2s1 _42984_inst ( .DIN1(_42866), .DIN2(_38017), .Q(_42408) );
  hi1s1 _42985_inst ( .DIN(_35534), .Q(_38017) );
  nor2s1 _42986_inst ( .DIN1(_37995), .DIN2(_36201), .Q(_42866) );
  nnd2s1 _42987_inst ( .DIN1(_42607), .DIN2(_42401), .Q(_42865) );
  hi1s1 _42988_inst ( .DIN(_42342), .Q(_42401) );
  hi1s1 _42989_inst ( .DIN(_42251), .Q(_42607) );
  nnd2s1 _42990_inst ( .DIN1(_36203), .DIN2(_42341), .Q(_42251) );
  hi1s1 _42991_inst ( .DIN(_42859), .Q(_42341) );
  nnd2s1 _42992_inst ( .DIN1(_42659), .DIN2(_42236), .Q(_42863) );
  nnd2s1 _42993_inst ( .DIN1(_42867), .DIN2(_42312), .Q(_42236) );
  nnd2s1 _42994_inst ( .DIN1(_42868), .DIN2(_42741), .Q(_42867) );
  nnd2s1 _42995_inst ( .DIN1(_42869), .DIN2(_42671), .Q(_42741) );
  nor2s1 _42996_inst ( .DIN1(_26279), .DIN2(_26539), .Q(_42671) );
  nor2s1 _42997_inst ( .DIN1(_42672), .DIN2(_42870), .Q(_42869) );
  xor2s1 _42998_inst ( .DIN1(_28860), .DIN2(_42550), .Q(_42868) );
  hi1s1 _42999_inst ( .DIN(_42106), .Q(_42550) );
  nnd2s1 _43000_inst ( .DIN1(_42599), .DIN2(_42603), .Q(_42106) );
  hi1s1 _43001_inst ( .DIN(_42598), .Q(_42603) );
  hi1s1 _43002_inst ( .DIN(_33214), .Q(_28860) );
  nnd2s1 _43003_inst ( .DIN1(_42871), .DIN2(_42872), .Q(_33214) );
  nor2s1 _43004_inst ( .DIN1(_42873), .DIN2(_42874), .Q(_42872) );
  nnd2s1 _43005_inst ( .DIN1(_42875), .DIN2(_40395), .Q(_42874) );
  nnd2s1 _43006_inst ( .DIN1(_42876), .DIN2(_42877), .Q(_42873) );
  nor2s1 _43007_inst ( .DIN1(_42878), .DIN2(_42879), .Q(_42871) );
  nnd2s1 _43008_inst ( .DIN1(_42880), .DIN2(_42881), .Q(_42879) );
  nnd2s1 _43009_inst ( .DIN1(_42882), .DIN2(_42883), .Q(_42659) );
  nor2s1 _43010_inst ( .DIN1(_42884), .DIN2(_35103), .Q(_42883) );
  nor2s1 _43011_inst ( .DIN1(_42338), .DIN2(_42387), .Q(_42882) );
  nor2s1 _43012_inst ( .DIN1(_42885), .DIN2(_42886), .Q(_42861) );
  nnd2s1 _43013_inst ( .DIN1(_42186), .DIN2(_42126), .Q(_42886) );
  nor2s1 _43014_inst ( .DIN1(_42651), .DIN2(_42887), .Q(_42126) );
  and2s1 _43015_inst ( .DIN1(_42231), .DIN2(_42471), .Q(_42887) );
  nnd2s1 _43016_inst ( .DIN1(_42888), .DIN2(_42406), .Q(_42471) );
  hi1s1 _43017_inst ( .DIN(_42407), .Q(_42231) );
  xnr2s1 _43018_inst ( .DIN1(_26321), .DIN2(_42889), .Q(_42651) );
  nor2s1 _43019_inst ( .DIN1(_42153), .DIN2(_42406), .Q(_42889) );
  nnd2s1 _43020_inst ( .DIN1(_35929), .DIN2(_42692), .Q(_42406) );
  nor2s1 _43021_inst ( .DIN1(_42842), .DIN2(_53425), .Q(_35929) );
  and2s1 _43022_inst ( .DIN1(_42890), .DIN2(_42891), .Q(_42186) );
  nor2s1 _43023_inst ( .DIN1(_42892), .DIN2(_42893), .Q(_42891) );
  nnd2s1 _43024_inst ( .DIN1(_42894), .DIN2(_42110), .Q(_42893) );
  nnd2s1 _43025_inst ( .DIN1(_42895), .DIN2(_42896), .Q(_42110) );
  hi1s1 _43026_inst ( .DIN(_42774), .Q(_42896) );
  nor2s1 _43027_inst ( .DIN1(_42387), .DIN2(_35270), .Q(_42895) );
  nnd2s1 _43028_inst ( .DIN1(_42054), .DIN2(_42312), .Q(_42894) );
  and2s1 _43029_inst ( .DIN1(_42897), .DIN2(_39317), .Q(_42054) );
  nor2s1 _43030_inst ( .DIN1(_37810), .DIN2(_36207), .Q(_42897) );
  nor2s1 _43031_inst ( .DIN1(_42190), .DIN2(_42250), .Q(_42892) );
  nnd2s1 _43032_inst ( .DIN1(_42898), .DIN2(_37467), .Q(_42250) );
  nor2s1 _43033_inst ( .DIN1(_35104), .DIN2(_28567), .Q(_42898) );
  hi1s1 _43034_inst ( .DIN(_28599), .Q(_28567) );
  nor2s1 _43035_inst ( .DIN1(_42481), .DIN2(_42085), .Q(_42890) );
  nnd2s1 _43036_inst ( .DIN1(_42899), .DIN2(_42900), .Q(_42085) );
  nnd2s1 _43037_inst ( .DIN1(_42901), .DIN2(_35113), .Q(_42900) );
  nor2s1 _43038_inst ( .DIN1(_42545), .DIN2(_42407), .Q(_42901) );
  nnd2s1 _43039_inst ( .DIN1(_42490), .DIN2(_42160), .Q(_42899) );
  hi1s1 _43040_inst ( .DIN(_42630), .Q(_42490) );
  nnd2s1 _43041_inst ( .DIN1(_42902), .DIN2(_35433), .Q(_42630) );
  hi1s1 _43042_inst ( .DIN(_42884), .Q(_35433) );
  nor2s1 _43043_inst ( .DIN1(_37810), .DIN2(_37323), .Q(_42902) );
  nnd2s1 _43044_inst ( .DIN1(_42903), .DIN2(_42904), .Q(_42481) );
  nnd2s1 _43045_inst ( .DIN1(_42905), .DIN2(_42371), .Q(_42904) );
  nor2s1 _43046_inst ( .DIN1(_36207), .DIN2(_42859), .Q(_42905) );
  nnd2s1 _43047_inst ( .DIN1(_28599), .DIN2(_37468), .Q(_42859) );
  nnd2s1 _43048_inst ( .DIN1(_42906), .DIN2(_42907), .Q(_36207) );
  nnd2s1 _43049_inst ( .DIN1(_42908), .DIN2(_41830), .Q(_42903) );
  hi1s1 _43050_inst ( .DIN(_42249), .Q(_41830) );
  nnd2s1 _43051_inst ( .DIN1(_42246), .DIN2(_42909), .Q(_42885) );
  nnd2s1 _43052_inst ( .DIN1(_42786), .DIN2(_42552), .Q(_42909) );
  nnd2s1 _43053_inst ( .DIN1(_41936), .DIN2(_42050), .Q(_42552) );
  nnd2s1 _43054_inst ( .DIN1(_42910), .DIN2(_42846), .Q(_42050) );
  nnd2s1 _43055_inst ( .DIN1(_42819), .DIN2(_37189), .Q(_41936) );
  hi1s1 _43056_inst ( .DIN(_41935), .Q(_42786) );
  xor2s1 _43057_inst ( .DIN1(_31269), .DIN2(_42911), .Q(_42246) );
  nor2s1 _43058_inst ( .DIN1(_42852), .DIN2(_42912), .Q(_42911) );
  nnd2s1 _43059_inst ( .DIN1(_42913), .DIN2(_42312), .Q(_42912) );
  nnd2s1 _43060_inst ( .DIN1(_42914), .DIN2(_42596), .Q(_42852) );
  nor2s1 _43061_inst ( .DIN1(_42000), .DIN2(_42392), .Q(_42860) );
  nnd2s1 _43062_inst ( .DIN1(_42702), .DIN2(_42915), .Q(_42392) );
  nnd2s1 _43063_inst ( .DIN1(_42771), .DIN2(_42371), .Q(_42915) );
  hi1s1 _43064_inst ( .DIN(_42714), .Q(_42771) );
  nnd2s1 _43065_inst ( .DIN1(_37671), .DIN2(_42916), .Q(_42714) );
  nnd2s1 _43066_inst ( .DIN1(_42917), .DIN2(_42918), .Q(_42916) );
  nnd2s1 _43067_inst ( .DIN1(_36456), .DIN2(_28596), .Q(_42917) );
  xor2s1 _43068_inst ( .DIN1(_31222), .DIN2(_36694), .Q(_37671) );
  nnd2s1 _43069_inst ( .DIN1(_42919), .DIN2(_42920), .Q(_31222) );
  nor2s1 _43070_inst ( .DIN1(_42921), .DIN2(_42922), .Q(_42920) );
  nnd2s1 _43071_inst ( .DIN1(_42923), .DIN2(_42924), .Q(_42922) );
  nor2s1 _43072_inst ( .DIN1(_42925), .DIN2(_42926), .Q(_42919) );
  nnd2s1 _43073_inst ( .DIN1(_42927), .DIN2(_42928), .Q(_42926) );
  nnd2s1 _43074_inst ( .DIN1(_42315), .DIN2(_41896), .Q(_42702) );
  nor2s1 _43075_inst ( .DIN1(_42388), .DIN2(_37034), .Q(_42315) );
  nnd2s1 _43076_inst ( .DIN1(_42929), .DIN2(_42906), .Q(_37034) );
  and2s1 _43077_inst ( .DIN1(_42930), .DIN2(_42479), .Q(_42000) );
  hi1s1 _43078_inst ( .DIN(_42837), .Q(_42479) );
  nnd2s1 _43079_inst ( .DIN1(_39317), .DIN2(_37468), .Q(_42837) );
  hi1s1 _43080_inst ( .DIN(_39042), .Q(_39317) );
  nor2s1 _43081_inst ( .DIN1(_36065), .DIN2(_42342), .Q(_42930) );
  nor2s1 _43082_inst ( .DIN1(_42931), .DIN2(_42932), .Q(_42800) );
  nnd2s1 _43083_inst ( .DIN1(_42933), .DIN2(_42934), .Q(_42932) );
  hi1s1 _43084_inst ( .DIN(_42464), .Q(_42934) );
  nnd2s1 _43085_inst ( .DIN1(_42935), .DIN2(_42936), .Q(_42464) );
  nor2s1 _43086_inst ( .DIN1(_42937), .DIN2(_42938), .Q(_42936) );
  nnd2s1 _43087_inst ( .DIN1(_42939), .DIN2(_42940), .Q(_42938) );
  nnd2s1 _43088_inst ( .DIN1(_41819), .DIN2(_42160), .Q(_42940) );
  hi1s1 _43089_inst ( .DIN(_42629), .Q(_41819) );
  nnd2s1 _43090_inst ( .DIN1(_42941), .DIN2(_42230), .Q(_42629) );
  hi1s1 _43091_inst ( .DIN(_35269), .Q(_42230) );
  nor2s1 _43092_inst ( .DIN1(_42677), .DIN2(_42942), .Q(_42939) );
  nor2s1 _43093_inst ( .DIN1(_41935), .DIN2(_42571), .Q(_42942) );
  nnd2s1 _43094_inst ( .DIN1(_42941), .DIN2(_36203), .Q(_42571) );
  nor2s1 _43095_inst ( .DIN1(_37810), .DIN2(_39042), .Q(_42941) );
  nnd2s1 _43096_inst ( .DIN1(_42943), .DIN2(_42944), .Q(_39042) );
  nnd2s1 _43097_inst ( .DIN1(_42312), .DIN2(_42945), .Q(_41935) );
  nnd2s1 _43098_inst ( .DIN1(_42946), .DIN2(______[29]), .Q(_42945) );
  nor2s1 _43099_inst ( .DIN1(______[11]), .DIN2(_39015), .Q(_42946) );
  nor2s1 _43100_inst ( .DIN1(_42947), .DIN2(_42330), .Q(_42677) );
  nnd2s1 _43101_inst ( .DIN1(_42312), .DIN2(_37334), .Q(_42947) );
  nnd2s1 _43102_inst ( .DIN1(_42948), .DIN2(_42719), .Q(_42937) );
  nnd2s1 _43103_inst ( .DIN1(_42949), .DIN2(_36063), .Q(_42719) );
  hi1s1 _43104_inst ( .DIN(_37320), .Q(_36063) );
  nnd2s1 _43105_inst ( .DIN1(_42791), .DIN2(_42950), .Q(_37320) );
  nor2s1 _43106_inst ( .DIN1(_42363), .DIN2(_42774), .Q(_42949) );
  nnd2s1 _43107_inst ( .DIN1(_28597), .DIN2(_37468), .Q(_42774) );
  nnd2s1 _43108_inst ( .DIN1(_42312), .DIN2(_42951), .Q(_42363) );
  nnd2s1 _43109_inst ( .DIN1(_42952), .DIN2(______[11]), .Q(_42951) );
  nor2s1 _43110_inst ( .DIN1(_41939), .DIN2(_42061), .Q(_42948) );
  nor2s1 _43111_inst ( .DIN1(_41944), .DIN2(_42224), .Q(_42061) );
  nnd2s1 _43112_inst ( .DIN1(_42819), .DIN2(_35114), .Q(_42224) );
  hi1s1 _43113_inst ( .DIN(_36202), .Q(_35114) );
  hi1s1 _43114_inst ( .DIN(_42388), .Q(_42819) );
  nnd2s1 _43115_inst ( .DIN1(_37673), .DIN2(_42846), .Q(_42388) );
  hi1s1 _43116_inst ( .DIN(_39312), .Q(_42846) );
  and2s1 _43117_inst ( .DIN1(_41831), .DIN2(_42953), .Q(_41939) );
  nnd2s1 _43118_inst ( .DIN1(_42190), .DIN2(_42249), .Q(_42953) );
  nnd2s1 _43119_inst ( .DIN1(_42312), .DIN2(_42954), .Q(_42249) );
  nnd2s1 _43120_inst ( .DIN1(_42955), .DIN2(______[11]), .Q(_42954) );
  nor2s1 _43121_inst ( .DIN1(______[7]), .DIN2(_39120), .Q(_42955) );
  nor2s1 _43122_inst ( .DIN1(_42649), .DIN2(_42293), .Q(_41831) );
  nnd2s1 _43123_inst ( .DIN1(_42956), .DIN2(_42929), .Q(_42649) );
  nor2s1 _43124_inst ( .DIN1(_42957), .DIN2(_42958), .Q(_42935) );
  or2s1 _43125_inst ( .DIN1(_42344), .DIN2(_42009), .Q(_42958) );
  nnd2s1 _43126_inst ( .DIN1(_41893), .DIN2(_42959), .Q(_42009) );
  nnd2s1 _43127_inst ( .DIN1(_42960), .DIN2(_42961), .Q(_42959) );
  nor2s1 _43128_inst ( .DIN1(_42687), .DIN2(_42342), .Q(_42960) );
  nnd2s1 _43129_inst ( .DIN1(_42257), .DIN2(_42292), .Q(_41893) );
  and2s1 _43130_inst ( .DIN1(_42962), .DIN2(_37467), .Q(_42257) );
  nor2s1 _43131_inst ( .DIN1(_42884), .DIN2(_36066), .Q(_42962) );
  hi1s1 _43132_inst ( .DIN(_36456), .Q(_36066) );
  nor2s1 _43133_inst ( .DIN1(_42597), .DIN2(_53425), .Q(_36456) );
  nnd2s1 _43134_inst ( .DIN1(_42631), .DIN2(_42963), .Q(_42344) );
  nnd2s1 _43135_inst ( .DIN1(_42964), .DIN2(_42857), .Q(_42963) );
  nor2s1 _43136_inst ( .DIN1(_37995), .DIN2(_35688), .Q(_42857) );
  nnd2s1 _43137_inst ( .DIN1(_42943), .DIN2(_42965), .Q(_35688) );
  nor2s1 _43138_inst ( .DIN1(_42104), .DIN2(_35930), .Q(_42964) );
  nnd2s1 _43139_inst ( .DIN1(_37328), .DIN2(_42950), .Q(_35930) );
  nnd2s1 _43140_inst ( .DIN1(_42966), .DIN2(_42967), .Q(_42104) );
  nnd2s1 _43141_inst ( .DIN1(_42908), .DIN2(_42114), .Q(_42631) );
  and2s1 _43142_inst ( .DIN1(_42968), .DIN2(_37189), .Q(_42908) );
  nor2s1 _43143_inst ( .DIN1(_39312), .DIN2(_37923), .Q(_42968) );
  nnd2s1 _43144_inst ( .DIN1(_42969), .DIN2(_42965), .Q(_39312) );
  nnd2s1 _43145_inst ( .DIN1(_42970), .DIN2(_42971), .Q(_42957) );
  hi1s1 _43146_inst ( .DIN(_42398), .Q(_42971) );
  nnd2s1 _43147_inst ( .DIN1(_42632), .DIN2(_42972), .Q(_42398) );
  nnd2s1 _43148_inst ( .DIN1(_42160), .DIN2(_42145), .Q(_42972) );
  hi1s1 _43149_inst ( .DIN(_42462), .Q(_42160) );
  nnd2s1 _43150_inst ( .DIN1(_42973), .DIN2(_42967), .Q(_42462) );
  nnd2s1 _43151_inst ( .DIN1(_42710), .DIN2(_42114), .Q(_42632) );
  nor2s1 _43152_inst ( .DIN1(_37211), .DIN2(_42293), .Q(_42710) );
  nnd2s1 _43153_inst ( .DIN1(_42974), .DIN2(_42907), .Q(_37211) );
  nor2s1 _43154_inst ( .DIN1(_42975), .DIN2(_42389), .Q(_42970) );
  nnd2s1 _43155_inst ( .DIN1(_42976), .DIN2(_42977), .Q(_42389) );
  nnd2s1 _43156_inst ( .DIN1(_41899), .DIN2(_42371), .Q(_42977) );
  hi1s1 _43157_inst ( .DIN(_42701), .Q(_41899) );
  nnd2s1 _43158_inst ( .DIN1(_42978), .DIN2(_37189), .Q(_42701) );
  nor2s1 _43159_inst ( .DIN1(_37670), .DIN2(_39040), .Q(_42978) );
  hi1s1 _43160_inst ( .DIN(_37673), .Q(_37670) );
  nor2s1 _43161_inst ( .DIN1(_42979), .DIN2(_53429), .Q(_37673) );
  nor2s1 _43162_inst ( .DIN1(_42980), .DIN2(_42981), .Q(_42976) );
  nor2s1 _43163_inst ( .DIN1(_42161), .DIN2(_42982), .Q(_42981) );
  nnd2s1 _43164_inst ( .DIN1(_42292), .DIN2(_37194), .Q(_42982) );
  hi1s1 _43165_inst ( .DIN(_36455), .Q(_37194) );
  nnd2s1 _43166_inst ( .DIN1(_42983), .DIN2(_42791), .Q(_36455) );
  hi1s1 _43167_inst ( .DIN(_42052), .Q(_42292) );
  nnd2s1 _43168_inst ( .DIN1(_28525), .DIN2(_37471), .Q(_42161) );
  hi1s1 _43169_inst ( .DIN(_37923), .Q(_37471) );
  hi1s1 _43170_inst ( .DIN(_42703), .Q(_42980) );
  nnd2s1 _43171_inst ( .DIN1(_42984), .DIN2(_36203), .Q(_42703) );
  nor2s1 _43172_inst ( .DIN1(_42985), .DIN2(_42986), .Q(_36203) );
  nnd2s1 _43173_inst ( .DIN1(_53425), .DIN2(_42929), .Q(_42985) );
  nor2s1 _43174_inst ( .DIN1(_42407), .DIN2(_42640), .Q(_42984) );
  nor2s1 _43175_inst ( .DIN1(_41903), .DIN2(_42023), .Q(_42975) );
  nnd2s1 _43176_inst ( .DIN1(_42987), .DIN2(_37197), .Q(_42023) );
  hi1s1 _43177_inst ( .DIN(_36201), .Q(_37197) );
  nnd2s1 _43178_inst ( .DIN1(_42929), .DIN2(_42950), .Q(_36201) );
  xnr2s1 _43179_inst ( .DIN1(_29049), .DIN2(_42621), .Q(_42987) );
  nor2s1 _43180_inst ( .DIN1(_35534), .DIN2(_37923), .Q(_42621) );
  nnd2s1 _43181_inst ( .DIN1(_42988), .DIN2(_53418), .Q(_37923) );
  nor2s1 _43182_inst ( .DIN1(_53419), .DIN2(_53429), .Q(_42988) );
  xor2s1 _43183_inst ( .DIN1(_42989), .DIN2(_28088), .Q(_42933) );
  nnd2s1 _43184_inst ( .DIN1(_42589), .DIN2(_42676), .Q(_42989) );
  nnd2s1 _43185_inst ( .DIN1(_42427), .DIN2(_42312), .Q(_42676) );
  hi1s1 _43186_inst ( .DIN(_42331), .Q(_42427) );
  nnd2s1 _43187_inst ( .DIN1(_42990), .DIN2(_28596), .Q(_42331) );
  nor2s1 _43188_inst ( .DIN1(_37445), .DIN2(_37318), .Q(_42990) );
  nnd2s1 _43189_inst ( .DIN1(_42302), .DIN2(_42991), .Q(_42589) );
  hi1s1 _43190_inst ( .DIN(_42379), .Q(_42991) );
  nnd2s1 _43191_inst ( .DIN1(_42992), .DIN2(_42596), .Q(_42379) );
  hi1s1 _43192_inst ( .DIN(_42993), .Q(_42596) );
  nor2s1 _43193_inst ( .DIN1(_42842), .DIN2(_42994), .Q(_42992) );
  hi1s1 _43194_inst ( .DIN(_41944), .Q(_42302) );
  nnd2s1 _43195_inst ( .DIN1(_42995), .DIN2(_42240), .Q(_42931) );
  and2s1 _43196_inst ( .DIN1(_42996), .DIN2(_42997), .Q(_42240) );
  nor2s1 _43197_inst ( .DIN1(_41934), .DIN2(_42998), .Q(_42997) );
  nnd2s1 _43198_inst ( .DIN1(_42011), .DIN2(_42174), .Q(_42998) );
  nnd2s1 _43199_inst ( .DIN1(_42504), .DIN2(_42258), .Q(_42174) );
  nor2s1 _43200_inst ( .DIN1(_42687), .DIN2(_42884), .Q(_42504) );
  nnd2s1 _43201_inst ( .DIN1(_42999), .DIN2(_42944), .Q(_42884) );
  nnd2s1 _43202_inst ( .DIN1(_35272), .DIN2(_36694), .Q(_42687) );
  hi1s1 _43203_inst ( .DIN(_36065), .Q(_35272) );
  nnd2s1 _43204_inst ( .DIN1(_42956), .DIN2(_42907), .Q(_36065) );
  nnd2s1 _43205_inst ( .DIN1(_42461), .DIN2(_42371), .Q(_42011) );
  hi1s1 _43206_inst ( .DIN(_42095), .Q(_42461) );
  nnd2s1 _43207_inst ( .DIN1(_43000), .DIN2(_43001), .Q(_42095) );
  nor2s1 _43208_inst ( .DIN1(_43002), .DIN2(_42613), .Q(_43001) );
  nor2s1 _43209_inst ( .DIN1(_42661), .DIN2(_42093), .Q(_41934) );
  nnd2s1 _43210_inst ( .DIN1(_42602), .DIN2(_42600), .Q(_42093) );
  nor2s1 _43211_inst ( .DIN1(_43003), .DIN2(_42817), .Q(_42602) );
  or2s1 _43212_inst ( .DIN1(_43002), .DIN2(_42613), .Q(_43003) );
  nor2s1 _43213_inst ( .DIN1(_41815), .DIN2(_42073), .Q(_42996) );
  nnd2s1 _43214_inst ( .DIN1(_43004), .DIN2(_43005), .Q(_42073) );
  nnd2s1 _43215_inst ( .DIN1(_42495), .DIN2(_41900), .Q(_43005) );
  nnd2s1 _43216_inst ( .DIN1(_42342), .DIN2(_42387), .Q(_41900) );
  nnd2s1 _43217_inst ( .DIN1(_42312), .DIN2(_43006), .Q(_42342) );
  nnd2s1 _43218_inst ( .DIN1(_42952), .DIN2(_43007), .Q(_43006) );
  nor2s1 _43219_inst ( .DIN1(______[7]), .DIN2(______[29]), .Q(_42952) );
  nor2s1 _43220_inst ( .DIN1(_42330), .DIN2(_37323), .Q(_42495) );
  nnd2s1 _43221_inst ( .DIN1(_42974), .DIN2(_37328), .Q(_37323) );
  nnd2s1 _43222_inst ( .DIN1(_28599), .DIN2(_36694), .Q(_42330) );
  nor2s1 _43223_inst ( .DIN1(_43008), .DIN2(_42207), .Q(_28599) );
  nnd2s1 _43224_inst ( .DIN1(_26538), .DIN2(_26275), .Q(_43008) );
  nnd2s1 _43225_inst ( .DIN1(_42371), .DIN2(_42402), .Q(_43004) );
  hi1s1 _43226_inst ( .DIN(_42489), .Q(_42402) );
  nnd2s1 _43227_inst ( .DIN1(_43009), .DIN2(_42914), .Q(_42489) );
  nor2s1 _43228_inst ( .DIN1(_43010), .DIN2(_42613), .Q(_42914) );
  nor2s1 _43229_inst ( .DIN1(_42817), .DIN2(_42994), .Q(_43009) );
  nnd2s1 _43230_inst ( .DIN1(_43011), .DIN2(_53425), .Q(_42817) );
  nor2s1 _43231_inst ( .DIN1(_26334), .DIN2(_42979), .Q(_43011) );
  hi1s1 _43232_inst ( .DIN(_42387), .Q(_42371) );
  nnd2s1 _43233_inst ( .DIN1(_43012), .DIN2(_43013), .Q(_42387) );
  nor2s1 _43234_inst ( .DIN1(_42533), .DIN2(_42423), .Q(_41815) );
  nnd2s1 _43235_inst ( .DIN1(_43000), .DIN2(_43014), .Q(_42423) );
  nor2s1 _43236_inst ( .DIN1(_43010), .DIN2(_42986), .Q(_43014) );
  nor2s1 _43237_inst ( .DIN1(_42598), .DIN2(_42993), .Q(_43000) );
  nnd2s1 _43238_inst ( .DIN1(_43015), .DIN2(_42944), .Q(_42598) );
  nor2s1 _43239_inst ( .DIN1(_43016), .DIN2(_42195), .Q(_42995) );
  nnd2s1 _43240_inst ( .DIN1(_42060), .DIN2(_43017), .Q(_42195) );
  nnd2s1 _43241_inst ( .DIN1(_41895), .DIN2(_42258), .Q(_43017) );
  hi1s1 _43242_inst ( .DIN(_42509), .Q(_41895) );
  nnd2s1 _43243_inst ( .DIN1(_43018), .DIN2(_28596), .Q(_42509) );
  nor2s1 _43244_inst ( .DIN1(_37810), .DIN2(_35103), .Q(_43018) );
  nnd2s1 _43245_inst ( .DIN1(_43019), .DIN2(_53425), .Q(_35103) );
  nor2s1 _43246_inst ( .DIN1(_43002), .DIN2(_37329), .Q(_43019) );
  nnd2s1 _43247_inst ( .DIN1(_43020), .DIN2(_43021), .Q(_42060) );
  hi1s1 _43248_inst ( .DIN(_42918), .Q(_43021) );
  nnd2s1 _43249_inst ( .DIN1(_42961), .DIN2(_37334), .Q(_42918) );
  hi1s1 _43250_inst ( .DIN(_37318), .Q(_37334) );
  hi1s1 _43251_inst ( .DIN(_39311), .Q(_42961) );
  nnd2s1 _43252_inst ( .DIN1(_43022), .DIN2(_42943), .Q(_39311) );
  nor2s1 _43253_inst ( .DIN1(_37445), .DIN2(_42407), .Q(_43020) );
  nnd2s1 _43254_inst ( .DIN1(_43012), .DIN2(_42967), .Q(_42407) );
  hi1s1 _43255_inst ( .DIN(_41920), .Q(_43016) );
  nor2s1 _43256_inst ( .DIN1(_43023), .DIN2(_41840), .Q(_41920) );
  nnd2s1 _43257_inst ( .DIN1(_43024), .DIN2(_43025), .Q(_41840) );
  nor2s1 _43258_inst ( .DIN1(_42063), .DIN2(_43026), .Q(_43025) );
  hi1s1 _43259_inst ( .DIN(_42662), .Q(_43026) );
  nnd2s1 _43260_inst ( .DIN1(_43027), .DIN2(_42692), .Q(_42662) );
  hi1s1 _43261_inst ( .DIN(_42779), .Q(_42692) );
  xor2s1 _43262_inst ( .DIN1(_43028), .DIN2(_30367), .Q(_43027) );
  hi1s1 _43263_inst ( .DIN(_30349), .Q(_30367) );
  nnd2s1 _43264_inst ( .DIN1(_27840), .DIN2(_43029), .Q(_30349) );
  hi1s1 _43265_inst ( .DIN(_32362), .Q(_27840) );
  nnd2s1 _43266_inst ( .DIN1(_43030), .DIN2(_33865), .Q(_32362) );
  nnd2s1 _43267_inst ( .DIN1(_36199), .DIN2(_42025), .Q(_43028) );
  hi1s1 _43268_inst ( .DIN(_42533), .Q(_42025) );
  nnd2s1 _43269_inst ( .DIN1(_43031), .DIN2(_43013), .Q(_42533) );
  hi1s1 _43270_inst ( .DIN(_35104), .Q(_36199) );
  nnd2s1 _43271_inst ( .DIN1(_42956), .DIN2(_37328), .Q(_35104) );
  nor2s1 _43272_inst ( .DIN1(_42986), .DIN2(_53425), .Q(_42956) );
  and2s1 _43273_inst ( .DIN1(_42725), .DIN2(_42258), .Q(_42063) );
  xor2s1 _43274_inst ( .DIN1(_43032), .DIN2(_27329), .Q(_42258) );
  nnd2s1 _43275_inst ( .DIN1(_42052), .DIN2(_42083), .Q(_43032) );
  nnd2s1 _43276_inst ( .DIN1(_42966), .DIN2(_43013), .Q(_42052) );
  nor2s1 _43277_inst ( .DIN1(______[11]), .DIN2(_39120), .Q(_42966) );
  hi1s1 _43278_inst ( .DIN(_42537), .Q(_42725) );
  nnd2s1 _43279_inst ( .DIN1(_42568), .DIN2(_42600), .Q(_42537) );
  and2s1 _43280_inst ( .DIN1(_43033), .DIN2(_43034), .Q(_42568) );
  nor2s1 _43281_inst ( .DIN1(_43035), .DIN2(_42993), .Q(_43033) );
  nor2s1 _43282_inst ( .DIN1(_42261), .DIN2(_43036), .Q(_43024) );
  nor2s1 _43283_inst ( .DIN1(_42650), .DIN2(_42219), .Q(_43036) );
  nnd2s1 _43284_inst ( .DIN1(_43037), .DIN2(_42600), .Q(_42219) );
  hi1s1 _43285_inst ( .DIN(_42853), .Q(_42600) );
  nnd2s1 _43286_inst ( .DIN1(_42969), .DIN2(_42944), .Q(_42853) );
  nor2s1 _43287_inst ( .DIN1(_53417), .DIN2(_53420), .Q(_42944) );
  nor2s1 _43288_inst ( .DIN1(_42842), .DIN2(_42993), .Q(_43037) );
  or2s1 _43289_inst ( .DIN1(_43035), .DIN2(_37329), .Q(_42842) );
  hi1s1 _43290_inst ( .DIN(_42541), .Q(_42650) );
  nnd2s1 _43291_inst ( .DIN1(_41944), .DIN2(_42225), .Q(_42541) );
  nnd2s1 _43292_inst ( .DIN1(_42312), .DIN2(_43038), .Q(_42225) );
  nnd2s1 _43293_inst ( .DIN1(_43039), .DIN2(______[11]), .Q(_43038) );
  nor2s1 _43294_inst ( .DIN1(______[29]), .DIN2(_39015), .Q(_43039) );
  nnd2s1 _43295_inst ( .DIN1(_43031), .DIN2(_42967), .Q(_41944) );
  nor2s1 _43296_inst ( .DIN1(_39015), .DIN2(_41903), .Q(_42967) );
  nor2s1 _43297_inst ( .DIN1(______[29]), .DIN2(_43007), .Q(_43031) );
  nor2s1 _43298_inst ( .DIN1(_41903), .DIN2(_42674), .Q(_42261) );
  nnd2s1 _43299_inst ( .DIN1(_42599), .DIN2(_42913), .Q(_42674) );
  hi1s1 _43300_inst ( .DIN(_42994), .Q(_42913) );
  nnd2s1 _43301_inst ( .DIN1(_43040), .DIN2(_42943), .Q(_42994) );
  nor2s1 _43302_inst ( .DIN1(_53421), .DIN2(_53422), .Q(_42943) );
  nor2s1 _43303_inst ( .DIN1(_42672), .DIN2(_42979), .Q(_42599) );
  nnd2s1 _43304_inst ( .DIN1(_26539), .DIN2(_26279), .Q(_42979) );
  nnd2s1 _43305_inst ( .DIN1(_43041), .DIN2(_43042), .Q(_42672) );
  nor2s1 _43306_inst ( .DIN1(_53425), .DIN2(_26334), .Q(_43042) );
  nor2s1 _43307_inst ( .DIN1(_37329), .DIN2(_43043), .Q(_43041) );
  or2s1 _43308_inst ( .DIN1(_42002), .DIN2(_41839), .Q(_43023) );
  nnd2s1 _43309_inst ( .DIN1(_43044), .DIN2(_43045), .Q(_41839) );
  nnd2s1 _43310_inst ( .DIN1(_42145), .DIN2(_42012), .Q(_43045) );
  hi1s1 _43311_inst ( .DIN(_42661), .Q(_42012) );
  nnd2s1 _43312_inst ( .DIN1(_42312), .DIN2(_43046), .Q(_42661) );
  nnd2s1 _43313_inst ( .DIN1(_43047), .DIN2(______[11]), .Q(_43046) );
  nor2s1 _43314_inst ( .DIN1(_39015), .DIN2(_39120), .Q(_43047) );
  and2s1 _43315_inst ( .DIN1(_42910), .DIN2(_28526), .Q(_42145) );
  hi1s1 _43316_inst ( .DIN(_39040), .Q(_28526) );
  nnd2s1 _43317_inst ( .DIN1(_43048), .DIN2(_53417), .Q(_39040) );
  nor2s1 _43318_inst ( .DIN1(_53422), .DIN2(_42207), .Q(_43048) );
  nor2s1 _43319_inst ( .DIN1(_36202), .DIN2(_37995), .Q(_42910) );
  nnd2s1 _43320_inst ( .DIN1(_42791), .DIN2(_42974), .Q(_36202) );
  and2s1 _43321_inst ( .DIN1(_43034), .DIN2(_53425), .Q(_42974) );
  nor2s1 _43322_inst ( .DIN1(_53416), .DIN2(_53460), .Q(_43034) );
  nnd2s1 _43323_inst ( .DIN1(_41896), .DIN2(_42146), .Q(_43044) );
  nnd2s1 _43324_inst ( .DIN1(_42536), .DIN2(_43049), .Q(_42146) );
  or2s1 _43325_inst ( .DIN1(_42293), .DIN2(_37199), .Q(_43049) );
  nnd2s1 _43326_inst ( .DIN1(_42950), .DIN2(_42907), .Q(_37199) );
  and2s1 _43327_inst ( .DIN1(_43050), .DIN2(_26585), .Q(_42950) );
  nor2s1 _43328_inst ( .DIN1(_53416), .DIN2(_53425), .Q(_43050) );
  nnd2s1 _43329_inst ( .DIN1(_28525), .DIN2(_36695), .Q(_42293) );
  hi1s1 _43330_inst ( .DIN(_37995), .Q(_36695) );
  hi1s1 _43331_inst ( .DIN(_39314), .Q(_28525) );
  nnd2s1 _43332_inst ( .DIN1(_43022), .DIN2(_42969), .Q(_39314) );
  nor2s1 _43333_inst ( .DIN1(_53417), .DIN2(_26298), .Q(_43022) );
  nnd2s1 _43334_inst ( .DIN1(_43051), .DIN2(_37189), .Q(_42536) );
  hi1s1 _43335_inst ( .DIN(_42255), .Q(_37189) );
  nnd2s1 _43336_inst ( .DIN1(_42790), .DIN2(_37328), .Q(_42255) );
  nor2s1 _43337_inst ( .DIN1(_37329), .DIN2(_26212), .Q(_42790) );
  nor2s1 _43338_inst ( .DIN1(_37995), .DIN2(_35534), .Q(_43051) );
  nnd2s1 _43339_inst ( .DIN1(_43052), .DIN2(_53417), .Q(_35534) );
  nor2s1 _43340_inst ( .DIN1(_42207), .DIN2(_26275), .Q(_43052) );
  nnd2s1 _43341_inst ( .DIN1(_43053), .DIN2(_53419), .Q(_37995) );
  nor2s1 _43342_inst ( .DIN1(_53418), .DIN2(_53429), .Q(_43053) );
  hi1s1 _43343_inst ( .DIN(_42090), .Q(_42002) );
  nnd2s1 _43344_inst ( .DIN1(_42732), .DIN2(_42114), .Q(_42090) );
  hi1s1 _43345_inst ( .DIN(_42190), .Q(_42114) );
  nnd2s1 _43346_inst ( .DIN1(_42973), .DIN2(_43013), .Q(_42190) );
  nor2s1 _43347_inst ( .DIN1(______[7]), .DIN2(_41903), .Q(_43013) );
  nor2s1 _43348_inst ( .DIN1(_39120), .DIN2(_43007), .Q(_42973) );
  hi1s1 _43349_inst ( .DIN(______[11]), .Q(_43007) );
  hi1s1 _43350_inst ( .DIN(______[29]), .Q(_39120) );
  nor2s1 _43351_inst ( .DIN1(_42986), .DIN2(_42612), .Q(_42732) );
  nnd2s1 _43352_inst ( .DIN1(_43054), .DIN2(_42567), .Q(_42612) );
  nor2s1 _43353_inst ( .DIN1(_43002), .DIN2(_42993), .Q(_43054) );
  nnd2s1 _43354_inst ( .DIN1(_43055), .DIN2(_43056), .Q(_42782) );
  nnd2s1 _43355_inst ( .DIN1(_42021), .DIN2(_43057), .Q(_43056) );
  nnd2s1 _43356_inst ( .DIN1(_43058), .DIN2(_43059), .Q(_43057) );
  nor2s1 _43357_inst ( .DIN1(_43060), .DIN2(_43061), .Q(_43059) );
  nor2s1 _43358_inst ( .DIN1(_35270), .DIN2(_43062), .Q(_43061) );
  nnd2s1 _43359_inst ( .DIN1(_42789), .DIN2(_26410), .Q(_43062) );
  hi1s1 _43360_inst ( .DIN(_42545), .Q(_42789) );
  nnd2s1 _43361_inst ( .DIN1(_28597), .DIN2(_36694), .Q(_42545) );
  hi1s1 _43362_inst ( .DIN(_35686), .Q(_28597) );
  nnd2s1 _43363_inst ( .DIN1(_43063), .DIN2(_53422), .Q(_35686) );
  nor2s1 _43364_inst ( .DIN1(_53417), .DIN2(_42207), .Q(_43063) );
  nnd2s1 _43365_inst ( .DIN1(_53420), .DIN2(_53421), .Q(_42207) );
  hi1s1 _43366_inst ( .DIN(_35113), .Q(_35270) );
  nor2s1 _43367_inst ( .DIN1(_43064), .DIN2(_37329), .Q(_35113) );
  nnd2s1 _43368_inst ( .DIN1(_53416), .DIN2(_53460), .Q(_37329) );
  nnd2s1 _43369_inst ( .DIN1(_26212), .DIN2(_42907), .Q(_43064) );
  hi1s1 _43370_inst ( .DIN(_43002), .Q(_42907) );
  nnd2s1 _43371_inst ( .DIN1(_53424), .DIN2(_26722), .Q(_43002) );
  hi1s1 _43372_inst ( .DIN(_42888), .Q(_43060) );
  nnd2s1 _43373_inst ( .DIN1(_42767), .DIN2(_36060), .Q(_42888) );
  xnr2s1 _43374_inst ( .DIN1(_37332), .DIN2(_35821), .Q(_36060) );
  hi1s1 _43375_inst ( .DIN(_42640), .Q(_42767) );
  nnd2s1 _43376_inst ( .DIN1(_37467), .DIN2(_28596), .Q(_42640) );
  hi1s1 _43377_inst ( .DIN(_39313), .Q(_28596) );
  nnd2s1 _43378_inst ( .DIN1(_43015), .DIN2(_42965), .Q(_39313) );
  nor2s1 _43379_inst ( .DIN1(_53422), .DIN2(_26626), .Q(_43015) );
  hi1s1 _43380_inst ( .DIN(_42338), .Q(_37467) );
  nnd2s1 _43381_inst ( .DIN1(_43065), .DIN2(_53418), .Q(_42338) );
  nor2s1 _43382_inst ( .DIN1(_53429), .DIN2(_26279), .Q(_43065) );
  nor2s1 _43383_inst ( .DIN1(_43066), .DIN2(_43067), .Q(_43058) );
  nor2s1 _43384_inst ( .DIN1(_42779), .DIN2(_37318), .Q(_43067) );
  nnd2s1 _43385_inst ( .DIN1(_42906), .DIN2(_37328), .Q(_37318) );
  hi1s1 _43386_inst ( .DIN(_43010), .Q(_37328) );
  nnd2s1 _43387_inst ( .DIN1(_53423), .DIN2(_26285), .Q(_43010) );
  nnd2s1 _43388_inst ( .DIN1(_38018), .DIN2(_36694), .Q(_42779) );
  hi1s1 _43389_inst ( .DIN(_37810), .Q(_36694) );
  nnd2s1 _43390_inst ( .DIN1(_43068), .DIN2(_53418), .Q(_37810) );
  nor2s1 _43391_inst ( .DIN1(_53419), .DIN2(_26334), .Q(_43068) );
  nor2s1 _43392_inst ( .DIN1(_35269), .DIN2(_42228), .Q(_43066) );
  nnd2s1 _43393_inst ( .DIN1(_42983), .DIN2(_42929), .Q(_35269) );
  hi1s1 _43394_inst ( .DIN(_43035), .Q(_42929) );
  nnd2s1 _43395_inst ( .DIN1(_26722), .DIN2(_26285), .Q(_43035) );
  nor2s1 _43396_inst ( .DIN1(_26212), .DIN2(_42613), .Q(_42983) );
  hi1s1 _43397_inst ( .DIN(_42153), .Q(_42021) );
  nnd2s1 _43398_inst ( .DIN1(_42312), .DIN2(_43069), .Q(_42153) );
  nnd2s1 _43399_inst ( .DIN1(_43012), .DIN2(______[7]), .Q(_43069) );
  nor2s1 _43400_inst ( .DIN1(______[29]), .DIN2(______[11]), .Q(_43012) );
  nnd2s1 _43401_inst ( .DIN1(_41896), .DIN2(_43070), .Q(_43055) );
  nnd2s1 _43402_inst ( .DIN1(_42084), .DIN2(_43071), .Q(_43070) );
  nnd2s1 _43403_inst ( .DIN1(_43072), .DIN2(_37332), .Q(_43071) );
  and2s1 _43404_inst ( .DIN1(_42791), .DIN2(_42906), .Q(_37332) );
  nor2s1 _43405_inst ( .DIN1(_42613), .DIN2(_53425), .Q(_42906) );
  nnd2s1 _43406_inst ( .DIN1(_53416), .DIN2(_26585), .Q(_42613) );
  hi1s1 _43407_inst ( .DIN(_43043), .Q(_42791) );
  hi1s1 _43408_inst ( .DIN(_42228), .Q(_43072) );
  nnd2s1 _43409_inst ( .DIN1(_38018), .DIN2(_37468), .Q(_42228) );
  hi1s1 _43410_inst ( .DIN(_37445), .Q(_37468) );
  nnd2s1 _43411_inst ( .DIN1(_43073), .DIN2(_53419), .Q(_37445) );
  nor2s1 _43412_inst ( .DIN1(_53418), .DIN2(_26334), .Q(_43073) );
  hi1s1 _43413_inst ( .DIN(_35533), .Q(_38018) );
  nnd2s1 _43414_inst ( .DIN1(_42999), .DIN2(_42965), .Q(_35533) );
  nor2s1 _43415_inst ( .DIN1(_26538), .DIN2(_53420), .Q(_42965) );
  nor2s1 _43416_inst ( .DIN1(_26626), .DIN2(_26275), .Q(_42999) );
  nnd2s1 _43417_inst ( .DIN1(_43074), .DIN2(_42567), .Q(_42084) );
  hi1s1 _43418_inst ( .DIN(_42870), .Q(_42567) );
  nnd2s1 _43419_inst ( .DIN1(_43040), .DIN2(_42969), .Q(_42870) );
  nor2s1 _43420_inst ( .DIN1(_26275), .DIN2(_53421), .Q(_42969) );
  nor2s1 _43421_inst ( .DIN1(_26298), .DIN2(_26538), .Q(_43040) );
  nor2s1 _43422_inst ( .DIN1(_42597), .DIN2(_42993), .Q(_43074) );
  nnd2s1 _43423_inst ( .DIN1(_43075), .DIN2(_43076), .Q(_42993) );
  nor2s1 _43424_inst ( .DIN1(_26334), .DIN2(_26279), .Q(_43076) );
  nor2s1 _43425_inst ( .DIN1(_26539), .DIN2(_26212), .Q(_43075) );
  or2s1 _43426_inst ( .DIN1(_43043), .DIN2(_42986), .Q(_42597) );
  nnd2s1 _43427_inst ( .DIN1(_53460), .DIN2(_26699), .Q(_42986) );
  nnd2s1 _43428_inst ( .DIN1(_53424), .DIN2(_53423), .Q(_43043) );
  hi1s1 _43429_inst ( .DIN(_42083), .Q(_41896) );
  nnd2s1 _43430_inst ( .DIN1(_42312), .DIN2(_43077), .Q(_42083) );
  nnd2s1 _43431_inst ( .DIN1(_43078), .DIN2(______[29]), .Q(_43077) );
  nor2s1 _43432_inst ( .DIN1(______[7]), .DIN2(______[11]), .Q(_43078) );
  nnd2s1 _43433_inst ( .DIN1(_43079), .DIN2(_43080), .Q(
        ____0____________9_____) );
  nnd2s1 _43434_inst ( .DIN1(_43081), .DIN2(_43082), .Q(_43080) );
  nnd2s1 _43435_inst ( .DIN1(_53444), .DIN2(_41806), .Q(_43081) );
  nnd2s1 _43436_inst ( .DIN1(_43083), .DIN2(_41807), .Q(_43079) );
  nor2s1 _43437_inst ( .DIN1(_43084), .DIN2(_43085), .Q(_43083) );
  nnd2s1 _43438_inst ( .DIN1(_43086), .DIN2(_43087), .Q(_43085) );
  nor2s1 _43439_inst ( .DIN1(_43088), .DIN2(_43089), .Q(_43087) );
  nnd2s1 _43440_inst ( .DIN1(_43090), .DIN2(_43091), .Q(_43089) );
  hi1s1 _43441_inst ( .DIN(_43092), .Q(_43090) );
  nnd2s1 _43442_inst ( .DIN1(_43093), .DIN2(_43094), .Q(_43088) );
  or2s1 _43443_inst ( .DIN1(_43095), .DIN2(_43096), .Q(_43094) );
  nor2s1 _43444_inst ( .DIN1(_43097), .DIN2(_43098), .Q(_43086) );
  nnd2s1 _43445_inst ( .DIN1(_43099), .DIN2(_43100), .Q(_43098) );
  nnd2s1 _43446_inst ( .DIN1(_43101), .DIN2(_43102), .Q(_43084) );
  nor2s1 _43447_inst ( .DIN1(_43103), .DIN2(_43104), .Q(_43102) );
  nnd2s1 _43448_inst ( .DIN1(_43105), .DIN2(_43106), .Q(_43104) );
  hi1s1 _43449_inst ( .DIN(_43107), .Q(_43106) );
  nnd2s1 _43450_inst ( .DIN1(_43108), .DIN2(_43109), .Q(_43105) );
  nnd2s1 _43451_inst ( .DIN1(_43110), .DIN2(_43111), .Q(_43109) );
  or2s1 _43452_inst ( .DIN1(_43112), .DIN2(_43113), .Q(_43103) );
  nor2s1 _43453_inst ( .DIN1(_43114), .DIN2(_43115), .Q(_43101) );
  nnd2s1 _43454_inst ( .DIN1(_43116), .DIN2(_43117), .Q(_43115) );
  nnd2s1 _43455_inst ( .DIN1(_43118), .DIN2(_43119), .Q(_43117) );
  or2s1 _43456_inst ( .DIN1(_43120), .DIN2(_43121), .Q(_43116) );
  nor2s1 _43457_inst ( .DIN1(_43122), .DIN2(_43123), .Q(_43114) );
  nnd2s1 _43458_inst ( .DIN1(_43124), .DIN2(_43125), .Q(
        ____0____________8_____) );
  nnd2s1 _43459_inst ( .DIN1(_43126), .DIN2(_41806), .Q(_43125) );
  xor2s1 _43460_inst ( .DIN1(_26215), .DIN2(_43127), .Q(_43126) );
  nnd2s1 _43461_inst ( .DIN1(_41807), .DIN2(_43128), .Q(_43124) );
  nnd2s1 _43462_inst ( .DIN1(_43129), .DIN2(_43130), .Q(_43128) );
  nor2s1 _43463_inst ( .DIN1(_43131), .DIN2(_43132), .Q(_43130) );
  nnd2s1 _43464_inst ( .DIN1(_43133), .DIN2(_43134), .Q(_43132) );
  nor2s1 _43465_inst ( .DIN1(_43135), .DIN2(_43136), .Q(_43134) );
  nor2s1 _43466_inst ( .DIN1(_43137), .DIN2(_43138), .Q(_43136) );
  nor2s1 _43467_inst ( .DIN1(_43139), .DIN2(_43140), .Q(_43135) );
  nor2s1 _43468_inst ( .DIN1(_43141), .DIN2(_43142), .Q(_43133) );
  nnd2s1 _43469_inst ( .DIN1(_43143), .DIN2(_43144), .Q(_43131) );
  nor2s1 _43470_inst ( .DIN1(_43145), .DIN2(_43146), .Q(_43144) );
  or2s1 _43471_inst ( .DIN1(_43147), .DIN2(_43148), .Q(_43146) );
  nor2s1 _43472_inst ( .DIN1(_43149), .DIN2(_43150), .Q(_43143) );
  nor2s1 _43473_inst ( .DIN1(_43151), .DIN2(_43152), .Q(_43150) );
  nor2s1 _43474_inst ( .DIN1(_43096), .DIN2(_43153), .Q(_43149) );
  nor2s1 _43475_inst ( .DIN1(_43154), .DIN2(_43155), .Q(_43129) );
  nnd2s1 _43476_inst ( .DIN1(_43156), .DIN2(_43157), .Q(_43155) );
  nor2s1 _43477_inst ( .DIN1(_43158), .DIN2(_43159), .Q(_43157) );
  nor2s1 _43478_inst ( .DIN1(_43160), .DIN2(_43161), .Q(_43156) );
  nnd2s1 _43479_inst ( .DIN1(_43162), .DIN2(_43163), .Q(_43154) );
  nor2s1 _43480_inst ( .DIN1(_43164), .DIN2(_43165), .Q(_43163) );
  nor2s1 _43481_inst ( .DIN1(_43166), .DIN2(_43167), .Q(_43164) );
  nor2s1 _43482_inst ( .DIN1(_43168), .DIN2(_43169), .Q(_43162) );
  nnd2s1 _43483_inst ( .DIN1(_43170), .DIN2(_43171), .Q(
        ____0____________7_____) );
  nor2s1 _43484_inst ( .DIN1(_43172), .DIN2(_43173), .Q(_43170) );
  nor2s1 _43485_inst ( .DIN1(_43174), .DIN2(_43175), .Q(_43173) );
  nnd2s1 _43486_inst ( .DIN1(_43176), .DIN2(_43177), .Q(_43175) );
  nor2s1 _43487_inst ( .DIN1(_43178), .DIN2(_43179), .Q(_43177) );
  nnd2s1 _43488_inst ( .DIN1(_43180), .DIN2(_43100), .Q(_43179) );
  hi1s1 _43489_inst ( .DIN(_43181), .Q(_43100) );
  nor2s1 _43490_inst ( .DIN1(_43182), .DIN2(_43183), .Q(_43180) );
  nnd2s1 _43491_inst ( .DIN1(_43184), .DIN2(_43185), .Q(_43178) );
  nnd2s1 _43492_inst ( .DIN1(_43186), .DIN2(_43187), .Q(_43185) );
  nnd2s1 _43493_inst ( .DIN1(_43188), .DIN2(_43189), .Q(_43187) );
  nor2s1 _43494_inst ( .DIN1(_43190), .DIN2(_43191), .Q(_43184) );
  nor2s1 _43495_inst ( .DIN1(_43192), .DIN2(_43193), .Q(_43176) );
  nnd2s1 _43496_inst ( .DIN1(_43194), .DIN2(_43195), .Q(_43193) );
  nor2s1 _43497_inst ( .DIN1(_43196), .DIN2(_43197), .Q(_43194) );
  nnd2s1 _43498_inst ( .DIN1(_43198), .DIN2(_43199), .Q(_43192) );
  hi1s1 _43499_inst ( .DIN(_43200), .Q(_43199) );
  nor2s1 _43500_inst ( .DIN1(_43201), .DIN2(_43202), .Q(_43198) );
  nor2s1 _43501_inst ( .DIN1(_43203), .DIN2(_43204), .Q(_43172) );
  nor2s1 _43502_inst ( .DIN1(_43205), .DIN2(_28646), .Q(_43204) );
  xor2s1 _43503_inst ( .DIN1(_26215), .DIN2(_53448), .Q(_43205) );
  nnd2s1 _43504_inst ( .DIN1(_43206), .DIN2(_43171), .Q(
        ____0____________6_____) );
  nor2s1 _43505_inst ( .DIN1(_43207), .DIN2(_43208), .Q(_43206) );
  nor2s1 _43506_inst ( .DIN1(_43174), .DIN2(_43209), .Q(_43208) );
  nnd2s1 _43507_inst ( .DIN1(_43210), .DIN2(_43211), .Q(_43209) );
  nor2s1 _43508_inst ( .DIN1(_43212), .DIN2(_43213), .Q(_43211) );
  nnd2s1 _43509_inst ( .DIN1(_43214), .DIN2(_43215), .Q(_43213) );
  nor2s1 _43510_inst ( .DIN1(_43216), .DIN2(_43217), .Q(_43215) );
  nor2s1 _43511_inst ( .DIN1(_43137), .DIN2(_43218), .Q(_43216) );
  nor2s1 _43512_inst ( .DIN1(_43219), .DIN2(_43220), .Q(_43214) );
  nnd2s1 _43513_inst ( .DIN1(_43221), .DIN2(_43222), .Q(_43212) );
  nor2s1 _43514_inst ( .DIN1(_43223), .DIN2(_43224), .Q(_43222) );
  nor2s1 _43515_inst ( .DIN1(_43225), .DIN2(_43226), .Q(_43224) );
  nor2s1 _43516_inst ( .DIN1(_43227), .DIN2(_43228), .Q(_43225) );
  nnd2s1 _43517_inst ( .DIN1(_43229), .DIN2(_43230), .Q(_43228) );
  nor2s1 _43518_inst ( .DIN1(_43231), .DIN2(_43232), .Q(_43221) );
  nor2s1 _43519_inst ( .DIN1(_43233), .DIN2(_43234), .Q(_43232) );
  nor2s1 _43520_inst ( .DIN1(_43235), .DIN2(_43236), .Q(_43210) );
  nnd2s1 _43521_inst ( .DIN1(_43237), .DIN2(_43238), .Q(_43236) );
  nor2s1 _43522_inst ( .DIN1(_43239), .DIN2(_43240), .Q(_43238) );
  nor2s1 _43523_inst ( .DIN1(_43241), .DIN2(_43242), .Q(_43237) );
  nnd2s1 _43524_inst ( .DIN1(_43243), .DIN2(_43244), .Q(_43235) );
  nor2s1 _43525_inst ( .DIN1(_43245), .DIN2(_43092), .Q(_43244) );
  nnd2s1 _43526_inst ( .DIN1(_43246), .DIN2(_43247), .Q(_43092) );
  nor2s1 _43527_inst ( .DIN1(_43248), .DIN2(_43249), .Q(_43247) );
  nor2s1 _43528_inst ( .DIN1(_43250), .DIN2(_43251), .Q(_43246) );
  nor2s1 _43529_inst ( .DIN1(_43252), .DIN2(_43253), .Q(_43250) );
  nor2s1 _43530_inst ( .DIN1(_43254), .DIN2(_43255), .Q(_43243) );
  nor2s1 _43531_inst ( .DIN1(_53449), .DIN2(_43203), .Q(_43207) );
  nnd2s1 _43532_inst ( .DIN1(_43256), .DIN2(_43257), .Q(
        ____0____________5_____) );
  nnd2s1 _43533_inst ( .DIN1(_43258), .DIN2(______[14]), .Q(_43257) );
  nor2s1 _43534_inst ( .DIN1(_43259), .DIN2(_43260), .Q(_43258) );
  xor2s1 _43535_inst ( .DIN1(_26262), .DIN2(_53429), .Q(_43260) );
  nnd2s1 _43536_inst ( .DIN1(_41807), .DIN2(_43261), .Q(_43256) );
  nnd2s1 _43537_inst ( .DIN1(_43262), .DIN2(_43263), .Q(_43261) );
  nor2s1 _43538_inst ( .DIN1(_43264), .DIN2(_43265), .Q(_43263) );
  nnd2s1 _43539_inst ( .DIN1(_43266), .DIN2(_43267), .Q(_43265) );
  nor2s1 _43540_inst ( .DIN1(_43268), .DIN2(_43269), .Q(_43267) );
  nor2s1 _43541_inst ( .DIN1(_43270), .DIN2(_43271), .Q(_43266) );
  nor2s1 _43542_inst ( .DIN1(_43137), .DIN2(_43272), .Q(_43270) );
  nnd2s1 _43543_inst ( .DIN1(_43273), .DIN2(_43274), .Q(_43264) );
  nor2s1 _43544_inst ( .DIN1(_43275), .DIN2(_43276), .Q(_43274) );
  hi1s1 _43545_inst ( .DIN(_43277), .Q(_43276) );
  nor2s1 _43546_inst ( .DIN1(_43278), .DIN2(_43279), .Q(_43273) );
  nor2s1 _43547_inst ( .DIN1(_43280), .DIN2(_43281), .Q(_43262) );
  nnd2s1 _43548_inst ( .DIN1(_43282), .DIN2(_43283), .Q(_43281) );
  nor2s1 _43549_inst ( .DIN1(_43284), .DIN2(_43285), .Q(_43282) );
  nnd2s1 _43550_inst ( .DIN1(_43286), .DIN2(_43287), .Q(_43280) );
  nor2s1 _43551_inst ( .DIN1(_43168), .DIN2(_43159), .Q(_43287) );
  nnd2s1 _43552_inst ( .DIN1(_43288), .DIN2(_43289), .Q(_43168) );
  nor2s1 _43553_inst ( .DIN1(_43248), .DIN2(_43290), .Q(_43289) );
  hi1s1 _43554_inst ( .DIN(_43291), .Q(_43290) );
  nor2s1 _43555_inst ( .DIN1(_43292), .DIN2(_43293), .Q(_43288) );
  nor2s1 _43556_inst ( .DIN1(_43233), .DIN2(_43294), .Q(_43293) );
  nor2s1 _43557_inst ( .DIN1(_43234), .DIN2(_43226), .Q(_43292) );
  nor2s1 _43558_inst ( .DIN1(_43295), .DIN2(_43296), .Q(_43286) );
  nnd2s1 _43559_inst ( .DIN1(_43297), .DIN2(_43298), .Q(
        ____0____________4_____) );
  nnd2s1 _43560_inst ( .DIN1(_43299), .DIN2(_43300), .Q(_43298) );
  xor2s1 _43561_inst ( .DIN1(_43301), .DIN2(_43302), .Q(_43300) );
  xor2s1 _43562_inst ( .DIN1(_53451), .DIN2(_53458), .Q(_43302) );
  nnd2s1 _43563_inst ( .DIN1(_43203), .DIN2(_43303), .Q(_43297) );
  nnd2s1 _43564_inst ( .DIN1(_43304), .DIN2(_43305), .Q(_43303) );
  nor2s1 _43565_inst ( .DIN1(_43306), .DIN2(_43307), .Q(_43305) );
  nnd2s1 _43566_inst ( .DIN1(_43308), .DIN2(_43309), .Q(_43307) );
  hi1s1 _43567_inst ( .DIN(_43310), .Q(_43309) );
  nor2s1 _43568_inst ( .DIN1(_43311), .DIN2(_43312), .Q(_43308) );
  nor2s1 _43569_inst ( .DIN1(_43166), .DIN2(_43313), .Q(_43311) );
  nnd2s1 _43570_inst ( .DIN1(_43314), .DIN2(_43315), .Q(_43306) );
  nor2s1 _43571_inst ( .DIN1(_43316), .DIN2(_43317), .Q(_43315) );
  nor2s1 _43572_inst ( .DIN1(_43318), .DIN2(_43319), .Q(_43314) );
  nor2s1 _43573_inst ( .DIN1(_43294), .DIN2(_43226), .Q(_43318) );
  nor2s1 _43574_inst ( .DIN1(_43320), .DIN2(_43321), .Q(_43304) );
  nnd2s1 _43575_inst ( .DIN1(_43322), .DIN2(_43323), .Q(_43321) );
  nor2s1 _43576_inst ( .DIN1(_43324), .DIN2(_43325), .Q(_43322) );
  nnd2s1 _43577_inst ( .DIN1(_43326), .DIN2(_43327), .Q(_43320) );
  nor2s1 _43578_inst ( .DIN1(_43328), .DIN2(_43169), .Q(_43327) );
  nnd2s1 _43579_inst ( .DIN1(_43329), .DIN2(_43330), .Q(_43169) );
  nor2s1 _43580_inst ( .DIN1(_43331), .DIN2(_43332), .Q(_43330) );
  nnd2s1 _43581_inst ( .DIN1(_43333), .DIN2(_43334), .Q(_43332) );
  nnd2s1 _43582_inst ( .DIN1(_43335), .DIN2(_43336), .Q(_43333) );
  nnd2s1 _43583_inst ( .DIN1(_43337), .DIN2(_43338), .Q(_43331) );
  nor2s1 _43584_inst ( .DIN1(_43339), .DIN2(_43340), .Q(_43329) );
  nnd2s1 _43585_inst ( .DIN1(_43341), .DIN2(_43342), .Q(_43340) );
  nor2s1 _43586_inst ( .DIN1(_43239), .DIN2(_43296), .Q(_43326) );
  nnd2s1 _43587_inst ( .DIN1(_43343), .DIN2(_43344), .Q(_43296) );
  nor2s1 _43588_inst ( .DIN1(_43345), .DIN2(_43346), .Q(_43344) );
  nnd2s1 _43589_inst ( .DIN1(_43347), .DIN2(_43348), .Q(_43346) );
  nnd2s1 _43590_inst ( .DIN1(_43186), .DIN2(_43349), .Q(_43348) );
  nnd2s1 _43591_inst ( .DIN1(_43350), .DIN2(_43351), .Q(_43349) );
  nnd2s1 _43592_inst ( .DIN1(_43352), .DIN2(_43119), .Q(_43347) );
  or2s1 _43593_inst ( .DIN1(_43353), .DIN2(_43354), .Q(_43345) );
  nor2s1 _43594_inst ( .DIN1(_43355), .DIN2(_43356), .Q(_43343) );
  or2s1 _43595_inst ( .DIN1(_43357), .DIN2(_43358), .Q(_43356) );
  nnd2s1 _43596_inst ( .DIN1(_43359), .DIN2(_43360), .Q(_43355) );
  xor2s1 _43597_inst ( .DIN1(_29579), .DIN2(_43361), .Q(_43360) );
  nnd2s1 _43598_inst ( .DIN1(_43362), .DIN2(_43363), .Q(_43361) );
  hi1s1 _43599_inst ( .DIN(_43364), .Q(_43359) );
  nnd2s1 _43600_inst ( .DIN1(_43365), .DIN2(_43366), .Q(_43239) );
  nnd2s1 _43601_inst ( .DIN1(_43119), .DIN2(_43367), .Q(_43366) );
  nnd2s1 _43602_inst ( .DIN1(_43368), .DIN2(_43369), .Q(_43367) );
  or2s1 _43603_inst ( .DIN1(_43370), .DIN2(_43371), .Q(_43365) );
  nnd2s1 _43604_inst ( .DIN1(_43372), .DIN2(_43373), .Q(
        ____0____________3_____) );
  nnd2s1 _43605_inst ( .DIN1(_43374), .DIN2(_43082), .Q(_43373) );
  nnd2s1 _43606_inst ( .DIN1(_43375), .DIN2(______[12]), .Q(_43374) );
  nor2s1 _43607_inst ( .DIN1(_43259), .DIN2(_43376), .Q(_43375) );
  xor2s1 _43608_inst ( .DIN1(_26387), .DIN2(_53448), .Q(_43376) );
  nnd2s1 _43609_inst ( .DIN1(_43377), .DIN2(_41807), .Q(_43372) );
  nor2s1 _43610_inst ( .DIN1(_43378), .DIN2(_43379), .Q(_43377) );
  nnd2s1 _43611_inst ( .DIN1(_43380), .DIN2(_43381), .Q(_43379) );
  nor2s1 _43612_inst ( .DIN1(_43382), .DIN2(_43383), .Q(_43381) );
  or2s1 _43613_inst ( .DIN1(_43384), .DIN2(_43385), .Q(_43383) );
  nnd2s1 _43614_inst ( .DIN1(_43386), .DIN2(_43341), .Q(_43382) );
  and2s1 _43615_inst ( .DIN1(_43387), .DIN2(_43388), .Q(_43341) );
  nnd2s1 _43616_inst ( .DIN1(_43389), .DIN2(_43390), .Q(_43388) );
  nor2s1 _43617_inst ( .DIN1(_26825), .DIN2(_30236), .Q(_43390) );
  nor2s1 _43618_inst ( .DIN1(_32080), .DIN2(_43392), .Q(_43389) );
  or2s1 _43619_inst ( .DIN1(_43123), .DIN2(_43122), .Q(_43387) );
  hi1s1 _43620_inst ( .DIN(_43255), .Q(_43386) );
  nnd2s1 _43621_inst ( .DIN1(_43393), .DIN2(_43394), .Q(_43255) );
  nnd2s1 _43622_inst ( .DIN1(_43395), .DIN2(_43396), .Q(_43394) );
  nor2s1 _43623_inst ( .DIN1(_43397), .DIN2(_43398), .Q(_43380) );
  or2s1 _43624_inst ( .DIN1(_43399), .DIN2(_43400), .Q(_43398) );
  nnd2s1 _43625_inst ( .DIN1(_43401), .DIN2(_43402), .Q(_43378) );
  nor2s1 _43626_inst ( .DIN1(_43403), .DIN2(_43404), .Q(_43402) );
  nnd2s1 _43627_inst ( .DIN1(_43405), .DIN2(_43406), .Q(_43404) );
  nnd2s1 _43628_inst ( .DIN1(_43407), .DIN2(_43408), .Q(_43403) );
  nor2s1 _43629_inst ( .DIN1(_43409), .DIN2(_43410), .Q(_43401) );
  nnd2s1 _43630_inst ( .DIN1(_43411), .DIN2(_43412), .Q(_43410) );
  nnd2s1 _43631_inst ( .DIN1(_43413), .DIN2(_43414), .Q(_43412) );
  or2s1 _43632_inst ( .DIN1(_43226), .DIN2(_43415), .Q(_43411) );
  nnd2s1 _43633_inst ( .DIN1(_43416), .DIN2(_43417), .Q(
        ____0____________2_____) );
  nnd2s1 _43634_inst ( .DIN1(_43418), .DIN2(______[22]), .Q(_43417) );
  nor2s1 _43635_inst ( .DIN1(_43259), .DIN2(_43419), .Q(_43418) );
  xor2s1 _43636_inst ( .DIN1(_43420), .DIN2(_26334), .Q(_43419) );
  hi1s1 _43637_inst ( .DIN(_41806), .Q(_43259) );
  nnd2s1 _43638_inst ( .DIN1(_43421), .DIN2(_43422), .Q(_41806) );
  nor2s1 _43639_inst ( .DIN1(_29433), .DIN2(_32807), .Q(_43421) );
  nnd2s1 _43640_inst ( .DIN1(_41807), .DIN2(_43423), .Q(_43416) );
  nnd2s1 _43641_inst ( .DIN1(_43424), .DIN2(_43425), .Q(_43423) );
  nor2s1 _43642_inst ( .DIN1(_43426), .DIN2(_43427), .Q(_43425) );
  nnd2s1 _43643_inst ( .DIN1(_43428), .DIN2(_43429), .Q(_43427) );
  nor2s1 _43644_inst ( .DIN1(_43430), .DIN2(_43431), .Q(_43429) );
  nor2s1 _43645_inst ( .DIN1(_43432), .DIN2(_43433), .Q(_43428) );
  nor2s1 _43646_inst ( .DIN1(_43434), .DIN2(_43435), .Q(_43432) );
  nnd2s1 _43647_inst ( .DIN1(_43436), .DIN2(_43437), .Q(_43426) );
  and2s1 _43648_inst ( .DIN1(_43438), .DIN2(_43439), .Q(_43437) );
  nor2s1 _43649_inst ( .DIN1(_43440), .DIN2(_43248), .Q(_43436) );
  nor2s1 _43650_inst ( .DIN1(_43441), .DIN2(_43233), .Q(_43248) );
  nor2s1 _43651_inst ( .DIN1(_43442), .DIN2(_43443), .Q(_43424) );
  nnd2s1 _43652_inst ( .DIN1(_43444), .DIN2(_43445), .Q(_43443) );
  hi1s1 _43653_inst ( .DIN(_43446), .Q(_43445) );
  nor2s1 _43654_inst ( .DIN1(_43447), .DIN2(_43448), .Q(_43444) );
  nnd2s1 _43655_inst ( .DIN1(_43449), .DIN2(_43450), .Q(_43442) );
  nor2s1 _43656_inst ( .DIN1(_43181), .DIN2(_43451), .Q(_43450) );
  nnd2s1 _43657_inst ( .DIN1(_43452), .DIN2(_43453), .Q(_43181) );
  nor2s1 _43658_inst ( .DIN1(_43454), .DIN2(_43455), .Q(_43453) );
  nnd2s1 _43659_inst ( .DIN1(_43456), .DIN2(_43457), .Q(_43455) );
  nnd2s1 _43660_inst ( .DIN1(_43458), .DIN2(_26770), .Q(_43457) );
  nor2s1 _43661_inst ( .DIN1(_43459), .DIN2(_43460), .Q(_43456) );
  nor2s1 _43662_inst ( .DIN1(_43461), .DIN2(_43462), .Q(_43460) );
  nor2s1 _43663_inst ( .DIN1(_26825), .DIN2(_43294), .Q(_43459) );
  hi1s1 _43664_inst ( .DIN(_43395), .Q(_43294) );
  nnd2s1 _43665_inst ( .DIN1(_43463), .DIN2(_43464), .Q(_43454) );
  nor2s1 _43666_inst ( .DIN1(_43465), .DIN2(_43466), .Q(_43463) );
  nor2s1 _43667_inst ( .DIN1(_43467), .DIN2(_43468), .Q(_43452) );
  nnd2s1 _43668_inst ( .DIN1(_43469), .DIN2(_43470), .Q(_43468) );
  xor2s1 _43669_inst ( .DIN1(_33865), .DIN2(_43471), .Q(_43470) );
  nor2s1 _43670_inst ( .DIN1(_43472), .DIN2(_43473), .Q(_43471) );
  and2s1 _43671_inst ( .DIN1(_43474), .DIN2(_43475), .Q(_43472) );
  nor2s1 _43672_inst ( .DIN1(_43476), .DIN2(_43477), .Q(_43469) );
  nnd2s1 _43673_inst ( .DIN1(_43478), .DIN2(_43479), .Q(_43467) );
  hi1s1 _43674_inst ( .DIN(_43271), .Q(_43479) );
  nnd2s1 _43675_inst ( .DIN1(_43480), .DIN2(_43481), .Q(_43271) );
  nor2s1 _43676_inst ( .DIN1(_43482), .DIN2(_43483), .Q(_43481) );
  hi1s1 _43677_inst ( .DIN(_43484), .Q(_43482) );
  nor2s1 _43678_inst ( .DIN1(_43485), .DIN2(_43486), .Q(_43480) );
  nor2s1 _43679_inst ( .DIN1(_43487), .DIN2(_43310), .Q(_43478) );
  nnd2s1 _43680_inst ( .DIN1(_43488), .DIN2(_43489), .Q(_43310) );
  nor2s1 _43681_inst ( .DIN1(_43490), .DIN2(_43491), .Q(_43487) );
  nor2s1 _43682_inst ( .DIN1(_43492), .DIN2(_43493), .Q(_43449) );
  hi1s1 _43683_inst ( .DIN(_43082), .Q(_41807) );
  nnd2s1 _43684_inst ( .DIN1(_43494), .DIN2(_43495), .Q(_43082) );
  nor2s1 _43685_inst ( .DIN1(_27310), .DIN2(_43496), .Q(_43495) );
  nnd2s1 _43686_inst ( .DIN1(_27441), .DIN2(_43497), .Q(_43496) );
  nor2s1 _43687_inst ( .DIN1(_27311), .DIN2(_43498), .Q(_43494) );
  nnd2s1 _43688_inst ( .DIN1(_43499), .DIN2(_43500), .Q(
        ____0____________1_____) );
  nnd2s1 _43689_inst ( .DIN1(_43501), .DIN2(_43299), .Q(_43500) );
  nor2s1 _43690_inst ( .DIN1(_43502), .DIN2(_43203), .Q(_43299) );
  nor2s1 _43691_inst ( .DIN1(_27039), .DIN2(_26353), .Q(_43501) );
  nnd2s1 _43692_inst ( .DIN1(_43203), .DIN2(_43503), .Q(_43499) );
  nnd2s1 _43693_inst ( .DIN1(_43504), .DIN2(_43505), .Q(_43503) );
  nor2s1 _43694_inst ( .DIN1(_43506), .DIN2(_43507), .Q(_43505) );
  nnd2s1 _43695_inst ( .DIN1(_43508), .DIN2(_43509), .Q(_43507) );
  nor2s1 _43696_inst ( .DIN1(_43510), .DIN2(_43511), .Q(_43509) );
  nor2s1 _43697_inst ( .DIN1(_43512), .DIN2(_43140), .Q(_43511) );
  nor2s1 _43698_inst ( .DIN1(_43513), .DIN2(_43514), .Q(_43510) );
  nor2s1 _43699_inst ( .DIN1(_43515), .DIN2(_43516), .Q(_43513) );
  nor2s1 _43700_inst ( .DIN1(_43517), .DIN2(_43518), .Q(_43508) );
  nor2s1 _43701_inst ( .DIN1(_43233), .DIN2(_43519), .Q(_43518) );
  nor2s1 _43702_inst ( .DIN1(_43520), .DIN2(_43521), .Q(_43517) );
  nnd2s1 _43703_inst ( .DIN1(_43522), .DIN2(_43523), .Q(_43506) );
  nor2s1 _43704_inst ( .DIN1(_43524), .DIN2(_43525), .Q(_43523) );
  or2s1 _43705_inst ( .DIN1(_43526), .DIN2(_43278), .Q(_43525) );
  nor2s1 _43706_inst ( .DIN1(_43527), .DIN2(_43353), .Q(_43522) );
  nor2s1 _43707_inst ( .DIN1(_43528), .DIN2(_43529), .Q(_43504) );
  nnd2s1 _43708_inst ( .DIN1(_43530), .DIN2(_43531), .Q(_43529) );
  nor2s1 _43709_inst ( .DIN1(_43532), .DIN2(_43533), .Q(_43531) );
  nor2s1 _43710_inst ( .DIN1(_43534), .DIN2(_43535), .Q(_43530) );
  nnd2s1 _43711_inst ( .DIN1(_43536), .DIN2(_43537), .Q(_43528) );
  nor2s1 _43712_inst ( .DIN1(_43538), .DIN2(_43158), .Q(_43537) );
  nnd2s1 _43713_inst ( .DIN1(_43539), .DIN2(_43540), .Q(_43158) );
  nor2s1 _43714_inst ( .DIN1(_43541), .DIN2(_43542), .Q(_43540) );
  nnd2s1 _43715_inst ( .DIN1(_43543), .DIN2(_43544), .Q(_43542) );
  hi1s1 _43716_inst ( .DIN(_43430), .Q(_43543) );
  nor2s1 _43717_inst ( .DIN1(_43166), .DIN2(_43545), .Q(_43541) );
  nor2s1 _43718_inst ( .DIN1(_43546), .DIN2(_43547), .Q(_43539) );
  nor2s1 _43719_inst ( .DIN1(_43252), .DIN2(_43548), .Q(_43547) );
  nor2s1 _43720_inst ( .DIN1(_43137), .DIN2(_43253), .Q(_43546) );
  nor2s1 _43721_inst ( .DIN1(_43549), .DIN2(_43400), .Q(_43536) );
  nnd2s1 _43722_inst ( .DIN1(_43550), .DIN2(_43551), .Q(_43400) );
  nor2s1 _43723_inst ( .DIN1(_43552), .DIN2(_43553), .Q(_43551) );
  or2s1 _43724_inst ( .DIN1(_43254), .DIN2(_43201), .Q(_43553) );
  nnd2s1 _43725_inst ( .DIN1(_43554), .DIN2(_43555), .Q(_43201) );
  nnd2s1 _43726_inst ( .DIN1(_43556), .DIN2(_43336), .Q(_43555) );
  nor2s1 _43727_inst ( .DIN1(_43557), .DIN2(_43141), .Q(_43554) );
  nor2s1 _43728_inst ( .DIN1(_43252), .DIN2(_43558), .Q(_43141) );
  nor2s1 _43729_inst ( .DIN1(_43151), .DIN2(_43559), .Q(_43557) );
  nnd2s1 _43730_inst ( .DIN1(_43484), .DIN2(_43560), .Q(_43254) );
  nnd2s1 _43731_inst ( .DIN1(_43561), .DIN2(_43562), .Q(_43560) );
  nnd2s1 _43732_inst ( .DIN1(_43563), .DIN2(_43564), .Q(_43484) );
  nor2s1 _43733_inst ( .DIN1(_43565), .DIN2(_43566), .Q(_43563) );
  nor2s1 _43734_inst ( .DIN1(_43567), .DIN2(_43568), .Q(_43566) );
  nnd2s1 _43735_inst ( .DIN1(_43569), .DIN2(_43570), .Q(_43552) );
  hi1s1 _43736_inst ( .DIN(_43159), .Q(_43569) );
  nnd2s1 _43737_inst ( .DIN1(_43571), .DIN2(_43572), .Q(_43159) );
  nnd2s1 _43738_inst ( .DIN1(_43573), .DIN2(_43574), .Q(_43572) );
  nor2s1 _43739_inst ( .DIN1(_43575), .DIN2(_43576), .Q(_43550) );
  or2s1 _43740_inst ( .DIN1(_43577), .DIN2(_43578), .Q(_43576) );
  xor2s1 _43741_inst ( .DIN1(_40991), .DIN2(_43579), .Q(_43575) );
  nor2s1 _43742_inst ( .DIN1(_43580), .DIN2(_43581), .Q(_43579) );
  nnd2s1 _43743_inst ( .DIN1(_43582), .DIN2(_43583), .Q(_43581) );
  hi1s1 _43744_inst ( .DIN(_43447), .Q(_43583) );
  nnd2s1 _43745_inst ( .DIN1(_43291), .DIN2(_43584), .Q(_43447) );
  nnd2s1 _43746_inst ( .DIN1(_43585), .DIN2(_43586), .Q(_43584) );
  nor2s1 _43747_inst ( .DIN1(_43587), .DIN2(_43588), .Q(_43582) );
  nnd2s1 _43748_inst ( .DIN1(_43589), .DIN2(_43590), .Q(_43580) );
  nor2s1 _43749_inst ( .DIN1(_43591), .DIN2(_43317), .Q(_43590) );
  nor2s1 _43750_inst ( .DIN1(_43592), .DIN2(_43593), .Q(_43589) );
  nor2s1 _43751_inst ( .DIN1(_43233), .DIN2(_43230), .Q(_43593) );
  nor2s1 _43752_inst ( .DIN1(_43565), .DIN2(_43594), .Q(_43592) );
  nnd2s1 _43753_inst ( .DIN1(_43595), .DIN2(_43596), .Q(
        ____0____________15_____) );
  nnd2s1 _43754_inst ( .DIN1(_43597), .DIN2(_35502), .Q(_43596) );
  hi1s1 _43755_inst ( .DIN(_27895), .Q(_35502) );
  nnd2s1 _43756_inst ( .DIN1(_43598), .DIN2(_35501), .Q(_43597) );
  or2s1 _43757_inst ( .DIN1(_43599), .DIN2(_33181), .Q(_35501) );
  xor2s1 _43758_inst ( .DIN1(_53069), .DIN2(_43600), .Q(_43598) );
  nor2s1 _43759_inst ( .DIN1(_53430), .DIN2(_26576), .Q(_43600) );
  nnd2s1 _43760_inst ( .DIN1(_43601), .DIN2(_27895), .Q(_43595) );
  nor2s1 _43761_inst ( .DIN1(_37702), .DIN2(_33696), .Q(_27895) );
  nnd2s1 _43762_inst ( .DIN1(_34488), .DIN2(_43602), .Q(_33696) );
  and2s1 _43763_inst ( .DIN1(_43603), .DIN2(_43604), .Q(_34488) );
  nor2s1 _43764_inst ( .DIN1(_38884), .DIN2(_43605), .Q(_43604) );
  nnd2s1 _43765_inst ( .DIN1(_34485), .DIN2(_30174), .Q(_43605) );
  nor2s1 _43766_inst ( .DIN1(_33182), .DIN2(_38853), .Q(_43603) );
  nor2s1 _43767_inst ( .DIN1(_43606), .DIN2(_43607), .Q(_43601) );
  nnd2s1 _43768_inst ( .DIN1(_43608), .DIN2(_43609), .Q(_43607) );
  nor2s1 _43769_inst ( .DIN1(_43610), .DIN2(_43611), .Q(_43609) );
  or2s1 _43770_inst ( .DIN1(_43202), .DIN2(_43165), .Q(_43611) );
  nnd2s1 _43771_inst ( .DIN1(_43612), .DIN2(_43613), .Q(_43165) );
  nor2s1 _43772_inst ( .DIN1(_43614), .DIN2(_43615), .Q(_43613) );
  nnd2s1 _43773_inst ( .DIN1(_43616), .DIN2(_43617), .Q(_43615) );
  nor2s1 _43774_inst ( .DIN1(_43618), .DIN2(_43619), .Q(_43616) );
  nor2s1 _43775_inst ( .DIN1(_43620), .DIN2(_43621), .Q(_43618) );
  nnd2s1 _43776_inst ( .DIN1(_43622), .DIN2(_43623), .Q(_43614) );
  nor2s1 _43777_inst ( .DIN1(_43278), .DIN2(_43624), .Q(_43623) );
  nor2s1 _43778_inst ( .DIN1(_43625), .DIN2(_43112), .Q(_43622) );
  nor2s1 _43779_inst ( .DIN1(_43626), .DIN2(_43627), .Q(_43612) );
  nnd2s1 _43780_inst ( .DIN1(_43628), .DIN2(_43629), .Q(_43627) );
  hi1s1 _43781_inst ( .DIN(_43451), .Q(_43629) );
  nor2s1 _43782_inst ( .DIN1(_43364), .DIN2(_43630), .Q(_43628) );
  nnd2s1 _43783_inst ( .DIN1(_43631), .DIN2(_43632), .Q(_43364) );
  nnd2s1 _43784_inst ( .DIN1(_43561), .DIN2(_43414), .Q(_43632) );
  nnd2s1 _43785_inst ( .DIN1(_43633), .DIN2(_43634), .Q(_43626) );
  hi1s1 _43786_inst ( .DIN(_43328), .Q(_43634) );
  nnd2s1 _43787_inst ( .DIN1(_43635), .DIN2(_43636), .Q(_43328) );
  nor2s1 _43788_inst ( .DIN1(_43465), .DIN2(_43637), .Q(_43636) );
  nor2s1 _43789_inst ( .DIN1(_43638), .DIN2(_43151), .Q(_43637) );
  nor2s1 _43790_inst ( .DIN1(_43413), .DIN2(_43639), .Q(_43638) );
  nor2s1 _43791_inst ( .DIN1(_43640), .DIN2(_43641), .Q(_43635) );
  nor2s1 _43792_inst ( .DIN1(_43514), .DIN2(_43475), .Q(_43640) );
  nor2s1 _43793_inst ( .DIN1(_43245), .DIN2(_43183), .Q(_43633) );
  xnr2s1 _43794_inst ( .DIN1(_31975), .DIN2(_43642), .Q(_43183) );
  nor2s1 _43795_inst ( .DIN1(_43643), .DIN2(_43644), .Q(_43642) );
  nnd2s1 _43796_inst ( .DIN1(_43645), .DIN2(_43646), .Q(_43644) );
  hi1s1 _43797_inst ( .DIN(_43647), .Q(_43646) );
  nor2s1 _43798_inst ( .DIN1(_43648), .DIN2(_43588), .Q(_43645) );
  nnd2s1 _43799_inst ( .DIN1(_43649), .DIN2(_43650), .Q(_43643) );
  nor2s1 _43800_inst ( .DIN1(_43651), .DIN2(_43527), .Q(_43650) );
  hi1s1 _43801_inst ( .DIN(_43652), .Q(_43527) );
  nor2s1 _43802_inst ( .DIN1(_43268), .DIN2(_43653), .Q(_43649) );
  nnd2s1 _43803_inst ( .DIN1(_43654), .DIN2(_43655), .Q(_43202) );
  nor2s1 _43804_inst ( .DIN1(_43656), .DIN2(_43657), .Q(_43655) );
  nor2s1 _43805_inst ( .DIN1(_43514), .DIN2(_43658), .Q(_43657) );
  nor2s1 _43806_inst ( .DIN1(_43565), .DIN2(_43659), .Q(_43656) );
  nor2s1 _43807_inst ( .DIN1(_43660), .DIN2(_43661), .Q(_43659) );
  nor2s1 _43808_inst ( .DIN1(_43662), .DIN2(_43663), .Q(_43654) );
  nor2s1 _43809_inst ( .DIN1(_43664), .DIN2(_43313), .Q(_43662) );
  nnd2s1 _43810_inst ( .DIN1(_43665), .DIN2(_43099), .Q(_43610) );
  and2s1 _43811_inst ( .DIN1(_43666), .DIN2(_43667), .Q(_43099) );
  nor2s1 _43812_inst ( .DIN1(_43668), .DIN2(_43669), .Q(_43667) );
  or2s1 _43813_inst ( .DIN1(_43354), .DIN2(_43670), .Q(_43669) );
  nnd2s1 _43814_inst ( .DIN1(_43671), .DIN2(_43439), .Q(_43668) );
  nor2s1 _43815_inst ( .DIN1(_43672), .DIN2(_43279), .Q(_43671) );
  nor2s1 _43816_inst ( .DIN1(_43673), .DIN2(_43674), .Q(_43666) );
  or2s1 _43817_inst ( .DIN1(_43433), .DIN2(_43312), .Q(_43674) );
  nnd2s1 _43818_inst ( .DIN1(_43675), .DIN2(_43676), .Q(_43312) );
  or2s1 _43819_inst ( .DIN1(_43229), .DIN2(_43233), .Q(_43676) );
  nnd2s1 _43820_inst ( .DIN1(_43677), .DIN2(_43678), .Q(_43433) );
  nor2s1 _43821_inst ( .DIN1(_43679), .DIN2(_43680), .Q(_43677) );
  nor2s1 _43822_inst ( .DIN1(_43252), .DIN2(_43681), .Q(_43680) );
  nnd2s1 _43823_inst ( .DIN1(_43682), .DIN2(_43683), .Q(_43673) );
  hi1s1 _43824_inst ( .DIN(_43220), .Q(_43683) );
  nnd2s1 _43825_inst ( .DIN1(_43684), .DIN2(_43685), .Q(_43220) );
  nnd2s1 _43826_inst ( .DIN1(_43686), .DIN2(_26770), .Q(_43685) );
  xor2s1 _43827_inst ( .DIN1(_43687), .DIN2(_43688), .Q(_43684) );
  nor2s1 _43828_inst ( .DIN1(_43689), .DIN2(_43690), .Q(_43688) );
  nor2s1 _43829_inst ( .DIN1(_43137), .DIN2(_43558), .Q(_43689) );
  nor2s1 _43830_inst ( .DIN1(_43691), .DIN2(_43692), .Q(_43682) );
  and2s1 _43831_inst ( .DIN1(_43414), .DIN2(_43516), .Q(_43692) );
  nor2s1 _43832_inst ( .DIN1(_43514), .DIN2(_43693), .Q(_43691) );
  nor2s1 _43833_inst ( .DIN1(_43694), .DIN2(_43695), .Q(_43608) );
  or2s1 _43834_inst ( .DIN1(_43532), .DIN2(_43284), .Q(_43695) );
  nnd2s1 _43835_inst ( .DIN1(_43696), .DIN2(_43697), .Q(_43284) );
  nor2s1 _43836_inst ( .DIN1(_43698), .DIN2(_43699), .Q(_43697) );
  nor2s1 _43837_inst ( .DIN1(_43700), .DIN2(_43701), .Q(_43696) );
  nnd2s1 _43838_inst ( .DIN1(_43702), .DIN2(_43703), .Q(_43532) );
  nnd2s1 _43839_inst ( .DIN1(_43704), .DIN2(_43705), .Q(_43703) );
  nnd2s1 _43840_inst ( .DIN1(_43706), .DIN2(_43707), .Q(_43702) );
  nnd2s1 _43841_inst ( .DIN1(_43708), .DIN2(_43709), .Q(_43606) );
  nor2s1 _43842_inst ( .DIN1(_43710), .DIN2(_43711), .Q(_43709) );
  nnd2s1 _43843_inst ( .DIN1(_43712), .DIN2(_43713), .Q(_43711) );
  nnd2s1 _43844_inst ( .DIN1(_43714), .DIN2(_43715), .Q(_43710) );
  hi1s1 _43845_inst ( .DIN(_43223), .Q(_43714) );
  nor2s1 _43846_inst ( .DIN1(_43716), .DIN2(_43717), .Q(_43708) );
  nnd2s1 _43847_inst ( .DIN1(_43489), .DIN2(_43718), .Q(_43717) );
  nnd2s1 _43848_inst ( .DIN1(_43719), .DIN2(_43720), .Q(_43718) );
  nor2s1 _43849_inst ( .DIN1(_43392), .DIN2(_43226), .Q(_43719) );
  nnd2s1 _43850_inst ( .DIN1(_43145), .DIN2(_39969), .Q(_43489) );
  nnd2s1 _43851_inst ( .DIN1(_43721), .DIN2(_43722), .Q(_43716) );
  nnd2s1 _43852_inst ( .DIN1(_43723), .DIN2(_43396), .Q(_43722) );
  nnd2s1 _43853_inst ( .DIN1(_43724), .DIN2(_43725), .Q(_43721) );
  nnd2s1 _43854_inst ( .DIN1(_43726), .DIN2(_27970), .Q(
        ____0____________14_____) );
  nnd2s1 _43855_inst ( .DIN1(_27913), .DIN2(_27973), .Q(_27970) );
  hi1s1 _43856_inst ( .DIN(_37213), .Q(_27913) );
  nnd2s1 _43857_inst ( .DIN1(_43727), .DIN2(_39745), .Q(_37213) );
  nor2s1 _43858_inst ( .DIN1(_43728), .DIN2(_43729), .Q(_43726) );
  nor2s1 _43859_inst ( .DIN1(_27973), .DIN2(_43730), .Q(_43729) );
  nnd2s1 _43860_inst ( .DIN1(_43731), .DIN2(_43732), .Q(_43730) );
  nor2s1 _43861_inst ( .DIN1(_43733), .DIN2(_43734), .Q(_43732) );
  nnd2s1 _43862_inst ( .DIN1(_43735), .DIN2(_43736), .Q(_43734) );
  nor2s1 _43863_inst ( .DIN1(_43737), .DIN2(_43738), .Q(_43736) );
  nnd2s1 _43864_inst ( .DIN1(_43739), .DIN2(_43740), .Q(_43738) );
  or2s1 _43865_inst ( .DIN1(_43475), .DIN2(_43514), .Q(_43740) );
  nnd2s1 _43866_inst ( .DIN1(_43741), .DIN2(_43742), .Q(_43739) );
  nor2s1 _43867_inst ( .DIN1(_43391), .DIN2(_43743), .Q(_43737) );
  nor2s1 _43868_inst ( .DIN1(_43744), .DIN2(_43486), .Q(_43735) );
  nnd2s1 _43869_inst ( .DIN1(_43745), .DIN2(_43746), .Q(_43486) );
  nnd2s1 _43870_inst ( .DIN1(_43747), .DIN2(_43119), .Q(_43746) );
  nnd2s1 _43871_inst ( .DIN1(_43748), .DIN2(_43749), .Q(_43745) );
  nor2s1 _43872_inst ( .DIN1(_43750), .DIN2(_43096), .Q(_43744) );
  nor2s1 _43873_inst ( .DIN1(_43751), .DIN2(_43352), .Q(_43750) );
  nnd2s1 _43874_inst ( .DIN1(_43752), .DIN2(_43753), .Q(_43733) );
  nor2s1 _43875_inst ( .DIN1(_43191), .DIN2(_43754), .Q(_43753) );
  nnd2s1 _43876_inst ( .DIN1(_43755), .DIN2(_43438), .Q(_43754) );
  hi1s1 _43877_inst ( .DIN(_43756), .Q(_43191) );
  nor2s1 _43878_inst ( .DIN1(_43757), .DIN2(_43758), .Q(_43752) );
  nor2s1 _43879_inst ( .DIN1(_42312), .DIN2(_43226), .Q(_43758) );
  nor2s1 _43880_inst ( .DIN1(_43371), .DIN2(_43759), .Q(_43757) );
  nor2s1 _43881_inst ( .DIN1(_43760), .DIN2(_43761), .Q(_43731) );
  nnd2s1 _43882_inst ( .DIN1(_43762), .DIN2(_43763), .Q(_43761) );
  nor2s1 _43883_inst ( .DIN1(_43694), .DIN2(_43764), .Q(_43763) );
  nnd2s1 _43884_inst ( .DIN1(_43765), .DIN2(_43766), .Q(_43764) );
  hi1s1 _43885_inst ( .DIN(_43533), .Q(_43765) );
  nnd2s1 _43886_inst ( .DIN1(_43767), .DIN2(_43768), .Q(_43533) );
  nor2s1 _43887_inst ( .DIN1(_43769), .DIN2(_43770), .Q(_43768) );
  nor2s1 _43888_inst ( .DIN1(_43771), .DIN2(_43772), .Q(_43767) );
  nor2s1 _43889_inst ( .DIN1(_43252), .DIN2(_43368), .Q(_43771) );
  nnd2s1 _43890_inst ( .DIN1(_43773), .DIN2(_43488), .Q(_43694) );
  and2s1 _43891_inst ( .DIN1(_43774), .DIN2(_43775), .Q(_43488) );
  nnd2s1 _43892_inst ( .DIN1(_43515), .DIN2(_26770), .Q(_43775) );
  nnd2s1 _43893_inst ( .DIN1(_43776), .DIN2(_43707), .Q(_43774) );
  nor2s1 _43894_inst ( .DIN1(_43777), .DIN2(_43778), .Q(_43773) );
  nor2s1 _43895_inst ( .DIN1(_43779), .DIN2(_43780), .Q(_43778) );
  nor2s1 _43896_inst ( .DIN1(_43781), .DIN2(_43782), .Q(_43777) );
  nnd2s1 _43897_inst ( .DIN1(_43564), .DIN2(_43108), .Q(_43782) );
  nor2s1 _43898_inst ( .DIN1(_43783), .DIN2(_43784), .Q(_43762) );
  nnd2s1 _43899_inst ( .DIN1(_43785), .DIN2(_43786), .Q(_43760) );
  nor2s1 _43900_inst ( .DIN1(_43325), .DIN2(_43787), .Q(_43786) );
  or2s1 _43901_inst ( .DIN1(_43240), .DIN2(_43160), .Q(_43787) );
  nnd2s1 _43902_inst ( .DIN1(_43788), .DIN2(_43789), .Q(_43160) );
  nnd2s1 _43903_inst ( .DIN1(_43660), .DIN2(_43790), .Q(_43789) );
  nor2s1 _43904_inst ( .DIN1(_43431), .DIN2(_43791), .Q(_43788) );
  nor2s1 _43905_inst ( .DIN1(_43461), .DIN2(_43434), .Q(_43791) );
  nor2s1 _43906_inst ( .DIN1(_43391), .DIN2(_43229), .Q(_43431) );
  nnd2s1 _43907_inst ( .DIN1(_43792), .DIN2(_43793), .Q(_43240) );
  nor2s1 _43908_inst ( .DIN1(_43142), .DIN2(_43794), .Q(_43793) );
  nnd2s1 _43909_inst ( .DIN1(_43795), .DIN2(_43337), .Q(_43794) );
  nor2s1 _43910_inst ( .DIN1(_43520), .DIN2(_43796), .Q(_43142) );
  nor2s1 _43911_inst ( .DIN1(_43797), .DIN2(_43798), .Q(_43792) );
  or2s1 _43912_inst ( .DIN1(_43485), .DIN2(_43799), .Q(_43798) );
  nnd2s1 _43913_inst ( .DIN1(_43570), .DIN2(_43405), .Q(_43485) );
  nnd2s1 _43914_inst ( .DIN1(_43706), .DIN2(_26770), .Q(_43405) );
  hi1s1 _43915_inst ( .DIN(_43800), .Q(_43706) );
  and2s1 _43916_inst ( .DIN1(_43712), .DIN2(_43801), .Q(_43570) );
  or2s1 _43917_inst ( .DIN1(_43620), .DIN2(_43565), .Q(_43801) );
  nnd2s1 _43918_inst ( .DIN1(_43802), .DIN2(_43803), .Q(_43712) );
  nor2s1 _43919_inst ( .DIN1(_43804), .DIN2(_43805), .Q(_43803) );
  nnd2s1 _43920_inst ( .DIN1(_43806), .DIN2(_26770), .Q(_43805) );
  and2s1 _43921_inst ( .DIN1(_43807), .DIN2(_43808), .Q(_43802) );
  xor2s1 _43922_inst ( .DIN1(_32005), .DIN2(_43809), .Q(_43797) );
  nor2s1 _43923_inst ( .DIN1(_43430), .DIN2(_43353), .Q(_43809) );
  and2s1 _43924_inst ( .DIN1(_43810), .DIN2(_29203), .Q(_43353) );
  nor2s1 _43925_inst ( .DIN1(_43811), .DIN2(_43151), .Q(_43810) );
  nor2s1 _43926_inst ( .DIN1(_43812), .DIN2(_43096), .Q(_43430) );
  nnd2s1 _43927_inst ( .DIN1(_43813), .DIN2(_43814), .Q(_43325) );
  nnd2s1 _43928_inst ( .DIN1(_43815), .DIN2(_43704), .Q(_43814) );
  nnd2s1 _43929_inst ( .DIN1(_43458), .DIN2(_43396), .Q(_43813) );
  hi1s1 _43930_inst ( .DIN(_43816), .Q(_43458) );
  nor2s1 _43931_inst ( .DIN1(_43817), .DIN2(_43818), .Q(_43785) );
  nor2s1 _43932_inst ( .DIN1(_53431), .DIN2(_27915), .Q(_43728) );
  hi1s1 _43933_inst ( .DIN(_27973), .Q(_27915) );
  nnd2s1 _43934_inst ( .DIN1(_43819), .DIN2(_43727), .Q(_27973) );
  nor2s1 _43935_inst ( .DIN1(_34490), .DIN2(_38884), .Q(_43727) );
  nor2s1 _43936_inst ( .DIN1(_36302), .DIN2(_37702), .Q(_43819) );
  nnd2s1 _43937_inst ( .DIN1(_39745), .DIN2(_34485), .Q(_36302) );
  nnd2s1 _43938_inst ( .DIN1(_43820), .DIN2(_43821), .Q(
        ____0____________13_____) );
  nnd2s1 _43939_inst ( .DIN1(_43822), .DIN2(_43823), .Q(_43821) );
  xor2s1 _43940_inst ( .DIN1(_52915), .DIN2(_53432), .Q(_43823) );
  hi1s1 _43941_inst ( .DIN(_28976), .Q(_43822) );
  nnd2s1 _43942_inst ( .DIN1(_27325), .DIN2(_43824), .Q(_43820) );
  nnd2s1 _43943_inst ( .DIN1(_43825), .DIN2(_43826), .Q(_43824) );
  nor2s1 _43944_inst ( .DIN1(_43827), .DIN2(_43828), .Q(_43826) );
  nnd2s1 _43945_inst ( .DIN1(_43829), .DIN2(_43830), .Q(_43828) );
  nor2s1 _43946_inst ( .DIN1(_43831), .DIN2(_43161), .Q(_43830) );
  nnd2s1 _43947_inst ( .DIN1(_43832), .DIN2(_43833), .Q(_43161) );
  nor2s1 _43948_inst ( .DIN1(_43834), .DIN2(_43835), .Q(_43833) );
  nor2s1 _43949_inst ( .DIN1(_43594), .DIN2(_43664), .Q(_43835) );
  nor2s1 _43950_inst ( .DIN1(_43799), .DIN2(_43836), .Q(_43832) );
  nor2s1 _43951_inst ( .DIN1(_43837), .DIN2(_43838), .Q(_43829) );
  nnd2s1 _43952_inst ( .DIN1(_43839), .DIN2(_43840), .Q(_43827) );
  and2s1 _43953_inst ( .DIN1(_43841), .DIN2(_43464), .Q(_43840) );
  hi1s1 _43954_inst ( .DIN(_43842), .Q(_43464) );
  nor2s1 _43955_inst ( .DIN1(_43591), .DIN2(_43843), .Q(_43839) );
  and2s1 _43956_inst ( .DIN1(_43414), .DIN2(_43844), .Q(_43843) );
  hi1s1 _43957_inst ( .DIN(_43755), .Q(_43591) );
  nnd2s1 _43958_inst ( .DIN1(_43845), .DIN2(_43586), .Q(_43755) );
  nor2s1 _43959_inst ( .DIN1(_43846), .DIN2(_43847), .Q(_43825) );
  nnd2s1 _43960_inst ( .DIN1(_43848), .DIN2(_43849), .Q(_43847) );
  hi1s1 _43961_inst ( .DIN(_43850), .Q(_43849) );
  nor2s1 _43962_inst ( .DIN1(_43534), .DIN2(_43851), .Q(_43848) );
  nnd2s1 _43963_inst ( .DIN1(_43852), .DIN2(_43853), .Q(_43534) );
  nor2s1 _43964_inst ( .DIN1(_43107), .DIN2(_43854), .Q(_43853) );
  nnd2s1 _43965_inst ( .DIN1(_43438), .DIN2(_43855), .Q(_43854) );
  nnd2s1 _43966_inst ( .DIN1(_43815), .DIN2(_43856), .Q(_43438) );
  nor2s1 _43967_inst ( .DIN1(_43857), .DIN2(_43858), .Q(_43852) );
  nnd2s1 _43968_inst ( .DIN1(_43859), .DIN2(_43860), .Q(_43846) );
  and2s1 _43969_inst ( .DIN1(_43323), .DIN2(_43861), .Q(_43860) );
  and2s1 _43970_inst ( .DIN1(_43862), .DIN2(_43795), .Q(_43323) );
  nnd2s1 _43971_inst ( .DIN1(_43863), .DIN2(_43186), .Q(_43795) );
  or2s1 _43972_inst ( .DIN1(_43759), .DIN2(_43864), .Q(_43862) );
  nor2s1 _43973_inst ( .DIN1(_43385), .DIN2(_43865), .Q(_43859) );
  nnd2s1 _43974_inst ( .DIN1(_43866), .DIN2(_43867), .Q(_43385) );
  nor2s1 _43975_inst ( .DIN1(_43868), .DIN2(_43869), .Q(_43867) );
  nnd2s1 _43976_inst ( .DIN1(_43870), .DIN2(_43871), .Q(_43869) );
  or2s1 _43977_inst ( .DIN1(_43658), .DIN2(_43514), .Q(_43871) );
  nor2s1 _43978_inst ( .DIN1(_43872), .DIN2(_43873), .Q(_43870) );
  nor2s1 _43979_inst ( .DIN1(_43096), .DIN2(_43218), .Q(_43873) );
  nor2s1 _43980_inst ( .DIN1(_43519), .DIN2(_43226), .Q(_43872) );
  nnd2s1 _43981_inst ( .DIN1(_43874), .DIN2(_43875), .Q(_43868) );
  hi1s1 _43982_inst ( .DIN(_43217), .Q(_43875) );
  nor2s1 _43983_inst ( .DIN1(_43876), .DIN2(_43461), .Q(_43217) );
  nor2s1 _43984_inst ( .DIN1(_43625), .DIN2(_43877), .Q(_43874) );
  hi1s1 _43985_inst ( .DIN(_43878), .Q(_43625) );
  nor2s1 _43986_inst ( .DIN1(_43879), .DIN2(_43880), .Q(_43866) );
  or2s1 _43987_inst ( .DIN1(_43881), .DIN2(_43882), .Q(_43880) );
  nnd2s1 _43988_inst ( .DIN1(_43883), .DIN2(_43884), .Q(_43879) );
  hi1s1 _43989_inst ( .DIN(_43251), .Q(_43884) );
  nnd2s1 _43990_inst ( .DIN1(_43885), .DIN2(_43886), .Q(_43251) );
  nnd2s1 _43991_inst ( .DIN1(_43639), .DIN2(_26770), .Q(_43885) );
  hi1s1 _43992_inst ( .DIN(_43887), .Q(_43639) );
  nor2s1 _43993_inst ( .DIN1(_43888), .DIN2(_43889), .Q(_43883) );
  nor2s1 _43994_inst ( .DIN1(_43890), .DIN2(_43891), .Q(_43888) );
  nor2s1 _43995_inst ( .DIN1(_43892), .DIN2(_43893), .Q(_43890) );
  nnd2s1 _43996_inst ( .DIN1(_43894), .DIN2(_43895), .Q(
        ____0____________12_____) );
  nnd2s1 _43997_inst ( .DIN1(_43896), .DIN2(_27779), .Q(_43895) );
  nnd2s1 _43998_inst ( .DIN1(_53433), .DIN2(_27780), .Q(_43896) );
  nnd2s1 _43999_inst ( .DIN1(_43897), .DIN2(_38919), .Q(_27780) );
  and2s1 _44000_inst ( .DIN1(_43898), .DIN2(_43899), .Q(_38919) );
  nor2s1 _44001_inst ( .DIN1(_37961), .DIN2(_39461), .Q(_43899) );
  nor2s1 _44002_inst ( .DIN1(_37418), .DIN2(_40867), .Q(_43898) );
  nor2s1 _44003_inst ( .DIN1(_43900), .DIN2(_40868), .Q(_43897) );
  nnd2s1 _44004_inst ( .DIN1(_43901), .DIN2(_27782), .Q(_43894) );
  hi1s1 _44005_inst ( .DIN(_27779), .Q(_27782) );
  nnd2s1 _44006_inst ( .DIN1(_43902), .DIN2(_40866), .Q(_27779) );
  nor2s1 _44007_inst ( .DIN1(_43900), .DIN2(_37961), .Q(_40866) );
  nor2s1 _44008_inst ( .DIN1(_40868), .DIN2(_39456), .Q(_43902) );
  nnd2s1 _44009_inst ( .DIN1(_43903), .DIN2(_37448), .Q(_39456) );
  nor2s1 _44010_inst ( .DIN1(_37417), .DIN2(_39461), .Q(_37448) );
  hi1s1 _44011_inst ( .DIN(_43904), .Q(_39461) );
  nor2s1 _44012_inst ( .DIN1(_40732), .DIN2(_43905), .Q(_43903) );
  hi1s1 _44013_inst ( .DIN(_43906), .Q(_40868) );
  nor2s1 _44014_inst ( .DIN1(_43907), .DIN2(_43908), .Q(_43901) );
  nnd2s1 _44015_inst ( .DIN1(_43909), .DIN2(_43910), .Q(_43908) );
  nor2s1 _44016_inst ( .DIN1(_43911), .DIN2(_43912), .Q(_43910) );
  or2s1 _44017_inst ( .DIN1(_43324), .DIN2(_43285), .Q(_43912) );
  nnd2s1 _44018_inst ( .DIN1(_43913), .DIN2(_43914), .Q(_43285) );
  nnd2s1 _44019_inst ( .DIN1(_43119), .DIN2(_43915), .Q(_43914) );
  nnd2s1 _44020_inst ( .DIN1(_43916), .DIN2(_43396), .Q(_43913) );
  nnd2s1 _44021_inst ( .DIN1(_43917), .DIN2(_43918), .Q(_43324) );
  nnd2s1 _44022_inst ( .DIN1(_43919), .DIN2(_43920), .Q(_43918) );
  nnd2s1 _44023_inst ( .DIN1(_43556), .DIN2(_43921), .Q(_43917) );
  nnd2s1 _44024_inst ( .DIN1(_43922), .DIN2(_43923), .Q(_43911) );
  hi1s1 _44025_inst ( .DIN(_43241), .Q(_43923) );
  nnd2s1 _44026_inst ( .DIN1(_43924), .DIN2(_43925), .Q(_43241) );
  nnd2s1 _44027_inst ( .DIN1(_43926), .DIN2(_43742), .Q(_43925) );
  hi1s1 _44028_inst ( .DIN(_43166), .Q(_43742) );
  nor2s1 _44029_inst ( .DIN1(_43927), .DIN2(_43928), .Q(_43924) );
  nor2s1 _44030_inst ( .DIN1(_43929), .DIN2(_43930), .Q(_43928) );
  hi1s1 _44031_inst ( .DIN(_43338), .Q(_43927) );
  nnd2s1 _44032_inst ( .DIN1(_43844), .DIN2(_43562), .Q(_43338) );
  nor2s1 _44033_inst ( .DIN1(_43836), .DIN2(_43200), .Q(_43922) );
  nnd2s1 _44034_inst ( .DIN1(_43931), .DIN2(_43932), .Q(_43200) );
  nor2s1 _44035_inst ( .DIN1(_43933), .DIN2(_43934), .Q(_43932) );
  nnd2s1 _44036_inst ( .DIN1(_43408), .DIN2(_43855), .Q(_43934) );
  hi1s1 _44037_inst ( .DIN(_43279), .Q(_43408) );
  nor2s1 _44038_inst ( .DIN1(_43252), .DIN2(_43812), .Q(_43279) );
  nor2s1 _44039_inst ( .DIN1(_43233), .DIN2(_43229), .Q(_43933) );
  nor2s1 _44040_inst ( .DIN1(_43935), .DIN2(_43936), .Q(_43931) );
  nnd2s1 _44041_inst ( .DIN1(_43937), .DIN2(_43938), .Q(_43936) );
  nnd2s1 _44042_inst ( .DIN1(_43118), .DIN2(_43939), .Q(_43938) );
  or2s1 _44043_inst ( .DIN1(_43940), .DIN2(_43461), .Q(_43937) );
  nnd2s1 _44044_inst ( .DIN1(_43941), .DIN2(_43942), .Q(_43836) );
  or2s1 _44045_inst ( .DIN1(_43351), .DIN2(_43891), .Q(_43942) );
  nnd2s1 _44046_inst ( .DIN1(_41903), .DIN2(_43336), .Q(_43941) );
  nor2s1 _44047_inst ( .DIN1(_43943), .DIN2(_43944), .Q(_43909) );
  or2s1 _44048_inst ( .DIN1(_43945), .DIN2(_43851), .Q(_43944) );
  nnd2s1 _44049_inst ( .DIN1(_43946), .DIN2(_43571), .Q(_43851) );
  xnr2s1 _44050_inst ( .DIN1(_31975), .DIN2(_43947), .Q(_43571) );
  nor2s1 _44051_inst ( .DIN1(_43864), .DIN2(_43370), .Q(_43947) );
  nnd2s1 _44052_inst ( .DIN1(_43948), .DIN2(_30163), .Q(_31975) );
  nor2s1 _44053_inst ( .DIN1(_43949), .DIN2(_41914), .Q(_43948) );
  nor2s1 _44054_inst ( .DIN1(_43619), .DIN2(_43950), .Q(_43946) );
  nor2s1 _44055_inst ( .DIN1(_43891), .DIN2(_43951), .Q(_43950) );
  nor2s1 _44056_inst ( .DIN1(_43743), .DIN2(_43226), .Q(_43619) );
  nnd2s1 _44057_inst ( .DIN1(_43952), .DIN2(_43953), .Q(_43943) );
  hi1s1 _44058_inst ( .DIN(_43783), .Q(_43953) );
  nnd2s1 _44059_inst ( .DIN1(_43954), .DIN2(_43955), .Q(_43783) );
  nor2s1 _44060_inst ( .DIN1(_43956), .DIN2(_43957), .Q(_43955) );
  nnd2s1 _44061_inst ( .DIN1(_43958), .DIN2(_43959), .Q(_43957) );
  nor2s1 _44062_inst ( .DIN1(_43145), .DIN2(_43249), .Q(_43958) );
  nor2s1 _44063_inst ( .DIN1(_43151), .DIN2(_43658), .Q(_43249) );
  hi1s1 _44064_inst ( .DIN(_43960), .Q(_43145) );
  nnd2s1 _44065_inst ( .DIN1(_43961), .DIN2(_43291), .Q(_43956) );
  nnd2s1 _44066_inst ( .DIN1(_43227), .DIN2(_43396), .Q(_43291) );
  nor2s1 _44067_inst ( .DIN1(_43465), .DIN2(_43624), .Q(_43961) );
  and2s1 _44068_inst ( .DIN1(_43962), .DIN2(_43963), .Q(_43624) );
  nor2s1 _44069_inst ( .DIN1(_43565), .DIN2(_26227), .Q(_43963) );
  nor2s1 _44070_inst ( .DIN1(_43964), .DIN2(_43965), .Q(_43962) );
  and2s1 _44071_inst ( .DIN1(_43966), .DIN2(_26770), .Q(_43465) );
  nor2s1 _44072_inst ( .DIN1(_43967), .DIN2(_43968), .Q(_43954) );
  or2s1 _44073_inst ( .DIN1(_43969), .DIN2(_43970), .Q(_43968) );
  nnd2s1 _44074_inst ( .DIN1(_43971), .DIN2(_43972), .Q(_43967) );
  hi1s1 _44075_inst ( .DIN(_43701), .Q(_43972) );
  nnd2s1 _44076_inst ( .DIN1(_43973), .DIN2(_43974), .Q(_43701) );
  or2s1 _44077_inst ( .DIN1(_43491), .DIN2(_43779), .Q(_43974) );
  nor2s1 _44078_inst ( .DIN1(_43466), .DIN2(_43975), .Q(_43973) );
  nor2s1 _44079_inst ( .DIN1(_43151), .DIN2(_43474), .Q(_43975) );
  and2s1 _44080_inst ( .DIN1(_43976), .DIN2(_43977), .Q(_43466) );
  nor2s1 _44081_inst ( .DIN1(_43512), .DIN2(_43978), .Q(_43976) );
  nor2s1 _44082_inst ( .DIN1(_43979), .DIN2(_43196), .Q(_43971) );
  nnd2s1 _44083_inst ( .DIN1(_43980), .DIN2(_43981), .Q(_43196) );
  nnd2s1 _44084_inst ( .DIN1(_43982), .DIN2(_43414), .Q(_43981) );
  or2s1 _44085_inst ( .DIN1(_43253), .DIN2(_43137), .Q(_43980) );
  nor2s1 _44086_inst ( .DIN1(_43882), .DIN2(_43399), .Q(_43952) );
  nnd2s1 _44087_inst ( .DIN1(_43983), .DIN2(_43984), .Q(_43399) );
  nor2s1 _44088_inst ( .DIN1(_43985), .DIN2(_43986), .Q(_43984) );
  nor2s1 _44089_inst ( .DIN1(_43864), .DIN2(_43987), .Q(_43986) );
  and2s1 _44090_inst ( .DIN1(_43759), .DIN2(_43988), .Q(_43987) );
  nor2s1 _44091_inst ( .DIN1(_43989), .DIN2(_43990), .Q(_43983) );
  nor2s1 _44092_inst ( .DIN1(_43096), .DIN2(_43368), .Q(_43989) );
  nnd2s1 _44093_inst ( .DIN1(_43713), .DIN2(_43991), .Q(_43882) );
  nnd2s1 _44094_inst ( .DIN1(_43992), .DIN2(_29203), .Q(_43991) );
  nor2s1 _44095_inst ( .DIN1(_43473), .DIN2(_43811), .Q(_43992) );
  nnd2s1 _44096_inst ( .DIN1(_43993), .DIN2(_43994), .Q(_43907) );
  nor2s1 _44097_inst ( .DIN1(_43995), .DIN2(_43996), .Q(_43994) );
  nnd2s1 _44098_inst ( .DIN1(_43997), .DIN2(_43998), .Q(_43996) );
  nnd2s1 _44099_inst ( .DIN1(_43515), .DIN2(_43414), .Q(_43998) );
  hi1s1 _44100_inst ( .DIN(_43152), .Q(_43515) );
  nnd2s1 _44101_inst ( .DIN1(_43999), .DIN2(_43977), .Q(_43152) );
  nor2s1 _44102_inst ( .DIN1(_27474), .DIN2(_43804), .Q(_43999) );
  nor2s1 _44103_inst ( .DIN1(_44000), .DIN2(_44001), .Q(_43997) );
  nor2s1 _44104_inst ( .DIN1(_43122), .DIN2(_43167), .Q(_44001) );
  hi1s1 _44105_inst ( .DIN(_43845), .Q(_43167) );
  nnd2s1 _44106_inst ( .DIN1(_44002), .DIN2(_44003), .Q(_43995) );
  nnd2s1 _44107_inst ( .DIN1(_43660), .DIN2(_43186), .Q(_44003) );
  nor2s1 _44108_inst ( .DIN1(_43526), .DIN2(_44004), .Q(_44002) );
  nor2s1 _44109_inst ( .DIN1(_44005), .DIN2(_44006), .Q(_43993) );
  nnd2s1 _44110_inst ( .DIN1(_43093), .DIN2(_44007), .Q(_44006) );
  hi1s1 _44111_inst ( .DIN(_43588), .Q(_44007) );
  xor2s1 _44112_inst ( .DIN1(_32753), .DIN2(_44008), .Q(_43093) );
  nor2s1 _44113_inst ( .DIN1(_44009), .DIN2(_44010), .Q(_44008) );
  nnd2s1 _44114_inst ( .DIN1(_44011), .DIN2(_44012), .Q(_44010) );
  nor2s1 _44115_inst ( .DIN1(_44013), .DIN2(_44014), .Q(_44012) );
  nor2s1 _44116_inst ( .DIN1(_43230), .DIN2(_43226), .Q(_44014) );
  nor2s1 _44117_inst ( .DIN1(_43514), .DIN2(_44015), .Q(_44013) );
  nor2s1 _44118_inst ( .DIN1(_43538), .DIN2(_43245), .Q(_44011) );
  nnd2s1 _44119_inst ( .DIN1(_44016), .DIN2(_44017), .Q(_43245) );
  nnd2s1 _44120_inst ( .DIN1(_44018), .DIN2(_43414), .Q(_44017) );
  or2s1 _44121_inst ( .DIN1(_43664), .DIN2(_43545), .Q(_44016) );
  nor2s1 _44122_inst ( .DIN1(_43252), .DIN2(_43272), .Q(_43538) );
  nnd2s1 _44123_inst ( .DIN1(_44019), .DIN2(_44020), .Q(_44009) );
  nor2s1 _44124_inst ( .DIN1(_44021), .DIN2(_43147), .Q(_44020) );
  nor2s1 _44125_inst ( .DIN1(_44022), .DIN2(_44023), .Q(_44019) );
  nor2s1 _44126_inst ( .DIN1(_43151), .DIN2(_44024), .Q(_44023) );
  nor2s1 _44127_inst ( .DIN1(_43350), .DIN2(_43520), .Q(_44022) );
  nor2s1 _44128_inst ( .DIN1(_44025), .DIN2(_44026), .Q(_43350) );
  nnd2s1 _44129_inst ( .DIN1(_44027), .DIN2(_44028), .Q(_32753) );
  nor2s1 _44130_inst ( .DIN1(_44029), .DIN2(_44030), .Q(_44028) );
  nor2s1 _44131_inst ( .DIN1(_44031), .DIN2(_44032), .Q(_44027) );
  nnd2s1 _44132_inst ( .DIN1(_44033), .DIN2(_44034), .Q(_44005) );
  nnd2s1 _44133_inst ( .DIN1(_43686), .DIN2(_43939), .Q(_44034) );
  hi1s1 _44134_inst ( .DIN(_43548), .Q(_43686) );
  nor2s1 _44135_inst ( .DIN1(_43483), .DIN2(_44035), .Q(_44033) );
  nor2s1 _44136_inst ( .DIN1(_43473), .DIN2(_43475), .Q(_44035) );
  nor2s1 _44137_inst ( .DIN1(_43490), .DIN2(_43780), .Q(_43483) );
  nnd2s1 _44138_inst ( .DIN1(_44036), .DIN2(_43171), .Q(
        ____0____________11_____) );
  nor2s1 _44139_inst ( .DIN1(_44037), .DIN2(_44038), .Q(_44036) );
  nor2s1 _44140_inst ( .DIN1(_43174), .DIN2(_44039), .Q(_44038) );
  nnd2s1 _44141_inst ( .DIN1(_44040), .DIN2(_44041), .Q(_44039) );
  nor2s1 _44142_inst ( .DIN1(_44042), .DIN2(_44043), .Q(_44041) );
  nnd2s1 _44143_inst ( .DIN1(_44044), .DIN2(_44045), .Q(_44043) );
  nor2s1 _44144_inst ( .DIN1(_43769), .DIN2(_43317), .Q(_44045) );
  and2s1 _44145_inst ( .DIN1(_44046), .DIN2(_44047), .Q(_43317) );
  hi1s1 _44146_inst ( .DIN(_43334), .Q(_43769) );
  nnd2s1 _44147_inst ( .DIN1(_43921), .DIN2(_43723), .Q(_43334) );
  hi1s1 _44148_inst ( .DIN(_43226), .Q(_43921) );
  nor2s1 _44149_inst ( .DIN1(_44048), .DIN2(_44049), .Q(_44044) );
  nor2s1 _44150_inst ( .DIN1(_43779), .DIN2(_43620), .Q(_44049) );
  nnd2s1 _44151_inst ( .DIN1(_44050), .DIN2(_44051), .Q(_43620) );
  nor2s1 _44152_inst ( .DIN1(_43978), .DIN2(_44052), .Q(_44050) );
  nnd2s1 _44153_inst ( .DIN1(_44053), .DIN2(_44054), .Q(_44042) );
  nor2s1 _44154_inst ( .DIN1(_43985), .DIN2(_43834), .Q(_44054) );
  and2s1 _44155_inst ( .DIN1(_44055), .DIN2(_43567), .Q(_43834) );
  hi1s1 _44156_inst ( .DIN(_43781), .Q(_43567) );
  nnd2s1 _44157_inst ( .DIN1(_43808), .DIN2(_44056), .Q(_43781) );
  nor2s1 _44158_inst ( .DIN1(_43151), .DIN2(_43964), .Q(_44055) );
  and2s1 _44159_inst ( .DIN1(_44057), .DIN2(_44058), .Q(_43985) );
  nor2s1 _44160_inst ( .DIN1(_27349), .DIN2(_43514), .Q(_44057) );
  nor2s1 _44161_inst ( .DIN1(_43670), .DIN2(_43842), .Q(_44053) );
  nor2s1 _44162_inst ( .DIN1(_43234), .DIN2(_43565), .Q(_43842) );
  nnd2s1 _44163_inst ( .DIN1(_43568), .DIN2(_44059), .Q(_43234) );
  nor2s1 _44164_inst ( .DIN1(_26227), .DIN2(_43965), .Q(_43568) );
  nor2s1 _44165_inst ( .DIN1(_44060), .DIN2(_44061), .Q(_44040) );
  nnd2s1 _44166_inst ( .DIN1(_44062), .DIN2(_44063), .Q(_44061) );
  nor2s1 _44167_inst ( .DIN1(_43242), .DIN2(_43357), .Q(_44063) );
  nnd2s1 _44168_inst ( .DIN1(_44064), .DIN2(_44065), .Q(_43357) );
  nor2s1 _44169_inst ( .DIN1(_44066), .DIN2(_44067), .Q(_44065) );
  nnd2s1 _44170_inst ( .DIN1(_43959), .DIN2(_44068), .Q(_44067) );
  hi1s1 _44171_inst ( .DIN(_43679), .Q(_44068) );
  nnd2s1 _44172_inst ( .DIN1(_43892), .DIN2(_43790), .Q(_43959) );
  nor2s1 _44173_inst ( .DIN1(_43096), .DIN2(_43558), .Q(_44066) );
  nor2s1 _44174_inst ( .DIN1(_43578), .DIN2(_44069), .Q(_44064) );
  xor2s1 _44175_inst ( .DIN1(_44070), .DIN2(_44071), .Q(_44069) );
  nor2s1 _44176_inst ( .DIN1(_44072), .DIN2(_43112), .Q(_44071) );
  nor2s1 _44177_inst ( .DIN1(_43189), .DIN2(_43864), .Q(_43112) );
  nor2s1 _44178_inst ( .DIN1(_43435), .DIN2(_44073), .Q(_44072) );
  nnd2s1 _44179_inst ( .DIN1(_44074), .DIN2(_43617), .Q(_43578) );
  nnd2s1 _44180_inst ( .DIN1(_43926), .DIN2(_44047), .Q(_43617) );
  hi1s1 _44181_inst ( .DIN(_44075), .Q(_43926) );
  xor2s1 _44182_inst ( .DIN1(_43439), .DIN2(_37195), .Q(_44074) );
  nnd2s1 _44183_inst ( .DIN1(_44076), .DIN2(_44077), .Q(_37195) );
  and2s1 _44184_inst ( .DIN1(_44078), .DIN2(_44079), .Q(_44076) );
  nnd2s1 _44185_inst ( .DIN1(_41903), .DIN2(_43396), .Q(_43439) );
  nnd2s1 _44186_inst ( .DIN1(_44080), .DIN2(_44081), .Q(_43242) );
  nor2s1 _44187_inst ( .DIN1(_44082), .DIN2(_44083), .Q(_44081) );
  nnd2s1 _44188_inst ( .DIN1(_44084), .DIN2(_43091), .Q(_44083) );
  nor2s1 _44189_inst ( .DIN1(_43889), .DIN2(_43319), .Q(_44084) );
  nor2s1 _44190_inst ( .DIN1(_43151), .DIN2(_43110), .Q(_43319) );
  nor2s1 _44191_inst ( .DIN1(_43780), .DIN2(_43621), .Q(_43889) );
  nnd2s1 _44192_inst ( .DIN1(_44085), .DIN2(_44086), .Q(_43780) );
  nnd2s1 _44193_inst ( .DIN1(_44087), .DIN2(_44088), .Q(_44082) );
  hi1s1 _44194_inst ( .DIN(_43190), .Q(_44088) );
  nor2s1 _44195_inst ( .DIN1(_44089), .DIN2(_43354), .Q(_44087) );
  nor2s1 _44196_inst ( .DIN1(_43415), .DIN2(_43233), .Q(_43354) );
  nor2s1 _44197_inst ( .DIN1(_44090), .DIN2(_44091), .Q(_44080) );
  or2s1 _44198_inst ( .DIN1(_44092), .DIN2(_43838), .Q(_44091) );
  nnd2s1 _44199_inst ( .DIN1(_44093), .DIN2(_44094), .Q(_43838) );
  nor2s1 _44200_inst ( .DIN1(_44095), .DIN2(_44096), .Q(_44094) );
  nor2s1 _44201_inst ( .DIN1(_43514), .DIN2(_43474), .Q(_44096) );
  nnd2s1 _44202_inst ( .DIN1(_44097), .DIN2(_43977), .Q(_43474) );
  nor2s1 _44203_inst ( .DIN1(_44098), .DIN2(_44099), .Q(_44097) );
  nor2s1 _44204_inst ( .DIN1(_43816), .DIN2(_43226), .Q(_44095) );
  nnd2s1 _44205_inst ( .DIN1(_44100), .DIN2(_44059), .Q(_43816) );
  nor2s1 _44206_inst ( .DIN1(_44101), .DIN2(_43804), .Q(_44059) );
  nor2s1 _44207_inst ( .DIN1(_44102), .DIN2(_44103), .Q(_44100) );
  nor2s1 _44208_inst ( .DIN1(_44104), .DIN2(_43477), .Q(_44093) );
  nnd2s1 _44209_inst ( .DIN1(_44105), .DIN2(_44106), .Q(_43477) );
  nnd2s1 _44210_inst ( .DIN1(_43574), .DIN2(_44107), .Q(_44106) );
  nnd2s1 _44211_inst ( .DIN1(_44108), .DIN2(_44109), .Q(_44107) );
  nnd2s1 _44212_inst ( .DIN1(_43977), .DIN2(_44110), .Q(_44109) );
  nnd2s1 _44213_inst ( .DIN1(_43573), .DIN2(_43707), .Q(_44105) );
  hi1s1 _44214_inst ( .DIN(_44108), .Q(_43573) );
  nnd2s1 _44215_inst ( .DIN1(_44111), .DIN2(_44085), .Q(_44108) );
  and2s1 _44216_inst ( .DIN1(_44112), .DIN2(_44113), .Q(_44085) );
  nor2s1 _44217_inst ( .DIN1(_53448), .DIN2(_27374), .Q(_44112) );
  nor2s1 _44218_inst ( .DIN1(_53457), .DIN2(_44114), .Q(_44111) );
  nor2s1 _44219_inst ( .DIN1(_43491), .DIN2(_43621), .Q(_44104) );
  nnd2s1 _44220_inst ( .DIN1(_44115), .DIN2(_44116), .Q(_44090) );
  hi1s1 _44221_inst ( .DIN(_43295), .Q(_44116) );
  nnd2s1 _44222_inst ( .DIN1(_44117), .DIN2(_44118), .Q(_43295) );
  nor2s1 _44223_inst ( .DIN1(_43770), .DIN2(_44119), .Q(_44118) );
  nor2s1 _44224_inst ( .DIN1(_43121), .DIN2(_43120), .Q(_44119) );
  nor2s1 _44225_inst ( .DIN1(_43473), .DIN2(_44015), .Q(_43770) );
  nor2s1 _44226_inst ( .DIN1(_43476), .DIN2(_44120), .Q(_44117) );
  xor2s1 _44227_inst ( .DIN1(_32716), .DIN2(_44121), .Q(_44120) );
  nnd2s1 _44228_inst ( .DIN1(_44122), .DIN2(_44123), .Q(_44121) );
  hi1s1 _44229_inst ( .DIN(_43877), .Q(_44123) );
  nor2s1 _44230_inst ( .DIN1(_43475), .DIN2(_43151), .Q(_43877) );
  nnd2s1 _44231_inst ( .DIN1(_44124), .DIN2(_44125), .Q(_43475) );
  nor2s1 _44232_inst ( .DIN1(_44126), .DIN2(_43148), .Q(_44122) );
  hi1s1 _44233_inst ( .DIN(_43406), .Q(_43148) );
  nnd2s1 _44234_inst ( .DIN1(_43704), .DIN2(_43920), .Q(_43406) );
  hi1s1 _44235_inst ( .DIN(_43462), .Q(_43704) );
  nnd2s1 _44236_inst ( .DIN1(_44127), .DIN2(_44128), .Q(_43462) );
  nor2s1 _44237_inst ( .DIN1(_27475), .DIN2(_44129), .Q(_44128) );
  nnd2s1 _44238_inst ( .DIN1(_44130), .DIN2(_26227), .Q(_44129) );
  nor2s1 _44239_inst ( .DIN1(_44131), .DIN2(_44132), .Q(_44127) );
  nnd2s1 _44240_inst ( .DIN1(_44056), .DIN2(_44133), .Q(_44132) );
  nnd2s1 _44241_inst ( .DIN1(_44134), .DIN2(_44135), .Q(_43476) );
  xor2s1 _44242_inst ( .DIN1(_27413), .DIN2(_44136), .Q(_44135) );
  nnd2s1 _44243_inst ( .DIN1(_43741), .DIN2(_26770), .Q(_44136) );
  hi1s1 _44244_inst ( .DIN(_43594), .Q(_43741) );
  nnd2s1 _44245_inst ( .DIN1(_44137), .DIN2(_44138), .Q(_43594) );
  nor2s1 _44246_inst ( .DIN1(_44139), .DIN2(_44140), .Q(_44138) );
  or2s1 _44247_inst ( .DIN1(_43804), .DIN2(_27474), .Q(_44140) );
  nor2s1 _44248_inst ( .DIN1(_44131), .DIN2(_44141), .Q(_44137) );
  nnd2s1 _44249_inst ( .DIN1(_53448), .DIN2(_44056), .Q(_44141) );
  hi1s1 _44250_inst ( .DIN(_43409), .Q(_44134) );
  nnd2s1 _44251_inst ( .DIN1(_44142), .DIN2(_44143), .Q(_43409) );
  nnd2s1 _44252_inst ( .DIN1(_44144), .DIN2(_43336), .Q(_44143) );
  nnd2s1 _44253_inst ( .DIN1(_44145), .DIN2(_26770), .Q(_44142) );
  nor2s1 _44254_inst ( .DIN1(_43339), .DIN2(_43549), .Q(_44115) );
  nnd2s1 _44255_inst ( .DIN1(_44146), .DIN2(_44147), .Q(_43549) );
  hi1s1 _44256_inst ( .DIN(_44148), .Q(_44147) );
  nor2s1 _44257_inst ( .DIN1(_44149), .DIN2(_44150), .Q(_44146) );
  nor2s1 _44258_inst ( .DIN1(_43461), .DIN2(_43940), .Q(_44150) );
  hi1s1 _44259_inst ( .DIN(_44151), .Q(_44149) );
  nnd2s1 _44260_inst ( .DIN1(_44152), .DIN2(_44153), .Q(_43339) );
  nor2s1 _44261_inst ( .DIN1(_43113), .DIN2(_44004), .Q(_44153) );
  hi1s1 _44262_inst ( .DIN(_44154), .Q(_44004) );
  nor2s1 _44263_inst ( .DIN1(_44155), .DIN2(_44156), .Q(_44152) );
  nor2s1 _44264_inst ( .DIN1(_43520), .DIN2(_44157), .Q(_44156) );
  nor2s1 _44265_inst ( .DIN1(_43137), .DIN2(_43095), .Q(_44155) );
  nor2s1 _44266_inst ( .DIN1(_44158), .DIN2(_44159), .Q(_44062) );
  hi1s1 _44267_inst ( .DIN(_43283), .Q(_44158) );
  nor2s1 _44268_inst ( .DIN1(_44160), .DIN2(_43630), .Q(_43283) );
  nnd2s1 _44269_inst ( .DIN1(_44161), .DIN2(_44162), .Q(_43630) );
  nnd2s1 _44270_inst ( .DIN1(_43556), .DIN2(_43396), .Q(_44162) );
  nor2s1 _44271_inst ( .DIN1(_44021), .DIN2(_43107), .Q(_44161) );
  nor2s1 _44272_inst ( .DIN1(_43520), .DIN2(_43988), .Q(_43107) );
  or2s1 _44273_inst ( .DIN1(_43524), .DIN2(_44163), .Q(_44160) );
  nor2s1 _44274_inst ( .DIN1(_43891), .DIN2(_43796), .Q(_44163) );
  nnd2s1 _44275_inst ( .DIN1(_44164), .DIN2(_44165), .Q(_44060) );
  nor2s1 _44276_inst ( .DIN1(_44166), .DIN2(_44167), .Q(_44165) );
  nor2s1 _44277_inst ( .DIN1(_43891), .DIN2(_44168), .Q(_44167) );
  nor2s1 _44278_inst ( .DIN1(_43197), .DIN2(_43858), .Q(_44164) );
  xor2s1 _44279_inst ( .DIN1(_44169), .DIN2(_34151), .Q(_43858) );
  nnd2s1 _44280_inst ( .DIN1(_44170), .DIN2(_44171), .Q(_44169) );
  nnd2s1 _44281_inst ( .DIN1(_43707), .DIN2(_43966), .Q(_44171) );
  and2s1 _44282_inst ( .DIN1(_44172), .DIN2(_44173), .Q(_43966) );
  nor2s1 _44283_inst ( .DIN1(_27474), .DIN2(_44174), .Q(_44173) );
  or2s1 _44284_inst ( .DIN1(_44175), .DIN2(_53448), .Q(_44174) );
  nor2s1 _44285_inst ( .DIN1(_26353), .DIN2(_44114), .Q(_44172) );
  hi1s1 _44286_inst ( .DIN(_43512), .Q(_43707) );
  nnd2s1 _44287_inst ( .DIN1(_43395), .DIN2(_43336), .Q(_44170) );
  nor2s1 _44288_inst ( .DIN1(_44176), .DIN2(_44052), .Q(_43395) );
  or2s1 _44289_inst ( .DIN1(_44114), .DIN2(_43978), .Q(_44176) );
  nnd2s1 _44290_inst ( .DIN1(_44177), .DIN2(_44178), .Q(_43197) );
  nor2s1 _44291_inst ( .DIN1(_44179), .DIN2(_44180), .Q(_44178) );
  nnd2s1 _44292_inst ( .DIN1(_43631), .DIN2(_43342), .Q(_44180) );
  nnd2s1 _44293_inst ( .DIN1(_43414), .DIN2(_44181), .Q(_43342) );
  and2s1 _44294_inst ( .DIN1(_44182), .DIN2(_44183), .Q(_43631) );
  nnd2s1 _44295_inst ( .DIN1(_44184), .DIN2(_43108), .Q(_44183) );
  nnd2s1 _44296_inst ( .DIN1(_43713), .DIN2(_44185), .Q(_44179) );
  hi1s1 _44297_inst ( .DIN(_43440), .Q(_43713) );
  nor2s1 _44298_inst ( .DIN1(_44186), .DIN2(_43891), .Q(_43440) );
  nor2s1 _44299_inst ( .DIN1(_44187), .DIN2(_44188), .Q(_44177) );
  or2s1 _44300_inst ( .DIN1(_43979), .DIN2(_43837), .Q(_44188) );
  nnd2s1 _44301_inst ( .DIN1(_44189), .DIN2(_44190), .Q(_43837) );
  nor2s1 _44302_inst ( .DIN1(_43278), .DIN2(_44191), .Q(_44190) );
  nor2s1 _44303_inst ( .DIN1(_43151), .DIN2(_43111), .Q(_44191) );
  nor2s1 _44304_inst ( .DIN1(_43930), .DIN2(_43121), .Q(_43278) );
  nor2s1 _44305_inst ( .DIN1(_43587), .DIN2(_43451), .Q(_44189) );
  nnd2s1 _44306_inst ( .DIN1(_44192), .DIN2(_44193), .Q(_43451) );
  nnd2s1 _44307_inst ( .DIN1(_44026), .DIN2(_43186), .Q(_44193) );
  nnd2s1 _44308_inst ( .DIN1(_43751), .DIN2(_43119), .Q(_44192) );
  hi1s1 _44309_inst ( .DIN(_43137), .Q(_43119) );
  hi1s1 _44310_inst ( .DIN(_43272), .Q(_43751) );
  nor2s1 _44311_inst ( .DIN1(_43441), .DIN2(_43226), .Q(_43587) );
  or2s1 _44312_inst ( .DIN1(_44194), .DIN2(_43700), .Q(_44187) );
  nnd2s1 _44313_inst ( .DIN1(_44195), .DIN2(_44196), .Q(_43700) );
  nnd2s1 _44314_inst ( .DIN1(_43815), .DIN2(_43919), .Q(_44196) );
  nnd2s1 _44315_inst ( .DIN1(_43335), .DIN2(_43396), .Q(_44195) );
  hi1s1 _44316_inst ( .DIN(_43233), .Q(_43396) );
  nor2s1 _44317_inst ( .DIN1(_43203), .DIN2(_44197), .Q(_44037) );
  nor2s1 _44318_inst ( .DIN1(_27241), .DIN2(_26243), .Q(_44197) );
  nnd2s1 _44319_inst ( .DIN1(_44198), .DIN2(_44199), .Q(
        ____0____________10_____) );
  nnd2s1 _44320_inst ( .DIN1(_44200), .DIN2(_53434), .Q(_44199) );
  nor2s1 _44321_inst ( .DIN1(_32183), .DIN2(_27241), .Q(_44200) );
  hi1s1 _44322_inst ( .DIN(_41984), .Q(_32183) );
  nnd2s1 _44323_inst ( .DIN1(_44201), .DIN2(_44202), .Q(_41984) );
  nor2s1 _44324_inst ( .DIN1(_38884), .DIN2(_39740), .Q(_44201) );
  nnd2s1 _44325_inst ( .DIN1(_28056), .DIN2(_44203), .Q(_44198) );
  nnd2s1 _44326_inst ( .DIN1(_44204), .DIN2(_44205), .Q(_44203) );
  nor2s1 _44327_inst ( .DIN1(_44206), .DIN2(_44207), .Q(_44205) );
  nnd2s1 _44328_inst ( .DIN1(_44208), .DIN2(_44209), .Q(_44207) );
  nor2s1 _44329_inst ( .DIN1(_44210), .DIN2(_44166), .Q(_44209) );
  nor2s1 _44330_inst ( .DIN1(_43139), .DIN2(_43800), .Q(_44166) );
  nnd2s1 _44331_inst ( .DIN1(_44211), .DIN2(_44086), .Q(_43800) );
  hi1s1 _44332_inst ( .DIN(_43965), .Q(_44086) );
  nnd2s1 _44333_inst ( .DIN1(_44212), .DIN2(_44213), .Q(_43965) );
  nor2s1 _44334_inst ( .DIN1(_44214), .DIN2(_44215), .Q(_44213) );
  nnd2s1 _44335_inst ( .DIN1(_26428), .DIN2(_26207), .Q(_44215) );
  nor2s1 _44336_inst ( .DIN1(_26624), .DIN2(_44216), .Q(_44212) );
  nnd2s1 _44337_inst ( .DIN1(_44217), .DIN2(_44218), .Q(_44216) );
  nor2s1 _44338_inst ( .DIN1(_53448), .DIN2(_43978), .Q(_44211) );
  hi1s1 _44339_inst ( .DIN(_44110), .Q(_43978) );
  nor2s1 _44340_inst ( .DIN1(_43804), .DIN2(_44099), .Q(_44110) );
  nor2s1 _44341_inst ( .DIN1(_44219), .DIN2(_43233), .Q(_44210) );
  nor2s1 _44342_inst ( .DIN1(_44144), .DIN2(_43723), .Q(_44219) );
  hi1s1 _44343_inst ( .DIN(_43743), .Q(_44144) );
  nnd2s1 _44344_inst ( .DIN1(_44220), .DIN2(_44051), .Q(_43743) );
  nor2s1 _44345_inst ( .DIN1(_43964), .DIN2(_44052), .Q(_44220) );
  nor2s1 _44346_inst ( .DIN1(_44221), .DIN2(_44222), .Q(_44208) );
  nor2s1 _44347_inst ( .DIN1(_43166), .DIN2(_43123), .Q(_44222) );
  nor2s1 _44348_inst ( .DIN1(_43812), .DIN2(_43137), .Q(_44221) );
  nnd2s1 _44349_inst ( .DIN1(_44223), .DIN2(_44224), .Q(_43812) );
  nor2s1 _44350_inst ( .DIN1(_44214), .DIN2(_44225), .Q(_44224) );
  nnd2s1 _44351_inst ( .DIN1(_26227), .DIN2(_26207), .Q(_44225) );
  nor2s1 _44352_inst ( .DIN1(_43964), .DIN2(_44226), .Q(_44223) );
  nnd2s1 _44353_inst ( .DIN1(_44227), .DIN2(_43807), .Q(_44226) );
  nnd2s1 _44354_inst ( .DIN1(_44228), .DIN2(_44229), .Q(_44206) );
  nor2s1 _44355_inst ( .DIN1(_43316), .DIN2(_44230), .Q(_44229) );
  nnd2s1 _44356_inst ( .DIN1(_44231), .DIN2(_43277), .Q(_44230) );
  nnd2s1 _44357_inst ( .DIN1(_43920), .DIN2(_43856), .Q(_43277) );
  hi1s1 _44358_inst ( .DIN(_43121), .Q(_43920) );
  nor2s1 _44359_inst ( .DIN1(_43690), .DIN2(_43679), .Q(_44228) );
  nor2s1 _44360_inst ( .DIN1(_43559), .DIN2(_43514), .Q(_43679) );
  nor2s1 _44361_inst ( .DIN1(_44232), .DIN2(_44233), .Q(_44204) );
  nnd2s1 _44362_inst ( .DIN1(_44234), .DIN2(_44235), .Q(_44233) );
  nor2s1 _44363_inst ( .DIN1(_43535), .DIN2(_43784), .Q(_44235) );
  nnd2s1 _44364_inst ( .DIN1(_44236), .DIN2(_44237), .Q(_43784) );
  nnd2s1 _44365_inst ( .DIN1(_43725), .DIN2(_44238), .Q(_44237) );
  nnd2s1 _44366_inst ( .DIN1(_43189), .DIN2(_43988), .Q(_44238) );
  nor2s1 _44367_inst ( .DIN1(_43672), .DIN2(_44239), .Q(_44236) );
  nor2s1 _44368_inst ( .DIN1(_44240), .DIN2(_43520), .Q(_44239) );
  nor2s1 _44369_inst ( .DIN1(_44145), .DIN2(_43724), .Q(_44240) );
  hi1s1 _44370_inst ( .DIN(_43951), .Q(_44145) );
  nnd2s1 _44371_inst ( .DIN1(_44241), .DIN2(_44242), .Q(_43951) );
  nor2s1 _44372_inst ( .DIN1(_53457), .DIN2(_44101), .Q(_44241) );
  nnd2s1 _44373_inst ( .DIN1(_44243), .DIN2(_44244), .Q(_43535) );
  nor2s1 _44374_inst ( .DIN1(_43275), .DIN2(_44245), .Q(_44244) );
  nor2s1 _44375_inst ( .DIN1(_43229), .DIN2(_43226), .Q(_44245) );
  nnd2s1 _44376_inst ( .DIN1(_44246), .DIN2(_43808), .Q(_43229) );
  hi1s1 _44377_inst ( .DIN(_44103), .Q(_43808) );
  nnd2s1 _44378_inst ( .DIN1(_44247), .DIN2(_44248), .Q(_44103) );
  nor2s1 _44379_inst ( .DIN1(_53448), .DIN2(_44139), .Q(_44247) );
  nor2s1 _44380_inst ( .DIN1(_44102), .DIN2(_43964), .Q(_44246) );
  nor2s1 _44381_inst ( .DIN1(_44249), .DIN2(_44250), .Q(_44243) );
  nor2s1 _44382_inst ( .DIN1(_43252), .DIN2(_43369), .Q(_44250) );
  nor2s1 _44383_inst ( .DIN1(_43779), .DIN2(_43491), .Q(_44249) );
  nnd2s1 _44384_inst ( .DIN1(_44251), .DIN2(_44242), .Q(_43491) );
  and2s1 _44385_inst ( .DIN1(_44252), .DIN2(_44051), .Q(_44242) );
  hi1s1 _44386_inst ( .DIN(_44253), .Q(_44051) );
  nor2s1 _44387_inst ( .DIN1(_53448), .DIN2(_43804), .Q(_44252) );
  nor2s1 _44388_inst ( .DIN1(_27474), .DIN2(_26353), .Q(_44251) );
  nor2s1 _44389_inst ( .DIN1(_43850), .DIN2(_43945), .Q(_44234) );
  nnd2s1 _44390_inst ( .DIN1(_44254), .DIN2(_44255), .Q(_43945) );
  nor2s1 _44391_inst ( .DIN1(_44048), .DIN2(_44256), .Q(_44254) );
  nor2s1 _44392_inst ( .DIN1(_43121), .DIN2(_44073), .Q(_44256) );
  nor2s1 _44393_inst ( .DIN1(_43887), .DIN2(_43514), .Q(_44048) );
  nnd2s1 _44394_inst ( .DIN1(_44257), .DIN2(_44258), .Q(_43850) );
  nor2s1 _44395_inst ( .DIN1(_44259), .DIN2(_44260), .Q(_44258) );
  nnd2s1 _44396_inst ( .DIN1(_44261), .DIN2(_43756), .Q(_44260) );
  nnd2s1 _44397_inst ( .DIN1(_44262), .DIN2(_43705), .Q(_43756) );
  or2s1 _44398_inst ( .DIN1(_26825), .DIN2(_44263), .Q(_44261) );
  nnd2s1 _44399_inst ( .DIN1(_44151), .DIN2(_44264), .Q(_44259) );
  nor2s1 _44400_inst ( .DIN1(_43448), .DIN2(_44265), .Q(_44257) );
  nnd2s1 _44401_inst ( .DIN1(_44266), .DIN2(_44267), .Q(_44265) );
  nnd2s1 _44402_inst ( .DIN1(_44018), .DIN2(_43108), .Q(_44267) );
  nnd2s1 _44403_inst ( .DIN1(_44268), .DIN2(_43939), .Q(_44266) );
  nnd2s1 _44404_inst ( .DIN1(_44269), .DIN2(_44270), .Q(_43448) );
  nor2s1 _44405_inst ( .DIN1(_44271), .DIN2(_44272), .Q(_44270) );
  nor2s1 _44406_inst ( .DIN1(_43137), .DIN2(_43548), .Q(_44272) );
  nor2s1 _44407_inst ( .DIN1(_43514), .DIN2(_44024), .Q(_44271) );
  hi1s1 _44408_inst ( .DIN(_44184), .Q(_44024) );
  nor2s1 _44409_inst ( .DIN1(_43588), .DIN2(_44148), .Q(_44269) );
  nnd2s1 _44410_inst ( .DIN1(_44273), .DIN2(_44274), .Q(_44148) );
  nnd2s1 _44411_inst ( .DIN1(_43747), .DIN2(_43939), .Q(_44274) );
  hi1s1 _44412_inst ( .DIN(_43153), .Q(_43747) );
  nnd2s1 _44413_inst ( .DIN1(_43977), .DIN2(_43564), .Q(_43153) );
  hi1s1 _44414_inst ( .DIN(_43964), .Q(_43564) );
  nnd2s1 _44415_inst ( .DIN1(_44113), .DIN2(_44130), .Q(_43964) );
  nor2s1 _44416_inst ( .DIN1(_43127), .DIN2(_44114), .Q(_43977) );
  nnd2s1 _44417_inst ( .DIN1(_43776), .DIN2(_43574), .Q(_44273) );
  hi1s1 _44418_inst ( .DIN(_43140), .Q(_43776) );
  nnd2s1 _44419_inst ( .DIN1(_44275), .DIN2(_44125), .Q(_43140) );
  nor2s1 _44420_inst ( .DIN1(_44175), .DIN2(_27474), .Q(_44125) );
  nor2s1 _44421_inst ( .DIN1(_43127), .DIN2(_44253), .Q(_44275) );
  nnd2s1 _44422_inst ( .DIN1(_44276), .DIN2(_44277), .Q(_44253) );
  nor2s1 _44423_inst ( .DIN1(_44139), .DIN2(_44278), .Q(_44277) );
  nnd2s1 _44424_inst ( .DIN1(_53449), .DIN2(_26207), .Q(_44278) );
  nor2s1 _44425_inst ( .DIN1(_26345), .DIN2(_44279), .Q(_44276) );
  nnd2s1 _44426_inst ( .DIN1(_53448), .DIN2(_53457), .Q(_43127) );
  xor2s1 _44427_inst ( .DIN1(_31842), .DIN2(_44280), .Q(_43588) );
  nor2s1 _44428_inst ( .DIN1(_43520), .DIN2(_44168), .Q(_44280) );
  nnd2s1 _44429_inst ( .DIN1(_44281), .DIN2(_44282), .Q(_31842) );
  nor2s1 _44430_inst ( .DIN1(_44283), .DIN2(_42925), .Q(_44281) );
  nnd2s1 _44431_inst ( .DIN1(_44284), .DIN2(_44285), .Q(_42925) );
  nor2s1 _44432_inst ( .DIN1(_44286), .DIN2(_42796), .Q(_44285) );
  nor2s1 _44433_inst ( .DIN1(_44287), .DIN2(_44288), .Q(_44284) );
  nnd2s1 _44434_inst ( .DIN1(_44289), .DIN2(_44290), .Q(_44232) );
  nor2s1 _44435_inst ( .DIN1(_43698), .DIN2(_43097), .Q(_44290) );
  nnd2s1 _44436_inst ( .DIN1(_44291), .DIN2(_44292), .Q(_43097) );
  nnd2s1 _44437_inst ( .DIN1(_43108), .DIN2(_44181), .Q(_44292) );
  hi1s1 _44438_inst ( .DIN(_44293), .Q(_44181) );
  nor2s1 _44439_inst ( .DIN1(_44294), .DIN2(_43641), .Q(_44291) );
  nor2s1 _44440_inst ( .DIN1(_43940), .DIN2(_43121), .Q(_43641) );
  nor2s1 _44441_inst ( .DIN1(_44295), .DIN2(_43166), .Q(_44294) );
  nor2s1 _44442_inst ( .DIN1(_43585), .DIN2(_43845), .Q(_44295) );
  hi1s1 _44443_inst ( .DIN(_43313), .Q(_43585) );
  nor2s1 _44444_inst ( .DIN1(_43252), .DIN2(_43095), .Q(_43698) );
  nor2s1 _44445_inst ( .DIN1(_43358), .DIN2(_43384), .Q(_44289) );
  nnd2s1 _44446_inst ( .DIN1(_44296), .DIN2(_43861), .Q(_43384) );
  nor2s1 _44447_inst ( .DIN1(_44297), .DIN2(_43653), .Q(_43861) );
  nor2s1 _44448_inst ( .DIN1(_43435), .DIN2(_43120), .Q(_43653) );
  nor2s1 _44449_inst ( .DIN1(_44298), .DIN2(_44092), .Q(_44296) );
  nnd2s1 _44450_inst ( .DIN1(_44299), .DIN2(_44300), .Q(_44092) );
  nnd2s1 _44451_inst ( .DIN1(_43748), .DIN2(_43939), .Q(_44300) );
  hi1s1 _44452_inst ( .DIN(_43138), .Q(_43748) );
  nnd2s1 _44453_inst ( .DIN1(_44124), .DIN2(_44301), .Q(_43138) );
  nor2s1 _44454_inst ( .DIN1(_44101), .DIN2(_27475), .Q(_44301) );
  nor2s1 _44455_inst ( .DIN1(_44114), .DIN2(_44052), .Q(_44124) );
  nnd2s1 _44456_inst ( .DIN1(_53448), .DIN2(_26353), .Q(_44052) );
  nnd2s1 _44457_inst ( .DIN1(_44302), .DIN2(_44248), .Q(_44114) );
  hi1s1 _44458_inst ( .DIN(_44131), .Q(_44248) );
  nnd2s1 _44459_inst ( .DIN1(_44303), .DIN2(_44227), .Q(_44131) );
  hi1s1 _44460_inst ( .DIN(_44279), .Q(_44227) );
  nnd2s1 _44461_inst ( .DIN1(_44304), .DIN2(_43420), .Q(_44279) );
  nor2s1 _44462_inst ( .DIN1(_26624), .DIN2(_26262), .Q(_43420) );
  nor2s1 _44463_inst ( .DIN1(_53451), .DIN2(_26387), .Q(_44304) );
  nor2s1 _44464_inst ( .DIN1(_53449), .DIN2(_26207), .Q(_44303) );
  nor2s1 _44465_inst ( .DIN1(_44305), .DIN2(_26345), .Q(_44302) );
  nnd2s1 _44466_inst ( .DIN1(_44025), .DIN2(_43363), .Q(_44299) );
  nnd2s1 _44467_inst ( .DIN1(_44306), .DIN2(_43678), .Q(_43358) );
  hi1s1 _44468_inst ( .DIN(_43990), .Q(_43678) );
  nnd2s1 _44469_inst ( .DIN1(_44307), .DIN2(_44308), .Q(_43990) );
  or2s1 _44470_inst ( .DIN1(_44309), .DIN2(_43779), .Q(_44308) );
  nnd2s1 _44471_inst ( .DIN1(_43863), .DIN2(_43790), .Q(_44307) );
  hi1s1 _44472_inst ( .DIN(_43520), .Q(_43790) );
  nor2s1 _44473_inst ( .DIN1(_43147), .DIN2(_43219), .Q(_44306) );
  xnr2s1 _44474_inst ( .DIN1(_34338), .DIN2(_43544), .Q(_43219) );
  nnd2s1 _44475_inst ( .DIN1(_44310), .DIN2(_44058), .Q(_43544) );
  nor2s1 _44476_inst ( .DIN1(_27349), .DIN2(_43151), .Q(_44310) );
  nnd2s1 _44477_inst ( .DIN1(_44311), .DIN2(_44312), .Q(_34338) );
  hi1s1 _44478_inst ( .DIN(_44313), .Q(_44312) );
  nor2s1 _44479_inst ( .DIN1(_44314), .DIN2(_42799), .Q(_44311) );
  nnd2s1 _44480_inst ( .DIN1(_44315), .DIN2(_44316), .Q(_42799) );
  nor2s1 _44481_inst ( .DIN1(_42921), .DIN2(_44317), .Q(_44315) );
  nor2s1 _44482_inst ( .DIN1(_43876), .DIN2(_43121), .Q(_43147) );
  nor2s1 _44483_inst ( .DIN1(_43599), .DIN2(_37702), .Q(_28056) );
  nnd2s1 _44484_inst ( .DIN1(_44318), .DIN2(_44202), .Q(_37702) );
  nor2s1 _44485_inst ( .DIN1(_34489), .DIN2(_37411), .Q(_44318) );
  hi1s1 _44486_inst ( .DIN(_44319), .Q(_34489) );
  nnd2s1 _44487_inst ( .DIN1(_44320), .DIN2(_38713), .Q(_43599) );
  nor2s1 _44488_inst ( .DIN1(_38884), .DIN2(_33182), .Q(_44320) );
  nnd2s1 _44489_inst ( .DIN1(_44321), .DIN2(_43171), .Q(
        ____0____________0_____) );
  nnd2s1 _44490_inst ( .DIN1(_43502), .DIN2(_43174), .Q(_43171) );
  nor2s1 _44491_inst ( .DIN1(_44322), .DIN2(_44323), .Q(_43502) );
  nnd2s1 _44492_inst ( .DIN1(_44324), .DIN2(_31399), .Q(_44322) );
  hi1s1 _44493_inst ( .DIN(_31404), .Q(_31399) );
  nnd2s1 _44494_inst ( .DIN1(_44325), .DIN2(_44326), .Q(_31404) );
  nor2s1 _44495_inst ( .DIN1(_42750), .DIN2(_27308), .Q(_44325) );
  nor2s1 _44496_inst ( .DIN1(_44327), .DIN2(_44328), .Q(_44321) );
  nor2s1 _44497_inst ( .DIN1(_43174), .DIN2(_44329), .Q(_44328) );
  nnd2s1 _44498_inst ( .DIN1(_44330), .DIN2(_44331), .Q(_44329) );
  nor2s1 _44499_inst ( .DIN1(_44332), .DIN2(_44333), .Q(_44331) );
  nnd2s1 _44500_inst ( .DIN1(_44334), .DIN2(_44335), .Q(_44333) );
  nor2s1 _44501_inst ( .DIN1(_44336), .DIN2(_44337), .Q(_44335) );
  nor2s1 _44502_inst ( .DIN1(_43490), .DIN2(_44309), .Q(_44337) );
  nnd2s1 _44503_inst ( .DIN1(_44338), .DIN2(_44339), .Q(_44309) );
  nor2s1 _44504_inst ( .DIN1(_30820), .DIN2(_27473), .Q(_44338) );
  and2s1 _44505_inst ( .DIN1(_43621), .DIN2(_43779), .Q(_43490) );
  nnd2s1 _44506_inst ( .DIN1(_44340), .DIN2(_44341), .Q(_43779) );
  nor2s1 _44507_inst ( .DIN1(_44342), .DIN2(_44343), .Q(_44340) );
  nnd2s1 _44508_inst ( .DIN1(_26770), .DIN2(_44344), .Q(_43621) );
  nnd2s1 _44509_inst ( .DIN1(_44345), .DIN2(______[1]), .Q(_44344) );
  nor2s1 _44510_inst ( .DIN1(_26773), .DIN2(_44342), .Q(_44345) );
  nor2s1 _44511_inst ( .DIN1(_44346), .DIN2(_43514), .Q(_44336) );
  nor2s1 _44512_inst ( .DIN1(_44347), .DIN2(_44348), .Q(_44346) );
  nnd2s1 _44513_inst ( .DIN1(_44349), .DIN2(_44350), .Q(_44348) );
  nnd2s1 _44514_inst ( .DIN1(_43516), .DIN2(_53221), .Q(_44350) );
  nnd2s1 _44515_inst ( .DIN1(_30965), .DIN2(_44351), .Q(_44349) );
  nnd2s1 _44516_inst ( .DIN1(_44352), .DIN2(_44353), .Q(_44347) );
  nnd2s1 _44517_inst ( .DIN1(_44354), .DIN2(_44355), .Q(_44352) );
  nor2s1 _44518_inst ( .DIN1(_43831), .DIN2(_44356), .Q(_44334) );
  nor2s1 _44519_inst ( .DIN1(_43252), .DIN2(_44357), .Q(_44356) );
  nor2s1 _44520_inst ( .DIN1(_39969), .DIN2(_43960), .Q(_43831) );
  nnd2s1 _44521_inst ( .DIN1(_44358), .DIN2(_32088), .Q(_43960) );
  nor2s1 _44522_inst ( .DIN1(_43565), .DIN2(_44359), .Q(_44358) );
  hi1s1 _44523_inst ( .DIN(_41312), .Q(_39969) );
  nor2s1 _44524_inst ( .DIN1(_39635), .DIN2(_40460), .Q(_41312) );
  hi1s1 _44525_inst ( .DIN(_39721), .Q(_40460) );
  nnd2s1 _44526_inst ( .DIN1(_44360), .DIN2(_40363), .Q(_39721) );
  nor2s1 _44527_inst ( .DIN1(_34359), .DIN2(_39976), .Q(_40363) );
  nnd2s1 _44528_inst ( .DIN1(_40425), .DIN2(_53443), .Q(_39976) );
  nor2s1 _44529_inst ( .DIN1(_53436), .DIN2(_53442), .Q(_40425) );
  nnd2s1 _44530_inst ( .DIN1(_53439), .DIN2(_53438), .Q(_34359) );
  nor2s1 _44531_inst ( .DIN1(_40138), .DIN2(_40150), .Q(_44360) );
  nnd2s1 _44532_inst ( .DIN1(_44361), .DIN2(_53435), .Q(_40150) );
  nor2s1 _44533_inst ( .DIN1(_53392), .DIN2(_26211), .Q(_44361) );
  nnd2s1 _44534_inst ( .DIN1(_40431), .DIN2(_26238), .Q(_40138) );
  nor2s1 _44535_inst ( .DIN1(_26228), .DIN2(_53437), .Q(_40431) );
  nor2s1 _44536_inst ( .DIN1(_40467), .DIN2(_40073), .Q(_39635) );
  nnd2s1 _44537_inst ( .DIN1(_40468), .DIN2(_26437), .Q(_40073) );
  nor2s1 _44538_inst ( .DIN1(_26211), .DIN2(_53435), .Q(_40468) );
  hi1s1 _44539_inst ( .DIN(_39795), .Q(_40467) );
  nor2s1 _44540_inst ( .DIN1(_40404), .DIN2(_40166), .Q(_39795) );
  nnd2s1 _44541_inst ( .DIN1(_40337), .DIN2(_44362), .Q(_40166) );
  nor2s1 _44542_inst ( .DIN1(_26286), .DIN2(_44363), .Q(_44362) );
  nnd2s1 _44543_inst ( .DIN1(_26238), .DIN2(_26587), .Q(_44363) );
  nor2s1 _44544_inst ( .DIN1(_26356), .DIN2(_26228), .Q(_40337) );
  nnd2s1 _44545_inst ( .DIN1(_44364), .DIN2(_53436), .Q(_40404) );
  nor2s1 _44546_inst ( .DIN1(_26288), .DIN2(_26466), .Q(_44364) );
  nnd2s1 _44547_inst ( .DIN1(_44365), .DIN2(_44366), .Q(_44332) );
  nor2s1 _44548_inst ( .DIN1(_44367), .DIN2(_44368), .Q(_44366) );
  nnd2s1 _44549_inst ( .DIN1(_44369), .DIN2(_43652), .Q(_44368) );
  nnd2s1 _44550_inst ( .DIN1(_43352), .DIN2(_43939), .Q(_43652) );
  hi1s1 _44551_inst ( .DIN(_43252), .Q(_43939) );
  hi1s1 _44552_inst ( .DIN(_43218), .Q(_43352) );
  nnd2s1 _44553_inst ( .DIN1(_44370), .DIN2(_44371), .Q(_43218) );
  nor2s1 _44554_inst ( .DIN1(_39069), .DIN2(_30875), .Q(_44370) );
  nnd2s1 _44555_inst ( .DIN1(_44372), .DIN2(_44373), .Q(_44369) );
  nor2s1 _44556_inst ( .DIN1(_28214), .DIN2(_43139), .Q(_44372) );
  hi1s1 _44557_inst ( .DIN(_43574), .Q(_43139) );
  xor2s1 _44558_inst ( .DIN1(_44374), .DIN2(_36757), .Q(_43574) );
  hi1s1 _44559_inst ( .DIN(_41367), .Q(_36757) );
  nnd2s1 _44560_inst ( .DIN1(_44375), .DIN2(_44376), .Q(_41367) );
  and2s1 _44561_inst ( .DIN1(_44377), .DIN2(_44378), .Q(_44375) );
  nnd2s1 _44562_inst ( .DIN1(_26770), .DIN2(_44379), .Q(_44374) );
  nnd2s1 _44563_inst ( .DIN1(_44380), .DIN2(______[1]), .Q(_44379) );
  nor2s1 _44564_inst ( .DIN1(______[28]), .DIN2(______[19]), .Q(_44380) );
  nor2s1 _44565_inst ( .DIN1(_43864), .DIN2(_44381), .Q(_44367) );
  nor2s1 _44566_inst ( .DIN1(_43362), .DIN2(_44382), .Q(_44381) );
  nnd2s1 _44567_inst ( .DIN1(_44383), .DIN2(_44186), .Q(_44382) );
  nnd2s1 _44568_inst ( .DIN1(_44384), .DIN2(_29997), .Q(_44186) );
  hi1s1 _44569_inst ( .DIN(_30820), .Q(_29997) );
  nor2s1 _44570_inst ( .DIN1(_44385), .DIN2(_31190), .Q(_44384) );
  xor2s1 _44571_inst ( .DIN1(_44386), .DIN2(_2064), .Q(_44385) );
  nnd2s1 _44572_inst ( .DIN1(_29499), .DIN2(_32801), .Q(_44386) );
  nor2s1 _44573_inst ( .DIN1(_27475), .DIN2(_27474), .Q(_29499) );
  hi1s1 _44574_inst ( .DIN(_43863), .Q(_44383) );
  nor2s1 _44575_inst ( .DIN1(_44359), .DIN2(_32080), .Q(_43863) );
  hi1s1 _44576_inst ( .DIN(_44168), .Q(_43362) );
  nnd2s1 _44577_inst ( .DIN1(_44387), .DIN2(_44388), .Q(_44168) );
  nor2s1 _44578_inst ( .DIN1(_30964), .DIN2(_28114), .Q(_44388) );
  nor2s1 _44579_inst ( .DIN1(_31702), .DIN2(_29481), .Q(_44387) );
  nor2s1 _44580_inst ( .DIN1(_44389), .DIN2(_44390), .Q(_44365) );
  nor2s1 _44581_inst ( .DIN1(_44391), .DIN2(_43520), .Q(_44390) );
  nor2s1 _44582_inst ( .DIN1(_44392), .DIN2(_44393), .Q(_44391) );
  nnd2s1 _44583_inst ( .DIN1(_44394), .DIN2(_44395), .Q(_44393) );
  nnd2s1 _44584_inst ( .DIN1(_44396), .DIN2(_30375), .Q(_44395) );
  hi1s1 _44585_inst ( .DIN(_32012), .Q(_30375) );
  nor2s1 _44586_inst ( .DIN1(_44397), .DIN2(_27359), .Q(_44396) );
  nnd2s1 _44587_inst ( .DIN1(_43893), .DIN2(_26528), .Q(_44394) );
  nnd2s1 _44588_inst ( .DIN1(_44398), .DIN2(_44399), .Q(_44392) );
  nor2s1 _44589_inst ( .DIN1(_44400), .DIN2(_43233), .Q(_44389) );
  nor2s1 _44590_inst ( .DIN1(_44401), .DIN2(_44402), .Q(_44400) );
  nnd2s1 _44591_inst ( .DIN1(_44403), .DIN2(_44404), .Q(_44402) );
  nnd2s1 _44592_inst ( .DIN1(_44405), .DIN2(_44355), .Q(_44404) );
  nnd2s1 _44593_inst ( .DIN1(_44354), .DIN2(_44406), .Q(_44403) );
  hi1s1 _44594_inst ( .DIN(_27473), .Q(_44406) );
  and2s1 _44595_inst ( .DIN1(_29325), .DIN2(_44058), .Q(_44401) );
  hi1s1 _44596_inst ( .DIN(_29482), .Q(_29325) );
  nor2s1 _44597_inst ( .DIN1(_44407), .DIN2(_44408), .Q(_44330) );
  nnd2s1 _44598_inst ( .DIN1(_44409), .DIN2(_44410), .Q(_44408) );
  nor2s1 _44599_inst ( .DIN1(_43881), .DIN2(_43397), .Q(_44410) );
  nnd2s1 _44600_inst ( .DIN1(_44411), .DIN2(_44412), .Q(_43397) );
  nor2s1 _44601_inst ( .DIN1(_43113), .DIN2(_44413), .Q(_44412) );
  nor2s1 _44602_inst ( .DIN1(_43565), .DIN2(_43548), .Q(_44413) );
  nnd2s1 _44603_inst ( .DIN1(_44414), .DIN2(_44415), .Q(_43548) );
  nor2s1 _44604_inst ( .DIN1(_31190), .DIN2(_44416), .Q(_44415) );
  nor2s1 _44605_inst ( .DIN1(_30848), .DIN2(_27492), .Q(_44414) );
  and2s1 _44606_inst ( .DIN1(_43856), .DIN2(_43705), .Q(_43113) );
  nor2s1 _44607_inst ( .DIN1(_27493), .DIN2(_43811), .Q(_43856) );
  nor2s1 _44608_inst ( .DIN1(_44417), .DIN2(_43857), .Q(_44411) );
  nnd2s1 _44609_inst ( .DIN1(_44418), .DIN2(_44419), .Q(_43857) );
  nor2s1 _44610_inst ( .DIN1(_44420), .DIN2(_44421), .Q(_44419) );
  nnd2s1 _44611_inst ( .DIN1(_44422), .DIN2(_44423), .Q(_44421) );
  nnd2s1 _44612_inst ( .DIN1(_43660), .DIN2(_26770), .Q(_44423) );
  and2s1 _44613_inst ( .DIN1(_44424), .DIN2(_27296), .Q(_43660) );
  hi1s1 _44614_inst ( .DIN(_43979), .Q(_44422) );
  nnd2s1 _44615_inst ( .DIN1(_44425), .DIN2(_44426), .Q(_43979) );
  nnd2s1 _44616_inst ( .DIN1(_44427), .DIN2(_44354), .Q(_44426) );
  nor2s1 _44617_inst ( .DIN1(_43151), .DIN2(_27466), .Q(_44427) );
  nnd2s1 _44618_inst ( .DIN1(_44428), .DIN2(_44429), .Q(_44425) );
  nor2s1 _44619_inst ( .DIN1(_43891), .DIN2(_44397), .Q(_44429) );
  nor2s1 _44620_inst ( .DIN1(_27359), .DIN2(_32012), .Q(_44428) );
  nnd2s1 _44621_inst ( .DIN1(_44231), .DIN2(_44430), .Q(_44420) );
  hi1s1 _44622_inst ( .DIN(_43672), .Q(_44430) );
  nor2s1 _44623_inst ( .DIN1(_44353), .DIN2(_43151), .Q(_43672) );
  nnd2s1 _44624_inst ( .DIN1(_44431), .DIN2(_44432), .Q(_44353) );
  nor2s1 _44625_inst ( .DIN1(_28985), .DIN2(_30849), .Q(_44432) );
  nor2s1 _44626_inst ( .DIN1(_28170), .DIN2(_27359), .Q(_44431) );
  or2s1 _44627_inst ( .DIN1(_44398), .DIN2(_43891), .Q(_44231) );
  nnd2s1 _44628_inst ( .DIN1(_44433), .DIN2(_44434), .Q(_44398) );
  nor2s1 _44629_inst ( .DIN1(_28985), .DIN2(_44416), .Q(_44434) );
  nor2s1 _44630_inst ( .DIN1(_32340), .DIN2(_27466), .Q(_44433) );
  nor2s1 _44631_inst ( .DIN1(_44435), .DIN2(_44436), .Q(_44418) );
  or2s1 _44632_inst ( .DIN1(_43493), .DIN2(_43817), .Q(_44436) );
  or2s1 _44633_inst ( .DIN1(_44437), .DIN2(_43492), .Q(_43817) );
  nnd2s1 _44634_inst ( .DIN1(_44438), .DIN2(_44439), .Q(_43492) );
  nor2s1 _44635_inst ( .DIN1(_43648), .DIN2(_44440), .Q(_44439) );
  nnd2s1 _44636_inst ( .DIN1(_43675), .DIN2(_44182), .Q(_44440) );
  nnd2s1 _44637_inst ( .DIN1(_44441), .DIN2(_44058), .Q(_44182) );
  nor2s1 _44638_inst ( .DIN1(_29482), .DIN2(_43226), .Q(_44441) );
  hi1s1 _44639_inst ( .DIN(_44089), .Q(_43675) );
  nor2s1 _44640_inst ( .DIN1(_44357), .DIN2(_43137), .Q(_44089) );
  nnd2s1 _44641_inst ( .DIN1(_44442), .DIN2(_44443), .Q(_44357) );
  nor2s1 _44642_inst ( .DIN1(_28985), .DIN2(_28170), .Q(_44443) );
  nor2s1 _44643_inst ( .DIN1(_32340), .DIN2(_29482), .Q(_44442) );
  nnd2s1 _44644_inst ( .DIN1(_44113), .DIN2(_44444), .Q(_29482) );
  nor2s1 _44645_inst ( .DIN1(_44073), .DIN2(_43565), .Q(_43648) );
  nnd2s1 _44646_inst ( .DIN1(_44373), .DIN2(_30821), .Q(_44073) );
  hi1s1 _44647_inst ( .DIN(_28170), .Q(_30821) );
  nor2s1 _44648_inst ( .DIN1(_44445), .DIN2(_43699), .Q(_44438) );
  nor2s1 _44649_inst ( .DIN1(_43473), .DIN2(_44293), .Q(_43699) );
  nnd2s1 _44650_inst ( .DIN1(_44446), .DIN2(_44447), .Q(_44293) );
  nor2s1 _44651_inst ( .DIN1(_44416), .DIN2(_27373), .Q(_44446) );
  nor2s1 _44652_inst ( .DIN1(_43096), .DIN2(_43095), .Q(_44445) );
  nnd2s1 _44653_inst ( .DIN1(_44448), .DIN2(_44449), .Q(_43095) );
  nor2s1 _44654_inst ( .DIN1(_32341), .DIN2(_27335), .Q(_44448) );
  hi1s1 _44655_inst ( .DIN(_44450), .Q(_27335) );
  or2s1 _44656_inst ( .DIN1(_43651), .DIN2(_43190), .Q(_44437) );
  nor2s1 _44657_inst ( .DIN1(_43351), .DIN2(_43520), .Q(_43190) );
  nnd2s1 _44658_inst ( .DIN1(_44451), .DIN2(_44452), .Q(_43351) );
  and2s1 _44659_inst ( .DIN1(_44453), .DIN2(_44405), .Q(_43651) );
  nor2s1 _44660_inst ( .DIN1(_27466), .DIN2(_43226), .Q(_44453) );
  nnd2s1 _44661_inst ( .DIN1(_44454), .DIN2(_44455), .Q(_43493) );
  nnd2s1 _44662_inst ( .DIN1(_43661), .DIN2(_26770), .Q(_44455) );
  hi1s1 _44663_inst ( .DIN(_43796), .Q(_43661) );
  nnd2s1 _44664_inst ( .DIN1(_44424), .DIN2(_29801), .Q(_43796) );
  nor2s1 _44665_inst ( .DIN1(_44021), .DIN2(_44000), .Q(_44454) );
  nor2s1 _44666_inst ( .DIN1(_43189), .DIN2(_43520), .Q(_44000) );
  nnd2s1 _44667_inst ( .DIN1(_44456), .DIN2(_44457), .Q(_43189) );
  nor2s1 _44668_inst ( .DIN1(_28114), .DIN2(_30677), .Q(_44457) );
  nor2s1 _44669_inst ( .DIN1(_30963), .DIN2(_27497), .Q(_44456) );
  nor2s1 _44670_inst ( .DIN1(_44399), .DIN2(_43891), .Q(_44021) );
  hi1s1 _44671_inst ( .DIN(_43725), .Q(_43891) );
  nnd2s1 _44672_inst ( .DIN1(_44458), .DIN2(_44459), .Q(_44399) );
  nor2s1 _44673_inst ( .DIN1(_28985), .DIN2(_27349), .Q(_44459) );
  nor2s1 _44674_inst ( .DIN1(_30849), .DIN2(_32081), .Q(_44458) );
  or2s1 _44675_inst ( .DIN1(_44159), .DIN2(_43935), .Q(_44435) );
  nnd2s1 _44676_inst ( .DIN1(_43715), .DIN2(_44460), .Q(_43935) );
  nnd2s1 _44677_inst ( .DIN1(_43724), .DIN2(_43363), .Q(_44460) );
  hi1s1 _44678_inst ( .DIN(_44157), .Q(_43724) );
  nnd2s1 _44679_inst ( .DIN1(_44461), .DIN2(_44449), .Q(_44157) );
  nor2s1 _44680_inst ( .DIN1(_30834), .DIN2(_27349), .Q(_44461) );
  nnd2s1 _44681_inst ( .DIN1(_44462), .DIN2(_43414), .Q(_43715) );
  and2s1 _44682_inst ( .DIN1(_44351), .DIN2(_30965), .Q(_44462) );
  nnd2s1 _44683_inst ( .DIN1(_44463), .DIN2(_44464), .Q(_44351) );
  nnd2s1 _44684_inst ( .DIN1(_44465), .DIN2(_30369), .Q(_44464) );
  nor2s1 _44685_inst ( .DIN1(_27349), .DIN2(_44416), .Q(_44465) );
  hi1s1 _44686_inst ( .DIN(_28215), .Q(_44416) );
  nor2s1 _44687_inst ( .DIN1(_44214), .DIN2(_26207), .Q(_28215) );
  nnd2s1 _44688_inst ( .DIN1(_44466), .DIN2(_53458), .Q(_44214) );
  nor2s1 _44689_inst ( .DIN1(_53446), .DIN2(_53449), .Q(_44466) );
  nnd2s1 _44690_inst ( .DIN1(_44467), .DIN2(_29354), .Q(_44463) );
  hi1s1 _44691_inst ( .DIN(_27336), .Q(_29354) );
  nor2s1 _44692_inst ( .DIN1(_32081), .DIN2(_30848), .Q(_44467) );
  nnd2s1 _44693_inst ( .DIN1(_44468), .DIN2(_44469), .Q(_44159) );
  nnd2s1 _44694_inst ( .DIN1(_43982), .DIN2(_26770), .Q(_44469) );
  hi1s1 _44695_inst ( .DIN(_43693), .Q(_43982) );
  nnd2s1 _44696_inst ( .DIN1(_44470), .DIN2(_44339), .Q(_43693) );
  nor2s1 _44697_inst ( .DIN1(_28170), .DIN2(_27358), .Q(_44470) );
  nnd2s1 _44698_inst ( .DIN1(_43516), .DIN2(_43414), .Q(_44468) );
  hi1s1 _44699_inst ( .DIN(_43151), .Q(_43414) );
  xor2s1 _44700_inst ( .DIN1(_27329), .DIN2(_44471), .Q(_43516) );
  nor2s1 _44701_inst ( .DIN1(_44472), .DIN2(_44473), .Q(_44471) );
  nnd2s1 _44702_inst ( .DIN1(_44450), .DIN2(_28849), .Q(_44473) );
  hi1s1 _44703_inst ( .DIN(_28985), .Q(_28849) );
  nor2s1 _44704_inst ( .DIN1(_43096), .DIN2(_43272), .Q(_44417) );
  nnd2s1 _44705_inst ( .DIN1(_44474), .DIN2(_29346), .Q(_43272) );
  nnd2s1 _44706_inst ( .DIN1(_43337), .DIN2(_44475), .Q(_43881) );
  nnd2s1 _44707_inst ( .DIN1(_43919), .DIN2(_43705), .Q(_44475) );
  hi1s1 _44708_inst ( .DIN(_43434), .Q(_43919) );
  nnd2s1 _44709_inst ( .DIN1(_44476), .DIN2(_30831), .Q(_43434) );
  hi1s1 _44710_inst ( .DIN(_44477), .Q(_30831) );
  nnd2s1 _44711_inst ( .DIN1(_43915), .DIN2(_26770), .Q(_43337) );
  hi1s1 _44712_inst ( .DIN(_43681), .Q(_43915) );
  nnd2s1 _44713_inst ( .DIN1(_44478), .DIN2(_44479), .Q(_43681) );
  nor2s1 _44714_inst ( .DIN1(_30964), .DIN2(_27493), .Q(_44479) );
  nnd2s1 _44715_inst ( .DIN1(_43806), .DIN2(_44480), .Q(_27493) );
  nor2s1 _44716_inst ( .DIN1(_32339), .DIN2(_44481), .Q(_44478) );
  nor2s1 _44717_inst ( .DIN1(_43446), .DIN2(_43969), .Q(_44409) );
  nnd2s1 _44718_inst ( .DIN1(_44482), .DIN2(_43195), .Q(_43969) );
  and2s1 _44719_inst ( .DIN1(_44151), .DIN2(_44483), .Q(_43195) );
  nnd2s1 _44720_inst ( .DIN1(_43561), .DIN2(_43108), .Q(_44483) );
  and2s1 _44721_inst ( .DIN1(_44484), .DIN2(_44485), .Q(_43561) );
  nor2s1 _44722_inst ( .DIN1(_44477), .DIN2(_28114), .Q(_44485) );
  nor2s1 _44723_inst ( .DIN1(_30963), .DIN2(_27348), .Q(_44484) );
  nnd2s1 _44724_inst ( .DIN1(_44486), .DIN2(_43720), .Q(_44151) );
  nor2s1 _44725_inst ( .DIN1(_43233), .DIN2(_43392), .Q(_44486) );
  hi1s1 _44726_inst ( .DIN(_44487), .Q(_43392) );
  nor2s1 _44727_inst ( .DIN1(_43231), .DIN2(_44488), .Q(_44482) );
  nor2s1 _44728_inst ( .DIN1(_43391), .DIN2(_43441), .Q(_44488) );
  nnd2s1 _44729_inst ( .DIN1(_44489), .DIN2(_29204), .Q(_43441) );
  hi1s1 _44730_inst ( .DIN(_29501), .Q(_29204) );
  nor2s1 _44731_inst ( .DIN1(_30834), .DIN2(_44490), .Q(_44489) );
  nor2s1 _44732_inst ( .DIN1(_43473), .DIN2(_43559), .Q(_43231) );
  nnd2s1 _44733_inst ( .DIN1(_44491), .DIN2(_44492), .Q(_43559) );
  nor2s1 _44734_inst ( .DIN1(_28985), .DIN2(_27359), .Q(_44492) );
  nor2s1 _44735_inst ( .DIN1(_30848), .DIN2(_29999), .Q(_44491) );
  nnd2s1 _44736_inst ( .DIN1(_44493), .DIN2(_44494), .Q(_43446) );
  nor2s1 _44737_inst ( .DIN1(_44495), .DIN2(_44496), .Q(_44494) );
  nnd2s1 _44738_inst ( .DIN1(_43886), .DIN2(_44497), .Q(_44496) );
  nnd2s1 _44739_inst ( .DIN1(_43413), .DIN2(_43108), .Q(_44497) );
  hi1s1 _44740_inst ( .DIN(_44015), .Q(_43413) );
  nnd2s1 _44741_inst ( .DIN1(_44476), .DIN2(_30526), .Q(_44015) );
  hi1s1 _44742_inst ( .DIN(_30236), .Q(_30526) );
  and2s1 _44743_inst ( .DIN1(_44498), .DIN2(_29902), .Q(_44476) );
  hi1s1 _44744_inst ( .DIN(_44481), .Q(_29902) );
  nor2s1 _44745_inst ( .DIN1(_39069), .DIN2(_31121), .Q(_44498) );
  nnd2s1 _44746_inst ( .DIN1(_43723), .DIN2(_43336), .Q(_43886) );
  and2s1 _44747_inst ( .DIN1(_44424), .DIN2(_39068), .Q(_43723) );
  and2s1 _44748_inst ( .DIN1(_28116), .DIN2(_44339), .Q(_44424) );
  nnd2s1 _44749_inst ( .DIN1(_44499), .DIN2(_44500), .Q(_44495) );
  hi1s1 _44750_inst ( .DIN(_43524), .Q(_44500) );
  nor2s1 _44751_inst ( .DIN1(_43658), .DIN2(_43473), .Q(_43524) );
  nnd2s1 _44752_inst ( .DIN1(_44501), .DIN2(_44502), .Q(_43658) );
  nor2s1 _44753_inst ( .DIN1(_31190), .DIN2(_27373), .Q(_44502) );
  hi1s1 _44754_inst ( .DIN(_39068), .Q(_27373) );
  nor2s1 _44755_inst ( .DIN1(_27475), .DIN2(_27374), .Q(_39068) );
  nor2s1 _44756_inst ( .DIN1(_32012), .DIN2(_30820), .Q(_44501) );
  nor2s1 _44757_inst ( .DIN1(_43670), .DIN2(_43690), .Q(_44499) );
  and2s1 _44758_inst ( .DIN1(_43892), .DIN2(_43363), .Q(_43690) );
  and2s1 _44759_inst ( .DIN1(_44503), .DIN2(_44504), .Q(_43892) );
  nor2s1 _44760_inst ( .DIN1(_32010), .DIN2(_27336), .Q(_44503) );
  nor2s1 _44761_inst ( .DIN1(_43370), .DIN2(_43520), .Q(_43670) );
  nnd2s1 _44762_inst ( .DIN1(_44505), .DIN2(_44506), .Q(_43370) );
  nor2s1 _44763_inst ( .DIN1(_44477), .DIN2(_32080), .Q(_44506) );
  nor2s1 _44764_inst ( .DIN1(_30963), .DIN2(_39069), .Q(_44505) );
  nnd2s1 _44765_inst ( .DIN1(_44507), .DIN2(_44130), .Q(_39069) );
  nor2s1 _44766_inst ( .DIN1(_44508), .DIN2(_44509), .Q(_44493) );
  nnd2s1 _44767_inst ( .DIN1(_43665), .DIN2(_43766), .Q(_44509) );
  and2s1 _44768_inst ( .DIN1(_44510), .DIN2(_44511), .Q(_43766) );
  nor2s1 _44769_inst ( .DIN1(_44512), .DIN2(_44513), .Q(_44511) );
  or2s1 _44770_inst ( .DIN1(_43268), .DIN2(_43526), .Q(_44513) );
  nor2s1 _44771_inst ( .DIN1(_43120), .DIN2(_43461), .Q(_43526) );
  nnd2s1 _44772_inst ( .DIN1(_44514), .DIN2(_44449), .Q(_43120) );
  nor2s1 _44773_inst ( .DIN1(_27358), .DIN2(_32012), .Q(_44514) );
  hi1s1 _44774_inst ( .DIN(_44264), .Q(_43268) );
  nnd2s1 _44775_inst ( .DIN1(_44046), .DIN2(_43586), .Q(_44264) );
  hi1s1 _44776_inst ( .DIN(_43664), .Q(_43586) );
  and2s1 _44777_inst ( .DIN1(_44515), .DIN2(_44487), .Q(_44046) );
  nor2s1 _44778_inst ( .DIN1(_30236), .DIN2(_44481), .Q(_44515) );
  nnd2s1 _44779_inst ( .DIN1(_44516), .DIN2(_43878), .Q(_44512) );
  nnd2s1 _44780_inst ( .DIN1(_43118), .DIN2(_43749), .Q(_43878) );
  hi1s1 _44781_inst ( .DIN(_43369), .Q(_43118) );
  nnd2s1 _44782_inst ( .DIN1(_44517), .DIN2(_29816), .Q(_43369) );
  hi1s1 _44783_inst ( .DIN(_29353), .Q(_29816) );
  nnd2s1 _44784_inst ( .DIN1(_43806), .DIN2(_44507), .Q(_29353) );
  and2s1 _44785_inst ( .DIN1(_29969), .DIN2(_44339), .Q(_44517) );
  nor2s1 _44786_inst ( .DIN1(_32012), .DIN2(_28985), .Q(_44339) );
  nor2s1 _44787_inst ( .DIN1(_44126), .DIN2(_44298), .Q(_44516) );
  nor2s1 _44788_inst ( .DIN1(_43930), .DIN2(_43461), .Q(_44298) );
  hi1s1 _44789_inst ( .DIN(_43705), .Q(_43461) );
  nnd2s1 _44790_inst ( .DIN1(_43435), .DIN2(_43121), .Q(_43705) );
  nnd2s1 _44791_inst ( .DIN1(_44518), .DIN2(______[1]), .Q(_43121) );
  nor2s1 _44792_inst ( .DIN1(_44519), .DIN2(_44342), .Q(_44518) );
  hi1s1 _44793_inst ( .DIN(_43815), .Q(_43435) );
  nnd2s1 _44794_inst ( .DIN1(_44405), .DIN2(_29801), .Q(_43930) );
  hi1s1 _44795_inst ( .DIN(_27492), .Q(_29801) );
  nnd2s1 _44796_inst ( .DIN1(_43806), .DIN2(_44520), .Q(_27492) );
  nor2s1 _44797_inst ( .DIN1(_44490), .DIN2(_32340), .Q(_44405) );
  hi1s1 _44798_inst ( .DIN(_43855), .Q(_44126) );
  nnd2s1 _44799_inst ( .DIN1(_44521), .DIN2(_44373), .Q(_43855) );
  and2s1 _44800_inst ( .DIN1(_44522), .DIN2(_27342), .Q(_44373) );
  nor2s1 _44801_inst ( .DIN1(_28985), .DIN2(_32010), .Q(_44522) );
  nor2s1 _44802_inst ( .DIN1(_43512), .DIN2(_28214), .Q(_44521) );
  nnd2s1 _44803_inst ( .DIN1(_44523), .DIN2(______[1]), .Q(_43512) );
  nor2s1 _44804_inst ( .DIN1(______[19]), .DIN2(_44519), .Q(_44523) );
  nor2s1 _44805_inst ( .DIN1(_44524), .DIN2(_44525), .Q(_44510) );
  nnd2s1 _44806_inst ( .DIN1(_44526), .DIN2(_44255), .Q(_44525) );
  and2s1 _44807_inst ( .DIN1(_44527), .DIN2(_44528), .Q(_44255) );
  or2s1 _44808_inst ( .DIN1(_43558), .DIN2(_43096), .Q(_44528) );
  nnd2s1 _44809_inst ( .DIN1(_44450), .DIN2(_44474), .Q(_43558) );
  and2s1 _44810_inst ( .DIN1(_44504), .DIN2(_31699), .Q(_44474) );
  hi1s1 _44811_inst ( .DIN(_32340), .Q(_31699) );
  nor2s1 _44812_inst ( .DIN1(_28864), .DIN2(_29999), .Q(_44504) );
  nor2s1 _44813_inst ( .DIN1(_44175), .DIN2(_44101), .Q(_44450) );
  nor2s1 _44814_inst ( .DIN1(_44529), .DIN2(_44530), .Q(_44527) );
  nor2s1 _44815_inst ( .DIN1(_43391), .DIN2(_43415), .Q(_44530) );
  nnd2s1 _44816_inst ( .DIN1(_44531), .DIN2(_44447), .Q(_43415) );
  nor2s1 _44817_inst ( .DIN1(_32081), .DIN2(_27358), .Q(_44531) );
  hi1s1 _44818_inst ( .DIN(_43393), .Q(_44529) );
  nnd2s1 _44819_inst ( .DIN1(_44532), .DIN2(_44354), .Q(_43393) );
  and2s1 _44820_inst ( .DIN1(_44449), .DIN2(_32801), .Q(_44354) );
  hi1s1 _44821_inst ( .DIN(_30849), .Q(_32801) );
  nor2s1 _44822_inst ( .DIN1(_29999), .DIN2(_31190), .Q(_44449) );
  hi1s1 _44823_inst ( .DIN(_29894), .Q(_29999) );
  nor2s1 _44824_inst ( .DIN1(_44305), .DIN2(_44533), .Q(_29894) );
  nor2s1 _44825_inst ( .DIN1(_27473), .DIN2(_43226), .Q(_44532) );
  nnd2s1 _44826_inst ( .DIN1(_44520), .DIN2(_44444), .Q(_27473) );
  hi1s1 _44827_inst ( .DIN(_43865), .Q(_44526) );
  nnd2s1 _44828_inst ( .DIN1(_44534), .DIN2(_44535), .Q(_43865) );
  nor2s1 _44829_inst ( .DIN1(_43223), .DIN2(_43182), .Q(_44535) );
  nor2s1 _44830_inst ( .DIN1(_43664), .DIN2(_44075), .Q(_43182) );
  nnd2s1 _44831_inst ( .DIN1(_44536), .DIN2(_44537), .Q(_44075) );
  nor2s1 _44832_inst ( .DIN1(_44477), .DIN2(_30872), .Q(_44536) );
  nor2s1 _44833_inst ( .DIN1(_43664), .DIN2(_43123), .Q(_43223) );
  nnd2s1 _44834_inst ( .DIN1(_44538), .DIN2(_44487), .Q(_43123) );
  nor2s1 _44835_inst ( .DIN1(_30677), .DIN2(_44481), .Q(_44538) );
  nor2s1 _44836_inst ( .DIN1(_44539), .DIN2(_43269), .Q(_44534) );
  nor2s1 _44837_inst ( .DIN1(_43929), .DIN2(_43940), .Q(_43269) );
  nnd2s1 _44838_inst ( .DIN1(_44371), .DIN2(_44540), .Q(_43940) );
  nor2s1 _44839_inst ( .DIN1(_27467), .DIN2(_32080), .Q(_44540) );
  nor2s1 _44840_inst ( .DIN1(_30963), .DIN2(_31702), .Q(_44371) );
  nor2s1 _44841_inst ( .DIN1(_43520), .DIN2(_43188), .Q(_44539) );
  hi1s1 _44842_inst ( .DIN(_44025), .Q(_43188) );
  xor2s1 _44843_inst ( .DIN1(_44541), .DIN2(_44542), .Q(_44025) );
  hi1s1 _44844_inst ( .DIN(_31569), .Q(_44542) );
  nnd2s1 _44845_inst ( .DIN1(_44543), .DIN2(_44544), .Q(_44541) );
  nor2s1 _44846_inst ( .DIN1(_30236), .DIN2(_29655), .Q(_44544) );
  nnd2s1 _44847_inst ( .DIN1(_29818), .DIN2(_44130), .Q(_29655) );
  nor2s1 _44848_inst ( .DIN1(_28114), .DIN2(_30963), .Q(_44543) );
  nnd2s1 _44849_inst ( .DIN1(_44545), .DIN2(_43091), .Q(_44524) );
  and2s1 _44850_inst ( .DIN1(_44546), .DIN2(_44547), .Q(_43091) );
  nnd2s1 _44851_inst ( .DIN1(_43893), .DIN2(_43186), .Q(_44547) );
  hi1s1 _44852_inst ( .DIN(_43521), .Q(_43893) );
  nnd2s1 _44853_inst ( .DIN1(_44548), .DIN2(_44549), .Q(_43521) );
  nor2s1 _44854_inst ( .DIN1(_31190), .DIN2(_30849), .Q(_44549) );
  nor2s1 _44855_inst ( .DIN1(_27336), .DIN2(_28214), .Q(_44548) );
  nnd2s1 _44856_inst ( .DIN1(_43806), .DIN2(_29818), .Q(_27336) );
  nnd2s1 _44857_inst ( .DIN1(_43916), .DIN2(_26770), .Q(_44546) );
  hi1s1 _44858_inst ( .DIN(_43519), .Q(_43916) );
  nnd2s1 _44859_inst ( .DIN1(_44550), .DIN2(_44551), .Q(_43519) );
  nor2s1 _44860_inst ( .DIN1(_28864), .DIN2(_32081), .Q(_44551) );
  nor2s1 _44861_inst ( .DIN1(_32012), .DIN2(_27466), .Q(_44550) );
  hi1s1 _44862_inst ( .DIN(_44355), .Q(_27466) );
  nor2s1 _44863_inst ( .DIN1(_27374), .DIN2(_44175), .Q(_44355) );
  nnd2s1 _44864_inst ( .DIN1(_44217), .DIN2(_44552), .Q(_32012) );
  nor2s1 _44865_inst ( .DIN1(_44553), .DIN2(_44554), .Q(_44545) );
  nor2s1 _44866_inst ( .DIN1(_43565), .DIN2(_43887), .Q(_44554) );
  nnd2s1 _44867_inst ( .DIN1(_44555), .DIN2(_44447), .Q(_43887) );
  nor2s1 _44868_inst ( .DIN1(_28985), .DIN2(_32341), .Q(_44447) );
  nor2s1 _44869_inst ( .DIN1(_30820), .DIN2(_29501), .Q(_44555) );
  nnd2s1 _44870_inst ( .DIN1(_44520), .DIN2(_44130), .Q(_29501) );
  nnd2s1 _44871_inst ( .DIN1(_44556), .DIN2(_53458), .Q(_30820) );
  nor2s1 _44872_inst ( .DIN1(_53446), .DIN2(_44557), .Q(_44556) );
  nor2s1 _44873_inst ( .DIN1(_44263), .DIN2(_43233), .Q(_44553) );
  nor2s1 _44874_inst ( .DIN1(_43556), .DIN2(_43335), .Q(_44263) );
  hi1s1 _44875_inst ( .DIN(_43230), .Q(_43335) );
  nnd2s1 _44876_inst ( .DIN1(_43720), .DIN2(_44537), .Q(_43230) );
  nor2s1 _44877_inst ( .DIN1(_30236), .DIN2(_32080), .Q(_43720) );
  nnd2s1 _44878_inst ( .DIN1(_44217), .DIN2(_44558), .Q(_30236) );
  nor2s1 _44879_inst ( .DIN1(_44359), .DIN2(_28114), .Q(_43556) );
  nnd2s1 _44880_inst ( .DIN1(_44559), .DIN2(_28850), .Q(_44359) );
  hi1s1 _44881_inst ( .DIN(_31121), .Q(_28850) );
  nor2s1 _44882_inst ( .DIN1(_30677), .DIN2(_27348), .Q(_44559) );
  xor2s1 _44883_inst ( .DIN1(_31569), .DIN2(_44560), .Q(_43665) );
  nor2s1 _44884_inst ( .DIN1(_44297), .DIN2(_44561), .Q(_44560) );
  hi1s1 _44885_inst ( .DIN(_44185), .Q(_44561) );
  nnd2s1 _44886_inst ( .DIN1(_44562), .DIN2(_29203), .Q(_44185) );
  hi1s1 _44887_inst ( .DIN(_29481), .Q(_29203) );
  nor2s1 _44888_inst ( .DIN1(_43811), .DIN2(_43514), .Q(_44562) );
  nor2s1 _44889_inst ( .DIN1(_43253), .DIN2(_43096), .Q(_44297) );
  hi1s1 _44890_inst ( .DIN(_43749), .Q(_43096) );
  nnd2s1 _44891_inst ( .DIN1(_44563), .DIN2(_44564), .Q(_43253) );
  nor2s1 _44892_inst ( .DIN1(_31190), .DIN2(_28170), .Q(_44564) );
  nnd2s1 _44893_inst ( .DIN1(_44565), .DIN2(_44566), .Q(_28170) );
  nor2s1 _44894_inst ( .DIN1(_53449), .DIN2(_53458), .Q(_44566) );
  nor2s1 _44895_inst ( .DIN1(_26215), .DIN2(_26207), .Q(_44565) );
  nor2s1 _44896_inst ( .DIN1(_27358), .DIN2(_30848), .Q(_44563) );
  nnd2s1 _44897_inst ( .DIN1(_44567), .DIN2(_42880), .Q(_31569) );
  hi1s1 _44898_inst ( .DIN(_40399), .Q(_42880) );
  nnd2s1 _44899_inst ( .DIN1(_44568), .DIN2(_44569), .Q(_40399) );
  nor2s1 _44900_inst ( .DIN1(_44570), .DIN2(_44571), .Q(_44569) );
  nnd2s1 _44901_inst ( .DIN1(_44572), .DIN2(_44573), .Q(_44571) );
  nor2s1 _44902_inst ( .DIN1(_44574), .DIN2(_44575), .Q(_44568) );
  nnd2s1 _44903_inst ( .DIN1(_44576), .DIN2(_44577), .Q(_44575) );
  nor2s1 _44904_inst ( .DIN1(_44578), .DIN2(_44579), .Q(_44567) );
  nnd2s1 _44905_inst ( .DIN1(_44580), .DIN2(_44581), .Q(_44508) );
  hi1s1 _44906_inst ( .DIN(_43663), .Q(_44581) );
  nnd2s1 _44907_inst ( .DIN1(_43407), .DIN2(_43841), .Q(_43663) );
  nnd2s1 _44908_inst ( .DIN1(_44582), .DIN2(_44058), .Q(_43841) );
  nor2s1 _44909_inst ( .DIN1(_44490), .DIN2(_32341), .Q(_44058) );
  nnd2s1 _44910_inst ( .DIN1(_43807), .DIN2(_44558), .Q(_32341) );
  hi1s1 _44911_inst ( .DIN(_44583), .Q(_44490) );
  nor2s1 _44912_inst ( .DIN1(_43473), .DIN2(_27349), .Q(_44582) );
  hi1s1 _44913_inst ( .DIN(_29346), .Q(_27349) );
  hi1s1 _44914_inst ( .DIN(_43562), .Q(_43473) );
  nnd2s1 _44915_inst ( .DIN1(_43844), .DIN2(_43108), .Q(_43407) );
  hi1s1 _44916_inst ( .DIN(_43514), .Q(_43108) );
  nor2s1 _44917_inst ( .DIN1(_27497), .DIN2(_43811), .Q(_43844) );
  nnd2s1 _44918_inst ( .DIN1(_44444), .DIN2(_29818), .Q(_27497) );
  hi1s1 _44919_inst ( .DIN(_27375), .Q(_29818) );
  nor2s1 _44920_inst ( .DIN1(_44584), .DIN2(_43647), .Q(_44580) );
  nnd2s1 _44921_inst ( .DIN1(_44585), .DIN2(_44586), .Q(_43647) );
  nnd2s1 _44922_inst ( .DIN1(_44268), .DIN2(_43749), .Q(_44586) );
  nnd2s1 _44923_inst ( .DIN1(_43252), .DIN2(_43137), .Q(_43749) );
  nnd2s1 _44924_inst ( .DIN1(_44587), .DIN2(_44341), .Q(_43137) );
  nnd2s1 _44925_inst ( .DIN1(_26770), .DIN2(_44588), .Q(_43252) );
  nnd2s1 _44926_inst ( .DIN1(_44587), .DIN2(______[28]), .Q(_44588) );
  nor2s1 _44927_inst ( .DIN1(______[1]), .DIN2(______[19]), .Q(_44587) );
  hi1s1 _44928_inst ( .DIN(_43368), .Q(_44268) );
  nnd2s1 _44929_inst ( .DIN1(_44589), .DIN2(_44590), .Q(_43368) );
  nor2s1 _44930_inst ( .DIN1(_28985), .DIN2(_27358), .Q(_44590) );
  hi1s1 _44931_inst ( .DIN(_27296), .Q(_27358) );
  nor2s1 _44932_inst ( .DIN1(_44099), .DIN2(_44175), .Q(_27296) );
  nnd2s1 _44933_inst ( .DIN1(_44591), .DIN2(_53459), .Q(_44175) );
  nnd2s1 _44934_inst ( .DIN1(_44592), .DIN2(_53444), .Q(_28985) );
  nor2s1 _44935_inst ( .DIN1(_26227), .DIN2(_26428), .Q(_44592) );
  nor2s1 _44936_inst ( .DIN1(_30848), .DIN2(_28214), .Q(_44589) );
  hi1s1 _44937_inst ( .DIN(_28116), .Q(_28214) );
  nor2s1 _44938_inst ( .DIN1(_44593), .DIN2(_44557), .Q(_28116) );
  nnd2s1 _44939_inst ( .DIN1(_26243), .DIN2(_53446), .Q(_44593) );
  xor2s1 _44940_inst ( .DIN1(_43275), .DIN2(_29490), .Q(_44585) );
  nor2s1 _44941_inst ( .DIN1(_43759), .DIN2(_43520), .Q(_43275) );
  nnd2s1 _44942_inst ( .DIN1(_44594), .DIN2(_44595), .Q(_43759) );
  nor2s1 _44943_inst ( .DIN1(_44477), .DIN2(_27467), .Q(_44595) );
  nor2s1 _44944_inst ( .DIN1(_30963), .DIN2(_44481), .Q(_44594) );
  xor2s1 _44945_inst ( .DIN1(_34151), .DIN2(_44596), .Q(_44584) );
  nor2s1 _44946_inst ( .DIN1(_43864), .DIN2(_43988), .Q(_44596) );
  nnd2s1 _44947_inst ( .DIN1(_44597), .DIN2(_29346), .Q(_43988) );
  nor2s1 _44948_inst ( .DIN1(_43804), .DIN2(_27374), .Q(_29346) );
  nnd2s1 _44949_inst ( .DIN1(_44598), .DIN2(_53454), .Q(_43804) );
  nor2s1 _44950_inst ( .DIN1(_53455), .DIN2(_53459), .Q(_44598) );
  nor2s1 _44951_inst ( .DIN1(_44397), .DIN2(_30834), .Q(_44597) );
  nnd2s1 _44952_inst ( .DIN1(_44218), .DIN2(_44056), .Q(_30834) );
  hi1s1 _44953_inst ( .DIN(_43363), .Q(_43864) );
  nnd2s1 _44954_inst ( .DIN1(_43030), .DIN2(_43029), .Q(_34151) );
  and2s1 _44955_inst ( .DIN1(_44599), .DIN2(_44600), .Q(_43030) );
  nor2s1 _44956_inst ( .DIN1(_44601), .DIN2(_44602), .Q(_44599) );
  nnd2s1 _44957_inst ( .DIN1(_44603), .DIN2(_44604), .Q(_44407) );
  nor2s1 _44958_inst ( .DIN1(_44605), .DIN2(_43799), .Q(_44604) );
  xnr2s1 _44959_inst ( .DIN1(_28088), .DIN2(_44606), .Q(_43799) );
  nor2s1 _44960_inst ( .DIN1(_43122), .DIN2(_43313), .Q(_44606) );
  nnd2s1 _44961_inst ( .DIN1(_44607), .DIN2(_44608), .Q(_43313) );
  nor2s1 _44962_inst ( .DIN1(_32080), .DIN2(_27348), .Q(_44607) );
  nnd2s1 _44963_inst ( .DIN1(_44507), .DIN2(_29819), .Q(_27348) );
  hi1s1 _44964_inst ( .DIN(_28115), .Q(_32080) );
  hi1s1 _44965_inst ( .DIN(_44047), .Q(_43122) );
  hi1s1 _44966_inst ( .DIN(_38848), .Q(_28088) );
  nnd2s1 _44967_inst ( .DIN1(_36606), .DIN2(_44376), .Q(_38848) );
  nor2s1 _44968_inst ( .DIN1(_43391), .DIN2(_42312), .Q(_44605) );
  nnd2s1 _44969_inst ( .DIN1(_44609), .DIN2(_44608), .Q(_42312) );
  nor2s1 _44970_inst ( .DIN1(_30964), .DIN2(_44477), .Q(_44608) );
  nor2s1 _44971_inst ( .DIN1(_28114), .DIN2(_27467), .Q(_44609) );
  nnd2s1 _44972_inst ( .DIN1(_44610), .DIN2(_44611), .Q(_28114) );
  nor2s1 _44973_inst ( .DIN1(_53445), .DIN2(_53458), .Q(_44611) );
  nor2s1 _44974_inst ( .DIN1(_26215), .DIN2(_26408), .Q(_44610) );
  nor2s1 _44975_inst ( .DIN1(_44194), .DIN2(_43577), .Q(_44603) );
  nnd2s1 _44976_inst ( .DIN1(_44612), .DIN2(_44613), .Q(_43577) );
  nor2s1 _44977_inst ( .DIN1(_44614), .DIN2(_44615), .Q(_44613) );
  nnd2s1 _44978_inst ( .DIN1(_44616), .DIN2(_44154), .Q(_44615) );
  nnd2s1 _44979_inst ( .DIN1(_44262), .DIN2(_43815), .Q(_44154) );
  xor2s1 _44980_inst ( .DIN1(_43929), .DIN2(_32005), .Q(_43815) );
  and2s1 _44981_inst ( .DIN1(_44617), .DIN2(_44618), .Q(_32005) );
  nor2s1 _44982_inst ( .DIN1(_44031), .DIN2(_44619), .Q(_44618) );
  nnd2s1 _44983_inst ( .DIN1(_40395), .DIN2(_44572), .Q(_44619) );
  nnd2s1 _44984_inst ( .DIN1(_42877), .DIN2(_44620), .Q(_44031) );
  nor2s1 _44985_inst ( .DIN1(_44579), .DIN2(_44621), .Q(_44617) );
  hi1s1 _44986_inst ( .DIN(_44622), .Q(_44621) );
  nnd2s1 _44987_inst ( .DIN1(_44623), .DIN2(_44624), .Q(_44579) );
  nor2s1 _44988_inst ( .DIN1(_44029), .DIN2(_44625), .Q(_44624) );
  hi1s1 _44989_inst ( .DIN(_44626), .Q(_44029) );
  nor2s1 _44990_inst ( .DIN1(_44627), .DIN2(_44628), .Q(_44623) );
  and2s1 _44991_inst ( .DIN1(_44629), .DIN2(_44537), .Q(_44262) );
  nor2s1 _44992_inst ( .DIN1(_31121), .DIN2(_27467), .Q(_44537) );
  nnd2s1 _44993_inst ( .DIN1(_44130), .DIN2(_44480), .Q(_27467) );
  hi1s1 _44994_inst ( .DIN(_44101), .Q(_44130) );
  nor2s1 _44995_inst ( .DIN1(_31702), .DIN2(_44481), .Q(_44629) );
  nnd2s1 _44996_inst ( .DIN1(_44630), .DIN2(_44631), .Q(_44481) );
  nor2s1 _44997_inst ( .DIN1(_53445), .DIN2(_53446), .Q(_44631) );
  nor2s1 _44998_inst ( .DIN1(_26408), .DIN2(_26243), .Q(_44630) );
  nnd2s1 _44999_inst ( .DIN1(_44552), .DIN2(_44056), .Q(_31702) );
  nnd2s1 _45000_inst ( .DIN1(_44018), .DIN2(_43562), .Q(_44616) );
  and2s1 _45001_inst ( .DIN1(_44632), .DIN2(_27342), .Q(_44018) );
  hi1s1 _45002_inst ( .DIN(_27494), .Q(_27342) );
  nnd2s1 _45003_inst ( .DIN1(_44113), .DIN2(_43806), .Q(_27494) );
  hi1s1 _45004_inst ( .DIN(_27474), .Q(_43806) );
  nnd2s1 _45005_inst ( .DIN1(_53453), .DIN2(_26297), .Q(_27474) );
  and2s1 _45006_inst ( .DIN1(_44633), .DIN2(_53455), .Q(_44113) );
  nor2s1 _45007_inst ( .DIN1(_53454), .DIN2(_26214), .Q(_44633) );
  nor2s1 _45008_inst ( .DIN1(_44397), .DIN2(_32340), .Q(_44632) );
  nnd2s1 _45009_inst ( .DIN1(_43807), .DIN2(_44552), .Q(_32340) );
  nnd2s1 _45010_inst ( .DIN1(_29969), .DIN2(_30965), .Q(_44397) );
  nor2s1 _45011_inst ( .DIN1(_43545), .DIN2(_43664), .Q(_44614) );
  nnd2s1 _45012_inst ( .DIN1(_44634), .DIN2(_44452), .Q(_43545) );
  and2s1 _45013_inst ( .DIN1(_44635), .DIN2(_32088), .Q(_44452) );
  nor2s1 _45014_inst ( .DIN1(_44101), .DIN2(_27375), .Q(_44635) );
  nnd2s1 _45015_inst ( .DIN1(_44636), .DIN2(_53454), .Q(_27375) );
  nor2s1 _45016_inst ( .DIN1(_53459), .DIN2(_26465), .Q(_44636) );
  nnd2s1 _45017_inst ( .DIN1(_53452), .DIN2(_26576), .Q(_44101) );
  nor2s1 _45018_inst ( .DIN1(_44477), .DIN2(_30963), .Q(_44634) );
  nnd2s1 _45019_inst ( .DIN1(_43807), .DIN2(_44218), .Q(_44477) );
  nor2s1 _45020_inst ( .DIN1(_26345), .DIN2(_53457), .Q(_43807) );
  nor2s1 _45021_inst ( .DIN1(_43818), .DIN2(_43970), .Q(_44612) );
  nnd2s1 _45022_inst ( .DIN1(_44637), .DIN2(_44638), .Q(_43970) );
  or2s1 _45023_inst ( .DIN1(_43111), .DIN2(_43565), .Q(_44638) );
  nnd2s1 _45024_inst ( .DIN1(_44639), .DIN2(_44583), .Q(_43111) );
  nor2s1 _45025_inst ( .DIN1(_27359), .DIN2(_30848), .Q(_44639) );
  nnd2s1 _45026_inst ( .DIN1(_44640), .DIN2(_44552), .Q(_30848) );
  nor2s1 _45027_inst ( .DIN1(_26387), .DIN2(_53456), .Q(_44552) );
  or2s1 _45028_inst ( .DIN1(_43110), .DIN2(_43514), .Q(_44637) );
  nnd2s1 _45029_inst ( .DIN1(_44641), .DIN2(_44642), .Q(_43110) );
  nor2s1 _45030_inst ( .DIN1(_30963), .DIN2(_44643), .Q(_44642) );
  nor2s1 _45031_inst ( .DIN1(_32339), .DIN2(_30872), .Q(_44641) );
  nnd2s1 _45032_inst ( .DIN1(_44644), .DIN2(_44645), .Q(_43818) );
  nnd2s1 _45033_inst ( .DIN1(_44184), .DIN2(_43562), .Q(_44645) );
  nnd2s1 _45034_inst ( .DIN1(_43151), .DIN2(_43514), .Q(_43562) );
  nnd2s1 _45035_inst ( .DIN1(_26770), .DIN2(_44646), .Q(_43514) );
  nnd2s1 _45036_inst ( .DIN1(_44647), .DIN2(______[19]), .Q(_44646) );
  nor2s1 _45037_inst ( .DIN1(______[1]), .DIN2(_26773), .Q(_44647) );
  nnd2s1 _45038_inst ( .DIN1(_44648), .DIN2(_44341), .Q(_43151) );
  nor2s1 _45039_inst ( .DIN1(______[1]), .DIN2(_44342), .Q(_44648) );
  nor2s1 _45040_inst ( .DIN1(_44649), .DIN2(_44472), .Q(_44184) );
  nnd2s1 _45041_inst ( .DIN1(_30369), .DIN2(_28212), .Q(_44472) );
  hi1s1 _45042_inst ( .DIN(_32081), .Q(_28212) );
  nnd2s1 _45043_inst ( .DIN1(_44650), .DIN2(_44133), .Q(_32081) );
  hi1s1 _45044_inst ( .DIN(_44305), .Q(_44133) );
  nor2s1 _45045_inst ( .DIN1(_53445), .DIN2(_26408), .Q(_44650) );
  hi1s1 _45046_inst ( .DIN(_32010), .Q(_30369) );
  nnd2s1 _45047_inst ( .DIN1(_44640), .DIN2(_44558), .Q(_32010) );
  nnd2s1 _45048_inst ( .DIN1(_30965), .DIN2(_27295), .Q(_44649) );
  hi1s1 _45049_inst ( .DIN(_27359), .Q(_27295) );
  hi1s1 _45050_inst ( .DIN(_31190), .Q(_30965) );
  nnd2s1 _45051_inst ( .DIN1(_44651), .DIN2(_53444), .Q(_31190) );
  nor2s1 _45052_inst ( .DIN1(_53448), .DIN2(_26428), .Q(_44651) );
  nnd2s1 _45053_inst ( .DIN1(_44026), .DIN2(_43363), .Q(_44644) );
  nnd2s1 _45054_inst ( .DIN1(_43371), .DIN2(_43520), .Q(_43363) );
  nnd2s1 _45055_inst ( .DIN1(_26770), .DIN2(_44652), .Q(_43520) );
  nnd2s1 _45056_inst ( .DIN1(_44653), .DIN2(_44342), .Q(_44652) );
  hi1s1 _45057_inst ( .DIN(_43186), .Q(_43371) );
  xnr2s1 _45058_inst ( .DIN1(_26321), .DIN2(_43725), .Q(_43186) );
  nor2s1 _45059_inst ( .DIN1(_44654), .DIN2(_44519), .Q(_43725) );
  nnd2s1 _45060_inst ( .DIN1(_44343), .DIN2(_44342), .Q(_44654) );
  and2s1 _45061_inst ( .DIN1(_44655), .DIN2(_44583), .Q(_44026) );
  xor2s1 _45062_inst ( .DIN1(_44656), .DIN2(_32548), .Q(_44583) );
  hi1s1 _45063_inst ( .DIN(_27413), .Q(_32548) );
  nnd2s1 _45064_inst ( .DIN1(_40991), .DIN2(_44657), .Q(_27413) );
  hi1s1 _45065_inst ( .DIN(_34235), .Q(_40991) );
  nnd2s1 _45066_inst ( .DIN1(_44658), .DIN2(_44078), .Q(_34235) );
  nnd2s1 _45067_inst ( .DIN1(_29969), .DIN2(_28909), .Q(_44656) );
  hi1s1 _45068_inst ( .DIN(_28864), .Q(_28909) );
  nnd2s1 _45069_inst ( .DIN1(_44659), .DIN2(_53451), .Q(_28864) );
  nor2s1 _45070_inst ( .DIN1(_53444), .DIN2(_26227), .Q(_44659) );
  hi1s1 _45071_inst ( .DIN(_28169), .Q(_29969) );
  nnd2s1 _45072_inst ( .DIN1(_44660), .DIN2(_53446), .Q(_28169) );
  nor2s1 _45073_inst ( .DIN1(_53458), .DIN2(_44533), .Q(_44660) );
  nor2s1 _45074_inst ( .DIN1(_30849), .DIN2(_27359), .Q(_44655) );
  nnd2s1 _45075_inst ( .DIN1(_44507), .DIN2(_44444), .Q(_27359) );
  hi1s1 _45076_inst ( .DIN(_44099), .Q(_44444) );
  and2s1 _45077_inst ( .DIN1(_44591), .DIN2(_26214), .Q(_44507) );
  nor2s1 _45078_inst ( .DIN1(_53454), .DIN2(_53455), .Q(_44591) );
  nnd2s1 _45079_inst ( .DIN1(_44056), .DIN2(_44558), .Q(_30849) );
  nor2s1 _45080_inst ( .DIN1(_26262), .DIN2(_53447), .Q(_44558) );
  nor2s1 _45081_inst ( .DIN1(_53457), .DIN2(_53450), .Q(_44056) );
  nnd2s1 _45082_inst ( .DIN1(_44661), .DIN2(_44662), .Q(_44194) );
  nnd2s1 _45083_inst ( .DIN1(_43845), .DIN2(_44047), .Q(_44662) );
  nnd2s1 _45084_inst ( .DIN1(_43664), .DIN2(_43166), .Q(_44047) );
  nnd2s1 _45085_inst ( .DIN1(_44663), .DIN2(_44341), .Q(_43166) );
  nor2s1 _45086_inst ( .DIN1(_26773), .DIN2(_43565), .Q(_44341) );
  nor2s1 _45087_inst ( .DIN1(______[19]), .DIN2(_44343), .Q(_44663) );
  hi1s1 _45088_inst ( .DIN(______[1]), .Q(_44343) );
  nnd2s1 _45089_inst ( .DIN1(_26770), .DIN2(_44664), .Q(_43664) );
  nnd2s1 _45090_inst ( .DIN1(_44665), .DIN2(______[1]), .Q(_44664) );
  nor2s1 _45091_inst ( .DIN1(______[19]), .DIN2(_26773), .Q(_44665) );
  nor2s1 _45092_inst ( .DIN1(_44643), .DIN2(_43811), .Q(_43845) );
  nnd2s1 _45093_inst ( .DIN1(_44451), .DIN2(_28115), .Q(_43811) );
  nor2s1 _45094_inst ( .DIN1(_44305), .DIN2(_44557), .Q(_28115) );
  nnd2s1 _45095_inst ( .DIN1(_53458), .DIN2(_53446), .Q(_44305) );
  nor2s1 _45096_inst ( .DIN1(_30964), .DIN2(_30677), .Q(_44451) );
  nnd2s1 _45097_inst ( .DIN1(_44666), .DIN2(_53448), .Q(_30964) );
  nor2s1 _45098_inst ( .DIN1(_53444), .DIN2(_53451), .Q(_44666) );
  hi1s1 _45099_inst ( .DIN(_29820), .Q(_44643) );
  nor2s1 _45100_inst ( .DIN1(_44099), .DIN2(_27475), .Q(_29820) );
  nnd2s1 _45101_inst ( .DIN1(_44667), .DIN2(_53454), .Q(_27475) );
  nor2s1 _45102_inst ( .DIN1(_53455), .DIN2(_26214), .Q(_44667) );
  nnd2s1 _45103_inst ( .DIN1(_53453), .DIN2(_53452), .Q(_44099) );
  nor2s1 _45104_inst ( .DIN1(_43316), .DIN2(_43772), .Q(_44661) );
  nor2s1 _45105_inst ( .DIN1(_43929), .DIN2(_43876), .Q(_43772) );
  nnd2s1 _45106_inst ( .DIN1(_44668), .DIN2(_44669), .Q(_43876) );
  nor2s1 _45107_inst ( .DIN1(_31121), .DIN2(_29351), .Q(_44669) );
  nnd2s1 _45108_inst ( .DIN1(_29819), .DIN2(_44480), .Q(_29351) );
  hi1s1 _45109_inst ( .DIN(_44098), .Q(_44480) );
  nnd2s1 _45110_inst ( .DIN1(_44670), .DIN2(_53454), .Q(_44098) );
  nor2s1 _45111_inst ( .DIN1(_26214), .DIN2(_26465), .Q(_44670) );
  nnd2s1 _45112_inst ( .DIN1(_44671), .DIN2(_53451), .Q(_31121) );
  nor2s1 _45113_inst ( .DIN1(_32339), .DIN2(_30875), .Q(_44668) );
  hi1s1 _45114_inst ( .DIN(_32088), .Q(_30875) );
  nor2s1 _45115_inst ( .DIN1(_44139), .DIN2(_44533), .Q(_32088) );
  nnd2s1 _45116_inst ( .DIN1(_26408), .DIN2(_26207), .Q(_44533) );
  nnd2s1 _45117_inst ( .DIN1(_44672), .DIN2(_44217), .Q(_32339) );
  nor2s1 _45118_inst ( .DIN1(_26353), .DIN2(_53450), .Q(_44217) );
  nor2s1 _45119_inst ( .DIN1(_26262), .DIN2(_26387), .Q(_44672) );
  nnd2s1 _45120_inst ( .DIN1(_26770), .DIN2(_44673), .Q(_43929) );
  nnd2s1 _45121_inst ( .DIN1(_44674), .DIN2(______[1]), .Q(_44673) );
  nor2s1 _45122_inst ( .DIN1(______[28]), .DIN2(_44342), .Q(_44674) );
  hi1s1 _45123_inst ( .DIN(______[19]), .Q(_44342) );
  and2s1 _45124_inst ( .DIN1(_43227), .DIN2(_43336), .Q(_43316) );
  hi1s1 _45125_inst ( .DIN(_43391), .Q(_43336) );
  xor2s1 _45126_inst ( .DIN1(_44675), .DIN2(_36606), .Q(_43391) );
  hi1s1 _45127_inst ( .DIN(_26998), .Q(_36606) );
  nnd2s1 _45128_inst ( .DIN1(_43233), .DIN2(_43226), .Q(_44675) );
  nnd2s1 _45129_inst ( .DIN1(_44676), .DIN2(______[19]), .Q(_43226) );
  nor2s1 _45130_inst ( .DIN1(______[1]), .DIN2(_44519), .Q(_44676) );
  nnd2s1 _45131_inst ( .DIN1(_26774), .DIN2(_26770), .Q(_44519) );
  nnd2s1 _45132_inst ( .DIN1(_26770), .DIN2(_44677), .Q(_43233) );
  nnd2s1 _45133_inst ( .DIN1(_44653), .DIN2(______[19]), .Q(_44677) );
  nor2s1 _45134_inst ( .DIN1(______[28]), .DIN2(______[1]), .Q(_44653) );
  and2s1 _45135_inst ( .DIN1(_44678), .DIN2(_44487), .Q(_43227) );
  nor2s1 _45136_inst ( .DIN1(_29481), .DIN2(_30963), .Q(_44487) );
  nnd2s1 _45137_inst ( .DIN1(_44671), .DIN2(_26428), .Q(_30963) );
  nor2s1 _45138_inst ( .DIN1(_53444), .DIN2(_53448), .Q(_44671) );
  nnd2s1 _45139_inst ( .DIN1(_44520), .DIN2(_29819), .Q(_29481) );
  hi1s1 _45140_inst ( .DIN(_27374), .Q(_29819) );
  nnd2s1 _45141_inst ( .DIN1(_26297), .DIN2(_26576), .Q(_27374) );
  and2s1 _45142_inst ( .DIN1(_44679), .DIN2(_53455), .Q(_44520) );
  nor2s1 _45143_inst ( .DIN1(_53454), .DIN2(_53459), .Q(_44679) );
  nor2s1 _45144_inst ( .DIN1(_30677), .DIN2(_30872), .Q(_44678) );
  hi1s1 _45145_inst ( .DIN(_27977), .Q(_30872) );
  nor2s1 _45146_inst ( .DIN1(_44139), .DIN2(_44557), .Q(_27977) );
  nnd2s1 _45147_inst ( .DIN1(_53445), .DIN2(_53449), .Q(_44557) );
  nnd2s1 _45148_inst ( .DIN1(_26215), .DIN2(_26243), .Q(_44139) );
  nnd2s1 _45149_inst ( .DIN1(_44218), .DIN2(_44640), .Q(_30677) );
  hi1s1 _45150_inst ( .DIN(_44102), .Q(_44640) );
  nnd2s1 _45151_inst ( .DIN1(_53450), .DIN2(_53457), .Q(_44102) );
  nor2s1 _45152_inst ( .DIN1(_53447), .DIN2(_53456), .Q(_44218) );
  nor2s1 _45153_inst ( .DIN1(_43203), .DIN2(_44680), .Q(_44327) );
  nor2s1 _45154_inst ( .DIN1(_27082), .DIN2(_44681), .Q(_44680) );
  nnd2s1 _45155_inst ( .DIN1(_44682), .DIN2(_44683), .Q(_44681) );
  nnd2s1 _45156_inst ( .DIN1(_44684), .DIN2(_26214), .Q(_44683) );
  nnd2s1 _45157_inst ( .DIN1(_53451), .DIN2(_53458), .Q(_44684) );
  nnd2s1 _45158_inst ( .DIN1(_43301), .DIN2(_53451), .Q(_44682) );
  nor2s1 _45159_inst ( .DIN1(_26243), .DIN2(_26214), .Q(_43301) );
  hi1s1 _45160_inst ( .DIN(_43174), .Q(_43203) );
  nnd2s1 _45161_inst ( .DIN1(_44685), .DIN2(_44686), .Q(_43174) );
  nor2s1 _45162_inst ( .DIN1(_27309), .DIN2(_31396), .Q(_44686) );
  nor2s1 _45163_inst ( .DIN1(_44687), .DIN2(_43498), .Q(_44685) );
  nnd2s1 _45164_inst ( .DIN1(_44688), .DIN2(_27445), .Q(_43498) );
  nor2s1 _45165_inst ( .DIN1(_27316), .DIN2(_42131), .Q(_44688) );
  nnd2s1 _45166_inst ( .DIN1(_44689), .DIN2(_44690), .Q(
        ____0___________0_9_____) );
  nnd2s1 _45167_inst ( .DIN1(_44691), .DIN2(_44692), .Q(_44690) );
  nor2s1 _45168_inst ( .DIN1(_44693), .DIN2(_28100), .Q(_44691) );
  xor2s1 _45169_inst ( .DIN1(_44694), .DIN2(_53478), .Q(_44693) );
  nnd2s1 _45170_inst ( .DIN1(_53477), .DIN2(_53472), .Q(_44694) );
  nnd2s1 _45171_inst ( .DIN1(_39842), .DIN2(_44695), .Q(_44689) );
  nnd2s1 _45172_inst ( .DIN1(_44696), .DIN2(_44697), .Q(_44695) );
  nor2s1 _45173_inst ( .DIN1(_44698), .DIN2(_44699), .Q(_44697) );
  nnd2s1 _45174_inst ( .DIN1(_44700), .DIN2(_44701), .Q(_44699) );
  hi1s1 _45175_inst ( .DIN(_44702), .Q(_44701) );
  nor2s1 _45176_inst ( .DIN1(_44703), .DIN2(_44704), .Q(_44700) );
  xor2s1 _45177_inst ( .DIN1(_33865), .DIN2(_44705), .Q(_44703) );
  nor2s1 _45178_inst ( .DIN1(_44706), .DIN2(_44707), .Q(_44705) );
  nnd2s1 _45179_inst ( .DIN1(_44708), .DIN2(_44709), .Q(_44698) );
  nor2s1 _45180_inst ( .DIN1(_44710), .DIN2(_44711), .Q(_44709) );
  nor2s1 _45181_inst ( .DIN1(_44712), .DIN2(_44713), .Q(_44708) );
  nor2s1 _45182_inst ( .DIN1(_26767), .DIN2(_44714), .Q(_44713) );
  nor2s1 _45183_inst ( .DIN1(_44715), .DIN2(_44716), .Q(_44712) );
  nor2s1 _45184_inst ( .DIN1(_44717), .DIN2(_44718), .Q(_44696) );
  nnd2s1 _45185_inst ( .DIN1(_44719), .DIN2(_44720), .Q(_44718) );
  nor2s1 _45186_inst ( .DIN1(_44721), .DIN2(_44722), .Q(_44720) );
  nor2s1 _45187_inst ( .DIN1(_44723), .DIN2(_44724), .Q(_44722) );
  nor2s1 _45188_inst ( .DIN1(_26805), .DIN2(_44726), .Q(_44721) );
  nor2s1 _45189_inst ( .DIN1(_44727), .DIN2(_44728), .Q(_44719) );
  xor2s1 _45190_inst ( .DIN1(_31752), .DIN2(_44729), .Q(_44728) );
  nor2s1 _45191_inst ( .DIN1(_44730), .DIN2(_44731), .Q(_44729) );
  hi1s1 _45192_inst ( .DIN(_29450), .Q(_31752) );
  nnd2s1 _45193_inst ( .DIN1(_44732), .DIN2(_44376), .Q(_29450) );
  nnd2s1 _45194_inst ( .DIN1(_44733), .DIN2(_44734), .Q(_44717) );
  nor2s1 _45195_inst ( .DIN1(_44735), .DIN2(_44736), .Q(_44734) );
  nor2s1 _45196_inst ( .DIN1(_44737), .DIN2(_44738), .Q(_44733) );
  nnd2s1 _45197_inst ( .DIN1(_44739), .DIN2(_44740), .Q(
        ____0___________0_8_____) );
  nnd2s1 _45198_inst ( .DIN1(_44741), .DIN2(_44692), .Q(_44740) );
  nor2s1 _45199_inst ( .DIN1(_44742), .DIN2(_26771), .Q(_44741) );
  xor2s1 _45200_inst ( .DIN1(_26585), .DIN2(_53472), .Q(_44742) );
  nnd2s1 _45201_inst ( .DIN1(_39842), .DIN2(_44743), .Q(_44739) );
  nnd2s1 _45202_inst ( .DIN1(_44744), .DIN2(_44745), .Q(_44743) );
  nor2s1 _45203_inst ( .DIN1(_44746), .DIN2(_44747), .Q(_44745) );
  nnd2s1 _45204_inst ( .DIN1(_44748), .DIN2(_44749), .Q(_44747) );
  nor2s1 _45205_inst ( .DIN1(_44750), .DIN2(_44737), .Q(_44749) );
  nnd2s1 _45206_inst ( .DIN1(_44751), .DIN2(_44752), .Q(_44737) );
  nor2s1 _45207_inst ( .DIN1(_44753), .DIN2(_44754), .Q(_44752) );
  nnd2s1 _45208_inst ( .DIN1(_44755), .DIN2(_44756), .Q(_44754) );
  nor2s1 _45209_inst ( .DIN1(_44757), .DIN2(_44758), .Q(_44751) );
  nor2s1 _45210_inst ( .DIN1(_26766), .DIN2(_44759), .Q(_44758) );
  nor2s1 _45211_inst ( .DIN1(_26845), .DIN2(_44761), .Q(_44750) );
  nor2s1 _45212_inst ( .DIN1(_44762), .DIN2(_44763), .Q(_44748) );
  nnd2s1 _45213_inst ( .DIN1(_44764), .DIN2(_44765), .Q(_44746) );
  nor2s1 _45214_inst ( .DIN1(_44766), .DIN2(_44767), .Q(_44765) );
  nor2s1 _45215_inst ( .DIN1(_44768), .DIN2(_44769), .Q(_44764) );
  nor2s1 _45216_inst ( .DIN1(_44770), .DIN2(_44771), .Q(_44769) );
  nor2s1 _45217_inst ( .DIN1(_44772), .DIN2(_44773), .Q(_44770) );
  nor2s1 _45218_inst ( .DIN1(_44774), .DIN2(_44775), .Q(_44744) );
  nnd2s1 _45219_inst ( .DIN1(_44776), .DIN2(_44777), .Q(_44775) );
  nor2s1 _45220_inst ( .DIN1(_44778), .DIN2(_44779), .Q(_44777) );
  nor2s1 _45221_inst ( .DIN1(_44780), .DIN2(_44781), .Q(_44776) );
  nnd2s1 _45222_inst ( .DIN1(_44782), .DIN2(_44783), .Q(_44781) );
  or2s1 _45223_inst ( .DIN1(_44784), .DIN2(_26766), .Q(_44783) );
  nnd2s1 _45224_inst ( .DIN1(_44785), .DIN2(_26766), .Q(_44782) );
  nnd2s1 _45225_inst ( .DIN1(_44786), .DIN2(_44787), .Q(_44774) );
  nor2s1 _45226_inst ( .DIN1(_44788), .DIN2(_44789), .Q(_44787) );
  nor2s1 _45227_inst ( .DIN1(_44790), .DIN2(_44791), .Q(_44786) );
  nor2s1 _45228_inst ( .DIN1(_44792), .DIN2(_27235), .Q(
        ____0___________0_7_____) );
  nor2s1 _45229_inst ( .DIN1(_44793), .DIN2(_44794), .Q(_44792) );
  nnd2s1 _45230_inst ( .DIN1(_44795), .DIN2(_44796), .Q(_44794) );
  nor2s1 _45231_inst ( .DIN1(_44797), .DIN2(_44798), .Q(_44796) );
  nnd2s1 _45232_inst ( .DIN1(_44799), .DIN2(_44800), .Q(_44798) );
  nnd2s1 _45233_inst ( .DIN1(_44801), .DIN2(_44802), .Q(_44797) );
  hi1s1 _45234_inst ( .DIN(_44803), .Q(_44802) );
  nor2s1 _45235_inst ( .DIN1(_44804), .DIN2(_26765), .Q(_44801) );
  nor2s1 _45236_inst ( .DIN1(_44715), .DIN2(_44805), .Q(_44804) );
  nor2s1 _45237_inst ( .DIN1(_44806), .DIN2(_44807), .Q(_44795) );
  nnd2s1 _45238_inst ( .DIN1(_44808), .DIN2(_44809), .Q(_44807) );
  hi1s1 _45239_inst ( .DIN(_44810), .Q(_44808) );
  or2s1 _45240_inst ( .DIN1(_44811), .DIN2(_44812), .Q(_44806) );
  nnd2s1 _45241_inst ( .DIN1(_44813), .DIN2(_44814), .Q(_44793) );
  nor2s1 _45242_inst ( .DIN1(_44815), .DIN2(_44816), .Q(_44814) );
  nnd2s1 _45243_inst ( .DIN1(_44817), .DIN2(_44818), .Q(_44816) );
  nnd2s1 _45244_inst ( .DIN1(_44819), .DIN2(_44820), .Q(_44815) );
  nor2s1 _45245_inst ( .DIN1(_44821), .DIN2(_44822), .Q(_44819) );
  nor2s1 _45246_inst ( .DIN1(_44823), .DIN2(_44824), .Q(_44813) );
  nnd2s1 _45247_inst ( .DIN1(_44825), .DIN2(_44826), .Q(_44824) );
  nnd2s1 _45248_inst ( .DIN1(_44827), .DIN2(_44828), .Q(_44823) );
  nor2s1 _45249_inst ( .DIN1(_44829), .DIN2(_27235), .Q(
        ____0___________0_6_____) );
  nor2s1 _45250_inst ( .DIN1(_44830), .DIN2(_44831), .Q(_44829) );
  nnd2s1 _45251_inst ( .DIN1(_44832), .DIN2(_44833), .Q(_44831) );
  nor2s1 _45252_inst ( .DIN1(_44834), .DIN2(_44835), .Q(_44833) );
  nnd2s1 _45253_inst ( .DIN1(_44836), .DIN2(_44837), .Q(_44835) );
  nor2s1 _45254_inst ( .DIN1(_44838), .DIN2(_44839), .Q(_44832) );
  nnd2s1 _45255_inst ( .DIN1(_44840), .DIN2(_44841), .Q(_44830) );
  nor2s1 _45256_inst ( .DIN1(_44842), .DIN2(_44843), .Q(_44841) );
  nnd2s1 _45257_inst ( .DIN1(_44844), .DIN2(_44845), .Q(_44843) );
  hi1s1 _45258_inst ( .DIN(_44738), .Q(_44845) );
  nnd2s1 _45259_inst ( .DIN1(_44846), .DIN2(_44847), .Q(_44738) );
  nor2s1 _45260_inst ( .DIN1(_44848), .DIN2(_44849), .Q(_44847) );
  nor2s1 _45261_inst ( .DIN1(_26767), .DIN2(_44850), .Q(_44849) );
  nor2s1 _45262_inst ( .DIN1(_44851), .DIN2(_26765), .Q(_44850) );
  nor2s1 _45263_inst ( .DIN1(_44852), .DIN2(_44853), .Q(_44846) );
  nor2s1 _45264_inst ( .DIN1(_44854), .DIN2(_26845), .Q(_44853) );
  nor2s1 _45265_inst ( .DIN1(_44715), .DIN2(_44855), .Q(_44852) );
  and2s1 _45266_inst ( .DIN1(_44856), .DIN2(_44857), .Q(_44855) );
  nor2s1 _45267_inst ( .DIN1(_44811), .DIN2(_44858), .Q(_44840) );
  nor2s1 _45268_inst ( .DIN1(_44859), .DIN2(_39166), .Q(
        ____0___________0_5_____) );
  nnd2s1 _45269_inst ( .DIN1(_35720), .DIN2(_35721), .Q(_39166) );
  nor2s1 _45270_inst ( .DIN1(_44860), .DIN2(_44861), .Q(_44859) );
  nnd2s1 _45271_inst ( .DIN1(_44862), .DIN2(_44863), .Q(_44861) );
  nor2s1 _45272_inst ( .DIN1(_44864), .DIN2(_44865), .Q(_44863) );
  nnd2s1 _45273_inst ( .DIN1(_44866), .DIN2(_44867), .Q(_44865) );
  hi1s1 _45274_inst ( .DIN(_44868), .Q(_44866) );
  nnd2s1 _45275_inst ( .DIN1(_44869), .DIN2(_44870), .Q(_44864) );
  nnd2s1 _45276_inst ( .DIN1(_44871), .DIN2(_26767), .Q(_44870) );
  hi1s1 _45277_inst ( .DIN(_44872), .Q(_44869) );
  nor2s1 _45278_inst ( .DIN1(_44873), .DIN2(_44874), .Q(_44862) );
  nnd2s1 _45279_inst ( .DIN1(_44875), .DIN2(_44876), .Q(_44874) );
  hi1s1 _45280_inst ( .DIN(_44877), .Q(_44876) );
  nnd2s1 _45281_inst ( .DIN1(_44878), .DIN2(_44879), .Q(_44873) );
  nnd2s1 _45282_inst ( .DIN1(_26805), .DIN2(_44880), .Q(_44879) );
  nnd2s1 _45283_inst ( .DIN1(_44881), .DIN2(_26804), .Q(_44878) );
  nnd2s1 _45284_inst ( .DIN1(_44882), .DIN2(_44883), .Q(_44881) );
  nor2s1 _45285_inst ( .DIN1(_44884), .DIN2(_44885), .Q(_44882) );
  nnd2s1 _45286_inst ( .DIN1(_44886), .DIN2(_44887), .Q(_44860) );
  nor2s1 _45287_inst ( .DIN1(_44888), .DIN2(_44889), .Q(_44887) );
  nnd2s1 _45288_inst ( .DIN1(_44890), .DIN2(_44891), .Q(_44889) );
  nnd2s1 _45289_inst ( .DIN1(_44892), .DIN2(_44893), .Q(_44888) );
  nor2s1 _45290_inst ( .DIN1(_44894), .DIN2(_44895), .Q(_44886) );
  nnd2s1 _45291_inst ( .DIN1(_44896), .DIN2(_44897), .Q(_44895) );
  nnd2s1 _45292_inst ( .DIN1(_44715), .DIN2(_44898), .Q(_44896) );
  nnd2s1 _45293_inst ( .DIN1(_44899), .DIN2(_44827), .Q(_44898) );
  nor2s1 _45294_inst ( .DIN1(_44900), .DIN2(_26845), .Q(_44894) );
  nor2s1 _45295_inst ( .DIN1(_44711), .DIN2(_44901), .Q(_44900) );
  nnd2s1 _45296_inst ( .DIN1(_44902), .DIN2(_28073), .Q(
        ____0___________0_4_____) );
  nnd2s1 _45297_inst ( .DIN1(_27235), .DIN2(_28976), .Q(_28073) );
  nor2s1 _45298_inst ( .DIN1(_44903), .DIN2(_44904), .Q(_44902) );
  nor2s1 _45299_inst ( .DIN1(_27235), .DIN2(_44905), .Q(_44904) );
  nnd2s1 _45300_inst ( .DIN1(_44906), .DIN2(_44907), .Q(_44905) );
  nor2s1 _45301_inst ( .DIN1(_44908), .DIN2(_44909), .Q(_44907) );
  nnd2s1 _45302_inst ( .DIN1(_26317), .DIN2(_44910), .Q(_44909) );
  nnd2s1 _45303_inst ( .DIN1(_26805), .DIN2(_44911), .Q(_44910) );
  nnd2s1 _45304_inst ( .DIN1(_44912), .DIN2(_44724), .Q(_44911) );
  nnd2s1 _45305_inst ( .DIN1(_44913), .DIN2(_44914), .Q(_44908) );
  nor2s1 _45306_inst ( .DIN1(_44915), .DIN2(_44916), .Q(_44906) );
  or2s1 _45307_inst ( .DIN1(_44917), .DIN2(_44918), .Q(_44916) );
  nnd2s1 _45308_inst ( .DIN1(_44919), .DIN2(_44867), .Q(_44915) );
  nor2s1 _45309_inst ( .DIN1(_44920), .DIN2(_44921), .Q(_44919) );
  xor2s1 _45310_inst ( .DIN1(_26998), .DIN2(_44922), .Q(_44920) );
  nor2s1 _45311_inst ( .DIN1(_44799), .DIN2(_44771), .Q(_44922) );
  nor2s1 _45312_inst ( .DIN1(_44923), .DIN2(_44924), .Q(_44799) );
  nnd2s1 _45313_inst ( .DIN1(_27093), .DIN2(_44925), .Q(_26998) );
  hi1s1 _45314_inst ( .DIN(_28613), .Q(_27093) );
  nnd2s1 _45315_inst ( .DIN1(_44926), .DIN2(_44732), .Q(_28613) );
  nor2s1 _45316_inst ( .DIN1(_44927), .DIN2(_44928), .Q(_44732) );
  and2s1 _45317_inst ( .DIN1(_44929), .DIN2(_44378), .Q(_44926) );
  nor2s1 _45318_inst ( .DIN1(_27325), .DIN2(_44930), .Q(_44903) );
  nor2s1 _45319_inst ( .DIN1(_44931), .DIN2(_28684), .Q(_44930) );
  xor2s1 _45320_inst ( .DIN1(_26507), .DIN2(_53501), .Q(_44931) );
  hi1s1 _45321_inst ( .DIN(_27235), .Q(_27325) );
  nnd2s1 _45322_inst ( .DIN1(_44932), .DIN2(_44933), .Q(
        ____0___________0_3_____) );
  nor2s1 _45323_inst ( .DIN1(_44934), .DIN2(_44935), .Q(_44933) );
  nor2s1 _45324_inst ( .DIN1(_28032), .DIN2(_44936), .Q(_44935) );
  nnd2s1 _45325_inst ( .DIN1(_44937), .DIN2(_44938), .Q(_44936) );
  nor2s1 _45326_inst ( .DIN1(_44939), .DIN2(_44940), .Q(_44938) );
  nnd2s1 _45327_inst ( .DIN1(_44941), .DIN2(_44942), .Q(_44940) );
  nor2s1 _45328_inst ( .DIN1(_44943), .DIN2(_44944), .Q(_44942) );
  nnd2s1 _45329_inst ( .DIN1(_44945), .DIN2(_44946), .Q(_44944) );
  nnd2s1 _45330_inst ( .DIN1(_44947), .DIN2(_44948), .Q(_44943) );
  nnd2s1 _45331_inst ( .DIN1(_44949), .DIN2(_26845), .Q(_44948) );
  nnd2s1 _45332_inst ( .DIN1(_44950), .DIN2(_44951), .Q(_44947) );
  nor2s1 _45333_inst ( .DIN1(_44727), .DIN2(_44952), .Q(_44941) );
  nnd2s1 _45334_inst ( .DIN1(_44953), .DIN2(_44954), .Q(_44727) );
  and2s1 _45335_inst ( .DIN1(_44955), .DIN2(_44893), .Q(_44954) );
  nor2s1 _45336_inst ( .DIN1(_44956), .DIN2(_44880), .Q(_44953) );
  nor2s1 _45337_inst ( .DIN1(_44957), .DIN2(_44958), .Q(_44956) );
  nnd2s1 _45338_inst ( .DIN1(_44959), .DIN2(_44960), .Q(_44939) );
  nor2s1 _45339_inst ( .DIN1(_44961), .DIN2(_44962), .Q(_44960) );
  nnd2s1 _45340_inst ( .DIN1(_44963), .DIN2(_44964), .Q(_44962) );
  nor2s1 _45341_inst ( .DIN1(_44965), .DIN2(_44966), .Q(_44959) );
  nor2s1 _45342_inst ( .DIN1(_44967), .DIN2(_44968), .Q(_44937) );
  nnd2s1 _45343_inst ( .DIN1(_44969), .DIN2(_44970), .Q(_44968) );
  nor2s1 _45344_inst ( .DIN1(_44834), .DIN2(_44971), .Q(_44970) );
  nnd2s1 _45345_inst ( .DIN1(_44972), .DIN2(_44973), .Q(_44834) );
  xor2s1 _45346_inst ( .DIN1(_44974), .DIN2(_29490), .Q(_44973) );
  hi1s1 _45347_inst ( .DIN(_27346), .Q(_29490) );
  nnd2s1 _45348_inst ( .DIN1(_44975), .DIN2(_44976), .Q(_27346) );
  nor2s1 _45349_inst ( .DIN1(_44286), .DIN2(_44977), .Q(_44976) );
  nor2s1 _45350_inst ( .DIN1(_44314), .DIN2(_42798), .Q(_44975) );
  nnd2s1 _45351_inst ( .DIN1(_44978), .DIN2(_44979), .Q(_42798) );
  nor2s1 _45352_inst ( .DIN1(_44980), .DIN2(_44981), .Q(_44979) );
  nor2s1 _45353_inst ( .DIN1(_44982), .DIN2(_44983), .Q(_44978) );
  nnd2s1 _45354_inst ( .DIN1(_44984), .DIN2(_44985), .Q(_44983) );
  nnd2s1 _45355_inst ( .DIN1(_44986), .DIN2(_44892), .Q(_44974) );
  nor2s1 _45356_inst ( .DIN1(_44987), .DIN2(_44885), .Q(_44986) );
  xor2s1 _45357_inst ( .DIN1(_44988), .DIN2(_29049), .Q(_44972) );
  nor2s1 _45358_inst ( .DIN1(_44989), .DIN2(_44032), .Q(_29049) );
  nnd2s1 _45359_inst ( .DIN1(_44990), .DIN2(_44991), .Q(_44032) );
  nor2s1 _45360_inst ( .DIN1(_44992), .DIN2(_44993), .Q(_44991) );
  nnd2s1 _45361_inst ( .DIN1(_44994), .DIN2(_42876), .Q(_44993) );
  nnd2s1 _45362_inst ( .DIN1(_44995), .DIN2(_44573), .Q(_44992) );
  nor2s1 _45363_inst ( .DIN1(_40398), .DIN2(_44996), .Q(_44990) );
  nnd2s1 _45364_inst ( .DIN1(_44997), .DIN2(_44998), .Q(_44996) );
  nnd2s1 _45365_inst ( .DIN1(_42881), .DIN2(_44999), .Q(_40398) );
  and2s1 _45366_inst ( .DIN1(_45000), .DIN2(_45001), .Q(_42881) );
  nnd2s1 _45367_inst ( .DIN1(_45002), .DIN2(_44576), .Q(_44989) );
  nnd2s1 _45368_inst ( .DIN1(_45003), .DIN2(_45004), .Q(_44988) );
  nnd2s1 _45369_inst ( .DIN1(_45005), .DIN2(_26845), .Q(_45004) );
  nor2s1 _45370_inst ( .DIN1(_45006), .DIN2(_45007), .Q(_44969) );
  nnd2s1 _45371_inst ( .DIN1(_45008), .DIN2(_45009), .Q(_44967) );
  nor2s1 _45372_inst ( .DIN1(_45010), .DIN2(_44812), .Q(_45009) );
  nor2s1 _45373_inst ( .DIN1(_45011), .DIN2(_45012), .Q(_45008) );
  nor2s1 _45374_inst ( .DIN1(_28037), .DIN2(_45013), .Q(_44934) );
  nnd2s1 _45375_inst ( .DIN1(_53462), .DIN2(_28040), .Q(_45013) );
  nor2s1 _45376_inst ( .DIN1(_28041), .DIN2(_45014), .Q(_44932) );
  nor2s1 _45377_inst ( .DIN1(_53462), .DIN2(_28043), .Q(_45014) );
  hi1s1 _45378_inst ( .DIN(_32954), .Q(_28043) );
  nor2s1 _45379_inst ( .DIN1(_28040), .DIN2(_28037), .Q(_32954) );
  hi1s1 _45380_inst ( .DIN(_28032), .Q(_28037) );
  nnd2s1 _45381_inst ( .DIN1(_53464), .DIN2(_53463), .Q(_28040) );
  hi1s1 _45382_inst ( .DIN(_30112), .Q(_28041) );
  nnd2s1 _45383_inst ( .DIN1(_28032), .DIN2(_28976), .Q(_30112) );
  nnd2s1 _45384_inst ( .DIN1(_28976), .DIN2(_29221), .Q(_28032) );
  nor2s1 _45385_inst ( .DIN1(_45015), .DIN2(_27235), .Q(
        ____0___________0_2_____) );
  nnd2s1 _45386_inst ( .DIN1(_27994), .DIN2(_28976), .Q(_27235) );
  xor2s1 _45387_inst ( .DIN1(_31768), .DIN2(_45016), .Q(_45015) );
  nor2s1 _45388_inst ( .DIN1(_45017), .DIN2(_45018), .Q(_45016) );
  nnd2s1 _45389_inst ( .DIN1(_45019), .DIN2(_45020), .Q(_45018) );
  nor2s1 _45390_inst ( .DIN1(_44918), .DIN2(_45021), .Q(_45020) );
  or2s1 _45391_inst ( .DIN1(_44762), .DIN2(_45022), .Q(_45021) );
  hi1s1 _45392_inst ( .DIN(_45023), .Q(_44762) );
  nnd2s1 _45393_inst ( .DIN1(_45024), .DIN2(_45025), .Q(_44918) );
  nor2s1 _45394_inst ( .DIN1(_45026), .DIN2(_45027), .Q(_45025) );
  nnd2s1 _45395_inst ( .DIN1(_45028), .DIN2(_45029), .Q(_45027) );
  nnd2s1 _45396_inst ( .DIN1(_45030), .DIN2(_44723), .Q(_45029) );
  nnd2s1 _45397_inst ( .DIN1(_45031), .DIN2(_45032), .Q(_45026) );
  nor2s1 _45398_inst ( .DIN1(_45033), .DIN2(_45034), .Q(_45024) );
  nnd2s1 _45399_inst ( .DIN1(_45035), .DIN2(_45036), .Q(_45034) );
  or2s1 _45400_inst ( .DIN1(_45037), .DIN2(_44789), .Q(_45033) );
  nnd2s1 _45401_inst ( .DIN1(_45038), .DIN2(_45039), .Q(_44789) );
  nor2s1 _45402_inst ( .DIN1(_45040), .DIN2(_44966), .Q(_45039) );
  nor2s1 _45403_inst ( .DIN1(_45041), .DIN2(_45042), .Q(_45038) );
  nor2s1 _45404_inst ( .DIN1(_44951), .DIN2(_45043), .Q(_45042) );
  nor2s1 _45405_inst ( .DIN1(_26851), .DIN2(_45045), .Q(_45041) );
  nor2s1 _45406_inst ( .DIN1(_45046), .DIN2(_45047), .Q(_45019) );
  nnd2s1 _45407_inst ( .DIN1(_45048), .DIN2(_45049), .Q(_45047) );
  hi1s1 _45408_inst ( .DIN(_45050), .Q(_45048) );
  nnd2s1 _45409_inst ( .DIN1(_45051), .DIN2(_45052), .Q(_45046) );
  nnd2s1 _45410_inst ( .DIN1(_44880), .DIN2(_44723), .Q(_45052) );
  nnd2s1 _45411_inst ( .DIN1(_45053), .DIN2(_26805), .Q(_45051) );
  nnd2s1 _45412_inst ( .DIN1(_45054), .DIN2(_45055), .Q(_45017) );
  nor2s1 _45413_inst ( .DIN1(_45056), .DIN2(_45057), .Q(_45055) );
  nnd2s1 _45414_inst ( .DIN1(_45058), .DIN2(_45059), .Q(_45057) );
  nor2s1 _45415_inst ( .DIN1(_26845), .DIN2(_45060), .Q(_45056) );
  nor2s1 _45416_inst ( .DIN1(_45061), .DIN2(_45062), .Q(_45054) );
  nnd2s1 _45417_inst ( .DIN1(_45063), .DIN2(_45064), .Q(_45062) );
  hi1s1 _45418_inst ( .DIN(_44731), .Q(_45063) );
  nnd2s1 _45419_inst ( .DIN1(_45065), .DIN2(_45066), .Q(_44731) );
  or2s1 _45420_inst ( .DIN1(_45067), .DIN2(_26805), .Q(_45066) );
  nnd2s1 _45421_inst ( .DIN1(_44884), .DIN2(_26805), .Q(_45065) );
  nnd2s1 _45422_inst ( .DIN1(_45068), .DIN2(_45069), .Q(_31768) );
  nor2s1 _45423_inst ( .DIN1(_44286), .DIN2(_42797), .Q(_45069) );
  nor2s1 _45424_inst ( .DIN1(_45070), .DIN2(_45071), .Q(_45068) );
  nnd2s1 _45425_inst ( .DIN1(_45072), .DIN2(_45073), .Q(
        ____0___________0_1_____) );
  nnd2s1 _45426_inst ( .DIN1(_45074), .DIN2(_27509), .Q(_45073) );
  nnd2s1 _45427_inst ( .DIN1(_27510), .DIN2(_45075), .Q(_45074) );
  xor2s1 _45428_inst ( .DIN1(_45076), .DIN2(_45077), .Q(_45075) );
  xor2s1 _45429_inst ( .DIN1(_53465), .DIN2(_53466), .Q(_45077) );
  and2s1 _45430_inst ( .DIN1(_26467), .DIN2(_53152), .Q(_45076) );
  nor2s1 _45431_inst ( .DIN1(_27039), .DIN2(_35873), .Q(_27510) );
  hi1s1 _45432_inst ( .DIN(_45078), .Q(_35873) );
  nnd2s1 _45433_inst ( .DIN1(_45079), .DIN2(_27512), .Q(_45072) );
  hi1s1 _45434_inst ( .DIN(_27509), .Q(_27512) );
  nnd2s1 _45435_inst ( .DIN1(_27606), .DIN2(_35994), .Q(_27509) );
  nor2s1 _45436_inst ( .DIN1(_45078), .DIN2(_35511), .Q(_27606) );
  nnd2s1 _45437_inst ( .DIN1(_35993), .DIN2(_45080), .Q(_45078) );
  nor2s1 _45438_inst ( .DIN1(_45081), .DIN2(_45082), .Q(_45079) );
  nnd2s1 _45439_inst ( .DIN1(_45083), .DIN2(_45084), .Q(_45082) );
  nor2s1 _45440_inst ( .DIN1(_45085), .DIN2(_45086), .Q(_45084) );
  nnd2s1 _45441_inst ( .DIN1(_45023), .DIN2(_45087), .Q(_45086) );
  nnd2s1 _45442_inst ( .DIN1(_44812), .DIN2(_44723), .Q(_45087) );
  nnd2s1 _45443_inst ( .DIN1(_44724), .DIN2(_45067), .Q(_44812) );
  xor2s1 _45444_inst ( .DIN1(_41043), .DIN2(_45088), .Q(_45023) );
  nor2s1 _45445_inst ( .DIN1(_45089), .DIN2(_45090), .Q(_45088) );
  nnd2s1 _45446_inst ( .DIN1(_45091), .DIN2(_45003), .Q(_45090) );
  nnd2s1 _45447_inst ( .DIN1(_45092), .DIN2(_44723), .Q(_45003) );
  nnd2s1 _45448_inst ( .DIN1(_44946), .DIN2(_44892), .Q(_45089) );
  nnd2s1 _45449_inst ( .DIN1(_45093), .DIN2(_26852), .Q(_44946) );
  hi1s1 _45450_inst ( .DIN(_44825), .Q(_45093) );
  nnd2s1 _45451_inst ( .DIN1(_45094), .DIN2(_45095), .Q(_41043) );
  nor2s1 _45452_inst ( .DIN1(_44288), .DIN2(_44313), .Q(_45094) );
  nnd2s1 _45453_inst ( .DIN1(_45096), .DIN2(_45097), .Q(_44288) );
  nor2s1 _45454_inst ( .DIN1(_45098), .DIN2(_44317), .Q(_45097) );
  nor2s1 _45455_inst ( .DIN1(_45099), .DIN2(_45070), .Q(_45096) );
  nnd2s1 _45456_inst ( .DIN1(_45100), .DIN2(_44985), .Q(_45070) );
  nnd2s1 _45457_inst ( .DIN1(_45101), .DIN2(_45102), .Q(_44985) );
  nor2s1 _45458_inst ( .DIN1(_45103), .DIN2(_45104), .Q(_45101) );
  nor2s1 _45459_inst ( .DIN1(_44977), .DIN2(_44980), .Q(_45100) );
  nnd2s1 _45460_inst ( .DIN1(_45105), .DIN2(_45106), .Q(_45085) );
  nor2s1 _45461_inst ( .DIN1(_44868), .DIN2(_45107), .Q(_45083) );
  nnd2s1 _45462_inst ( .DIN1(_44809), .DIN2(_45108), .Q(_45107) );
  and2s1 _45463_inst ( .DIN1(_45109), .DIN2(_45110), .Q(_44809) );
  nor2s1 _45464_inst ( .DIN1(_45111), .DIN2(_45112), .Q(_45110) );
  nnd2s1 _45465_inst ( .DIN1(_45113), .DIN2(_44897), .Q(_45112) );
  and2s1 _45466_inst ( .DIN1(_45114), .DIN2(_45115), .Q(_45113) );
  nnd2s1 _45467_inst ( .DIN1(_45116), .DIN2(_45117), .Q(_45111) );
  nor2s1 _45468_inst ( .DIN1(_44773), .DIN2(_45118), .Q(_45117) );
  and2s1 _45469_inst ( .DIN1(_45032), .DIN2(_44955), .Q(_45116) );
  nor2s1 _45470_inst ( .DIN1(_45119), .DIN2(_45120), .Q(_45109) );
  nnd2s1 _45471_inst ( .DIN1(_45121), .DIN2(_45122), .Q(_45120) );
  hi1s1 _45472_inst ( .DIN(_45030), .Q(_45122) );
  nnd2s1 _45473_inst ( .DIN1(_44883), .DIN2(_45123), .Q(_45030) );
  nor2s1 _45474_inst ( .DIN1(_44790), .DIN2(_44952), .Q(_45121) );
  nnd2s1 _45475_inst ( .DIN1(_45124), .DIN2(_45125), .Q(_44952) );
  nnd2s1 _45476_inst ( .DIN1(_44767), .DIN2(_26845), .Q(_45125) );
  nnd2s1 _45477_inst ( .DIN1(_45126), .DIN2(_45127), .Q(_44790) );
  nor2s1 _45478_inst ( .DIN1(_45128), .DIN2(_45129), .Q(_45127) );
  nnd2s1 _45479_inst ( .DIN1(_45130), .DIN2(_45131), .Q(_45129) );
  or2s1 _45480_inst ( .DIN1(_45132), .DIN2(_26804), .Q(_45130) );
  nor2s1 _45481_inst ( .DIN1(_44715), .DIN2(_45133), .Q(_45128) );
  nor2s1 _45482_inst ( .DIN1(_44842), .DIN2(_45134), .Q(_45126) );
  xor2s1 _45483_inst ( .DIN1(_41072), .DIN2(_45135), .Q(_45134) );
  nor2s1 _45484_inst ( .DIN1(_45136), .DIN2(_44949), .Q(_45135) );
  nnd2s1 _45485_inst ( .DIN1(_44714), .DIN2(_45137), .Q(_44842) );
  nnd2s1 _45486_inst ( .DIN1(_45138), .DIN2(_26799), .Q(_45137) );
  nnd2s1 _45487_inst ( .DIN1(_45139), .DIN2(_45140), .Q(_45119) );
  nor2s1 _45488_inst ( .DIN1(_45141), .DIN2(_45142), .Q(_45140) );
  nor2s1 _45489_inst ( .DIN1(_26805), .DIN2(_44912), .Q(_45141) );
  nor2s1 _45490_inst ( .DIN1(_45143), .DIN2(_45144), .Q(_45139) );
  nnd2s1 _45491_inst ( .DIN1(_45145), .DIN2(_45146), .Q(_44868) );
  nor2s1 _45492_inst ( .DIN1(_44965), .DIN2(_45147), .Q(_45146) );
  nnd2s1 _45493_inst ( .DIN1(_44805), .DIN2(_45031), .Q(_45147) );
  hi1s1 _45494_inst ( .DIN(_44753), .Q(_45031) );
  nor2s1 _45495_inst ( .DIN1(_45148), .DIN2(_44811), .Q(_45145) );
  nnd2s1 _45496_inst ( .DIN1(_45149), .DIN2(_45150), .Q(_44811) );
  nor2s1 _45497_inst ( .DIN1(_45151), .DIN2(_45152), .Q(_45150) );
  nnd2s1 _45498_inst ( .DIN1(_45153), .DIN2(_45060), .Q(_45152) );
  nnd2s1 _45499_inst ( .DIN1(_45154), .DIN2(_26845), .Q(_45153) );
  nnd2s1 _45500_inst ( .DIN1(_26770), .DIN2(_45043), .Q(_45154) );
  nnd2s1 _45501_inst ( .DIN1(_44913), .DIN2(_45155), .Q(_45151) );
  nor2s1 _45502_inst ( .DIN1(_45156), .DIN2(_45157), .Q(_44913) );
  hi1s1 _45503_inst ( .DIN(_44755), .Q(_45156) );
  nor2s1 _45504_inst ( .DIN1(_45158), .DIN2(_45159), .Q(_45149) );
  or2s1 _45505_inst ( .DIN1(_45037), .DIN2(_45010), .Q(_45159) );
  nnd2s1 _45506_inst ( .DIN1(_45160), .DIN2(_45161), .Q(_45010) );
  nor2s1 _45507_inst ( .DIN1(_45162), .DIN2(_45163), .Q(_45161) );
  nor2s1 _45508_inst ( .DIN1(_26851), .DIN2(_45164), .Q(_45163) );
  nor2s1 _45509_inst ( .DIN1(_26766), .DIN2(_45165), .Q(_45162) );
  nor2s1 _45510_inst ( .DIN1(_45166), .DIN2(_45167), .Q(_45160) );
  nor2s1 _45511_inst ( .DIN1(_45168), .DIN2(_45169), .Q(_45167) );
  or2s1 _45512_inst ( .DIN1(_44736), .DIN2(_45170), .Q(_45158) );
  nnd2s1 _45513_inst ( .DIN1(_45171), .DIN2(_45172), .Q(_44736) );
  nor2s1 _45514_inst ( .DIN1(_45173), .DIN2(_45174), .Q(_45172) );
  nor2s1 _45515_inst ( .DIN1(_45175), .DIN2(_45176), .Q(_45171) );
  nor2s1 _45516_inst ( .DIN1(_44715), .DIN2(_44828), .Q(_45148) );
  nnd2s1 _45517_inst ( .DIN1(_45177), .DIN2(_45178), .Q(_45081) );
  nor2s1 _45518_inst ( .DIN1(_45179), .DIN2(_45180), .Q(_45178) );
  nnd2s1 _45519_inst ( .DIN1(_44964), .DIN2(_44899), .Q(_45180) );
  nnd2s1 _45520_inst ( .DIN1(_45181), .DIN2(_45182), .Q(_45179) );
  nor2s1 _45521_inst ( .DIN1(_45183), .DIN2(_45184), .Q(_45177) );
  nnd2s1 _45522_inst ( .DIN1(_45185), .DIN2(_45186), .Q(_45184) );
  nnd2s1 _45523_inst ( .DIN1(_45187), .DIN2(_45188), .Q(
        ____0___________0_13_____) );
  nnd2s1 _45524_inst ( .DIN1(_45189), .DIN2(_27520), .Q(_45188) );
  nnd2s1 _45525_inst ( .DIN1(_45190), .DIN2(_45191), .Q(_45189) );
  xnr2s1 _45526_inst ( .DIN1(_52896), .DIN2(_29710), .Q(_45191) );
  nor2s1 _45527_inst ( .DIN1(_53467), .DIN2(_53471), .Q(_29710) );
  nor2s1 _45528_inst ( .DIN1(_27522), .DIN2(_27614), .Q(_45190) );
  and2s1 _45529_inst ( .DIN1(_45192), .DIN2(_45193), .Q(_27522) );
  nor2s1 _45530_inst ( .DIN1(_45194), .DIN2(_45195), .Q(_45193) );
  or2s1 _45531_inst ( .DIN1(_45196), .DIN2(_27742), .Q(_45195) );
  nor2s1 _45532_inst ( .DIN1(_45197), .DIN2(_45198), .Q(_45192) );
  nnd2s1 _45533_inst ( .DIN1(_45199), .DIN2(_27524), .Q(_45187) );
  hi1s1 _45534_inst ( .DIN(_27520), .Q(_27524) );
  nnd2s1 _45535_inst ( .DIN1(_45200), .DIN2(_45201), .Q(_27520) );
  nor2s1 _45536_inst ( .DIN1(_27744), .DIN2(_45202), .Q(_45201) );
  nnd2s1 _45537_inst ( .DIN1(_45203), .DIN2(_45204), .Q(_45202) );
  nnd2s1 _45538_inst ( .DIN1(_45205), .DIN2(_45206), .Q(_27744) );
  nnd2s1 _45539_inst ( .DIN1(_45207), .DIN2(_45208), .Q(_45206) );
  nor2s1 _45540_inst ( .DIN1(_39518), .DIN2(_45209), .Q(_45200) );
  nnd2s1 _45541_inst ( .DIN1(_45210), .DIN2(_45211), .Q(_39518) );
  nor2s1 _45542_inst ( .DIN1(_45212), .DIN2(_45197), .Q(_45210) );
  nor2s1 _45543_inst ( .DIN1(_45213), .DIN2(_45214), .Q(_45199) );
  nnd2s1 _45544_inst ( .DIN1(_45215), .DIN2(_45216), .Q(_45214) );
  nor2s1 _45545_inst ( .DIN1(_45217), .DIN2(_45218), .Q(_45216) );
  nnd2s1 _45546_inst ( .DIN1(_44837), .DIN2(_45091), .Q(_45218) );
  and2s1 _45547_inst ( .DIN1(_45219), .DIN2(_45220), .Q(_45091) );
  nnd2s1 _45548_inst ( .DIN1(_26765), .DIN2(_26851), .Q(_45219) );
  and2s1 _45549_inst ( .DIN1(_45123), .DIN2(_45221), .Q(_44837) );
  nnd2s1 _45550_inst ( .DIN1(_45136), .DIN2(_26805), .Q(_45221) );
  hi1s1 _45551_inst ( .DIN(_45222), .Q(_45136) );
  nnd2s1 _45552_inst ( .DIN1(_45223), .DIN2(_45224), .Q(_45123) );
  nnd2s1 _45553_inst ( .DIN1(_45225), .DIN2(_45226), .Q(_45217) );
  nor2s1 _45554_inst ( .DIN1(_45227), .DIN2(_45228), .Q(_45225) );
  nor2s1 _45555_inst ( .DIN1(_26805), .DIN2(_45229), .Q(_45227) );
  nor2s1 _45556_inst ( .DIN1(_45230), .DIN2(_45231), .Q(_45215) );
  nnd2s1 _45557_inst ( .DIN1(_45232), .DIN2(_45233), .Q(_45231) );
  nnd2s1 _45558_inst ( .DIN1(_45234), .DIN2(_44867), .Q(_45230) );
  and2s1 _45559_inst ( .DIN1(_45235), .DIN2(_45236), .Q(_44867) );
  nnd2s1 _45560_inst ( .DIN1(_45237), .DIN2(_26851), .Q(_45236) );
  nnd2s1 _45561_inst ( .DIN1(_26805), .DIN2(_45238), .Q(_45235) );
  hi1s1 _45562_inst ( .DIN(_44971), .Q(_45234) );
  nnd2s1 _45563_inst ( .DIN1(_45239), .DIN2(_45240), .Q(_44971) );
  nor2s1 _45564_inst ( .DIN1(_45241), .DIN2(_45242), .Q(_45240) );
  nnd2s1 _45565_inst ( .DIN1(_45243), .DIN2(_45244), .Q(_45242) );
  nor2s1 _45566_inst ( .DIN1(_44791), .DIN2(_44810), .Q(_45243) );
  nnd2s1 _45567_inst ( .DIN1(_45245), .DIN2(_45246), .Q(_44810) );
  nnd2s1 _45568_inst ( .DIN1(_45183), .DIN2(_26845), .Q(_45246) );
  nnd2s1 _45569_inst ( .DIN1(_45247), .DIN2(_45248), .Q(_44791) );
  nor2s1 _45570_inst ( .DIN1(_45249), .DIN2(_45250), .Q(_45248) );
  nnd2s1 _45571_inst ( .DIN1(_45251), .DIN2(_45252), .Q(_45250) );
  nnd2s1 _45572_inst ( .DIN1(_44851), .DIN2(_26766), .Q(_45252) );
  nnd2s1 _45573_inst ( .DIN1(_45253), .DIN2(_26805), .Q(_45251) );
  nnd2s1 _45574_inst ( .DIN1(_45254), .DIN2(_45060), .Q(_45249) );
  hi1s1 _45575_inst ( .DIN(_45255), .Q(_45060) );
  nor2s1 _45576_inst ( .DIN1(_45256), .DIN2(_45174), .Q(_45254) );
  and2s1 _45577_inst ( .DIN1(_45257), .DIN2(_26766), .Q(_45174) );
  nor2s1 _45578_inst ( .DIN1(_45258), .DIN2(_45259), .Q(_45247) );
  nnd2s1 _45579_inst ( .DIN1(_45260), .DIN2(_45261), .Q(_45259) );
  hi1s1 _45580_inst ( .DIN(_45144), .Q(_45260) );
  nnd2s1 _45581_inst ( .DIN1(_45262), .DIN2(_45263), .Q(_45144) );
  nor2s1 _45582_inst ( .DIN1(_45264), .DIN2(_45265), .Q(_45263) );
  nnd2s1 _45583_inst ( .DIN1(_45266), .DIN2(_45267), .Q(_45265) );
  nor2s1 _45584_inst ( .DIN1(_45268), .DIN2(_45061), .Q(_45262) );
  nnd2s1 _45585_inst ( .DIN1(_45269), .DIN2(_45270), .Q(_45061) );
  nnd2s1 _45586_inst ( .DIN1(_45271), .DIN2(_45272), .Q(_45270) );
  nor2s1 _45587_inst ( .DIN1(_45168), .DIN2(_26845), .Q(_45271) );
  or2s1 _45588_inst ( .DIN1(_45273), .DIN2(_26799), .Q(_45269) );
  nnd2s1 _45589_inst ( .DIN1(_45274), .DIN2(_45108), .Q(_45258) );
  and2s1 _45590_inst ( .DIN1(_45275), .DIN2(_45276), .Q(_45108) );
  nnd2s1 _45591_inst ( .DIN1(_45277), .DIN2(_44771), .Q(_45276) );
  nor2s1 _45592_inst ( .DIN1(_45278), .DIN2(_44803), .Q(_45274) );
  nor2s1 _45593_inst ( .DIN1(_44951), .DIN2(_45279), .Q(_45278) );
  nnd2s1 _45594_inst ( .DIN1(_45280), .DIN2(_45281), .Q(_45241) );
  hi1s1 _45595_inst ( .DIN(_45282), .Q(_45281) );
  nor2s1 _45596_inst ( .DIN1(_44773), .DIN2(_45283), .Q(_45280) );
  nor2s1 _45597_inst ( .DIN1(_45284), .DIN2(_45285), .Q(_45239) );
  nnd2s1 _45598_inst ( .DIN1(_45286), .DIN2(_45287), .Q(_45285) );
  nor2s1 _45599_inst ( .DIN1(_45288), .DIN2(_45289), .Q(_45287) );
  nor2s1 _45600_inst ( .DIN1(_44771), .DIN2(_45290), .Q(_45289) );
  nor2s1 _45601_inst ( .DIN1(_44715), .DIN2(_45291), .Q(_45288) );
  nor2s1 _45602_inst ( .DIN1(_45292), .DIN2(_45293), .Q(_45286) );
  nor2s1 _45603_inst ( .DIN1(_26852), .DIN2(_45294), .Q(_45293) );
  nor2s1 _45604_inst ( .DIN1(_26767), .DIN2(_45295), .Q(_45292) );
  nnd2s1 _45605_inst ( .DIN1(_45296), .DIN2(_45297), .Q(_45284) );
  nor2s1 _45606_inst ( .DIN1(_45298), .DIN2(_45299), .Q(_45297) );
  nor2s1 _45607_inst ( .DIN1(_26845), .DIN2(_45300), .Q(_45299) );
  nor2s1 _45608_inst ( .DIN1(_44951), .DIN2(_45301), .Q(_45298) );
  nor2s1 _45609_inst ( .DIN1(_44858), .DIN2(_45302), .Q(_45296) );
  nnd2s1 _45610_inst ( .DIN1(_45303), .DIN2(_45304), .Q(_44858) );
  nnd2s1 _45611_inst ( .DIN1(_45305), .DIN2(_26845), .Q(_45304) );
  nnd2s1 _45612_inst ( .DIN1(_44761), .DIN2(_45114), .Q(_45305) );
  nnd2s1 _45613_inst ( .DIN1(_45053), .DIN2(_44723), .Q(_45303) );
  hi1s1 _45614_inst ( .DIN(_44897), .Q(_45053) );
  nnd2s1 _45615_inst ( .DIN1(_45306), .DIN2(_45307), .Q(_45213) );
  nor2s1 _45616_inst ( .DIN1(_45308), .DIN2(_45309), .Q(_45307) );
  nnd2s1 _45617_inst ( .DIN1(_45310), .DIN2(_45311), .Q(_45309) );
  nnd2s1 _45618_inst ( .DIN1(_45312), .DIN2(_45313), .Q(_45308) );
  and2s1 _45619_inst ( .DIN1(_44755), .DIN2(_44818), .Q(_45312) );
  nnd2s1 _45620_inst ( .DIN1(_26767), .DIN2(_45314), .Q(_44755) );
  nor2s1 _45621_inst ( .DIN1(_45315), .DIN2(_45316), .Q(_45306) );
  nnd2s1 _45622_inst ( .DIN1(_45317), .DIN2(_45318), .Q(_45316) );
  nnd2s1 _45623_inst ( .DIN1(_45319), .DIN2(_45064), .Q(_45315) );
  nnd2s1 _45624_inst ( .DIN1(_45320), .DIN2(_26767), .Q(_45064) );
  nnd2s1 _45625_inst ( .DIN1(_44951), .DIN2(_45321), .Q(_45319) );
  nnd2s1 _45626_inst ( .DIN1(_45322), .DIN2(_45323), .Q(
        ____0___________0_12_____) );
  nnd2s1 _45627_inst ( .DIN1(_39842), .DIN2(_45324), .Q(_45323) );
  nnd2s1 _45628_inst ( .DIN1(_45325), .DIN2(_45326), .Q(_45324) );
  nor2s1 _45629_inst ( .DIN1(_45327), .DIN2(_45328), .Q(_45326) );
  nnd2s1 _45630_inst ( .DIN1(_45329), .DIN2(_45330), .Q(_45328) );
  nor2s1 _45631_inst ( .DIN1(_44778), .DIN2(_44877), .Q(_45329) );
  nnd2s1 _45632_inst ( .DIN1(_45331), .DIN2(_45332), .Q(_44877) );
  nor2s1 _45633_inst ( .DIN1(_45333), .DIN2(_45334), .Q(_45332) );
  nnd2s1 _45634_inst ( .DIN1(_45133), .DIN2(_44964), .Q(_45334) );
  hi1s1 _45635_inst ( .DIN(_45335), .Q(_44964) );
  hi1s1 _45636_inst ( .DIN(_45058), .Q(_45333) );
  nor2s1 _45637_inst ( .DIN1(_45336), .DIN2(_45337), .Q(_45331) );
  nnd2s1 _45638_inst ( .DIN1(_45338), .DIN2(_45339), .Q(_45337) );
  nnd2s1 _45639_inst ( .DIN1(_44848), .DIN2(_44723), .Q(_45339) );
  hi1s1 _45640_inst ( .DIN(_45124), .Q(_44848) );
  nnd2s1 _45641_inst ( .DIN1(_44715), .DIN2(_44923), .Q(_45338) );
  nnd2s1 _45642_inst ( .DIN1(_45340), .DIN2(_45341), .Q(_44778) );
  nor2s1 _45643_inst ( .DIN1(_45342), .DIN2(_45343), .Q(_45341) );
  nnd2s1 _45644_inst ( .DIN1(_45344), .DIN2(_44912), .Q(_45343) );
  nnd2s1 _45645_inst ( .DIN1(_45345), .DIN2(_45346), .Q(_45342) );
  nnd2s1 _45646_inst ( .DIN1(_45157), .DIN2(_26852), .Q(_45346) );
  nor2s1 _45647_inst ( .DIN1(_45347), .DIN2(_45348), .Q(_45345) );
  nor2s1 _45648_inst ( .DIN1(_44951), .DIN2(_44914), .Q(_45348) );
  nor2s1 _45649_inst ( .DIN1(_44771), .DIN2(_44856), .Q(_45347) );
  nor2s1 _45650_inst ( .DIN1(_45349), .DIN2(_45350), .Q(_45340) );
  nnd2s1 _45651_inst ( .DIN1(_45351), .DIN2(_44844), .Q(_45350) );
  and2s1 _45652_inst ( .DIN1(_45032), .DIN2(_45352), .Q(_44844) );
  or2s1 _45653_inst ( .DIN1(_44724), .DIN2(_26805), .Q(_45352) );
  nnd2s1 _45654_inst ( .DIN1(_45353), .DIN2(_44771), .Q(_45032) );
  nor2s1 _45655_inst ( .DIN1(_45354), .DIN2(_45355), .Q(_45351) );
  nor2s1 _45656_inst ( .DIN1(_26805), .DIN2(_45067), .Q(_45354) );
  nnd2s1 _45657_inst ( .DIN1(_44800), .DIN2(_45028), .Q(_45349) );
  and2s1 _45658_inst ( .DIN1(_45356), .DIN2(_45311), .Q(_45028) );
  nor2s1 _45659_inst ( .DIN1(_45173), .DIN2(_44961), .Q(_45356) );
  nor2s1 _45660_inst ( .DIN1(_45357), .DIN2(_44723), .Q(_45173) );
  and2s1 _45661_inst ( .DIN1(_45358), .DIN2(_45359), .Q(_44800) );
  nnd2s1 _45662_inst ( .DIN1(_44965), .DIN2(_44723), .Q(_45359) );
  nor2s1 _45663_inst ( .DIN1(_45360), .DIN2(_45361), .Q(_45358) );
  nor2s1 _45664_inst ( .DIN1(_44771), .DIN2(_44899), .Q(_45361) );
  nor2s1 _45665_inst ( .DIN1(_26766), .DIN2(_45105), .Q(_45360) );
  nnd2s1 _45666_inst ( .DIN1(_45362), .DIN2(_45363), .Q(_45327) );
  nor2s1 _45667_inst ( .DIN1(_45364), .DIN2(_44901), .Q(_45363) );
  nor2s1 _45668_inst ( .DIN1(_45365), .DIN2(_44706), .Q(_45362) );
  nnd2s1 _45669_inst ( .DIN1(_45366), .DIN2(_45367), .Q(_44706) );
  nor2s1 _45670_inst ( .DIN1(_45228), .DIN2(_45368), .Q(_45367) );
  nnd2s1 _45671_inst ( .DIN1(_45369), .DIN2(_44883), .Q(_45368) );
  nnd2s1 _45672_inst ( .DIN1(_45370), .DIN2(_26766), .Q(_45369) );
  nor2s1 _45673_inst ( .DIN1(_44723), .DIN2(_44826), .Q(_45228) );
  nor2s1 _45674_inst ( .DIN1(_45371), .DIN2(_44921), .Q(_45366) );
  nnd2s1 _45675_inst ( .DIN1(_45372), .DIN2(_45373), .Q(_44921) );
  nnd2s1 _45676_inst ( .DIN1(_45374), .DIN2(_26851), .Q(_45373) );
  xor2s1 _45677_inst ( .DIN1(_45375), .DIN2(_36445), .Q(_45372) );
  hi1s1 _45678_inst ( .DIN(_34026), .Q(_36445) );
  nnd2s1 _45679_inst ( .DIN1(_37792), .DIN2(_44658), .Q(_34026) );
  nnd2s1 _45680_inst ( .DIN1(_45290), .DIN2(_45376), .Q(_45375) );
  nnd2s1 _45681_inst ( .DIN1(_43565), .DIN2(_44951), .Q(_45376) );
  hi1s1 _45682_inst ( .DIN(_26770), .Q(_43565) );
  nor2s1 _45683_inst ( .DIN1(_26805), .DIN2(_45377), .Q(_45365) );
  nor2s1 _45684_inst ( .DIN1(_44966), .DIN2(_45378), .Q(_45377) );
  nnd2s1 _45685_inst ( .DIN1(_45379), .DIN2(_45222), .Q(_45378) );
  nor2s1 _45686_inst ( .DIN1(_45380), .DIN2(_45381), .Q(_45325) );
  nnd2s1 _45687_inst ( .DIN1(_45382), .DIN2(_45383), .Q(_45381) );
  nor2s1 _45688_inst ( .DIN1(_45384), .DIN2(_45385), .Q(_45383) );
  and2s1 _45689_inst ( .DIN1(_26845), .DIN2(_45386), .Q(_45385) );
  nor2s1 _45690_inst ( .DIN1(_26845), .DIN2(_45387), .Q(_45384) );
  nor2s1 _45691_inst ( .DIN1(_45388), .DIN2(_45389), .Q(_45382) );
  nnd2s1 _45692_inst ( .DIN1(_45390), .DIN2(_45391), .Q(_45389) );
  nnd2s1 _45693_inst ( .DIN1(_45392), .DIN2(_26852), .Q(_45390) );
  nnd2s1 _45694_inst ( .DIN1(_45393), .DIN2(_45045), .Q(_45392) );
  nnd2s1 _45695_inst ( .DIN1(_45394), .DIN2(_45395), .Q(_45388) );
  nnd2s1 _45696_inst ( .DIN1(_45396), .DIN2(_44771), .Q(_45395) );
  nnd2s1 _45697_inst ( .DIN1(_45397), .DIN2(_44715), .Q(_45394) );
  nnd2s1 _45698_inst ( .DIN1(_45398), .DIN2(_45399), .Q(_45380) );
  nor2s1 _45699_inst ( .DIN1(_44917), .DIN2(_45006), .Q(_45398) );
  nnd2s1 _45700_inst ( .DIN1(_45400), .DIN2(_45401), .Q(_45006) );
  nnd2s1 _45701_inst ( .DIN1(_30081), .DIN2(_44714), .Q(_45401) );
  nor2s1 _45702_inst ( .DIN1(_45402), .DIN2(_45403), .Q(_45400) );
  nor2s1 _45703_inst ( .DIN1(_26767), .DIN2(_45404), .Q(_45403) );
  nor2s1 _45704_inst ( .DIN1(_44871), .DIN2(_30081), .Q(_45404) );
  nor2s1 _45705_inst ( .DIN1(_26851), .DIN2(_45405), .Q(_45402) );
  nnd2s1 _45706_inst ( .DIN1(_45237), .DIN2(_44070), .Q(_45405) );
  hi1s1 _45707_inst ( .DIN(_30081), .Q(_44070) );
  nnd2s1 _45708_inst ( .DIN1(_45406), .DIN2(_27924), .Q(_30081) );
  hi1s1 _45709_inst ( .DIN(_32716), .Q(_27924) );
  nnd2s1 _45710_inst ( .DIN1(_43029), .DIN2(_33865), .Q(_32716) );
  and2s1 _45711_inst ( .DIN1(_45407), .DIN2(_44600), .Q(_45406) );
  hi1s1 _45712_inst ( .DIN(_44714), .Q(_45237) );
  nnd2s1 _45713_inst ( .DIN1(_45408), .DIN2(_45409), .Q(_44917) );
  nor2s1 _45714_inst ( .DIN1(_45410), .DIN2(_45411), .Q(_45409) );
  nnd2s1 _45715_inst ( .DIN1(_45295), .DIN2(_45059), .Q(_45411) );
  nor2s1 _45716_inst ( .DIN1(_45412), .DIN2(_45413), .Q(_45408) );
  nor2s1 _45717_inst ( .DIN1(_26766), .DIN2(_45414), .Q(_45413) );
  nor2s1 _45718_inst ( .DIN1(_26845), .DIN2(_44890), .Q(_45412) );
  nnd2s1 _45719_inst ( .DIN1(_53477), .DIN2(_44692), .Q(_45322) );
  hi1s1 _45720_inst ( .DIN(_39841), .Q(_44692) );
  nnd2s1 _45721_inst ( .DIN1(_45415), .DIN2(_39947), .Q(_39841) );
  hi1s1 _45722_inst ( .DIN(_39842), .Q(_39947) );
  nor2s1 _45723_inst ( .DIN1(_42748), .DIN2(_27431), .Q(_39842) );
  nnd2s1 _45724_inst ( .DIN1(_45416), .DIN2(_32826), .Q(_27431) );
  nor2s1 _45725_inst ( .DIN1(_45417), .DIN2(_31396), .Q(_45416) );
  hi1s1 _45726_inst ( .DIN(_44324), .Q(_31396) );
  nnd2s1 _45727_inst ( .DIN1(_45418), .DIN2(_45419), .Q(_42748) );
  nor2s1 _45728_inst ( .DIN1(_32807), .DIN2(_45420), .Q(_45419) );
  nnd2s1 _45729_inst ( .DIN1(_27442), .DIN2(_29741), .Q(_45420) );
  nor2s1 _45730_inst ( .DIN1(_45421), .DIN2(_44323), .Q(_45418) );
  nnd2s1 _45731_inst ( .DIN1(_45422), .DIN2(_45423), .Q(_44323) );
  nor2s1 _45732_inst ( .DIN1(_29767), .DIN2(_45424), .Q(_45422) );
  nnd2s1 _45733_inst ( .DIN1(_42130), .DIN2(_32826), .Q(_45415) );
  hi1s1 _45734_inst ( .DIN(_27443), .Q(_42130) );
  nnd2s1 _45735_inst ( .DIN1(_45425), .DIN2(_45426), .Q(_27443) );
  nor2s1 _45736_inst ( .DIN1(_42753), .DIN2(_32813), .Q(_45426) );
  hi1s1 _45737_inst ( .DIN(_29741), .Q(_42753) );
  nor2s1 _45738_inst ( .DIN1(_45421), .DIN2(_44687), .Q(_45425) );
  nnd2s1 _45739_inst ( .DIN1(_45427), .DIN2(_45428), .Q(_44687) );
  nor2s1 _45740_inst ( .DIN1(_27308), .DIN2(_29767), .Q(_45428) );
  nor2s1 _45741_inst ( .DIN1(_27311), .DIN2(_27432), .Q(_45427) );
  nnd2s1 _45742_inst ( .DIN1(_45423), .DIN2(_43497), .Q(_27432) );
  and2s1 _45743_inst ( .DIN1(_32825), .DIN2(_45429), .Q(_45423) );
  nnd2s1 _45744_inst ( .DIN1(_45430), .DIN2(_45431), .Q(_45429) );
  or2s1 _45745_inst ( .DIN1(_32815), .DIN2(_27430), .Q(_27311) );
  nnd2s1 _45746_inst ( .DIN1(_45432), .DIN2(_45433), .Q(_32815) );
  nor2s1 _45747_inst ( .DIN1(_45417), .DIN2(_32807), .Q(_45433) );
  hi1s1 _45748_inst ( .DIN(_45434), .Q(_32807) );
  hi1s1 _45749_inst ( .DIN(_45435), .Q(_45417) );
  nor2s1 _45750_inst ( .DIN1(_45424), .DIN2(_32810), .Q(_45432) );
  hi1s1 _45751_inst ( .DIN(_45436), .Q(_32810) );
  nnd2s1 _45752_inst ( .DIN1(_27994), .DIN2(_45437), .Q(
        ____0___________0_11_____) );
  nnd2s1 _45753_inst ( .DIN1(_45438), .DIN2(_45439), .Q(_45437) );
  nor2s1 _45754_inst ( .DIN1(_45440), .DIN2(_45441), .Q(_45439) );
  nnd2s1 _45755_inst ( .DIN1(_45442), .DIN2(_45049), .Q(_45441) );
  and2s1 _45756_inst ( .DIN1(_44945), .DIN2(_45443), .Q(_45049) );
  nnd2s1 _45757_inst ( .DIN1(_44711), .DIN2(_44951), .Q(_45443) );
  hi1s1 _45758_inst ( .DIN(_45114), .Q(_44711) );
  nnd2s1 _45759_inst ( .DIN1(_45444), .DIN2(_45445), .Q(_45114) );
  nnd2s1 _45760_inst ( .DIN1(_45374), .DIN2(_26767), .Q(_44945) );
  hi1s1 _45761_inst ( .DIN(_45155), .Q(_45374) );
  nor2s1 _45762_inst ( .DIN1(_44707), .DIN2(_44779), .Q(_45442) );
  nnd2s1 _45763_inst ( .DIN1(_45446), .DIN2(_45447), .Q(_44779) );
  and2s1 _45764_inst ( .DIN1(_45106), .DIN2(_26770), .Q(_45447) );
  nor2s1 _45765_inst ( .DIN1(_44871), .DIN2(_45448), .Q(_45446) );
  nnd2s1 _45766_inst ( .DIN1(_45449), .DIN2(_45450), .Q(_45448) );
  nnd2s1 _45767_inst ( .DIN1(_44885), .DIN2(_44723), .Q(_45450) );
  or2s1 _45768_inst ( .DIN1(_45451), .DIN2(_26804), .Q(_45449) );
  nnd2s1 _45769_inst ( .DIN1(_45452), .DIN2(_45453), .Q(_44707) );
  nor2s1 _45770_inst ( .DIN1(_45454), .DIN2(_45455), .Q(_45453) );
  nor2s1 _45771_inst ( .DIN1(_26852), .DIN2(_45295), .Q(_45455) );
  hi1s1 _45772_inst ( .DIN(_45267), .Q(_45454) );
  nnd2s1 _45773_inst ( .DIN1(_45456), .DIN2(_45457), .Q(_45267) );
  nor2s1 _45774_inst ( .DIN1(_45458), .DIN2(_45459), .Q(_45457) );
  nor2s1 _45775_inst ( .DIN1(_45460), .DIN2(_45461), .Q(_45456) );
  nor2s1 _45776_inst ( .DIN1(_45462), .DIN2(_45463), .Q(_45452) );
  nnd2s1 _45777_inst ( .DIN1(_45464), .DIN2(_45465), .Q(_45463) );
  nnd2s1 _45778_inst ( .DIN1(_44961), .DIN2(_44951), .Q(_45465) );
  nnd2s1 _45779_inst ( .DIN1(_45466), .DIN2(_26845), .Q(_45464) );
  nnd2s1 _45780_inst ( .DIN1(_45467), .DIN2(_44891), .Q(_45466) );
  nor2s1 _45781_inst ( .DIN1(_26805), .DIN2(_45266), .Q(_45462) );
  nnd2s1 _45782_inst ( .DIN1(_45468), .DIN2(_45469), .Q(_45440) );
  nnd2s1 _45783_inst ( .DIN1(_45138), .DIN2(_44715), .Q(_45469) );
  hi1s1 _45784_inst ( .DIN(_45290), .Q(_45138) );
  nor2s1 _45785_inst ( .DIN1(_45470), .DIN2(_45471), .Q(_45468) );
  xor2s1 _45786_inst ( .DIN1(_31307), .DIN2(_45472), .Q(_45471) );
  nor2s1 _45787_inst ( .DIN1(_44723), .DIN2(_45067), .Q(_45472) );
  nor2s1 _45788_inst ( .DIN1(_45473), .DIN2(_45474), .Q(_45438) );
  nnd2s1 _45789_inst ( .DIN1(_45475), .DIN2(_45476), .Q(_45474) );
  nor2s1 _45790_inst ( .DIN1(_45477), .DIN2(_45478), .Q(_45476) );
  nor2s1 _45791_inst ( .DIN1(_44951), .DIN2(_45479), .Q(_45478) );
  nor2s1 _45792_inst ( .DIN1(_45183), .DIN2(_44949), .Q(_45479) );
  nor2s1 _45793_inst ( .DIN1(_26845), .DIN2(_44818), .Q(_45477) );
  nor2s1 _45794_inst ( .DIN1(_45480), .DIN2(_45481), .Q(_45475) );
  nnd2s1 _45795_inst ( .DIN1(_45482), .DIN2(_45483), .Q(_45481) );
  nnd2s1 _45796_inst ( .DIN1(_45410), .DIN2(_26852), .Q(_45483) );
  hi1s1 _45797_inst ( .DIN(_45294), .Q(_45410) );
  nnd2s1 _45798_inst ( .DIN1(_45318), .DIN2(_45220), .Q(_45480) );
  nnd2s1 _45799_inst ( .DIN1(_44923), .DIN2(_44771), .Q(_45220) );
  nnd2s1 _45800_inst ( .DIN1(_45353), .DIN2(_44715), .Q(_45318) );
  hi1s1 _45801_inst ( .DIN(_45484), .Q(_45353) );
  nnd2s1 _45802_inst ( .DIN1(_45485), .DIN2(_45486), .Q(_45473) );
  xnr2s1 _45803_inst ( .DIN1(_45487), .DIN2(_37577), .Q(_45486) );
  nnd2s1 _45804_inst ( .DIN1(_45036), .DIN2(_45488), .Q(_45487) );
  hi1s1 _45805_inst ( .DIN(_44838), .Q(_45488) );
  nnd2s1 _45806_inst ( .DIN1(_45391), .DIN2(_45489), .Q(_44838) );
  nnd2s1 _45807_inst ( .DIN1(_45283), .DIN2(_44951), .Q(_45489) );
  nnd2s1 _45808_inst ( .DIN1(_45490), .DIN2(_26766), .Q(_45391) );
  and2s1 _45809_inst ( .DIN1(_45491), .DIN2(_45492), .Q(_45036) );
  nor2s1 _45810_inst ( .DIN1(_45493), .DIN2(_45494), .Q(_45492) );
  nnd2s1 _45811_inst ( .DIN1(_45495), .DIN2(_45393), .Q(_45494) );
  nor2s1 _45812_inst ( .DIN1(_45496), .DIN2(_44768), .Q(_45495) );
  nnd2s1 _45813_inst ( .DIN1(_45497), .DIN2(_45379), .Q(_45493) );
  nor2s1 _45814_inst ( .DIN1(_45321), .DIN2(_45498), .Q(_45497) );
  nor2s1 _45815_inst ( .DIN1(_45499), .DIN2(_45500), .Q(_45491) );
  nnd2s1 _45816_inst ( .DIN1(_45501), .DIN2(_45330), .Q(_45500) );
  and2s1 _45817_inst ( .DIN1(_45502), .DIN2(_45503), .Q(_45330) );
  nor2s1 _45818_inst ( .DIN1(_45504), .DIN2(_45505), .Q(_45503) );
  nnd2s1 _45819_inst ( .DIN1(_45300), .DIN2(_45506), .Q(_45505) );
  nnd2s1 _45820_inst ( .DIN1(_44857), .DIN2(_45301), .Q(_45504) );
  nor2s1 _45821_inst ( .DIN1(_45507), .DIN2(_45508), .Q(_45502) );
  nnd2s1 _45822_inst ( .DIN1(_44963), .DIN2(_45509), .Q(_45508) );
  nor2s1 _45823_inst ( .DIN1(_44704), .DIN2(_45386), .Q(_45501) );
  nnd2s1 _45824_inst ( .DIN1(_44761), .DIN2(_45510), .Q(_45386) );
  nnd2s1 _45825_inst ( .DIN1(_45511), .DIN2(_45512), .Q(_44704) );
  nor2s1 _45826_inst ( .DIN1(_45513), .DIN2(_45396), .Q(_45512) );
  hi1s1 _45827_inst ( .DIN(_45514), .Q(_45396) );
  nor2s1 _45828_inst ( .DIN1(_45397), .DIN2(_45142), .Q(_45511) );
  nnd2s1 _45829_inst ( .DIN1(_45515), .DIN2(_45516), .Q(_45499) );
  nor2s1 _45830_inst ( .DIN1(_44757), .DIN2(_45517), .Q(_45515) );
  nor2s1 _45831_inst ( .DIN1(_26845), .DIN2(_45279), .Q(_45517) );
  nor2s1 _45832_inst ( .DIN1(_44805), .DIN2(_44771), .Q(_44757) );
  nor2s1 _45833_inst ( .DIN1(_45518), .DIN2(_45519), .Q(_45485) );
  xor2s1 _45834_inst ( .DIN1(_29599), .DIN2(_45520), .Q(_45519) );
  nnd2s1 _45835_inst ( .DIN1(_45521), .DIN2(_45522), .Q(_45520) );
  nor2s1 _45836_inst ( .DIN1(_45364), .DIN2(_45092), .Q(_45522) );
  hi1s1 _45837_inst ( .DIN(_44826), .Q(_45092) );
  nor2s1 _45838_inst ( .DIN1(_45320), .DIN2(_45523), .Q(_45521) );
  nor2s1 _45839_inst ( .DIN1(_44771), .DIN2(_44817), .Q(_45523) );
  hi1s1 _45840_inst ( .DIN(_27500), .Q(_27994) );
  nnd2s1 _45841_inst ( .DIN1(_37006), .DIN2(_29221), .Q(_27500) );
  nnd2s1 _45842_inst ( .DIN1(_45524), .DIN2(_45525), .Q(
        ____0___________0_10_____) );
  nnd2s1 _45843_inst ( .DIN1(_45526), .DIN2(_35902), .Q(_45525) );
  nnd2s1 _45844_inst ( .DIN1(_45527), .DIN2(______[30]), .Q(_45526) );
  nor2s1 _45845_inst ( .DIN1(_30866), .DIN2(_45528), .Q(_45527) );
  xor2s1 _45846_inst ( .DIN1(_26592), .DIN2(_53468), .Q(_45528) );
  hi1s1 _45847_inst ( .DIN(_29082), .Q(_30866) );
  nnd2s1 _45848_inst ( .DIN1(_45529), .DIN2(_45530), .Q(_29082) );
  nor2s1 _45849_inst ( .DIN1(_45194), .DIN2(_45531), .Q(_45530) );
  nnd2s1 _45850_inst ( .DIN1(_45532), .DIN2(_45533), .Q(_45531) );
  nor2s1 _45851_inst ( .DIN1(_45197), .DIN2(_27740), .Q(_45529) );
  nnd2s1 _45852_inst ( .DIN1(_45534), .DIN2(_29083), .Q(_45524) );
  hi1s1 _45853_inst ( .DIN(_35902), .Q(_29083) );
  nnd2s1 _45854_inst ( .DIN1(_45535), .DIN2(_45536), .Q(_35902) );
  nor2s1 _45855_inst ( .DIN1(_45537), .DIN2(_39523), .Q(_45536) );
  nor2s1 _45856_inst ( .DIN1(_27746), .DIN2(_28857), .Q(_45535) );
  nnd2s1 _45857_inst ( .DIN1(_45538), .DIN2(_45539), .Q(_28857) );
  nor2s1 _45858_inst ( .DIN1(_39521), .DIN2(_45540), .Q(_45539) );
  and2s1 _45859_inst ( .DIN1(_45541), .DIN2(_39516), .Q(_45538) );
  nnd2s1 _45860_inst ( .DIN1(_45542), .DIN2(_45543), .Q(_27746) );
  nor2s1 _45861_inst ( .DIN1(_45544), .DIN2(_45545), .Q(_45543) );
  nnd2s1 _45862_inst ( .DIN1(_45546), .DIN2(_45532), .Q(_45545) );
  nnd2s1 _45863_inst ( .DIN1(_45547), .DIN2(_45533), .Q(_45544) );
  nor2s1 _45864_inst ( .DIN1(_45548), .DIN2(_45549), .Q(_45542) );
  nnd2s1 _45865_inst ( .DIN1(_45550), .DIN2(_45551), .Q(_45549) );
  nnd2s1 _45866_inst ( .DIN1(_45552), .DIN2(_45553), .Q(_45548) );
  nor2s1 _45867_inst ( .DIN1(_45554), .DIN2(_45555), .Q(_45534) );
  nnd2s1 _45868_inst ( .DIN1(_45556), .DIN2(_45557), .Q(_45555) );
  nor2s1 _45869_inst ( .DIN1(_45558), .DIN2(_45559), .Q(_45557) );
  nnd2s1 _45870_inst ( .DIN1(_45035), .DIN2(_45560), .Q(_45559) );
  hi1s1 _45871_inst ( .DIN(_44839), .Q(_45560) );
  nnd2s1 _45872_inst ( .DIN1(_45561), .DIN2(_45562), .Q(_44839) );
  nor2s1 _45873_inst ( .DIN1(_45563), .DIN2(_45564), .Q(_45562) );
  nnd2s1 _45874_inst ( .DIN1(_45565), .DIN2(_45058), .Q(_45564) );
  nnd2s1 _45875_inst ( .DIN1(_45183), .DIN2(_44951), .Q(_45058) );
  hi1s1 _45876_inst ( .DIN(_44756), .Q(_45183) );
  nnd2s1 _45877_inst ( .DIN1(_45566), .DIN2(_45567), .Q(_44756) );
  nor2s1 _45878_inst ( .DIN1(_45459), .DIN2(_45568), .Q(_45567) );
  nnd2s1 _45879_inst ( .DIN1(_45569), .DIN2(_45570), .Q(_45568) );
  nor2s1 _45880_inst ( .DIN1(_45571), .DIN2(_45572), .Q(_45566) );
  nnd2s1 _45881_inst ( .DIN1(_45573), .DIN2(_45574), .Q(_45572) );
  nnd2s1 _45882_inst ( .DIN1(_44773), .DIN2(_44771), .Q(_45565) );
  nnd2s1 _45883_inst ( .DIN1(_45300), .DIN2(_45106), .Q(_45563) );
  nnd2s1 _45884_inst ( .DIN1(_44924), .DIN2(_44771), .Q(_45106) );
  hi1s1 _45885_inst ( .DIN(_44893), .Q(_44924) );
  nnd2s1 _45886_inst ( .DIN1(_45575), .DIN2(_45576), .Q(_44893) );
  xor2s1 _45887_inst ( .DIN1(_31658), .DIN2(_45577), .Q(_45576) );
  hi1s1 _45888_inst ( .DIN(_30186), .Q(_31658) );
  nnd2s1 _45889_inst ( .DIN1(_45578), .DIN2(_45579), .Q(_30186) );
  nor2s1 _45890_inst ( .DIN1(_44578), .DIN2(_45580), .Q(_45579) );
  nnd2s1 _45891_inst ( .DIN1(_44626), .DIN2(_44573), .Q(_45580) );
  nor2s1 _45892_inst ( .DIN1(_42878), .DIN2(_45581), .Q(_45578) );
  nnd2s1 _45893_inst ( .DIN1(_44622), .DIN2(_44577), .Q(_45581) );
  nor2s1 _45894_inst ( .DIN1(_45582), .DIN2(_44574), .Q(_44622) );
  nnd2s1 _45895_inst ( .DIN1(_44997), .DIN2(_45583), .Q(_44574) );
  nnd2s1 _45896_inst ( .DIN1(_45584), .DIN2(_45585), .Q(_45583) );
  nnd2s1 _45897_inst ( .DIN1(_45002), .DIN2(_44995), .Q(_45582) );
  nnd2s1 _45898_inst ( .DIN1(_45586), .DIN2(_45587), .Q(_42878) );
  nnd2s1 _45899_inst ( .DIN1(_44030), .DIN2(_45588), .Q(_45586) );
  nor2s1 _45900_inst ( .DIN1(_45589), .DIN2(_45590), .Q(_45575) );
  nor2s1 _45901_inst ( .DIN1(_45591), .DIN2(_45592), .Q(_45561) );
  nnd2s1 _45902_inst ( .DIN1(_45593), .DIN2(_45594), .Q(_45592) );
  xor2s1 _45903_inst ( .DIN1(_45595), .DIN2(_31269), .Q(_45594) );
  hi1s1 _45904_inst ( .DIN(_43687), .Q(_31269) );
  nnd2s1 _45905_inst ( .DIN1(_30787), .DIN2(_45596), .Q(_43687) );
  hi1s1 _45906_inst ( .DIN(_29518), .Q(_30787) );
  nnd2s1 _45907_inst ( .DIN1(_44376), .DIN2(_44925), .Q(_29518) );
  nnd2s1 _45908_inst ( .DIN1(_45597), .DIN2(_45245), .Q(_45595) );
  nnd2s1 _45909_inst ( .DIN1(_44884), .DIN2(_44723), .Q(_45245) );
  hi1s1 _45910_inst ( .DIN(_45185), .Q(_44884) );
  nnd2s1 _45911_inst ( .DIN1(_45598), .DIN2(_45599), .Q(_45185) );
  nor2s1 _45912_inst ( .DIN1(_45459), .DIN2(_45577), .Q(_45599) );
  nor2s1 _45913_inst ( .DIN1(_45600), .DIN2(_45601), .Q(_45598) );
  nor2s1 _45914_inst ( .DIN1(_44785), .DIN2(_44767), .Q(_45597) );
  hi1s1 _45915_inst ( .DIN(_45602), .Q(_44785) );
  nor2s1 _45916_inst ( .DIN1(_45470), .DIN2(_45603), .Q(_45593) );
  nor2s1 _45917_inst ( .DIN1(_44912), .DIN2(_44723), .Q(_45603) );
  nor2s1 _45918_inst ( .DIN1(_26805), .DIN2(_44955), .Q(_45470) );
  nnd2s1 _45919_inst ( .DIN1(_45604), .DIN2(_45244), .Q(_45591) );
  and2s1 _45920_inst ( .DIN1(_45115), .DIN2(_45605), .Q(_45244) );
  nnd2s1 _45921_inst ( .DIN1(_45513), .DIN2(_26851), .Q(_45605) );
  nnd2s1 _45922_inst ( .DIN1(_45606), .DIN2(_45607), .Q(_45115) );
  nor2s1 _45923_inst ( .DIN1(_45590), .DIN2(_26852), .Q(_45606) );
  hi1s1 _45924_inst ( .DIN(_45011), .Q(_45604) );
  nnd2s1 _45925_inst ( .DIN1(_45608), .DIN2(_45609), .Q(_45011) );
  nnd2s1 _45926_inst ( .DIN1(_45320), .DIN2(_26852), .Q(_45609) );
  hi1s1 _45927_inst ( .DIN(_45105), .Q(_45320) );
  nnd2s1 _45928_inst ( .DIN1(_45610), .DIN2(_45611), .Q(_45105) );
  nnd2s1 _45929_inst ( .DIN1(_44710), .DIN2(_44771), .Q(_45608) );
  hi1s1 _45930_inst ( .DIN(_44828), .Q(_44710) );
  nnd2s1 _45931_inst ( .DIN1(_45612), .DIN2(_45613), .Q(_44828) );
  nor2s1 _45932_inst ( .DIN1(_38865), .DIN2(_45614), .Q(_45613) );
  nor2s1 _45933_inst ( .DIN1(_45615), .DIN2(_45601), .Q(_45612) );
  and2s1 _45934_inst ( .DIN1(_45616), .DIN2(_45617), .Q(_45035) );
  nnd2s1 _45935_inst ( .DIN1(_45335), .DIN2(_26767), .Q(_45617) );
  nnd2s1 _45936_inst ( .DIN1(_44965), .DIN2(_26805), .Q(_45616) );
  hi1s1 _45937_inst ( .DIN(_45618), .Q(_44965) );
  nnd2s1 _45938_inst ( .DIN1(_45261), .DIN2(_45619), .Q(_45558) );
  hi1s1 _45939_inst ( .DIN(_44735), .Q(_45619) );
  nnd2s1 _45940_inst ( .DIN1(_45620), .DIN2(_45621), .Q(_44735) );
  nor2s1 _45941_inst ( .DIN1(_45622), .DIN2(_45623), .Q(_45621) );
  nnd2s1 _45942_inst ( .DIN1(_45482), .DIN2(_45624), .Q(_45623) );
  nnd2s1 _45943_inst ( .DIN1(_45625), .DIN2(_44715), .Q(_45624) );
  nnd2s1 _45944_inst ( .DIN1(_45157), .DIN2(_26766), .Q(_45482) );
  nnd2s1 _45945_inst ( .DIN1(_45626), .DIN2(_45627), .Q(_45622) );
  nnd2s1 _45946_inst ( .DIN1(_44951), .DIN2(_45628), .Q(_45627) );
  nnd2s1 _45947_inst ( .DIN1(_45629), .DIN2(_44914), .Q(_45628) );
  nor2s1 _45948_inst ( .DIN1(_44821), .DIN2(_45630), .Q(_45629) );
  nor2s1 _45949_inst ( .DIN1(_45166), .DIN2(_45631), .Q(_45626) );
  hi1s1 _45950_inst ( .DIN(_44892), .Q(_45631) );
  nnd2s1 _45951_inst ( .DIN1(_45632), .DIN2(_44771), .Q(_44892) );
  and2s1 _45952_inst ( .DIN1(_26805), .DIN2(_45633), .Q(_45166) );
  nnd2s1 _45953_inst ( .DIN1(_45451), .DIN2(_45634), .Q(_45633) );
  nnd2s1 _45954_inst ( .DIN1(_45635), .DIN2(_45636), .Q(_45634) );
  nor2s1 _45955_inst ( .DIN1(_53477), .DIN2(_26219), .Q(_45636) );
  nor2s1 _45956_inst ( .DIN1(_45637), .DIN2(_45638), .Q(_45620) );
  or2s1 _45957_inst ( .DIN1(_45264), .DIN2(_45143), .Q(_45638) );
  nnd2s1 _45958_inst ( .DIN1(_45639), .DIN2(_45640), .Q(_45143) );
  nor2s1 _45959_inst ( .DIN1(_45641), .DIN2(_44885), .Q(_45640) );
  nor2s1 _45960_inst ( .DIN1(_45642), .DIN2(_45282), .Q(_45639) );
  nnd2s1 _45961_inst ( .DIN1(_44784), .DIN2(_45643), .Q(_45282) );
  nnd2s1 _45962_inst ( .DIN1(_45644), .DIN2(_45645), .Q(_45643) );
  nor2s1 _45963_inst ( .DIN1(_26767), .DIN2(_45313), .Q(_45642) );
  nnd2s1 _45964_inst ( .DIN1(_45646), .DIN2(_45647), .Q(_45264) );
  nnd2s1 _45965_inst ( .DIN1(_45648), .DIN2(_45645), .Q(_45647) );
  nor2s1 _45966_inst ( .DIN1(_44723), .DIN2(_45649), .Q(_45648) );
  nnd2s1 _45967_inst ( .DIN1(_45650), .DIN2(_45226), .Q(_45637) );
  and2s1 _45968_inst ( .DIN1(_45651), .DIN2(_45652), .Q(_45226) );
  or2s1 _45969_inst ( .DIN1(_45510), .DIN2(_26845), .Q(_45652) );
  nnd2s1 _45970_inst ( .DIN1(_45653), .DIN2(_26805), .Q(_45651) );
  nor2s1 _45971_inst ( .DIN1(_44803), .DIN2(_45170), .Q(_45650) );
  nnd2s1 _45972_inst ( .DIN1(_45654), .DIN2(_45516), .Q(_45170) );
  nnd2s1 _45973_inst ( .DIN1(_45644), .DIN2(_45655), .Q(_45516) );
  nor2s1 _45974_inst ( .DIN1(_45256), .DIN2(_45040), .Q(_45654) );
  nor2s1 _45975_inst ( .DIN1(_45656), .DIN2(_44957), .Q(_45040) );
  nnd2s1 _45976_inst ( .DIN1(_45657), .DIN2(_45658), .Q(_44803) );
  nnd2s1 _45977_inst ( .DIN1(_45659), .DIN2(_26767), .Q(_45658) );
  and2s1 _45978_inst ( .DIN1(_45660), .DIN2(_45661), .Q(_45261) );
  xor2s1 _45979_inst ( .DIN1(_27338), .DIN2(_45662), .Q(_45661) );
  nor2s1 _45980_inst ( .DIN1(_44771), .DIN2(_44857), .Q(_45662) );
  nnd2s1 _45981_inst ( .DIN1(_45663), .DIN2(_44929), .Q(_27329) );
  nor2s1 _45982_inst ( .DIN1(_45664), .DIN2(_44928), .Q(_45663) );
  nor2s1 _45983_inst ( .DIN1(_44822), .DIN2(_45665), .Q(_45660) );
  nor2s1 _45984_inst ( .DIN1(_45666), .DIN2(_26851), .Q(_45665) );
  nor2s1 _45985_inst ( .DIN1(_45667), .DIN2(_45175), .Q(_45666) );
  nor2s1 _45986_inst ( .DIN1(_45668), .DIN2(_45669), .Q(_45556) );
  nnd2s1 _45987_inst ( .DIN1(_44716), .DIN2(_45670), .Q(_45669) );
  hi1s1 _45988_inst ( .DIN(_45518), .Q(_45670) );
  nnd2s1 _45989_inst ( .DIN1(_45671), .DIN2(_45672), .Q(_45518) );
  nor2s1 _45990_inst ( .DIN1(_45673), .DIN2(_45674), .Q(_45672) );
  nor2s1 _45991_inst ( .DIN1(_26852), .DIN2(_44714), .Q(_45674) );
  nnd2s1 _45992_inst ( .DIN1(_45675), .DIN2(_45676), .Q(_44714) );
  nor2s1 _45993_inst ( .DIN1(_26219), .DIN2(_45168), .Q(_45675) );
  nor2s1 _45994_inst ( .DIN1(_45677), .DIN2(_44723), .Q(_45673) );
  nor2s1 _45995_inst ( .DIN1(_44966), .DIN2(_45678), .Q(_45677) );
  nnd2s1 _45996_inst ( .DIN1(_44883), .DIN2(_45124), .Q(_45678) );
  nnd2s1 _45997_inst ( .DIN1(_45679), .DIN2(_45680), .Q(_45124) );
  nor2s1 _45998_inst ( .DIN1(_45458), .DIN2(_45681), .Q(_45680) );
  nnd2s1 _45999_inst ( .DIN1(_53471), .DIN2(_26558), .Q(_45681) );
  nor2s1 _46000_inst ( .DIN1(_45682), .DIN2(_45683), .Q(_45679) );
  nor2s1 _46001_inst ( .DIN1(_44788), .DIN2(_45684), .Q(_45671) );
  nnd2s1 _46002_inst ( .DIN1(_45685), .DIN2(_45686), .Q(_45684) );
  nnd2s1 _46003_inst ( .DIN1(_44950), .DIN2(_26845), .Q(_45686) );
  hi1s1 _46004_inst ( .DIN(_45311), .Q(_44950) );
  nnd2s1 _46005_inst ( .DIN1(_45687), .DIN2(_45688), .Q(_45311) );
  nor2s1 _46006_inst ( .DIN1(_53474), .DIN2(_45689), .Q(_45688) );
  nor2s1 _46007_inst ( .DIN1(_45690), .DIN2(_45691), .Q(_45687) );
  nnd2s1 _46008_inst ( .DIN1(_45255), .DIN2(_44951), .Q(_45685) );
  nnd2s1 _46009_inst ( .DIN1(_44726), .DIN2(_45692), .Q(_44788) );
  nnd2s1 _46010_inst ( .DIN1(_45005), .DIN2(_44951), .Q(_45692) );
  hi1s1 _46011_inst ( .DIN(_45059), .Q(_45005) );
  nnd2s1 _46012_inst ( .DIN1(_45693), .DIN2(_45224), .Q(_44726) );
  nor2s1 _46013_inst ( .DIN1(_45496), .DIN2(_45277), .Q(_44716) );
  hi1s1 _46014_inst ( .DIN(_44827), .Q(_45277) );
  nnd2s1 _46015_inst ( .DIN1(_45694), .DIN2(_45695), .Q(_44827) );
  or2s1 _46016_inst ( .DIN1(_45007), .DIN2(_45302), .Q(_45668) );
  nnd2s1 _46017_inst ( .DIN1(_45696), .DIN2(_45697), .Q(_45302) );
  nor2s1 _46018_inst ( .DIN1(_45118), .DIN2(_45498), .Q(_45697) );
  hi1s1 _46019_inst ( .DIN(_44856), .Q(_45498) );
  nnd2s1 _46020_inst ( .DIN1(_45698), .DIN2(_45699), .Q(_44856) );
  nor2s1 _46021_inst ( .DIN1(_44958), .DIN2(_45700), .Q(_45699) );
  nor2s1 _46022_inst ( .DIN1(_45701), .DIN2(_45702), .Q(_45696) );
  nor2s1 _46023_inst ( .DIN1(_44951), .DIN2(_26770), .Q(_45702) );
  nor2s1 _46024_inst ( .DIN1(_44715), .DIN2(_45703), .Q(_45701) );
  nnd2s1 _46025_inst ( .DIN1(_45704), .DIN2(_45705), .Q(_45007) );
  nor2s1 _46026_inst ( .DIN1(_45321), .DIN2(_45490), .Q(_45705) );
  nor2s1 _46027_inst ( .DIN1(_44923), .DIN2(_45706), .Q(_45704) );
  nnd2s1 _46028_inst ( .DIN1(_45707), .DIN2(_45708), .Q(_45706) );
  nnd2s1 _46029_inst ( .DIN1(_45176), .DIN2(_26852), .Q(_45708) );
  hi1s1 _46030_inst ( .DIN(_45045), .Q(_45176) );
  nnd2s1 _46031_inst ( .DIN1(_26765), .DIN2(_26766), .Q(_45707) );
  nnd2s1 _46032_inst ( .DIN1(_45709), .DIN2(_45710), .Q(_45554) );
  nor2s1 _46033_inst ( .DIN1(_45711), .DIN2(_45712), .Q(_45710) );
  nnd2s1 _46034_inst ( .DIN1(_45713), .DIN2(_44897), .Q(_45712) );
  nnd2s1 _46035_inst ( .DIN1(_45714), .DIN2(_45444), .Q(_44897) );
  nor2s1 _46036_inst ( .DIN1(_38865), .DIN2(_45715), .Q(_45714) );
  nnd2s1 _46037_inst ( .DIN1(_44951), .DIN2(_45716), .Q(_45713) );
  nnd2s1 _46038_inst ( .DIN1(_45717), .DIN2(_45043), .Q(_45716) );
  nnd2s1 _46039_inst ( .DIN1(_45718), .DIN2(_44761), .Q(_45711) );
  nnd2s1 _46040_inst ( .DIN1(_45719), .DIN2(_45720), .Q(_44761) );
  nor2s1 _46041_inst ( .DIN1(_45690), .DIN2(_44958), .Q(_45719) );
  nor2s1 _46042_inst ( .DIN1(_44851), .DIN2(_44901), .Q(_45718) );
  nor2s1 _46043_inst ( .DIN1(_45721), .DIN2(_45722), .Q(_45709) );
  nnd2s1 _46044_inst ( .DIN1(_45317), .DIN2(_45723), .Q(_45722) );
  hi1s1 _46045_inst ( .DIN(_44763), .Q(_45723) );
  nnd2s1 _46046_inst ( .DIN1(_45724), .DIN2(_45725), .Q(_44763) );
  nnd2s1 _46047_inst ( .DIN1(_45507), .DIN2(_26851), .Q(_45725) );
  nnd2s1 _46048_inst ( .DIN1(_45726), .DIN2(_26767), .Q(_45724) );
  and2s1 _46049_inst ( .DIN1(_45727), .DIN2(_45728), .Q(_45317) );
  nnd2s1 _46050_inst ( .DIN1(_44987), .DIN2(_44771), .Q(_45728) );
  hi1s1 _46051_inst ( .DIN(_44805), .Q(_44987) );
  nnd2s1 _46052_inst ( .DIN1(_45729), .DIN2(_45730), .Q(_44805) );
  nor2s1 _46053_inst ( .DIN1(_45459), .DIN2(_45731), .Q(_45730) );
  nnd2s1 _46054_inst ( .DIN1(_45569), .DIN2(_53478), .Q(_45731) );
  nor2s1 _46055_inst ( .DIN1(_45571), .DIN2(_45732), .Q(_45729) );
  nnd2s1 _46056_inst ( .DIN1(_45573), .DIN2(_45676), .Q(_45732) );
  nnd2s1 _46057_inst ( .DIN1(_44715), .DIN2(_45733), .Q(_45727) );
  nnd2s1 _46058_inst ( .DIN1(_44963), .DIN2(_45514), .Q(_45733) );
  nnd2s1 _46059_inst ( .DIN1(_45734), .DIN2(_45735), .Q(_45721) );
  nnd2s1 _46060_inst ( .DIN1(_26766), .DIN2(_45736), .Q(_45735) );
  nnd2s1 _46061_inst ( .DIN1(_45165), .DIN2(_44825), .Q(_45736) );
  nnd2s1 _46062_inst ( .DIN1(_29221), .DIN2(_45737), .Q(
        ____0___________0_0_____) );
  nnd2s1 _46063_inst ( .DIN1(_45738), .DIN2(_45739), .Q(_45737) );
  nor2s1 _46064_inst ( .DIN1(_45740), .DIN2(_45741), .Q(_45739) );
  nnd2s1 _46065_inst ( .DIN1(_45742), .DIN2(_45743), .Q(_45741) );
  nor2s1 _46066_inst ( .DIN1(_45744), .DIN2(_45745), .Q(_45743) );
  nnd2s1 _46067_inst ( .DIN1(_45746), .DIN2(_45747), .Q(_45745) );
  nnd2s1 _46068_inst ( .DIN1(_45224), .DIN2(_45748), .Q(_45747) );
  nnd2s1 _46069_inst ( .DIN1(_45656), .DIN2(_45460), .Q(_45748) );
  nnd2s1 _46070_inst ( .DIN1(_45749), .DIN2(_53095), .Q(_45746) );
  nor2s1 _46071_inst ( .DIN1(_26463), .DIN2(_45181), .Q(_45744) );
  nor2s1 _46072_inst ( .DIN1(_45371), .DIN2(_45750), .Q(_45742) );
  nnd2s1 _46073_inst ( .DIN1(_45751), .DIN2(_45752), .Q(_45750) );
  or2s1 _46074_inst ( .DIN1(_45182), .DIN2(_26362), .Q(_45752) );
  hi1s1 _46075_inst ( .DIN(_44880), .Q(_45751) );
  nnd2s1 _46076_inst ( .DIN1(_44912), .DIN2(_45222), .Q(_44880) );
  nnd2s1 _46077_inst ( .DIN1(_45753), .DIN2(_45754), .Q(_45222) );
  nor2s1 _46078_inst ( .DIN1(_26219), .DIN2(_45755), .Q(_45754) );
  nnd2s1 _46079_inst ( .DIN1(_31888), .DIN2(_26325), .Q(_45755) );
  nor2s1 _46080_inst ( .DIN1(_38912), .DIN2(_45756), .Q(_45753) );
  xor2s1 _46081_inst ( .DIN1(_45757), .DIN2(_31462), .Q(_44912) );
  nnd2s1 _46082_inst ( .DIN1(_45758), .DIN2(_53476), .Q(_45757) );
  nor2s1 _46083_inst ( .DIN1(_38528), .DIN2(_45759), .Q(_45758) );
  nnd2s1 _46084_inst ( .DIN1(_44825), .DIN2(_45760), .Q(_45371) );
  nnd2s1 _46085_inst ( .DIN1(_44768), .DIN2(_26845), .Q(_45760) );
  hi1s1 _46086_inst ( .DIN(_45717), .Q(_44768) );
  nnd2s1 _46087_inst ( .DIN1(_45761), .DIN2(_45762), .Q(_45717) );
  nor2s1 _46088_inst ( .DIN1(_45763), .DIN2(_45764), .Q(_45762) );
  nor2s1 _46089_inst ( .DIN1(_45765), .DIN2(_45766), .Q(_45761) );
  nnd2s1 _46090_inst ( .DIN1(_45767), .DIN2(_45768), .Q(_44825) );
  xor2s1 _46091_inst ( .DIN1(_45769), .DIN2(_35821), .Q(_45768) );
  nnd2s1 _46092_inst ( .DIN1(_38345), .DIN2(_45770), .Q(_45769) );
  nor2s1 _46093_inst ( .DIN1(_45614), .DIN2(_45689), .Q(_45767) );
  nnd2s1 _46094_inst ( .DIN1(_45771), .DIN2(_45772), .Q(_45740) );
  nor2s1 _46095_inst ( .DIN1(_45257), .DIN2(_45773), .Q(_45772) );
  nnd2s1 _46096_inst ( .DIN1(_45357), .DIN2(_45273), .Q(_45773) );
  nnd2s1 _46097_inst ( .DIN1(_45635), .DIN2(_45774), .Q(_45273) );
  nor2s1 _46098_inst ( .DIN1(_45756), .DIN2(_45775), .Q(_45635) );
  or2s1 _46099_inst ( .DIN1(_45776), .DIN2(_45777), .Q(_45357) );
  and2s1 _46100_inst ( .DIN1(_45778), .DIN2(_45779), .Q(_45257) );
  nor2s1 _46101_inst ( .DIN1(_45775), .DIN2(_45780), .Q(_45778) );
  nor2s1 _46102_inst ( .DIN1(_45255), .DIN2(_45781), .Q(_45771) );
  nnd2s1 _46103_inst ( .DIN1(_45506), .DIN2(_44857), .Q(_45781) );
  nnd2s1 _46104_inst ( .DIN1(_45782), .DIN2(_45783), .Q(_44857) );
  hi1s1 _46105_inst ( .DIN(_44851), .Q(_45506) );
  nor2s1 _46106_inst ( .DIN1(_45784), .DIN2(_45785), .Q(_44851) );
  nnd2s1 _46107_inst ( .DIN1(_45676), .DIN2(_45783), .Q(_45784) );
  hi1s1 _46108_inst ( .DIN(_45786), .Q(_45676) );
  nor2s1 _46109_inst ( .DIN1(_45787), .DIN2(_45766), .Q(_45255) );
  nnd2s1 _46110_inst ( .DIN1(_45788), .DIN2(_45645), .Q(_45787) );
  nor2s1 _46111_inst ( .DIN1(_45789), .DIN2(_45790), .Q(_45738) );
  nnd2s1 _46112_inst ( .DIN1(_45791), .DIN2(_45792), .Q(_45790) );
  nor2s1 _46113_inst ( .DIN1(_45238), .DIN2(_45793), .Q(_45792) );
  nnd2s1 _46114_inst ( .DIN1(_45399), .DIN2(_45232), .Q(_45793) );
  and2s1 _46115_inst ( .DIN1(_45794), .DIN2(_45795), .Q(_45232) );
  nor2s1 _46116_inst ( .DIN1(_45632), .DIN2(_45796), .Q(_45795) );
  nnd2s1 _46117_inst ( .DIN1(_45045), .DIN2(_45059), .Q(_45796) );
  nnd2s1 _46118_inst ( .DIN1(_45797), .DIN2(_45798), .Q(_45059) );
  nor2s1 _46119_inst ( .DIN1(_45690), .DIN2(_45700), .Q(_45798) );
  nnd2s1 _46120_inst ( .DIN1(_53479), .DIN2(_26364), .Q(_45700) );
  nor2s1 _46121_inst ( .DIN1(_45764), .DIN2(_45799), .Q(_45797) );
  nnd2s1 _46122_inst ( .DIN1(_45800), .DIN2(_45801), .Q(_45045) );
  nor2s1 _46123_inst ( .DIN1(_45802), .DIN2(_45780), .Q(_45800) );
  hi1s1 _46124_inst ( .DIN(_44817), .Q(_45632) );
  nnd2s1 _46125_inst ( .DIN1(_45803), .DIN2(_45804), .Q(_44817) );
  nor2s1 _46126_inst ( .DIN1(_45802), .DIN2(_38528), .Q(_45804) );
  nor2s1 _46127_inst ( .DIN1(_45601), .DIN2(_45805), .Q(_45803) );
  xor2s1 _46128_inst ( .DIN1(_35821), .DIN2(_45806), .Q(_45805) );
  nor2s1 _46129_inst ( .DIN1(_53500), .DIN2(_45807), .Q(_45806) );
  and2s1 _46130_inst ( .DIN1(_45808), .DIN2(_45809), .Q(_35821) );
  nor2s1 _46131_inst ( .DIN1(_45810), .DIN2(_45811), .Q(_45809) );
  nnd2s1 _46132_inst ( .DIN1(_45812), .DIN2(_42924), .Q(_45811) );
  nnd2s1 _46133_inst ( .DIN1(_45813), .DIN2(_45814), .Q(_45810) );
  nor2s1 _46134_inst ( .DIN1(_44313), .DIN2(_45815), .Q(_45808) );
  or2s1 _46135_inst ( .DIN1(_44982), .DIN2(_44287), .Q(_45815) );
  nnd2s1 _46136_inst ( .DIN1(_45816), .DIN2(_45817), .Q(_44313) );
  nor2s1 _46137_inst ( .DIN1(_45818), .DIN2(_45819), .Q(_45817) );
  and2s1 _46138_inst ( .DIN1(_42927), .DIN2(_44282), .Q(_45816) );
  nor2s1 _46139_inst ( .DIN1(_45820), .DIN2(_45821), .Q(_44282) );
  nnd2s1 _46140_inst ( .DIN1(_45822), .DIN2(_45823), .Q(_45820) );
  nor2s1 _46141_inst ( .DIN1(_45037), .DIN2(_45824), .Q(_45794) );
  nnd2s1 _46142_inst ( .DIN1(_45825), .DIN2(_45826), .Q(_45824) );
  nnd2s1 _46143_inst ( .DIN1(_44885), .DIN2(_26805), .Q(_45826) );
  and2s1 _46144_inst ( .DIN1(_45827), .DIN2(_45779), .Q(_44885) );
  nnd2s1 _46145_inst ( .DIN1(_44961), .DIN2(_26845), .Q(_45825) );
  and2s1 _46146_inst ( .DIN1(_45828), .DIN2(_45829), .Q(_44961) );
  nor2s1 _46147_inst ( .DIN1(_53503), .DIN2(_45830), .Q(_45828) );
  nnd2s1 _46148_inst ( .DIN1(_45831), .DIN2(_45832), .Q(_45037) );
  nnd2s1 _46149_inst ( .DIN1(_45833), .DIN2(_45834), .Q(_45832) );
  nor2s1 _46150_inst ( .DIN1(_44958), .DIN2(_45775), .Q(_45833) );
  nnd2s1 _46151_inst ( .DIN1(_45644), .DIN2(_45801), .Q(_45831) );
  hi1s1 _46152_inst ( .DIN(_45835), .Q(_45801) );
  and2s1 _46153_inst ( .DIN1(_45043), .DIN2(_45836), .Q(_45399) );
  nnd2s1 _46154_inst ( .DIN1(_44767), .DIN2(_44951), .Q(_45836) );
  hi1s1 _46155_inst ( .DIN(_44891), .Q(_44767) );
  nnd2s1 _46156_inst ( .DIN1(_45837), .DIN2(_45574), .Q(_44891) );
  nnd2s1 _46157_inst ( .DIN1(_45838), .DIN2(_45611), .Q(_45043) );
  hi1s1 _46158_inst ( .DIN(_45839), .Q(_45838) );
  nnd2s1 _46159_inst ( .DIN1(_45067), .DIN2(_45132), .Q(_45238) );
  nnd2s1 _46160_inst ( .DIN1(_45840), .DIN2(_45841), .Q(_45132) );
  nor2s1 _46161_inst ( .DIN1(_38912), .DIN2(_45842), .Q(_45841) );
  nor2s1 _46162_inst ( .DIN1(_44958), .DIN2(_45843), .Q(_45840) );
  nnd2s1 _46163_inst ( .DIN1(_45844), .DIN2(_45845), .Q(_45067) );
  nor2s1 _46164_inst ( .DIN1(_45169), .DIN2(_45839), .Q(_45844) );
  nnd2s1 _46165_inst ( .DIN1(_45846), .DIN2(_45573), .Q(_45839) );
  nor2s1 _46166_inst ( .DIN1(_38528), .DIN2(_37403), .Q(_45846) );
  nor2s1 _46167_inst ( .DIN1(_45847), .DIN2(_45848), .Q(_45791) );
  nnd2s1 _46168_inst ( .DIN1(_45849), .DIN2(_45850), .Q(_45848) );
  nnd2s1 _46169_inst ( .DIN1(_44966), .DIN2(_26805), .Q(_45850) );
  hi1s1 _46170_inst ( .DIN(_45229), .Q(_44966) );
  nnd2s1 _46171_inst ( .DIN1(_45851), .DIN2(_45852), .Q(_45229) );
  nor2s1 _46172_inst ( .DIN1(_53471), .DIN2(_53472), .Q(_45852) );
  nor2s1 _46173_inst ( .DIN1(_45656), .DIN2(_45853), .Q(_45851) );
  nnd2s1 _46174_inst ( .DIN1(_45854), .DIN2(_44723), .Q(_45849) );
  nnd2s1 _46175_inst ( .DIN1(_45451), .DIN2(_45855), .Q(_45854) );
  nnd2s1 _46176_inst ( .DIN1(_45645), .DIN2(_45856), .Q(_45855) );
  nnd2s1 _46177_inst ( .DIN1(_45857), .DIN2(_45774), .Q(_45451) );
  nor2s1 _46178_inst ( .DIN1(_53478), .DIN2(_26325), .Q(_45774) );
  nor2s1 _46179_inst ( .DIN1(_45756), .DIN2(_45835), .Q(_45857) );
  hi1s1 _46180_inst ( .DIN(_45788), .Q(_45756) );
  xor2s1 _46181_inst ( .DIN1(_31307), .DIN2(_45858), .Q(_45847) );
  nnd2s1 _46182_inst ( .DIN1(_45859), .DIN2(_45860), .Q(_45858) );
  nnd2s1 _46183_inst ( .DIN1(_45861), .DIN2(_26851), .Q(_45860) );
  nnd2s1 _46184_inst ( .DIN1(_45862), .DIN2(_45863), .Q(_45861) );
  nnd2s1 _46185_inst ( .DIN1(_45659), .DIN2(_26534), .Q(_45863) );
  hi1s1 _46186_inst ( .DIN(_45186), .Q(_45659) );
  nnd2s1 _46187_inst ( .DIN1(_45864), .DIN2(_45865), .Q(_45186) );
  nor2s1 _46188_inst ( .DIN1(_45777), .DIN2(_45656), .Q(_45864) );
  nnd2s1 _46189_inst ( .DIN1(_45866), .DIN2(_45770), .Q(_45777) );
  hi1s1 _46190_inst ( .DIN(_45458), .Q(_45770) );
  nor2s1 _46191_inst ( .DIN1(_45314), .DIN2(_45370), .Q(_45862) );
  hi1s1 _46192_inst ( .DIN(_45164), .Q(_45370) );
  nnd2s1 _46193_inst ( .DIN1(_45607), .DIN2(_45867), .Q(_45164) );
  and2s1 _46194_inst ( .DIN1(_45868), .DIN2(_45645), .Q(_45607) );
  and2s1 _46195_inst ( .DIN1(_45869), .DIN2(_45870), .Q(_45314) );
  nor2s1 _46196_inst ( .DIN1(_45786), .DIN2(_45871), .Q(_45869) );
  nor2s1 _46197_inst ( .DIN1(_44730), .DIN2(_45872), .Q(_45859) );
  nor2s1 _46198_inst ( .DIN1(_45871), .DIN2(_45873), .Q(_45872) );
  nnd2s1 _46199_inst ( .DIN1(_45655), .DIN2(_45874), .Q(_45873) );
  nor2s1 _46200_inst ( .DIN1(_45300), .DIN2(_44951), .Q(_44730) );
  nnd2s1 _46201_inst ( .DIN1(_45875), .DIN2(_45876), .Q(_45300) );
  nor2s1 _46202_inst ( .DIN1(_53474), .DIN2(_53503), .Q(_45876) );
  nor2s1 _46203_inst ( .DIN1(_45877), .DIN2(_45766), .Q(_45875) );
  nnd2s1 _46204_inst ( .DIN1(_26325), .DIN2(_26219), .Q(_45766) );
  nnd2s1 _46205_inst ( .DIN1(_45878), .DIN2(_30163), .Q(_31307) );
  nor2s1 _46206_inst ( .DIN1(_41912), .DIN2(_41914), .Q(_45878) );
  nnd2s1 _46207_inst ( .DIN1(_45879), .DIN2(_45880), .Q(_45789) );
  nor2s1 _46208_inst ( .DIN1(_44923), .DIN2(_45881), .Q(_45880) );
  nnd2s1 _46209_inst ( .DIN1(_45344), .DIN2(_45882), .Q(_45881) );
  hi1s1 _46210_inst ( .DIN(_44780), .Q(_45882) );
  nnd2s1 _46211_inst ( .DIN1(_45155), .DIN2(_45883), .Q(_44780) );
  nnd2s1 _46212_inst ( .DIN1(_45321), .DIN2(_26845), .Q(_45883) );
  hi1s1 _46213_inst ( .DIN(_44854), .Q(_45321) );
  nnd2s1 _46214_inst ( .DIN1(_45884), .DIN2(_45885), .Q(_44854) );
  nnd2s1 _46215_inst ( .DIN1(_45886), .DIN2(_45887), .Q(_45155) );
  nor2s1 _46216_inst ( .DIN1(_31459), .DIN2(_45802), .Q(_45887) );
  nor2s1 _46217_inst ( .DIN1(_45842), .DIN2(_36898), .Q(_45886) );
  and2s1 _46218_inst ( .DIN1(_45888), .DIN2(_45889), .Q(_45344) );
  or2s1 _46219_inst ( .DIN1(_45165), .DIN2(_26767), .Q(_45889) );
  nnd2s1 _46220_inst ( .DIN1(_45890), .DIN2(_45891), .Q(_45165) );
  nor2s1 _46221_inst ( .DIN1(_45682), .DIN2(_45892), .Q(_45891) );
  nnd2s1 _46222_inst ( .DIN1(_45569), .DIN2(_45893), .Q(_45892) );
  nor2s1 _46223_inst ( .DIN1(_45571), .DIN2(_45601), .Q(_45890) );
  nnd2s1 _46224_inst ( .DIN1(_45513), .DIN2(_26766), .Q(_45888) );
  and2s1 _46225_inst ( .DIN1(_45894), .DIN2(_45895), .Q(_45513) );
  nor2s1 _46226_inst ( .DIN1(_45764), .DIN2(_45896), .Q(_45895) );
  nor2s1 _46227_inst ( .DIN1(_45656), .DIN2(_45765), .Q(_45894) );
  xnr2s1 _46228_inst ( .DIN1(_26321), .DIN2(_45897), .Q(_44923) );
  nor2s1 _46229_inst ( .DIN1(_45898), .DIN2(_45899), .Q(_45897) );
  nnd2s1 _46230_inst ( .DIN1(_45900), .DIN2(_45901), .Q(_45899) );
  nnd2s1 _46231_inst ( .DIN1(_45902), .DIN2(_45903), .Q(_45898) );
  hi1s1 _46232_inst ( .DIN(_45802), .Q(_45903) );
  nor2s1 _46233_inst ( .DIN1(_45904), .DIN2(_38865), .Q(_45902) );
  nor2s1 _46234_inst ( .DIN1(_45050), .DIN2(_45905), .Q(_45879) );
  nnd2s1 _46235_inst ( .DIN1(_44875), .DIN2(_44836), .Q(_45905) );
  and2s1 _46236_inst ( .DIN1(_45906), .DIN2(_45907), .Q(_44836) );
  nor2s1 _46237_inst ( .DIN1(_45908), .DIN2(_45909), .Q(_45907) );
  nnd2s1 _46238_inst ( .DIN1(_45910), .DIN2(_44883), .Q(_45909) );
  hi1s1 _46239_inst ( .DIN(_45253), .Q(_44883) );
  nor2s1 _46240_inst ( .DIN1(_45911), .DIN2(_45799), .Q(_45253) );
  or2s1 _46241_inst ( .DIN1(_45590), .DIN2(_45683), .Q(_45911) );
  nor2s1 _46242_inst ( .DIN1(_44871), .DIN2(_45496), .Q(_45910) );
  hi1s1 _46243_inst ( .DIN(_45291), .Q(_45496) );
  nnd2s1 _46244_inst ( .DIN1(_45912), .DIN2(_45913), .Q(_45291) );
  hi1s1 _46245_inst ( .DIN(_45313), .Q(_44871) );
  nnd2s1 _46246_inst ( .DIN1(_45914), .DIN2(_45915), .Q(_45313) );
  nor2s1 _46247_inst ( .DIN1(_45577), .DIN2(_45600), .Q(_45914) );
  nnd2s1 _46248_inst ( .DIN1(_45916), .DIN2(_45901), .Q(_45577) );
  nor2s1 _46249_inst ( .DIN1(_45917), .DIN2(_38865), .Q(_45916) );
  nnd2s1 _46250_inst ( .DIN1(_45918), .DIN2(_45919), .Q(_45908) );
  nor2s1 _46251_inst ( .DIN1(_45630), .DIN2(_44753), .Q(_45919) );
  nor2s1 _46252_inst ( .DIN1(_44818), .DIN2(_44951), .Q(_44753) );
  nnd2s1 _46253_inst ( .DIN1(_45694), .DIN2(_38345), .Q(_44818) );
  and2s1 _46254_inst ( .DIN1(_45920), .DIN2(_45611), .Q(_45694) );
  nor2s1 _46255_inst ( .DIN1(_45715), .DIN2(_45571), .Q(_45920) );
  hi1s1 _46256_inst ( .DIN(_45301), .Q(_45630) );
  nnd2s1 _46257_inst ( .DIN1(_45921), .DIN2(_45720), .Q(_45301) );
  hi1s1 _46258_inst ( .DIN(_45853), .Q(_45720) );
  nor2s1 _46259_inst ( .DIN1(_45690), .DIN2(_45799), .Q(_45921) );
  nor2s1 _46260_inst ( .DIN1(_44766), .DIN2(_45397), .Q(_45918) );
  hi1s1 _46261_inst ( .DIN(_45703), .Q(_45397) );
  nnd2s1 _46262_inst ( .DIN1(_45922), .DIN2(_45923), .Q(_45703) );
  nor2s1 _46263_inst ( .DIN1(_53472), .DIN2(_26222), .Q(_45923) );
  nor2s1 _46264_inst ( .DIN1(_45924), .DIN2(_45691), .Q(_45922) );
  hi1s1 _46265_inst ( .DIN(_44820), .Q(_44766) );
  nnd2s1 _46266_inst ( .DIN1(_45335), .DIN2(_26852), .Q(_44820) );
  nor2s1 _46267_inst ( .DIN1(_45925), .DIN2(_45759), .Q(_45335) );
  nnd2s1 _46268_inst ( .DIN1(_26233), .DIN2(_45569), .Q(_45925) );
  hi1s1 _46269_inst ( .DIN(_38865), .Q(_45569) );
  nor2s1 _46270_inst ( .DIN1(_45926), .DIN2(_45927), .Q(_45906) );
  nnd2s1 _46271_inst ( .DIN1(_45928), .DIN2(_45929), .Q(_45927) );
  hi1s1 _46272_inst ( .DIN(_45012), .Q(_45929) );
  nnd2s1 _46273_inst ( .DIN1(_45930), .DIN2(_45931), .Q(_45012) );
  nor2s1 _46274_inst ( .DIN1(_45653), .DIN2(_45932), .Q(_45931) );
  nnd2s1 _46275_inst ( .DIN1(_45514), .DIN2(_45510), .Q(_45932) );
  nnd2s1 _46276_inst ( .DIN1(_45782), .DIN2(_45933), .Q(_45510) );
  nor2s1 _46277_inst ( .DIN1(_53477), .DIN2(_45763), .Q(_45782) );
  nnd2s1 _46278_inst ( .DIN1(_45934), .DIN2(_45913), .Q(_45514) );
  nor2s1 _46279_inst ( .DIN1(_53503), .DIN2(_26416), .Q(_45934) );
  hi1s1 _46280_inst ( .DIN(_45379), .Q(_45653) );
  nnd2s1 _46281_inst ( .DIN1(_45935), .DIN2(_45913), .Q(_45379) );
  nor2s1 _46282_inst ( .DIN1(_45936), .DIN2(_45937), .Q(_45930) );
  nnd2s1 _46283_inst ( .DIN1(_45938), .DIN2(_45939), .Q(_45937) );
  nnd2s1 _46284_inst ( .DIN1(_45726), .DIN2(_26851), .Q(_45939) );
  hi1s1 _46285_inst ( .DIN(_45393), .Q(_45726) );
  nnd2s1 _46286_inst ( .DIN1(_45940), .DIN2(_45941), .Q(_45393) );
  nor2s1 _46287_inst ( .DIN1(_53478), .DIN2(_45924), .Q(_45941) );
  nor2s1 _46288_inst ( .DIN1(_45785), .DIN2(_45853), .Q(_45940) );
  nnd2s1 _46289_inst ( .DIN1(_45935), .DIN2(_45942), .Q(_45853) );
  nor2s1 _46290_inst ( .DIN1(_53479), .DIN2(_26364), .Q(_45935) );
  nnd2s1 _46291_inst ( .DIN1(_45507), .DIN2(_26767), .Q(_45938) );
  hi1s1 _46292_inst ( .DIN(_45310), .Q(_45507) );
  nnd2s1 _46293_inst ( .DIN1(_45943), .DIN2(_45829), .Q(_45310) );
  hi1s1 _46294_inst ( .DIN(_45877), .Q(_45829) );
  nnd2s1 _46295_inst ( .DIN1(_45944), .DIN2(_45945), .Q(_45877) );
  nor2s1 _46296_inst ( .DIN1(_26231), .DIN2(_45946), .Q(_45945) );
  nnd2s1 _46297_inst ( .DIN1(_26416), .DIN2(_26222), .Q(_45946) );
  nor2s1 _46298_inst ( .DIN1(_45601), .DIN2(_45947), .Q(_45944) );
  nnd2s1 _46299_inst ( .DIN1(_45948), .DIN2(_53473), .Q(_45947) );
  nor2s1 _46300_inst ( .DIN1(_26364), .DIN2(_45830), .Q(_45943) );
  nnd2s1 _46301_inst ( .DIN1(_45949), .DIN2(_45950), .Q(_45936) );
  nnd2s1 _46302_inst ( .DIN1(_45625), .DIN2(_44771), .Q(_45950) );
  hi1s1 _46303_inst ( .DIN(_45133), .Q(_45625) );
  nnd2s1 _46304_inst ( .DIN1(_45951), .DIN2(_38345), .Q(_45133) );
  nor2s1 _46305_inst ( .DIN1(_53476), .DIN2(_45759), .Q(_45951) );
  nnd2s1 _46306_inst ( .DIN1(_45952), .DIN2(_45953), .Q(_45759) );
  nor2s1 _46307_inst ( .DIN1(_45917), .DIN2(_45954), .Q(_45953) );
  nnd2s1 _46308_inst ( .DIN1(_53500), .DIN2(_26369), .Q(_45954) );
  nor2s1 _46309_inst ( .DIN1(_45589), .DIN2(_45955), .Q(_45952) );
  nnd2s1 _46310_inst ( .DIN1(_45956), .DIN2(_45957), .Q(_45955) );
  nnd2s1 _46311_inst ( .DIN1(_45749), .DIN2(_44715), .Q(_45949) );
  hi1s1 _46312_inst ( .DIN(_44899), .Q(_45749) );
  nnd2s1 _46313_inst ( .DIN1(_45958), .DIN2(_45223), .Q(_44899) );
  nor2s1 _46314_inst ( .DIN1(_45022), .DIN2(_44872), .Q(_45928) );
  nnd2s1 _46315_inst ( .DIN1(_45959), .DIN2(_45960), .Q(_44872) );
  nnd2s1 _46316_inst ( .DIN1(_45641), .DIN2(_44951), .Q(_45960) );
  hi1s1 _46317_inst ( .DIN(_45279), .Q(_45641) );
  nnd2s1 _46318_inst ( .DIN1(_45961), .DIN2(_45693), .Q(_45279) );
  hi1s1 _46319_inst ( .DIN(_45169), .Q(_45693) );
  nor2s1 _46320_inst ( .DIN1(_45842), .DIN2(_45775), .Q(_45961) );
  or2s1 _46321_inst ( .DIN1(_45266), .DIN2(_26804), .Q(_45959) );
  nnd2s1 _46322_inst ( .DIN1(_45962), .DIN2(_45963), .Q(_45266) );
  nor2s1 _46323_inst ( .DIN1(_31459), .DIN2(_45590), .Q(_45963) );
  nnd2s1 _46324_inst ( .DIN1(_45964), .DIN2(_45957), .Q(_45590) );
  hi1s1 _46325_inst ( .DIN(_45459), .Q(_45957) );
  nor2s1 _46326_inst ( .DIN1(_45682), .DIN2(_36898), .Q(_45962) );
  nnd2s1 _46327_inst ( .DIN1(_45965), .DIN2(_45966), .Q(_45022) );
  nnd2s1 _46328_inst ( .DIN1(_45118), .DIN2(_26766), .Q(_45966) );
  hi1s1 _46329_inst ( .DIN(_44759), .Q(_45118) );
  nnd2s1 _46330_inst ( .DIN1(_45967), .DIN2(_45958), .Q(_44759) );
  nor2s1 _46331_inst ( .DIN1(_45968), .DIN2(_45780), .Q(_45958) );
  or2s1 _46332_inst ( .DIN1(_31459), .DIN2(_36898), .Q(_45968) );
  nor2s1 _46333_inst ( .DIN1(_26219), .DIN2(_45786), .Q(_45967) );
  nnd2s1 _46334_inst ( .DIN1(_45574), .DIN2(_26565), .Q(_45786) );
  hi1s1 _46335_inst ( .DIN(_45589), .Q(_45574) );
  nnd2s1 _46336_inst ( .DIN1(_53475), .DIN2(_26325), .Q(_45589) );
  and2s1 _46337_inst ( .DIN1(_45295), .DIN2(_45294), .Q(_45965) );
  nnd2s1 _46338_inst ( .DIN1(_45969), .DIN2(_45783), .Q(_45294) );
  hi1s1 _46339_inst ( .DIN(_45970), .Q(_45783) );
  nnd2s1 _46340_inst ( .DIN1(_45913), .DIN2(_45885), .Q(_45295) );
  and2s1 _46341_inst ( .DIN1(_45698), .DIN2(_45868), .Q(_45913) );
  nor2s1 _46342_inst ( .DIN1(_53475), .DIN2(_45830), .Q(_45868) );
  nor2s1 _46343_inst ( .DIN1(_45764), .DIN2(_45785), .Q(_45698) );
  nnd2s1 _46344_inst ( .DIN1(_53472), .DIN2(_26222), .Q(_45785) );
  nnd2s1 _46345_inst ( .DIN1(_45971), .DIN2(_45972), .Q(_45926) );
  nor2s1 _46346_inst ( .DIN1(_45973), .DIN2(_45336), .Q(_45972) );
  nor2s1 _46347_inst ( .DIN1(_26851), .DIN2(_44784), .Q(_45336) );
  nnd2s1 _46348_inst ( .DIN1(_45974), .DIN2(_45975), .Q(_44784) );
  nor2s1 _46349_inst ( .DIN1(_53474), .DIN2(_45683), .Q(_45975) );
  nor2s1 _46350_inst ( .DIN1(_45871), .DIN2(_45600), .Q(_45974) );
  and2s1 _46351_inst ( .DIN1(_45645), .DIN2(_45644), .Q(_45973) );
  nor2s1 _46352_inst ( .DIN1(_45976), .DIN2(_45871), .Q(_45644) );
  nnd2s1 _46353_inst ( .DIN1(_26805), .DIN2(_45874), .Q(_45976) );
  nor2s1 _46354_inst ( .DIN1(_45977), .DIN2(_44702), .Q(_45971) );
  nnd2s1 _46355_inst ( .DIN1(_45978), .DIN2(_45979), .Q(_44702) );
  nnd2s1 _46356_inst ( .DIN1(_44772), .DIN2(_44771), .Q(_45979) );
  hi1s1 _46357_inst ( .DIN(_44963), .Q(_44772) );
  nnd2s1 _46358_inst ( .DIN1(_45912), .DIN2(_45884), .Q(_44963) );
  and2s1 _46359_inst ( .DIN1(_45980), .DIN2(_45981), .Q(_45884) );
  nor2s1 _46360_inst ( .DIN1(_26222), .DIN2(_45982), .Q(_45981) );
  nnd2s1 _46361_inst ( .DIN1(_26231), .DIN2(_26369), .Q(_45982) );
  nor2s1 _46362_inst ( .DIN1(_45830), .DIN2(_45764), .Q(_45980) );
  hi1s1 _46363_inst ( .DIN(_45765), .Q(_45912) );
  nnd2s1 _46364_inst ( .DIN1(_53479), .DIN2(_53503), .Q(_45765) );
  nnd2s1 _46365_inst ( .DIN1(_45667), .DIN2(_26851), .Q(_45978) );
  hi1s1 _46366_inst ( .DIN(_45509), .Q(_45667) );
  nnd2s1 _46367_inst ( .DIN1(_45983), .DIN2(_45984), .Q(_45509) );
  nor2s1 _46368_inst ( .DIN1(_53474), .DIN2(_45896), .Q(_45984) );
  nnd2s1 _46369_inst ( .DIN1(_26369), .DIN2(_26222), .Q(_45896) );
  nor2s1 _46370_inst ( .DIN1(_45689), .DIN2(_45970), .Q(_45983) );
  nnd2s1 _46371_inst ( .DIN1(_45985), .DIN2(_45942), .Q(_45970) );
  hi1s1 _46372_inst ( .DIN(_45764), .Q(_45942) );
  and2s1 _46373_inst ( .DIN1(_26219), .DIN2(_45885), .Q(_45985) );
  nor2s1 _46374_inst ( .DIN1(_53479), .DIN2(_53503), .Q(_45885) );
  nor2s1 _46375_inst ( .DIN1(_26805), .DIN2(_45618), .Q(_45977) );
  nnd2s1 _46376_inst ( .DIN1(_45837), .DIN2(_45986), .Q(_45618) );
  and2s1 _46377_inst ( .DIN1(_45987), .DIN2(_45573), .Q(_45837) );
  nor2s1 _46378_inst ( .DIN1(_45614), .DIN2(_37922), .Q(_45987) );
  and2s1 _46379_inst ( .DIN1(_45988), .DIN2(_45989), .Q(_44875) );
  nor2s1 _46380_inst ( .DIN1(_45990), .DIN2(_45991), .Q(_45989) );
  nnd2s1 _46381_inst ( .DIN1(_45484), .DIN2(_44826), .Q(_45991) );
  nnd2s1 _46382_inst ( .DIN1(_45992), .DIN2(_45993), .Q(_44826) );
  nor2s1 _46383_inst ( .DIN1(_45614), .DIN2(_38528), .Q(_45993) );
  hi1s1 _46384_inst ( .DIN(_45994), .Q(_45614) );
  and2s1 _46385_inst ( .DIN1(_45573), .DIN2(_45995), .Q(_45992) );
  nnd2s1 _46386_inst ( .DIN1(_45996), .DIN2(_45610), .Q(_45484) );
  and2s1 _46387_inst ( .DIN1(_45997), .DIN2(_45900), .Q(_45610) );
  hi1s1 _46388_inst ( .DIN(_45601), .Q(_45900) );
  nor2s1 _46389_inst ( .DIN1(_37922), .DIN2(_45571), .Q(_45997) );
  nor2s1 _46390_inst ( .DIN1(_45998), .DIN2(_45689), .Q(_45996) );
  nnd2s1 _46391_inst ( .DIN1(_45999), .DIN2(_44724), .Q(_45990) );
  nnd2s1 _46392_inst ( .DIN1(_46000), .DIN2(_46001), .Q(_44724) );
  nor2s1 _46393_inst ( .DIN1(_45459), .DIN2(_46002), .Q(_46001) );
  nnd2s1 _46394_inst ( .DIN1(_45445), .DIN2(_45570), .Q(_46002) );
  nor2s1 _46395_inst ( .DIN1(_45571), .DIN2(_45600), .Q(_46000) );
  and2s1 _46396_inst ( .DIN1(_45290), .DIN2(_45646), .Q(_45999) );
  nnd2s1 _46397_inst ( .DIN1(_46003), .DIN2(_46004), .Q(_45646) );
  nor2s1 _46398_inst ( .DIN1(_45843), .DIN2(_46005), .Q(_46004) );
  nnd2s1 _46399_inst ( .DIN1(_46006), .DIN2(_45867), .Q(_46005) );
  nor2s1 _46400_inst ( .DIN1(_26852), .DIN2(_45169), .Q(_46003) );
  nnd2s1 _46401_inst ( .DIN1(_46007), .DIN2(_45994), .Q(_45290) );
  nor2s1 _46402_inst ( .DIN1(_46008), .DIN2(_46009), .Q(_45988) );
  or2s1 _46403_inst ( .DIN1(_45142), .DIN2(_26765), .Q(_46009) );
  nor2s1 _46404_inst ( .DIN1(_46011), .DIN2(_46012), .Q(_46010) );
  nnd2s1 _46405_inst ( .DIN1(_46013), .DIN2(_45573), .Q(_46012) );
  nor2s1 _46406_inst ( .DIN1(_26233), .DIN2(_53472), .Q(_45573) );
  xnr2s1 _46407_inst ( .DIN1(_37577), .DIN2(_45807), .Q(_46013) );
  nnd2s1 _46408_inst ( .DIN1(_45893), .DIN2(_34289), .Q(_45807) );
  nnd2s1 _46409_inst ( .DIN1(_46014), .DIN2(_46015), .Q(_37577) );
  nor2s1 _46410_inst ( .DIN1(_44287), .DIN2(_44981), .Q(_46015) );
  nnd2s1 _46411_inst ( .DIN1(_45822), .DIN2(_46016), .Q(_44981) );
  nor2s1 _46412_inst ( .DIN1(_44317), .DIN2(_45071), .Q(_46014) );
  nnd2s1 _46413_inst ( .DIN1(_46017), .DIN2(_46018), .Q(_45071) );
  nor2s1 _46414_inst ( .DIN1(_46019), .DIN2(_46020), .Q(_46018) );
  nnd2s1 _46415_inst ( .DIN1(_46021), .DIN2(_46022), .Q(_46020) );
  nor2s1 _46416_inst ( .DIN1(_44982), .DIN2(_45821), .Q(_46017) );
  nnd2s1 _46417_inst ( .DIN1(_46023), .DIN2(_44984), .Q(_45821) );
  nnd2s1 _46418_inst ( .DIN1(_46024), .DIN2(_46025), .Q(_44984) );
  nor2s1 _46419_inst ( .DIN1(_46026), .DIN2(_46027), .Q(_46023) );
  nnd2s1 _46420_inst ( .DIN1(_45095), .DIN2(_46028), .Q(_44982) );
  nor2s1 _46421_inst ( .DIN1(_46029), .DIN2(_46030), .Q(_45095) );
  nnd2s1 _46422_inst ( .DIN1(_46031), .DIN2(_38345), .Q(_46011) );
  hi1s1 _46423_inst ( .DIN(_37922), .Q(_38345) );
  nor2s1 _46424_inst ( .DIN1(_26241), .DIN2(_45682), .Q(_46031) );
  nnd2s1 _46425_inst ( .DIN1(_45874), .DIN2(_53478), .Q(_45682) );
  hi1s1 _46426_inst ( .DIN(_45924), .Q(_45874) );
  xor2s1 _46427_inst ( .DIN1(_29599), .DIN2(_46032), .Q(_45142) );
  nor2s1 _46428_inst ( .DIN1(_26766), .DIN2(_45602), .Q(_46032) );
  nnd2s1 _46429_inst ( .DIN1(_46033), .DIN2(_46007), .Q(_45602) );
  and2s1 _46430_inst ( .DIN1(_46034), .DIN2(_45995), .Q(_46007) );
  nor2s1 _46431_inst ( .DIN1(_45715), .DIN2(_37922), .Q(_46034) );
  nnd2s1 _46432_inst ( .DIN1(_46035), .DIN2(_53503), .Q(_37922) );
  nor2s1 _46433_inst ( .DIN1(_53501), .DIN2(_26467), .Q(_46035) );
  nor2s1 _46434_inst ( .DIN1(_45998), .DIN2(_37403), .Q(_46033) );
  hi1s1 _46435_inst ( .DIN(_37792), .Q(_29599) );
  nor2s1 _46436_inst ( .DIN1(_29579), .DIN2(_41914), .Q(_37792) );
  nnd2s1 _46437_inst ( .DIN1(_46036), .DIN2(_44079), .Q(_29579) );
  nor2s1 _46438_inst ( .DIN1(_43949), .DIN2(_41912), .Q(_46036) );
  nnd2s1 _46439_inst ( .DIN1(_45275), .DIN2(_46037), .Q(_46008) );
  nnd2s1 _46440_inst ( .DIN1(_46038), .DIN2(_45223), .Q(_46037) );
  nor2s1 _46441_inst ( .DIN1(_26805), .DIN2(_45168), .Q(_46038) );
  nnd2s1 _46442_inst ( .DIN1(_44821), .DIN2(_26845), .Q(_45275) );
  hi1s1 _46443_inst ( .DIN(_45387), .Q(_44821) );
  nnd2s1 _46444_inst ( .DIN1(_46039), .DIN2(_46040), .Q(_45387) );
  nor2s1 _46445_inst ( .DIN1(_45571), .DIN2(_46041), .Q(_46040) );
  nnd2s1 _46446_inst ( .DIN1(_45695), .DIN2(_45570), .Q(_46041) );
  hi1s1 _46447_inst ( .DIN(_38528), .Q(_45695) );
  nnd2s1 _46448_inst ( .DIN1(_45956), .DIN2(_26241), .Q(_45571) );
  nor2s1 _46449_inst ( .DIN1(_45780), .DIN2(_45600), .Q(_46039) );
  nnd2s1 _46450_inst ( .DIN1(_46042), .DIN2(_46043), .Q(_45050) );
  nor2s1 _46451_inst ( .DIN1(_46044), .DIN2(_46045), .Q(_46043) );
  nnd2s1 _46452_inst ( .DIN1(_46046), .DIN2(_45657), .Q(_46045) );
  hi1s1 _46453_inst ( .DIN(_45364), .Q(_45657) );
  nor2s1 _46454_inst ( .DIN1(_45182), .DIN2(_44723), .Q(_45364) );
  nnd2s1 _46455_inst ( .DIN1(_46047), .DIN2(_46048), .Q(_45182) );
  nor2s1 _46456_inst ( .DIN1(_38864), .DIN2(_45924), .Q(_46048) );
  nnd2s1 _46457_inst ( .DIN1(_45986), .DIN2(_26565), .Q(_45924) );
  hi1s1 _46458_inst ( .DIN(_45615), .Q(_45986) );
  nor2s1 _46459_inst ( .DIN1(_45843), .DIN2(_45871), .Q(_46047) );
  nnd2s1 _46460_inst ( .DIN1(_45867), .DIN2(_26219), .Q(_45871) );
  nor2s1 _46461_inst ( .DIN1(_45175), .DIN2(_45157), .Q(_46046) );
  and2s1 _46462_inst ( .DIN1(_46049), .DIN2(_45915), .Q(_45157) );
  nor2s1 _46463_inst ( .DIN1(_45904), .DIN2(_45715), .Q(_45915) );
  nor2s1 _46464_inst ( .DIN1(_45656), .DIN2(_45835), .Q(_46049) );
  nnd2s1 _46465_inst ( .DIN1(_46006), .DIN2(_31888), .Q(_45835) );
  hi1s1 _46466_inst ( .DIN(_31459), .Q(_31888) );
  hi1s1 _46467_inst ( .DIN(_45414), .Q(_45175) );
  nnd2s1 _46468_inst ( .DIN1(_46050), .DIN2(_45856), .Q(_45414) );
  hi1s1 _46469_inst ( .DIN(_45649), .Q(_45856) );
  nor2s1 _46470_inst ( .DIN1(_38912), .DIN2(_45843), .Q(_46050) );
  nnd2s1 _46471_inst ( .DIN1(_46051), .DIN2(_26770), .Q(_46044) );
  and2s1 _46472_inst ( .DIN1(_45445), .DIN2(_45994), .Q(_46052) );
  nor2s1 _46473_inst ( .DIN1(_46054), .DIN2(_45998), .Q(_45994) );
  nnd2s1 _46474_inst ( .DIN1(_53500), .DIN2(_45956), .Q(_46054) );
  xnr2s1 _46475_inst ( .DIN1(_34289), .DIN2(_41072), .Q(_45956) );
  hi1s1 _46476_inst ( .DIN(_32330), .Q(_41072) );
  nnd2s1 _46477_inst ( .DIN1(_30163), .DIN2(_44077), .Q(_32330) );
  hi1s1 _46478_inst ( .DIN(_28521), .Q(_30163) );
  nnd2s1 _46479_inst ( .DIN1(_44658), .DIN2(_44079), .Q(_28521) );
  nor2s1 _46480_inst ( .DIN1(_26416), .DIN2(_53499), .Q(_34289) );
  nor2s1 _46481_inst ( .DIN1(_45458), .DIN2(_38865), .Q(_45445) );
  nnd2s1 _46482_inst ( .DIN1(_46055), .DIN2(_53502), .Q(_38865) );
  nor2s1 _46483_inst ( .DIN1(_53501), .DIN2(_53503), .Q(_46055) );
  nor2s1 _46484_inst ( .DIN1(_45256), .DIN2(_44822), .Q(_46051) );
  nor2s1 _46485_inst ( .DIN1(_45181), .DIN2(_26851), .Q(_44822) );
  nnd2s1 _46486_inst ( .DIN1(_46056), .DIN2(_46057), .Q(_45181) );
  nor2s1 _46487_inst ( .DIN1(_45904), .DIN2(_45802), .Q(_46057) );
  nor2s1 _46488_inst ( .DIN1(_45715), .DIN2(_45775), .Q(_46056) );
  and2s1 _46489_inst ( .DIN1(_46058), .DIN2(_45834), .Q(_45256) );
  and2s1 _46490_inst ( .DIN1(_46059), .DIN2(_26767), .Q(_45834) );
  nor2s1 _46491_inst ( .DIN1(_45904), .DIN2(_45458), .Q(_46059) );
  nor2s1 _46492_inst ( .DIN1(_45461), .DIN2(_45799), .Q(_46058) );
  nnd2s1 _46493_inst ( .DIN1(_45995), .DIN2(_46060), .Q(_45799) );
  hi1s1 _46494_inst ( .DIN(_45645), .Q(_45461) );
  nor2s1 _46495_inst ( .DIN1(_46061), .DIN2(_46062), .Q(_46042) );
  nnd2s1 _46496_inst ( .DIN1(_46063), .DIN2(_45233), .Q(_46062) );
  and2s1 _46497_inst ( .DIN1(_46064), .DIN2(_46065), .Q(_45233) );
  or2s1 _46498_inst ( .DIN1(_45169), .DIN2(_44957), .Q(_46065) );
  nnd2s1 _46499_inst ( .DIN1(_26805), .DIN2(_45224), .Q(_44957) );
  hi1s1 _46500_inst ( .DIN(_45168), .Q(_45224) );
  nnd2s1 _46501_inst ( .DIN1(_45865), .DIN2(_45867), .Q(_45168) );
  nor2s1 _46502_inst ( .DIN1(_31459), .DIN2(_38912), .Q(_45865) );
  nnd2s1 _46503_inst ( .DIN1(_46066), .DIN2(_26241), .Q(_31459) );
  hi1s1 _46504_inst ( .DIN(_44723), .Q(_44725) );
  nnd2s1 _46505_inst ( .DIN1(_46067), .DIN2(_45995), .Q(_45169) );
  hi1s1 _46506_inst ( .DIN(_45600), .Q(_45995) );
  nnd2s1 _46507_inst ( .DIN1(_53477), .DIN2(_53475), .Q(_45600) );
  nnd2s1 _46508_inst ( .DIN1(_45490), .DIN2(_26852), .Q(_46064) );
  hi1s1 _46509_inst ( .DIN(_45131), .Q(_45490) );
  nnd2s1 _46510_inst ( .DIN1(_45827), .DIN2(_45272), .Q(_45131) );
  nor2s1 _46511_inst ( .DIN1(_46068), .DIN2(_45842), .Q(_45827) );
  nor2s1 _46512_inst ( .DIN1(_45355), .DIN2(_45268), .Q(_46063) );
  nnd2s1 _46513_inst ( .DIN1(_45734), .DIN2(_46069), .Q(_45268) );
  nnd2s1 _46514_inst ( .DIN1(_44901), .DIN2(_26845), .Q(_46069) );
  hi1s1 _46515_inst ( .DIN(_45467), .Q(_44901) );
  nnd2s1 _46516_inst ( .DIN1(_46070), .DIN2(_45444), .Q(_45467) );
  and2s1 _46517_inst ( .DIN1(_45611), .DIN2(_45901), .Q(_45444) );
  hi1s1 _46518_inst ( .DIN(_37403), .Q(_45901) );
  nnd2s1 _46519_inst ( .DIN1(_46071), .DIN2(_53499), .Q(_37403) );
  nor2s1 _46520_inst ( .DIN1(_53479), .DIN2(_53500), .Q(_46071) );
  nor2s1 _46521_inst ( .DIN1(_45615), .DIN2(_45998), .Q(_45611) );
  nnd2s1 _46522_inst ( .DIN1(_45570), .DIN2(_45893), .Q(_45998) );
  hi1s1 _46523_inst ( .DIN(_45904), .Q(_45893) );
  nnd2s1 _46524_inst ( .DIN1(_53473), .DIN2(_53471), .Q(_45904) );
  hi1s1 _46525_inst ( .DIN(_45917), .Q(_45570) );
  nnd2s1 _46526_inst ( .DIN1(_53474), .DIN2(_26219), .Q(_45917) );
  nnd2s1 _46527_inst ( .DIN1(_26325), .DIN2(_26231), .Q(_45615) );
  nor2s1 _46528_inst ( .DIN1(_38528), .DIN2(_45601), .Q(_46070) );
  nnd2s1 _46529_inst ( .DIN1(_53476), .DIN2(_53472), .Q(_45601) );
  nnd2s1 _46530_inst ( .DIN1(_46072), .DIN2(_53501), .Q(_38528) );
  nor2s1 _46531_inst ( .DIN1(_53502), .DIN2(_26364), .Q(_46072) );
  nnd2s1 _46532_inst ( .DIN1(_45867), .DIN2(_46073), .Q(_45734) );
  nnd2s1 _46533_inst ( .DIN1(_45776), .DIN2(_46074), .Q(_46073) );
  nnd2s1 _46534_inst ( .DIN1(_46075), .DIN2(_45645), .Q(_46074) );
  nor2s1 _46535_inst ( .DIN1(_36898), .DIN2(_35291), .Q(_45645) );
  nor2s1 _46536_inst ( .DIN1(_44958), .DIN2(_26852), .Q(_46075) );
  hi1s1 _46537_inst ( .DIN(_45223), .Q(_44958) );
  nor2s1 _46538_inst ( .DIN1(_45830), .DIN2(_26231), .Q(_45223) );
  nnd2s1 _46539_inst ( .DIN1(_46060), .DIN2(_26325), .Q(_45830) );
  nnd2s1 _46540_inst ( .DIN1(_45272), .DIN2(_45655), .Q(_45776) );
  hi1s1 _46541_inst ( .DIN(_45683), .Q(_45655) );
  hi1s1 _46542_inst ( .DIN(_45460), .Q(_45272) );
  nnd2s1 _46543_inst ( .DIN1(_46060), .DIN2(_46053), .Q(_45460) );
  nor2s1 _46544_inst ( .DIN1(_26565), .DIN2(_26219), .Q(_46060) );
  hi1s1 _46545_inst ( .DIN(_45842), .Q(_45867) );
  nnd2s1 _46546_inst ( .DIN1(_45866), .DIN2(_45964), .Q(_45842) );
  nor2s1 _46547_inst ( .DIN1(_53471), .DIN2(_26558), .Q(_45866) );
  nor2s1 _46548_inst ( .DIN1(_44723), .DIN2(_44955), .Q(_45355) );
  nnd2s1 _46549_inst ( .DIN1(_46076), .DIN2(_46077), .Q(_44955) );
  nor2s1 _46550_inst ( .DIN1(_45458), .DIN2(_46068), .Q(_46077) );
  nnd2s1 _46551_inst ( .DIN1(_38344), .DIN2(_32681), .Q(_46068) );
  hi1s1 _46552_inst ( .DIN(_38912), .Q(_38344) );
  nnd2s1 _46553_inst ( .DIN1(_46078), .DIN2(_26364), .Q(_38912) );
  nnd2s1 _46554_inst ( .DIN1(_53472), .DIN2(_26233), .Q(_45458) );
  nor2s1 _46555_inst ( .DIN1(_45459), .DIN2(_45802), .Q(_46076) );
  nnd2s1 _46556_inst ( .DIN1(_46067), .DIN2(_46053), .Q(_45802) );
  nor2s1 _46557_inst ( .DIN1(_53474), .DIN2(_26219), .Q(_46067) );
  nnd2s1 _46558_inst ( .DIN1(_26558), .DIN2(_26222), .Q(_45459) );
  nnd2s1 _46559_inst ( .DIN1(______[28]), .DIN2(_39015), .Q(_44723) );
  nnd2s1 _46560_inst ( .DIN1(_46079), .DIN2(_46080), .Q(_46061) );
  nnd2s1 _46561_inst ( .DIN1(_44773), .DIN2(_44715), .Q(_46080) );
  nnd2s1 _46562_inst ( .DIN1(______[7]), .DIN2(______[28]), .Q(_44771) );
  nor2s1 _46563_inst ( .DIN1(_45649), .DIN2(_45775), .Q(_44773) );
  hi1s1 _46564_inst ( .DIN(_45870), .Q(_45775) );
  nor2s1 _46565_inst ( .DIN1(_36898), .DIN2(_45843), .Q(_45870) );
  nnd2s1 _46566_inst ( .DIN1(_46081), .DIN2(_53479), .Q(_45843) );
  and2s1 _46567_inst ( .DIN1(_26241), .DIN2(_53499), .Q(_46081) );
  nnd2s1 _46568_inst ( .DIN1(_46082), .DIN2(_53501), .Q(_36898) );
  nor2s1 _46569_inst ( .DIN1(_53502), .DIN2(_53503), .Q(_46082) );
  nnd2s1 _46570_inst ( .DIN1(_46083), .DIN2(_45788), .Q(_45649) );
  nor2s1 _46571_inst ( .DIN1(_46084), .DIN2(_45763), .Q(_45788) );
  nnd2s1 _46572_inst ( .DIN1(_26233), .DIN2(_53473), .Q(_46084) );
  nor2s1 _46573_inst ( .DIN1(_26219), .DIN2(_26325), .Q(_46083) );
  nor2s1 _46574_inst ( .DIN1(_45283), .DIN2(_44949), .Q(_46079) );
  hi1s1 _46575_inst ( .DIN(_44890), .Q(_44949) );
  nnd2s1 _46576_inst ( .DIN1(_46085), .DIN2(_45779), .Q(_44890) );
  hi1s1 _46577_inst ( .DIN(_45656), .Q(_45779) );
  nnd2s1 _46578_inst ( .DIN1(_46086), .DIN2(_46053), .Q(_45656) );
  hi1s1 _46579_inst ( .DIN(_45689), .Q(_46053) );
  nnd2s1 _46580_inst ( .DIN1(_53477), .DIN2(_26231), .Q(_45689) );
  nor2s1 _46581_inst ( .DIN1(_53474), .DIN2(_53478), .Q(_46086) );
  nor2s1 _46582_inst ( .DIN1(_45683), .DIN2(_45780), .Q(_46085) );
  nnd2s1 _46583_inst ( .DIN1(_45845), .DIN2(_45964), .Q(_45780) );
  hi1s1 _46584_inst ( .DIN(_45715), .Q(_45964) );
  nnd2s1 _46585_inst ( .DIN1(_26233), .DIN2(_26369), .Q(_45715) );
  nor2s1 _46586_inst ( .DIN1(_53473), .DIN2(_26222), .Q(_45845) );
  nnd2s1 _46587_inst ( .DIN1(_46006), .DIN2(_32681), .Q(_45683) );
  hi1s1 _46588_inst ( .DIN(_35291), .Q(_32681) );
  nnd2s1 _46589_inst ( .DIN1(_46066), .DIN2(_53500), .Q(_35291) );
  nor2s1 _46590_inst ( .DIN1(_53479), .DIN2(_53499), .Q(_46066) );
  hi1s1 _46591_inst ( .DIN(_38864), .Q(_46006) );
  nnd2s1 _46592_inst ( .DIN1(_46078), .DIN2(_53503), .Q(_38864) );
  nor2s1 _46593_inst ( .DIN1(_53501), .DIN2(_53502), .Q(_46078) );
  hi1s1 _46594_inst ( .DIN(_44914), .Q(_45283) );
  nnd2s1 _46595_inst ( .DIN1(_45969), .DIN2(_45933), .Q(_44914) );
  hi1s1 _46596_inst ( .DIN(_45691), .Q(_45933) );
  nnd2s1 _46597_inst ( .DIN1(_46087), .DIN2(_46088), .Q(_45691) );
  nor2s1 _46598_inst ( .DIN1(_53478), .DIN2(_53503), .Q(_46088) );
  nor2s1 _46599_inst ( .DIN1(_26416), .DIN2(_45764), .Q(_46087) );
  nnd2s1 _46600_inst ( .DIN1(_46089), .DIN2(_45948), .Q(_45764) );
  and2s1 _46601_inst ( .DIN1(_46090), .DIN2(_28502), .Q(_45948) );
  and2s1 _46602_inst ( .DIN1(_53499), .DIN2(_53501), .Q(_28502) );
  nor2s1 _46603_inst ( .DIN1(_26241), .DIN2(_26467), .Q(_46090) );
  nor2s1 _46604_inst ( .DIN1(_53473), .DIN2(_26233), .Q(_46089) );
  nor2s1 _46605_inst ( .DIN1(_26325), .DIN2(_45763), .Q(_45969) );
  nnd2s1 _46606_inst ( .DIN1(_46091), .DIN2(_46092), .Q(_45763) );
  hi1s1 _46607_inst ( .DIN(_45690), .Q(_46092) );
  nnd2s1 _46608_inst ( .DIN1(_53472), .DIN2(_53471), .Q(_45690) );
  nor2s1 _46609_inst ( .DIN1(_53474), .DIN2(_26231), .Q(_46091) );
  hi1s1 _46610_inst ( .DIN(_32702), .Q(_14172) );
  xnr2s1 _46611_inst ( .DIN1(_46093), .DIN2(_32799), .Q(_32702) );
  nnd2s1 _46612_inst ( .DIN1(_46094), .DIN2(_46095), .Q(_32799) );
  nnd2s1 _46613_inst ( .DIN1(_53507), .DIN2(_46096), .Q(_46095) );
  or2s1 _46614_inst ( .DIN1(_26723), .DIN2(_32779), .Q(_46096) );
  nnd2s1 _46615_inst ( .DIN1(_32779), .DIN2(_26723), .Q(_46094) );
  nnd2s1 _46616_inst ( .DIN1(_46097), .DIN2(_46098), .Q(_32779) );
  nnd2s1 _46617_inst ( .DIN1(_46099), .DIN2(_26542), .Q(_46098) );
  nnd2s1 _46618_inst ( .DIN1(_26551), .DIN2(_32778), .Q(_46099) );
  or2s1 _46619_inst ( .DIN1(_26551), .DIN2(_32778), .Q(_46097) );
  nnd2s1 _46620_inst ( .DIN1(_46100), .DIN2(_46101), .Q(_32778) );
  nnd2s1 _46621_inst ( .DIN1(_53134), .DIN2(_46102), .Q(_46101) );
  or2s1 _46622_inst ( .DIN1(_32775), .DIN2(_53506), .Q(_46102) );
  nnd2s1 _46623_inst ( .DIN1(_53506), .DIN2(_32775), .Q(_46100) );
  nnd2s1 _46624_inst ( .DIN1(_46103), .DIN2(_46104), .Q(_32775) );
  nnd2s1 _46625_inst ( .DIN1(_52844), .DIN2(_46105), .Q(_46104) );
  nnd2s1 _46626_inst ( .DIN1(_53511), .DIN2(_32772), .Q(_46105) );
  or2s1 _46627_inst ( .DIN1(_32772), .DIN2(_53511), .Q(_46103) );
  or2s1 _46628_inst ( .DIN1(_26562), .DIN2(_53135), .Q(_32772) );
  xor2s1 _46629_inst ( .DIN1(_26559), .DIN2(_53513), .Q(_46093) );
  nnd2s1 _46630_inst ( .DIN1(_46106), .DIN2(_46107), .Q(____3___________[9])
         );
  nor2s1 _46631_inst ( .DIN1(_46108), .DIN2(_46109), .Q(_46107) );
  nnd2s1 _46632_inst ( .DIN1(_46110), .DIN2(_46111), .Q(_46109) );
  nnd2s1 _46633_inst ( .DIN1(_26840), .DIN2(_46113), .Q(_46111) );
  nnd2s1 _46634_inst ( .DIN1(_46114), .DIN2(_46115), .Q(_46113) );
  nor2s1 _46635_inst ( .DIN1(_46116), .DIN2(_46117), .Q(_46114) );
  nnd2s1 _46636_inst ( .DIN1(_46118), .DIN2(_46119), .Q(_46110) );
  nnd2s1 _46637_inst ( .DIN1(_46120), .DIN2(_46121), .Q(_46119) );
  nor2s1 _46638_inst ( .DIN1(_46122), .DIN2(_46123), .Q(_46120) );
  nnd2s1 _46639_inst ( .DIN1(_46124), .DIN2(_46125), .Q(_46108) );
  nnd2s1 _46640_inst ( .DIN1(_46126), .DIN2(_46127), .Q(_46124) );
  nnd2s1 _46641_inst ( .DIN1(_46128), .DIN2(_46129), .Q(_46126) );
  nor2s1 _46642_inst ( .DIN1(_46130), .DIN2(_46131), .Q(_46106) );
  nnd2s1 _46643_inst ( .DIN1(_46132), .DIN2(_46133), .Q(_46131) );
  hi1s1 _46644_inst ( .DIN(_46134), .Q(_46133) );
  nnd2s1 _46645_inst ( .DIN1(_46135), .DIN2(_46136), .Q(_46130) );
  hi1s1 _46646_inst ( .DIN(_46137), .Q(_46135) );
  nnd2s1 _46647_inst ( .DIN1(_46138), .DIN2(_46139), .Q(____3___________[8])
         );
  nor2s1 _46648_inst ( .DIN1(_46140), .DIN2(_46141), .Q(_46139) );
  nnd2s1 _46649_inst ( .DIN1(_46142), .DIN2(_46143), .Q(_46141) );
  nnd2s1 _46650_inst ( .DIN1(_46144), .DIN2(_46145), .Q(_46143) );
  nnd2s1 _46651_inst ( .DIN1(_26840), .DIN2(_46146), .Q(_46142) );
  nnd2s1 _46652_inst ( .DIN1(_46147), .DIN2(_46148), .Q(_46146) );
  nor2s1 _46653_inst ( .DIN1(_46149), .DIN2(_46150), .Q(_46148) );
  nnd2s1 _46654_inst ( .DIN1(_46151), .DIN2(_46152), .Q(_46150) );
  nnd2s1 _46655_inst ( .DIN1(_46153), .DIN2(_46154), .Q(_46149) );
  nor2s1 _46656_inst ( .DIN1(_46155), .DIN2(_46156), .Q(_46147) );
  nnd2s1 _46657_inst ( .DIN1(_46157), .DIN2(_46158), .Q(_46156) );
  nnd2s1 _46658_inst ( .DIN1(_46159), .DIN2(_46160), .Q(_46140) );
  nnd2s1 _46659_inst ( .DIN1(_46227), .DIN2(_46161), .Q(_46159) );
  nnd2s1 _46660_inst ( .DIN1(_46162), .DIN2(_46163), .Q(_46161) );
  nor2s1 _46661_inst ( .DIN1(_46164), .DIN2(_46165), .Q(_46162) );
  nor2s1 _46662_inst ( .DIN1(_46166), .DIN2(_46167), .Q(_46138) );
  or2s1 _46663_inst ( .DIN1(_46168), .DIN2(_46169), .Q(_46167) );
  nnd2s1 _46664_inst ( .DIN1(_46170), .DIN2(_46171), .Q(_46166) );
  hi1s1 _46665_inst ( .DIN(_46172), .Q(_46171) );
  nnd2s1 _46666_inst ( .DIN1(_46173), .DIN2(_46174), .Q(____3___________[7])
         );
  nor2s1 _46667_inst ( .DIN1(_46175), .DIN2(_46176), .Q(_46174) );
  nnd2s1 _46668_inst ( .DIN1(_46177), .DIN2(_46178), .Q(_46176) );
  nnd2s1 _46669_inst ( .DIN1(_46118), .DIN2(_46179), .Q(_46178) );
  nnd2s1 _46670_inst ( .DIN1(_46180), .DIN2(_46181), .Q(_46179) );
  nor2s1 _46671_inst ( .DIN1(_46116), .DIN2(_46182), .Q(_46181) );
  nnd2s1 _46672_inst ( .DIN1(_46183), .DIN2(_46184), .Q(_46182) );
  hi1s1 _46673_inst ( .DIN(_46185), .Q(_46116) );
  nor2s1 _46674_inst ( .DIN1(_46186), .DIN2(_46187), .Q(_46180) );
  nnd2s1 _46675_inst ( .DIN1(_46188), .DIN2(_46189), .Q(_46187) );
  hi1s1 _46676_inst ( .DIN(_46190), .Q(_46188) );
  hi1s1 _46677_inst ( .DIN(_46191), .Q(_46177) );
  nnd2s1 _46678_inst ( .DIN1(_46192), .DIN2(_46193), .Q(_46175) );
  nnd2s1 _46679_inst ( .DIN1(_26840), .DIN2(_46194), .Q(_46192) );
  nnd2s1 _46680_inst ( .DIN1(_46195), .DIN2(_46196), .Q(_46194) );
  nor2s1 _46681_inst ( .DIN1(_46197), .DIN2(_46198), .Q(_46195) );
  nor2s1 _46682_inst ( .DIN1(_46199), .DIN2(_46200), .Q(_46173) );
  nnd2s1 _46683_inst ( .DIN1(_46201), .DIN2(_46202), .Q(_46200) );
  nnd2s1 _46684_inst ( .DIN1(_46203), .DIN2(_46204), .Q(____3___________[6])
         );
  nor2s1 _46685_inst ( .DIN1(_46205), .DIN2(_46206), .Q(_46204) );
  nnd2s1 _46686_inst ( .DIN1(_46207), .DIN2(_46208), .Q(_46206) );
  nnd2s1 _46687_inst ( .DIN1(_46209), .DIN2(_45194), .Q(_46208) );
  nnd2s1 _46688_inst ( .DIN1(_46210), .DIN2(_46127), .Q(_46207) );
  nnd2s1 _46689_inst ( .DIN1(_46211), .DIN2(_46212), .Q(_46205) );
  nnd2s1 _46690_inst ( .DIN1(_46213), .DIN2(_46145), .Q(_46212) );
  nnd2s1 _46691_inst ( .DIN1(_46214), .DIN2(_46215), .Q(_46213) );
  nor2s1 _46692_inst ( .DIN1(_46216), .DIN2(_46217), .Q(_46215) );
  nnd2s1 _46693_inst ( .DIN1(_46218), .DIN2(_46219), .Q(_46217) );
  nor2s1 _46694_inst ( .DIN1(_46220), .DIN2(_46221), .Q(_46214) );
  nnd2s1 _46695_inst ( .DIN1(_46222), .DIN2(_46223), .Q(_46221) );
  nor2s1 _46696_inst ( .DIN1(_46224), .DIN2(_46225), .Q(_46211) );
  nor2s1 _46697_inst ( .DIN1(_46226), .DIN2(_26782), .Q(_46225) );
  nor2s1 _46698_inst ( .DIN1(_46228), .DIN2(_46229), .Q(_46226) );
  nnd2s1 _46699_inst ( .DIN1(_46230), .DIN2(_46231), .Q(_46229) );
  hi1s1 _46700_inst ( .DIN(_46232), .Q(_46224) );
  nor2s1 _46701_inst ( .DIN1(_46233), .DIN2(_46234), .Q(_46203) );
  nnd2s1 _46702_inst ( .DIN1(_46235), .DIN2(_46236), .Q(_46234) );
  nnd2s1 _46703_inst ( .DIN1(_46237), .DIN2(_46238), .Q(_46233) );
  nor2s1 _46704_inst ( .DIN1(_46239), .DIN2(_46169), .Q(_46237) );
  nnd2s1 _46705_inst ( .DIN1(_46240), .DIN2(_46241), .Q(_46169) );
  nor2s1 _46706_inst ( .DIN1(_46242), .DIN2(_46243), .Q(_46241) );
  nnd2s1 _46707_inst ( .DIN1(_46244), .DIN2(_46245), .Q(_46243) );
  nnd2s1 _46708_inst ( .DIN1(_26840), .DIN2(_46246), .Q(_46244) );
  nnd2s1 _46709_inst ( .DIN1(_46247), .DIN2(_46248), .Q(_46246) );
  nnd2s1 _46710_inst ( .DIN1(_46249), .DIN2(_46250), .Q(_46242) );
  nor2s1 _46711_inst ( .DIN1(_46251), .DIN2(_46252), .Q(_46240) );
  nnd2s1 _46712_inst ( .DIN1(_46202), .DIN2(_46253), .Q(_46252) );
  hi1s1 _46713_inst ( .DIN(_46254), .Q(_46253) );
  nor2s1 _46714_inst ( .DIN1(_46255), .DIN2(_46256), .Q(_46202) );
  nor2s1 _46715_inst ( .DIN1(_46257), .DIN2(_46258), .Q(_46256) );
  nnd2s1 _46716_inst ( .DIN1(_46259), .DIN2(_46260), .Q(_46251) );
  nnd2s1 _46717_inst ( .DIN1(_46227), .DIN2(_46261), .Q(_46260) );
  nnd2s1 _46718_inst ( .DIN1(_46262), .DIN2(_46263), .Q(_46261) );
  nnd2s1 _46719_inst ( .DIN1(_46264), .DIN2(_46265), .Q(____3___________[5])
         );
  nor2s1 _46720_inst ( .DIN1(_46266), .DIN2(_46267), .Q(_46265) );
  nnd2s1 _46721_inst ( .DIN1(_46268), .DIN2(_46269), .Q(_46267) );
  nnd2s1 _46722_inst ( .DIN1(_46118), .DIN2(_46270), .Q(_46269) );
  nnd2s1 _46723_inst ( .DIN1(_46271), .DIN2(_46272), .Q(_46270) );
  nnd2s1 _46724_inst ( .DIN1(_26840), .DIN2(_46273), .Q(_46268) );
  nnd2s1 _46725_inst ( .DIN1(_46274), .DIN2(_46275), .Q(_46273) );
  hi1s1 _46726_inst ( .DIN(_46220), .Q(_46275) );
  nnd2s1 _46727_inst ( .DIN1(_46276), .DIN2(_46151), .Q(_46220) );
  nor2s1 _46728_inst ( .DIN1(_46277), .DIN2(_46228), .Q(_46274) );
  nnd2s1 _46729_inst ( .DIN1(_46278), .DIN2(_46279), .Q(_46228) );
  hi1s1 _46730_inst ( .DIN(_46280), .Q(_46277) );
  nnd2s1 _46731_inst ( .DIN1(_46281), .DIN2(_46282), .Q(_46266) );
  nor2s1 _46732_inst ( .DIN1(_46283), .DIN2(_46284), .Q(_46264) );
  or2s1 _46733_inst ( .DIN1(_46285), .DIN2(_46286), .Q(_46284) );
  nnd2s1 _46734_inst ( .DIN1(_46287), .DIN2(_46288), .Q(_46283) );
  nnd2s1 _46735_inst ( .DIN1(_46289), .DIN2(_46145), .Q(_46288) );
  nnd2s1 _46736_inst ( .DIN1(_46290), .DIN2(_46291), .Q(____3___________[4])
         );
  nor2s1 _46737_inst ( .DIN1(_46292), .DIN2(_46293), .Q(_46291) );
  nnd2s1 _46738_inst ( .DIN1(_46294), .DIN2(_46295), .Q(_46293) );
  nnd2s1 _46739_inst ( .DIN1(_46296), .DIN2(_46127), .Q(_46295) );
  nnd2s1 _46740_inst ( .DIN1(_46297), .DIN2(_46298), .Q(_46296) );
  and2s1 _46741_inst ( .DIN1(_46262), .DIN2(_46299), .Q(_46298) );
  nor2s1 _46742_inst ( .DIN1(_46300), .DIN2(_46301), .Q(_46297) );
  nor2s1 _46743_inst ( .DIN1(_46302), .DIN2(_46303), .Q(_46294) );
  nor2s1 _46744_inst ( .DIN1(_46304), .DIN2(_46305), .Q(_46303) );
  nor2s1 _46745_inst ( .DIN1(_46306), .DIN2(_46307), .Q(_46304) );
  nnd2s1 _46746_inst ( .DIN1(_46271), .DIN2(_46219), .Q(_46307) );
  nor2s1 _46747_inst ( .DIN1(_46308), .DIN2(_26782), .Q(_46302) );
  and2s1 _46748_inst ( .DIN1(_46158), .DIN2(_46309), .Q(_46308) );
  nnd2s1 _46749_inst ( .DIN1(_46310), .DIN2(_46282), .Q(_46292) );
  nnd2s1 _46750_inst ( .DIN1(_46311), .DIN2(_46312), .Q(_46282) );
  nor2s1 _46751_inst ( .DIN1(_26782), .DIN2(_46313), .Q(_46311) );
  nor2s1 _46752_inst ( .DIN1(_46314), .DIN2(_46315), .Q(_46310) );
  nor2s1 _46753_inst ( .DIN1(_46316), .DIN2(_46317), .Q(_46290) );
  nnd2s1 _46754_inst ( .DIN1(_46318), .DIN2(_46319), .Q(_46317) );
  hi1s1 _46755_inst ( .DIN(_46320), .Q(_46319) );
  nor2s1 _46756_inst ( .DIN1(_46321), .DIN2(_46322), .Q(_46318) );
  nnd2s1 _46757_inst ( .DIN1(_46323), .DIN2(_46235), .Q(_46316) );
  and2s1 _46758_inst ( .DIN1(_46324), .DIN2(_46325), .Q(_46235) );
  nor2s1 _46759_inst ( .DIN1(_46326), .DIN2(_46327), .Q(_46325) );
  nnd2s1 _46760_inst ( .DIN1(_46328), .DIN2(_46281), .Q(_46327) );
  nnd2s1 _46761_inst ( .DIN1(_46329), .DIN2(_46145), .Q(_46281) );
  nnd2s1 _46762_inst ( .DIN1(_26840), .DIN2(_46330), .Q(_46328) );
  nnd2s1 _46763_inst ( .DIN1(_46331), .DIN2(_46332), .Q(_46330) );
  nor2s1 _46764_inst ( .DIN1(_26782), .DIN2(_46333), .Q(_46326) );
  nor2s1 _46765_inst ( .DIN1(_46334), .DIN2(_46335), .Q(_46324) );
  nor2s1 _46766_inst ( .DIN1(_46336), .DIN2(_46254), .Q(_46323) );
  nnd2s1 _46767_inst ( .DIN1(_46337), .DIN2(_46338), .Q(_46254) );
  nnd2s1 _46768_inst ( .DIN1(_46227), .DIN2(_46339), .Q(_46338) );
  nnd2s1 _46769_inst ( .DIN1(_46280), .DIN2(_46340), .Q(_46339) );
  nnd2s1 _46770_inst ( .DIN1(_46341), .DIN2(_46342), .Q(_46340) );
  nnd2s1 _46771_inst ( .DIN1(_26840), .DIN2(_46343), .Q(_46337) );
  nnd2s1 _46772_inst ( .DIN1(_46344), .DIN2(_46345), .Q(_46343) );
  nor2s1 _46773_inst ( .DIN1(_46346), .DIN2(_46347), .Q(_46344) );
  nnd2s1 _46774_inst ( .DIN1(_46348), .DIN2(_46349), .Q(____3___________[3])
         );
  nor2s1 _46775_inst ( .DIN1(_46350), .DIN2(_46351), .Q(_46349) );
  nnd2s1 _46776_inst ( .DIN1(_46352), .DIN2(_46353), .Q(_46351) );
  nor2s1 _46777_inst ( .DIN1(_46354), .DIN2(_46355), .Q(_46352) );
  nor2s1 _46778_inst ( .DIN1(_46356), .DIN2(_26782), .Q(_46355) );
  nor2s1 _46779_inst ( .DIN1(_46357), .DIN2(_46358), .Q(_46356) );
  nnd2s1 _46780_inst ( .DIN1(_46359), .DIN2(_46360), .Q(_46358) );
  hi1s1 _46781_inst ( .DIN(_46300), .Q(_46359) );
  nnd2s1 _46782_inst ( .DIN1(_46279), .DIN2(_46154), .Q(_46300) );
  nnd2s1 _46783_inst ( .DIN1(_46361), .DIN2(_46362), .Q(_46357) );
  nor2s1 _46784_inst ( .DIN1(_46363), .DIN2(_46364), .Q(_46354) );
  nor2s1 _46785_inst ( .DIN1(_46365), .DIN2(_46366), .Q(_46364) );
  nnd2s1 _46786_inst ( .DIN1(_46280), .DIN2(_46367), .Q(_46366) );
  nor2s1 _46787_inst ( .DIN1(_46368), .DIN2(_45553), .Q(_46365) );
  nnd2s1 _46788_inst ( .DIN1(_46369), .DIN2(_46370), .Q(_46350) );
  nnd2s1 _46789_inst ( .DIN1(_46371), .DIN2(_46127), .Q(_46370) );
  nnd2s1 _46790_inst ( .DIN1(_46257), .DIN2(_46372), .Q(_46371) );
  nor2s1 _46791_inst ( .DIN1(_46373), .DIN2(_46374), .Q(_46369) );
  nor2s1 _46792_inst ( .DIN1(_45205), .DIN2(_46375), .Q(_46374) );
  nnd2s1 _46793_inst ( .DIN1(_46376), .DIN2(_26840), .Q(_46375) );
  hi1s1 _46794_inst ( .DIN(_46377), .Q(_46373) );
  nor2s1 _46795_inst ( .DIN1(_46378), .DIN2(_46379), .Q(_46348) );
  nnd2s1 _46796_inst ( .DIN1(_46380), .DIN2(_46381), .Q(_46379) );
  nor2s1 _46797_inst ( .DIN1(_46286), .DIN2(_46320), .Q(_46380) );
  nnd2s1 _46798_inst ( .DIN1(_46382), .DIN2(_46383), .Q(_46320) );
  nor2s1 _46799_inst ( .DIN1(_46384), .DIN2(_46385), .Q(_46383) );
  nnd2s1 _46800_inst ( .DIN1(_46386), .DIN2(_46387), .Q(_46385) );
  nnd2s1 _46801_inst ( .DIN1(_46388), .DIN2(_46127), .Q(_46387) );
  nnd2s1 _46802_inst ( .DIN1(_46389), .DIN2(_46145), .Q(_46386) );
  nnd2s1 _46803_inst ( .DIN1(_46390), .DIN2(_46391), .Q(_46384) );
  nnd2s1 _46804_inst ( .DIN1(_46209), .DIN2(_45197), .Q(_46391) );
  nor2s1 _46805_inst ( .DIN1(_46392), .DIN2(_46255), .Q(_46390) );
  nor2s1 _46806_inst ( .DIN1(_46393), .DIN2(_46394), .Q(_46382) );
  nnd2s1 _46807_inst ( .DIN1(_46395), .DIN2(_46396), .Q(_46394) );
  hi1s1 _46808_inst ( .DIN(_46397), .Q(_46396) );
  nnd2s1 _46809_inst ( .DIN1(_46398), .DIN2(_46399), .Q(_46393) );
  nnd2s1 _46810_inst ( .DIN1(_46400), .DIN2(_46118), .Q(_46399) );
  nnd2s1 _46811_inst ( .DIN1(_46401), .DIN2(_46402), .Q(_46286) );
  nor2s1 _46812_inst ( .DIN1(_46403), .DIN2(_46404), .Q(_46402) );
  nor2s1 _46813_inst ( .DIN1(_46363), .DIN2(_46405), .Q(_46404) );
  nor2s1 _46814_inst ( .DIN1(_46216), .DIN2(_46347), .Q(_46405) );
  hi1s1 _46815_inst ( .DIN(_46406), .Q(_46347) );
  nor2s1 _46816_inst ( .DIN1(_46407), .DIN2(_46305), .Q(_46403) );
  nor2s1 _46817_inst ( .DIN1(_46408), .DIN2(_46409), .Q(_46407) );
  or2s1 _46818_inst ( .DIN1(_46165), .DIN2(_46410), .Q(_46409) );
  hi1s1 _46819_inst ( .DIN(_46183), .Q(_46165) );
  hi1s1 _46820_inst ( .DIN(_46222), .Q(_46408) );
  nor2s1 _46821_inst ( .DIN1(_46411), .DIN2(_46322), .Q(_46401) );
  nnd2s1 _46822_inst ( .DIN1(_46412), .DIN2(_46413), .Q(_46322) );
  nnd2s1 _46823_inst ( .DIN1(_46118), .DIN2(_46414), .Q(_46413) );
  nnd2s1 _46824_inst ( .DIN1(_46415), .DIN2(_46416), .Q(_46414) );
  and2s1 _46825_inst ( .DIN1(_46417), .DIN2(_46223), .Q(_46415) );
  nor2s1 _46826_inst ( .DIN1(_46418), .DIN2(_46419), .Q(_46412) );
  nor2s1 _46827_inst ( .DIN1(_26839), .DIN2(_46420), .Q(_46419) );
  hi1s1 _46828_inst ( .DIN(_46245), .Q(_46418) );
  nnd2s1 _46829_inst ( .DIN1(_46227), .DIN2(_46421), .Q(_46245) );
  nnd2s1 _46830_inst ( .DIN1(_46422), .DIN2(_46423), .Q(_46421) );
  nor2s1 _46831_inst ( .DIN1(_46424), .DIN2(_26782), .Q(_46411) );
  nor2s1 _46832_inst ( .DIN1(_46425), .DIN2(_46426), .Q(_46424) );
  nnd2s1 _46833_inst ( .DIN1(_46427), .DIN2(_46428), .Q(_46378) );
  hi1s1 _46834_inst ( .DIN(_46429), .Q(_46428) );
  nor2s1 _46835_inst ( .DIN1(_46134), .DIN2(_46172), .Q(_46427) );
  nnd2s1 _46836_inst ( .DIN1(_46430), .DIN2(_46431), .Q(_46172) );
  nnd2s1 _46837_inst ( .DIN1(_46432), .DIN2(_46118), .Q(_46431) );
  nnd2s1 _46838_inst ( .DIN1(_46433), .DIN2(_46434), .Q(_46134) );
  nor2s1 _46839_inst ( .DIN1(_46435), .DIN2(_46436), .Q(_46434) );
  nnd2s1 _46840_inst ( .DIN1(_46437), .DIN2(_46438), .Q(_46436) );
  nnd2s1 _46841_inst ( .DIN1(_46439), .DIN2(_46440), .Q(_46437) );
  nor2s1 _46842_inst ( .DIN1(_26782), .DIN2(_39517), .Q(_46439) );
  hi1s1 _46843_inst ( .DIN(_46441), .Q(_39517) );
  nor2s1 _46844_inst ( .DIN1(_46363), .DIN2(_46442), .Q(_46435) );
  nor2s1 _46845_inst ( .DIN1(_46289), .DIN2(_46443), .Q(_46442) );
  nor2s1 _46846_inst ( .DIN1(_46444), .DIN2(_46445), .Q(_46433) );
  nnd2s1 _46847_inst ( .DIN1(_46446), .DIN2(_46447), .Q(_46445) );
  nnd2s1 _46848_inst ( .DIN1(_46164), .DIN2(_46127), .Q(_46447) );
  hi1s1 _46849_inst ( .DIN(_46448), .Q(_46164) );
  nnd2s1 _46850_inst ( .DIN1(_46449), .DIN2(_26840), .Q(_46446) );
  nnd2s1 _46851_inst ( .DIN1(_46450), .DIN2(_46451), .Q(____3___________[2])
         );
  nor2s1 _46852_inst ( .DIN1(_46452), .DIN2(_46453), .Q(_46451) );
  nnd2s1 _46853_inst ( .DIN1(_46454), .DIN2(_46455), .Q(_46453) );
  nnd2s1 _46854_inst ( .DIN1(_46118), .DIN2(_46456), .Q(_46455) );
  nnd2s1 _46855_inst ( .DIN1(_46457), .DIN2(_46458), .Q(_46456) );
  nor2s1 _46856_inst ( .DIN1(_46459), .DIN2(_46449), .Q(_46457) );
  nnd2s1 _46857_inst ( .DIN1(_46443), .DIN2(_46145), .Q(_46454) );
  nnd2s1 _46858_inst ( .DIN1(_46460), .DIN2(_46377), .Q(_46452) );
  nnd2s1 _46859_inst ( .DIN1(_26840), .DIN2(_46461), .Q(_46377) );
  nnd2s1 _46860_inst ( .DIN1(_46309), .DIN2(_46462), .Q(_46461) );
  nnd2s1 _46861_inst ( .DIN1(_26840), .DIN2(_46463), .Q(_46460) );
  nnd2s1 _46862_inst ( .DIN1(_46464), .DIN2(_46465), .Q(_46463) );
  hi1s1 _46863_inst ( .DIN(_46186), .Q(_46465) );
  nnd2s1 _46864_inst ( .DIN1(_46466), .DIN2(_46467), .Q(_46186) );
  nor2s1 _46865_inst ( .DIN1(_46432), .DIN2(_46468), .Q(_46467) );
  nnd2s1 _46866_inst ( .DIN1(_46280), .DIN2(_46406), .Q(_46468) );
  hi1s1 _46867_inst ( .DIN(_46469), .Q(_46432) );
  nor2s1 _46868_inst ( .DIN1(_46470), .DIN2(_46471), .Q(_46466) );
  hi1s1 _46869_inst ( .DIN(_46115), .Q(_46471) );
  nor2s1 _46870_inst ( .DIN1(_46472), .DIN2(_46473), .Q(_46464) );
  nor2s1 _46871_inst ( .DIN1(_46474), .DIN2(_46475), .Q(_46450) );
  nnd2s1 _46872_inst ( .DIN1(_46476), .DIN2(_46395), .Q(_46475) );
  and2s1 _46873_inst ( .DIN1(_46477), .DIN2(_46478), .Q(_46395) );
  nor2s1 _46874_inst ( .DIN1(_46479), .DIN2(_46480), .Q(_46478) );
  nnd2s1 _46875_inst ( .DIN1(_46481), .DIN2(_46160), .Q(_46480) );
  nor2s1 _46876_inst ( .DIN1(_46482), .DIN2(_46305), .Q(_46479) );
  nor2s1 _46877_inst ( .DIN1(_46483), .DIN2(_46484), .Q(_46482) );
  nnd2s1 _46878_inst ( .DIN1(_46361), .DIN2(_46485), .Q(_46484) );
  hi1s1 _46879_inst ( .DIN(_46276), .Q(_46483) );
  nor2s1 _46880_inst ( .DIN1(_46486), .DIN2(_46487), .Q(_46477) );
  nor2s1 _46881_inst ( .DIN1(_26782), .DIN2(_46248), .Q(_46486) );
  nnd2s1 _46882_inst ( .DIN1(_46236), .DIN2(_46488), .Q(_46474) );
  hi1s1 _46883_inst ( .DIN(_46199), .Q(_46488) );
  nnd2s1 _46884_inst ( .DIN1(_46489), .DIN2(_46490), .Q(_46199) );
  nor2s1 _46885_inst ( .DIN1(_46491), .DIN2(_46492), .Q(_46490) );
  nnd2s1 _46886_inst ( .DIN1(_46493), .DIN2(_46494), .Q(_46492) );
  nnd2s1 _46887_inst ( .DIN1(_46495), .DIN2(_46145), .Q(_46494) );
  nnd2s1 _46888_inst ( .DIN1(_26840), .DIN2(_46496), .Q(_46493) );
  nnd2s1 _46889_inst ( .DIN1(_46497), .DIN2(_46498), .Q(_46496) );
  nor2s1 _46890_inst ( .DIN1(_46425), .DIN2(_46289), .Q(_46497) );
  hi1s1 _46891_inst ( .DIN(_46499), .Q(_46425) );
  nnd2s1 _46892_inst ( .DIN1(_46500), .DIN2(_46501), .Q(_46491) );
  nor2s1 _46893_inst ( .DIN1(_46429), .DIN2(_46502), .Q(_46489) );
  nnd2s1 _46894_inst ( .DIN1(_46430), .DIN2(_46503), .Q(_46502) );
  nnd2s1 _46895_inst ( .DIN1(_46227), .DIN2(_46504), .Q(_46503) );
  nnd2s1 _46896_inst ( .DIN1(_46505), .DIN2(_46158), .Q(_46504) );
  nor2s1 _46897_inst ( .DIN1(_46506), .DIN2(_46122), .Q(_46505) );
  hi1s1 _46898_inst ( .DIN(_46334), .Q(_46430) );
  nnd2s1 _46899_inst ( .DIN1(_46507), .DIN2(_46508), .Q(_46429) );
  nnd2s1 _46900_inst ( .DIN1(_46118), .DIN2(_46509), .Q(_46508) );
  nor2s1 _46901_inst ( .DIN1(_46510), .DIN2(_46511), .Q(_46507) );
  nor2s1 _46902_inst ( .DIN1(_26839), .DIN2(_46512), .Q(_46511) );
  and2s1 _46903_inst ( .DIN1(_46513), .DIN2(_46514), .Q(_46236) );
  nor2s1 _46904_inst ( .DIN1(_46515), .DIN2(_46516), .Q(_46514) );
  nnd2s1 _46905_inst ( .DIN1(_46517), .DIN2(_46518), .Q(_46516) );
  nnd2s1 _46906_inst ( .DIN1(_26840), .DIN2(_46519), .Q(_46518) );
  nnd2s1 _46907_inst ( .DIN1(_46520), .DIN2(_46521), .Q(_46519) );
  and2s1 _46908_inst ( .DIN1(_46230), .DIN2(_46183), .Q(_46520) );
  nnd2s1 _46909_inst ( .DIN1(_46227), .DIN2(_46522), .Q(_46517) );
  nnd2s1 _46910_inst ( .DIN1(_46523), .DIN2(_46416), .Q(_46522) );
  and2s1 _46911_inst ( .DIN1(_46524), .DIN2(_46184), .Q(_46416) );
  nor2s1 _46912_inst ( .DIN1(_46525), .DIN2(_46526), .Q(_46523) );
  nnd2s1 _46913_inst ( .DIN1(_46125), .DIN2(_46438), .Q(_46515) );
  or2s1 _46914_inst ( .DIN1(_46527), .DIN2(_26782), .Q(_46438) );
  nnd2s1 _46915_inst ( .DIN1(_46528), .DIN2(_46529), .Q(_46125) );
  nor2s1 _46916_inst ( .DIN1(_45551), .DIN2(_26782), .Q(_46528) );
  nor2s1 _46917_inst ( .DIN1(_46530), .DIN2(_46531), .Q(_46513) );
  nnd2s1 _46918_inst ( .DIN1(_46532), .DIN2(_46533), .Q(_46531) );
  nnd2s1 _46919_inst ( .DIN1(_46534), .DIN2(_46127), .Q(_46533) );
  or2s1 _46920_inst ( .DIN1(_46362), .DIN2(_46363), .Q(_46532) );
  nnd2s1 _46921_inst ( .DIN1(_46535), .DIN2(_46536), .Q(____3___________[1])
         );
  nor2s1 _46922_inst ( .DIN1(_46537), .DIN2(_46538), .Q(_46536) );
  nnd2s1 _46923_inst ( .DIN1(_46539), .DIN2(_46540), .Q(_46538) );
  nnd2s1 _46924_inst ( .DIN1(_46118), .DIN2(_46541), .Q(_46539) );
  nnd2s1 _46925_inst ( .DIN1(_46542), .DIN2(_46543), .Q(_46541) );
  hi1s1 _46926_inst ( .DIN(_46144), .Q(_46543) );
  and2s1 _46927_inst ( .DIN1(_46362), .DIN2(_46544), .Q(_46542) );
  nnd2s1 _46928_inst ( .DIN1(_46232), .DIN2(_46160), .Q(_46537) );
  nnd2s1 _46929_inst ( .DIN1(_46545), .DIN2(_46546), .Q(_46160) );
  nor2s1 _46930_inst ( .DIN1(_26249), .DIN2(_46305), .Q(_46546) );
  nor2s1 _46931_inst ( .DIN1(_29221), .DIN2(_46547), .Q(_46545) );
  nnd2s1 _46932_inst ( .DIN1(_26840), .DIN2(_46548), .Q(_46232) );
  nnd2s1 _46933_inst ( .DIN1(_46272), .DIN2(_46448), .Q(_46548) );
  nor2s1 _46934_inst ( .DIN1(_46549), .DIN2(_46550), .Q(_46535) );
  nnd2s1 _46935_inst ( .DIN1(_46476), .DIN2(_46551), .Q(_46550) );
  nnd2s1 _46936_inst ( .DIN1(_46346), .DIN2(_46145), .Q(_46551) );
  and2s1 _46937_inst ( .DIN1(_46552), .DIN2(_46553), .Q(_46476) );
  nnd2s1 _46938_inst ( .DIN1(_46554), .DIN2(_46127), .Q(_46553) );
  nnd2s1 _46939_inst ( .DIN1(_46555), .DIN2(_46556), .Q(_46554) );
  nor2s1 _46940_inst ( .DIN1(_46557), .DIN2(_46558), .Q(_46556) );
  nnd2s1 _46941_inst ( .DIN1(_46345), .DIN2(_46278), .Q(_46558) );
  nor2s1 _46942_inst ( .DIN1(______[21]), .DIN2(_46257), .Q(_46557) );
  nor2s1 _46943_inst ( .DIN1(_46559), .DIN2(_46560), .Q(_46555) );
  or2s1 _46944_inst ( .DIN1(_46123), .DIN2(_46198), .Q(_46560) );
  nnd2s1 _46945_inst ( .DIN1(_46561), .DIN2(_46562), .Q(_46549) );
  nnd2s1 _46946_inst ( .DIN1(_46563), .DIN2(_46127), .Q(_46562) );
  nnd2s1 _46947_inst ( .DIN1(_46564), .DIN2(_46565), .Q(_46563) );
  nor2s1 _46948_inst ( .DIN1(_46459), .DIN2(_46472), .Q(_46565) );
  hi1s1 _46949_inst ( .DIN(_46417), .Q(_46472) );
  nor2s1 _46950_inst ( .DIN1(_46388), .DIN2(_46301), .Q(_46564) );
  nnd2s1 _46951_inst ( .DIN1(_46566), .DIN2(_46567), .Q(_46301) );
  nor2s1 _46952_inst ( .DIN1(_46568), .DIN2(_46569), .Q(_46567) );
  or2s1 _46953_inst ( .DIN1(_46525), .DIN2(_46449), .Q(_46569) );
  hi1s1 _46954_inst ( .DIN(_46263), .Q(_46449) );
  nor2s1 _46955_inst ( .DIN1(_46470), .DIN2(_46155), .Q(_46566) );
  hi1s1 _46956_inst ( .DIN(_46570), .Q(_46155) );
  nnd2s1 _46957_inst ( .DIN1(_46117), .DIN2(_26840), .Q(_46561) );
  nnd2s1 _46958_inst ( .DIN1(_46571), .DIN2(_46572), .Q(____3___________[10])
         );
  nor2s1 _46959_inst ( .DIN1(_46573), .DIN2(_46574), .Q(_46572) );
  nnd2s1 _46960_inst ( .DIN1(_46575), .DIN2(_46576), .Q(_46574) );
  nor2s1 _46961_inst ( .DIN1(_46577), .DIN2(_46578), .Q(_46576) );
  nor2s1 _46962_inst ( .DIN1(_46363), .DIN2(_46579), .Q(_46578) );
  nor2s1 _46963_inst ( .DIN1(_46580), .DIN2(_46581), .Q(_46579) );
  nnd2s1 _46964_inst ( .DIN1(_46527), .DIN2(_46230), .Q(_46581) );
  nor2s1 _46965_inst ( .DIN1(_46582), .DIN2(_26782), .Q(_46577) );
  nor2s1 _46966_inst ( .DIN1(_46329), .DIN2(_46210), .Q(_46582) );
  nor2s1 _46967_inst ( .DIN1(_46583), .DIN2(_46584), .Q(_46575) );
  nor2s1 _46968_inst ( .DIN1(_46258), .DIN2(_46271), .Q(_46584) );
  nor2s1 _46969_inst ( .DIN1(_46585), .DIN2(_46305), .Q(_46583) );
  nor2s1 _46970_inst ( .DIN1(_46144), .DIN2(_46586), .Q(_46585) );
  nnd2s1 _46971_inst ( .DIN1(_46189), .DIN2(_46121), .Q(_46586) );
  nor2s1 _46972_inst ( .DIN1(_46197), .DIN2(_46568), .Q(_46121) );
  and2s1 _46973_inst ( .DIN1(_46587), .DIN2(_46588), .Q(_46189) );
  nor2s1 _46974_inst ( .DIN1(_46443), .DIN2(_46117), .Q(_46588) );
  hi1s1 _46975_inst ( .DIN(_46272), .Q(_46443) );
  nor2s1 _46976_inst ( .DIN1(_46589), .DIN2(_46590), .Q(_46587) );
  nor2s1 _46977_inst ( .DIN1(_46591), .DIN2(_46592), .Q(_46590) );
  hi1s1 _46978_inst ( .DIN(_46423), .Q(_46589) );
  nnd2s1 _46979_inst ( .DIN1(_46593), .DIN2(_46223), .Q(_46144) );
  nor2s1 _46980_inst ( .DIN1(_46495), .DIN2(_46594), .Q(_46593) );
  nnd2s1 _46981_inst ( .DIN1(_46595), .DIN2(_46596), .Q(_46573) );
  nor2s1 _46982_inst ( .DIN1(_46315), .DIN2(_46597), .Q(_46596) );
  hi1s1 _46983_inst ( .DIN(_46481), .Q(_46597) );
  nnd2s1 _46984_inst ( .DIN1(_46598), .DIN2(_39514), .Q(_46481) );
  and2s1 _46985_inst ( .DIN1(_46599), .DIN2(_27747), .Q(_46315) );
  nor2s1 _46986_inst ( .DIN1(_26782), .DIN2(_46600), .Q(_46599) );
  nor2s1 _46987_inst ( .DIN1(_46601), .DIN2(_46602), .Q(_46595) );
  hi1s1 _46988_inst ( .DIN(_46250), .Q(_46602) );
  nnd2s1 _46989_inst ( .DIN1(_46603), .DIN2(_46604), .Q(_46250) );
  nor2s1 _46990_inst ( .DIN1(_46605), .DIN2(_46606), .Q(_46571) );
  nnd2s1 _46991_inst ( .DIN1(_46607), .DIN2(_46381), .Q(_46606) );
  and2s1 _46992_inst ( .DIN1(_46608), .DIN2(_46609), .Q(_46381) );
  nnd2s1 _46993_inst ( .DIN1(_46227), .DIN2(_46610), .Q(_46609) );
  nnd2s1 _46994_inst ( .DIN1(_46152), .DIN2(_46611), .Q(_46610) );
  nnd2s1 _46995_inst ( .DIN1(_46525), .DIN2(_26840), .Q(_46608) );
  nor2s1 _46996_inst ( .DIN1(_46285), .DIN2(_46397), .Q(_46607) );
  nnd2s1 _46997_inst ( .DIN1(_46612), .DIN2(_46613), .Q(_46397) );
  nnd2s1 _46998_inst ( .DIN1(_46614), .DIN2(_46615), .Q(_46613) );
  nnd2s1 _46999_inst ( .DIN1(_46616), .DIN2(_46145), .Q(_46612) );
  nnd2s1 _47000_inst ( .DIN1(_46617), .DIN2(_46618), .Q(_46285) );
  nor2s1 _47001_inst ( .DIN1(_46619), .DIN2(_46620), .Q(_46618) );
  nnd2s1 _47002_inst ( .DIN1(_46621), .DIN2(_46622), .Q(_46620) );
  nnd2s1 _47003_inst ( .DIN1(_46623), .DIN2(_46127), .Q(_46622) );
  nnd2s1 _47004_inst ( .DIN1(_46624), .DIN2(_46448), .Q(_46623) );
  nnd2s1 _47005_inst ( .DIN1(_26840), .DIN2(_46625), .Q(_46621) );
  nnd2s1 _47006_inst ( .DIN1(_46626), .DIN2(_46627), .Q(_46625) );
  nor2s1 _47007_inst ( .DIN1(_46628), .DIN2(_46629), .Q(_46626) );
  nnd2s1 _47008_inst ( .DIN1(_46630), .DIN2(_46631), .Q(_46619) );
  nnd2s1 _47009_inst ( .DIN1(_46118), .DIN2(_46632), .Q(_46630) );
  nnd2s1 _47010_inst ( .DIN1(_46521), .DIN2(_46633), .Q(_46632) );
  hi1s1 _47011_inst ( .DIN(_46388), .Q(_46521) );
  nnd2s1 _47012_inst ( .DIN1(_46128), .DIN2(_46185), .Q(_46388) );
  nor2s1 _47013_inst ( .DIN1(_46321), .DIN2(_46634), .Q(_46617) );
  nnd2s1 _47014_inst ( .DIN1(_46635), .DIN2(_46636), .Q(_46634) );
  nnd2s1 _47015_inst ( .DIN1(_46506), .DIN2(_46145), .Q(_46636) );
  hi1s1 _47016_inst ( .DIN(_46637), .Q(_46635) );
  nnd2s1 _47017_inst ( .DIN1(_46500), .DIN2(_46638), .Q(_46321) );
  or2s1 _47018_inst ( .DIN1(_46153), .DIN2(_26839), .Q(_46638) );
  hi1s1 _47019_inst ( .DIN(_46639), .Q(_46500) );
  nnd2s1 _47020_inst ( .DIN1(_46640), .DIN2(_46641), .Q(_46605) );
  nor2s1 _47021_inst ( .DIN1(_46444), .DIN2(_46137), .Q(_46641) );
  nnd2s1 _47022_inst ( .DIN1(_46642), .DIN2(_46643), .Q(_46137) );
  or2s1 _47023_inst ( .DIN1(_46279), .DIN2(_46258), .Q(_46643) );
  nor2s1 _47024_inst ( .DIN1(_46644), .DIN2(_46645), .Q(_46642) );
  nor2s1 _47025_inst ( .DIN1(_46646), .DIN2(_46305), .Q(_46645) );
  and2s1 _47026_inst ( .DIN1(_46154), .DIN2(_46406), .Q(_46646) );
  nor2s1 _47027_inst ( .DIN1(_46647), .DIN2(_46648), .Q(_46644) );
  nnd2s1 _47028_inst ( .DIN1(_46649), .DIN2(_46118), .Q(_46648) );
  nnd2s1 _47029_inst ( .DIN1(_46650), .DIN2(_46651), .Q(_46444) );
  nnd2s1 _47030_inst ( .DIN1(_46346), .DIN2(_46227), .Q(_46651) );
  nor2s1 _47031_inst ( .DIN1(_46652), .DIN2(_46653), .Q(_46650) );
  nor2s1 _47032_inst ( .DIN1(_26839), .DIN2(_46218), .Q(_46653) );
  hi1s1 _47033_inst ( .DIN(_46540), .Q(_46652) );
  nnd2s1 _47034_inst ( .DIN1(_46654), .DIN2(_46655), .Q(_46540) );
  nor2s1 _47035_inst ( .DIN1(_46305), .DIN2(_45546), .Q(_46654) );
  nor2s1 _47036_inst ( .DIN1(_46168), .DIN2(_46335), .Q(_46640) );
  nnd2s1 _47037_inst ( .DIN1(_46656), .DIN2(_46657), .Q(_46335) );
  nnd2s1 _47038_inst ( .DIN1(_46289), .DIN2(_46118), .Q(_46657) );
  nnd2s1 _47039_inst ( .DIN1(_46122), .DIN2(_26840), .Q(_46656) );
  hi1s1 _47040_inst ( .DIN(_46372), .Q(_46122) );
  nnd2s1 _47041_inst ( .DIN1(_46658), .DIN2(_46659), .Q(_46168) );
  nor2s1 _47042_inst ( .DIN1(_46660), .DIN2(_46661), .Q(_46659) );
  nnd2s1 _47043_inst ( .DIN1(_46193), .DIN2(_46501), .Q(_46661) );
  nor2s1 _47044_inst ( .DIN1(_46662), .DIN2(_46305), .Q(_46660) );
  nor2s1 _47045_inst ( .DIN1(_46663), .DIN2(_46664), .Q(_46662) );
  nor2s1 _47046_inst ( .DIN1(_46665), .DIN2(_46666), .Q(_46658) );
  nnd2s1 _47047_inst ( .DIN1(_46667), .DIN2(_46668), .Q(_46666) );
  nnd2s1 _47048_inst ( .DIN1(_46227), .DIN2(_46669), .Q(_46668) );
  nnd2s1 _47049_inst ( .DIN1(_46670), .DIN2(_46671), .Q(_46669) );
  nnd2s1 _47050_inst ( .DIN1(_45540), .DIN2(_46376), .Q(_46671) );
  nnd2s1 _47051_inst ( .DIN1(_46672), .DIN2(_46127), .Q(_46667) );
  nnd2s1 _47052_inst ( .DIN1(_46417), .DIN2(_46333), .Q(_46672) );
  nor2s1 _47053_inst ( .DIN1(_46363), .DIN2(_46276), .Q(_46665) );
  nnd2s1 _47054_inst ( .DIN1(_46673), .DIN2(_46674), .Q(____3___________[0])
         );
  nor2s1 _47055_inst ( .DIN1(_46675), .DIN2(_46676), .Q(_46674) );
  nnd2s1 _47056_inst ( .DIN1(_46677), .DIN2(_46678), .Q(_46676) );
  nnd2s1 _47057_inst ( .DIN1(_46118), .DIN2(_46679), .Q(_46678) );
  nnd2s1 _47058_inst ( .DIN1(_46680), .DIN2(_46681), .Q(_46679) );
  nor2s1 _47059_inst ( .DIN1(_46682), .DIN2(_46683), .Q(_46681) );
  nnd2s1 _47060_inst ( .DIN1(_46684), .DIN2(_46685), .Q(_46683) );
  nnd2s1 _47061_inst ( .DIN1(_46686), .DIN2(_46687), .Q(_46685) );
  nor2s1 _47062_inst ( .DIN1(_26540), .DIN2(_45552), .Q(_46686) );
  nnd2s1 _47063_inst ( .DIN1(_46441), .DIN2(_46688), .Q(_46684) );
  nnd2s1 _47064_inst ( .DIN1(_46689), .DIN2(_46690), .Q(_46682) );
  nnd2s1 _47065_inst ( .DIN1(_46691), .DIN2(_46692), .Q(_46690) );
  nor2s1 _47066_inst ( .DIN1(_53044), .DIN2(_45541), .Q(_46691) );
  nor2s1 _47067_inst ( .DIN1(_46117), .DIN2(_46216), .Q(_46689) );
  hi1s1 _47068_inst ( .DIN(_46158), .Q(_46216) );
  nnd2s1 _47069_inst ( .DIN1(_46693), .DIN2(_46694), .Q(_46158) );
  nor2s1 _47070_inst ( .DIN1(_28976), .DIN2(_45203), .Q(_46693) );
  hi1s1 _47071_inst ( .DIN(_46524), .Q(_46117) );
  nnd2s1 _47072_inst ( .DIN1(_46695), .DIN2(_46696), .Q(_46524) );
  nor2s1 _47073_inst ( .DIN1(_26249), .DIN2(_28976), .Q(_46695) );
  nor2s1 _47074_inst ( .DIN1(_46697), .DIN2(_46698), .Q(_46680) );
  nnd2s1 _47075_inst ( .DIN1(_46699), .DIN2(_46196), .Q(_46698) );
  nor2s1 _47076_inst ( .DIN1(_46663), .DIN2(_46700), .Q(_46196) );
  and2s1 _47077_inst ( .DIN1(_46701), .DIN2(_45194), .Q(_46700) );
  nnd2s1 _47078_inst ( .DIN1(_46702), .DIN2(_46703), .Q(_46697) );
  hi1s1 _47079_inst ( .DIN(_46704), .Q(_46703) );
  nor2s1 _47080_inst ( .DIN1(_46705), .DIN2(_46706), .Q(_46702) );
  nnd2s1 _47081_inst ( .DIN1(_46614), .DIN2(_45209), .Q(_46677) );
  hi1s1 _47082_inst ( .DIN(_46707), .Q(_45209) );
  nnd2s1 _47083_inst ( .DIN1(_46708), .DIN2(_46709), .Q(_46675) );
  nnd2s1 _47084_inst ( .DIN1(_26840), .DIN2(_46710), .Q(_46709) );
  nnd2s1 _47085_inst ( .DIN1(_46711), .DIN2(_46712), .Q(_46710) );
  nor2s1 _47086_inst ( .DIN1(_46713), .DIN2(_46714), .Q(_46712) );
  nnd2s1 _47087_inst ( .DIN1(_46544), .DIN2(_46715), .Q(_46714) );
  nor2s1 _47088_inst ( .DIN1(_46473), .DIN2(_46329), .Q(_46544) );
  hi1s1 _47089_inst ( .DIN(_46512), .Q(_46329) );
  nnd2s1 _47090_inst ( .DIN1(_46716), .DIN2(_46717), .Q(_46512) );
  nnd2s1 _47091_inst ( .DIN1(_46469), .DIN2(_46223), .Q(_46713) );
  nnd2s1 _47092_inst ( .DIN1(_45196), .DIN2(_46655), .Q(_46223) );
  nor2s1 _47093_inst ( .DIN1(_46718), .DIN2(_46719), .Q(_46711) );
  or2s1 _47094_inst ( .DIN1(_46720), .DIN2(_46509), .Q(_46719) );
  nnd2s1 _47095_inst ( .DIN1(_46670), .DIN2(_46721), .Q(_46509) );
  nnd2s1 _47096_inst ( .DIN1(_46688), .DIN2(_45197), .Q(_46721) );
  nor2s1 _47097_inst ( .DIN1(_46639), .DIN2(_46722), .Q(_46708) );
  nor2s1 _47098_inst ( .DIN1(_46363), .DIN2(_46723), .Q(_46722) );
  nor2s1 _47099_inst ( .DIN1(_46724), .DIN2(_46725), .Q(_46723) );
  nnd2s1 _47100_inst ( .DIN1(_46115), .DIN2(_46406), .Q(_46725) );
  nnd2s1 _47101_inst ( .DIN1(_45537), .DIN2(_46688), .Q(_46406) );
  nor2s1 _47102_inst ( .DIN1(_46389), .DIN2(_46616), .Q(_46115) );
  hi1s1 _47103_inst ( .DIN(_46151), .Q(_46616) );
  nnd2s1 _47104_inst ( .DIN1(_46692), .DIN2(_46726), .Q(_46151) );
  nnd2s1 _47105_inst ( .DIN1(_46153), .DIN2(_46184), .Q(_46724) );
  nnd2s1 _47106_inst ( .DIN1(_46687), .DIN2(_45198), .Q(_46184) );
  nnd2s1 _47107_inst ( .DIN1(_46376), .DIN2(_46441), .Q(_46153) );
  nor2s1 _47108_inst ( .DIN1(_46367), .DIN2(_26782), .Q(_46639) );
  nnd2s1 _47109_inst ( .DIN1(_46727), .DIN2(_46694), .Q(_46367) );
  nor2s1 _47110_inst ( .DIN1(_28976), .DIN2(_46728), .Q(_46727) );
  nor2s1 _47111_inst ( .DIN1(_46729), .DIN2(_46730), .Q(_46673) );
  nnd2s1 _47112_inst ( .DIN1(_46201), .DIN2(_46170), .Q(_46730) );
  and2s1 _47113_inst ( .DIN1(_46731), .DIN2(_46732), .Q(_46170) );
  nor2s1 _47114_inst ( .DIN1(_46733), .DIN2(_46734), .Q(_46732) );
  nnd2s1 _47115_inst ( .DIN1(_46735), .DIN2(_46736), .Q(_46734) );
  nnd2s1 _47116_inst ( .DIN1(_46737), .DIN2(_46127), .Q(_46736) );
  nnd2s1 _47117_inst ( .DIN1(_46372), .DIN2(_46185), .Q(_46737) );
  nnd2s1 _47118_inst ( .DIN1(_46738), .DIN2(_46342), .Q(_46185) );
  nnd2s1 _47119_inst ( .DIN1(_46604), .DIN2(_46701), .Q(_46372) );
  nnd2s1 _47120_inst ( .DIN1(_46289), .DIN2(_26840), .Q(_46735) );
  and2s1 _47121_inst ( .DIN1(_46717), .DIN2(_46739), .Q(_46289) );
  nor2s1 _47122_inst ( .DIN1(_26782), .DIN2(_46272), .Q(_46733) );
  nnd2s1 _47123_inst ( .DIN1(_39522), .DIN2(_46739), .Q(_46272) );
  nor2s1 _47124_inst ( .DIN1(_46637), .DIN2(_46740), .Q(_46731) );
  nnd2s1 _47125_inst ( .DIN1(_46132), .DIN2(_46552), .Q(_46740) );
  nnd2s1 _47126_inst ( .DIN1(_46197), .DIN2(_46145), .Q(_46552) );
  hi1s1 _47127_inst ( .DIN(_46331), .Q(_46197) );
  nnd2s1 _47128_inst ( .DIN1(_46741), .DIN2(_46342), .Q(_46331) );
  and2s1 _47129_inst ( .DIN1(_46742), .DIN2(_46743), .Q(_46132) );
  nor2s1 _47130_inst ( .DIN1(_46314), .DIN2(_46510), .Q(_46743) );
  and2s1 _47131_inst ( .DIN1(_46598), .DIN2(_39521), .Q(_46510) );
  nor2s1 _47132_inst ( .DIN1(_46305), .DIN2(_46744), .Q(_46598) );
  and2s1 _47133_inst ( .DIN1(_46745), .DIN2(_46701), .Q(_46314) );
  nor2s1 _47134_inst ( .DIN1(_46746), .DIN2(_46747), .Q(_46742) );
  nor2s1 _47135_inst ( .DIN1(_46258), .DIN2(_46748), .Q(_46747) );
  nor2s1 _47136_inst ( .DIN1(_46459), .DIN2(_46400), .Q(_46748) );
  hi1s1 _47137_inst ( .DIN(_46278), .Q(_46400) );
  nnd2s1 _47138_inst ( .DIN1(_46749), .DIN2(_45207), .Q(_46278) );
  hi1s1 _47139_inst ( .DIN(_46420), .Q(_46459) );
  nnd2s1 _47140_inst ( .DIN1(_46342), .DIN2(_46750), .Q(_46420) );
  nor2s1 _47141_inst ( .DIN1(_46751), .DIN2(_26782), .Q(_46746) );
  nor2s1 _47142_inst ( .DIN1(_46752), .DIN2(_46506), .Q(_46751) );
  hi1s1 _47143_inst ( .DIN(_46219), .Q(_46506) );
  nnd2s1 _47144_inst ( .DIN1(_39514), .DIN2(_46529), .Q(_46219) );
  nor2s1 _47145_inst ( .DIN1(_45552), .DIN2(_46753), .Q(_46752) );
  nnd2s1 _47146_inst ( .DIN1(_46754), .DIN2(_46755), .Q(_46637) );
  nnd2s1 _47147_inst ( .DIN1(_26840), .DIN2(_46756), .Q(_46755) );
  nnd2s1 _47148_inst ( .DIN1(_46462), .DIN2(_46422), .Q(_46756) );
  nnd2s1 _47149_inst ( .DIN1(_45196), .DIN2(_46757), .Q(_46422) );
  nnd2s1 _47150_inst ( .DIN1(_46758), .DIN2(_46127), .Q(_46754) );
  nnd2s1 _47151_inst ( .DIN1(_46309), .DIN2(_46759), .Q(_46758) );
  nnd2s1 _47152_inst ( .DIN1(_46440), .DIN2(_46441), .Q(_46759) );
  nnd2s1 _47153_inst ( .DIN1(_27743), .DIN2(_46440), .Q(_46309) );
  and2s1 _47154_inst ( .DIN1(_46238), .DIN2(_46760), .Q(_46201) );
  nnd2s1 _47155_inst ( .DIN1(_46761), .DIN2(_46127), .Q(_46760) );
  nnd2s1 _47156_inst ( .DIN1(_46762), .DIN2(_46763), .Q(_46761) );
  nor2s1 _47157_inst ( .DIN1(_46764), .DIN2(_46765), .Q(_46763) );
  nnd2s1 _47158_inst ( .DIN1(_46766), .DIN2(_46128), .Q(_46765) );
  and2s1 _47159_inst ( .DIN1(_46767), .DIN2(_46768), .Q(_46128) );
  nnd2s1 _47160_inst ( .DIN1(_46769), .DIN2(_46750), .Q(_46768) );
  nnd2s1 _47161_inst ( .DIN1(_46770), .DIN2(_46771), .Q(_46767) );
  hi1s1 _47162_inst ( .DIN(_46123), .Q(_46766) );
  nnd2s1 _47163_inst ( .DIN1(_46417), .DIN2(_46154), .Q(_46764) );
  nnd2s1 _47164_inst ( .DIN1(_45198), .DIN2(_46772), .Q(_46154) );
  nnd2s1 _47165_inst ( .DIN1(_46312), .DIN2(_46750), .Q(_46417) );
  nor2s1 _47166_inst ( .DIN1(_46773), .DIN2(_46774), .Q(_46762) );
  nnd2s1 _47167_inst ( .DIN1(_46775), .DIN2(_46624), .Q(_46774) );
  and2s1 _47168_inst ( .DIN1(_46263), .DIN2(_46485), .Q(_46624) );
  nnd2s1 _47169_inst ( .DIN1(_46726), .DIN2(_46772), .Q(_46485) );
  nnd2s1 _47170_inst ( .DIN1(_46776), .DIN2(_46342), .Q(_46263) );
  hi1s1 _47171_inst ( .DIN(_46559), .Q(_46775) );
  nnd2s1 _47172_inst ( .DIN1(_46777), .DIN2(_46129), .Q(_46559) );
  nnd2s1 _47173_inst ( .DIN1(_46341), .DIN2(_46771), .Q(_46129) );
  and2s1 _47174_inst ( .DIN1(_46333), .DIN2(_46279), .Q(_46777) );
  nnd2s1 _47175_inst ( .DIN1(_46341), .DIN2(_46769), .Q(_46279) );
  nnd2s1 _47176_inst ( .DIN1(_46770), .DIN2(_46769), .Q(_46333) );
  nnd2s1 _47177_inst ( .DIN1(_46778), .DIN2(_46779), .Q(_46773) );
  nnd2s1 _47178_inst ( .DIN1(______[21]), .DIN2(_46780), .Q(_46779) );
  nnd2s1 _47179_inst ( .DIN1(_46781), .DIN2(_46782), .Q(_46780) );
  nor2s1 _47180_inst ( .DIN1(_46783), .DIN2(_46784), .Q(_46782) );
  nnd2s1 _47181_inst ( .DIN1(_46448), .DIN2(_46230), .Q(_46784) );
  nnd2s1 _47182_inst ( .DIN1(_46785), .DIN2(_46529), .Q(_46230) );
  nnd2s1 _47183_inst ( .DIN1(_39522), .DIN2(_46649), .Q(_46448) );
  hi1s1 _47184_inst ( .DIN(_46218), .Q(_46783) );
  nnd2s1 _47185_inst ( .DIN1(_46786), .DIN2(_46785), .Q(_46218) );
  nor2s1 _47186_inst ( .DIN1(_29221), .DIN2(_46787), .Q(_46786) );
  nor2s1 _47187_inst ( .DIN1(_46788), .DIN2(_46789), .Q(_46781) );
  nnd2s1 _47188_inst ( .DIN1(_46633), .DIN2(_46458), .Q(_46789) );
  hi1s1 _47189_inst ( .DIN(_46790), .Q(_46458) );
  and2s1 _47190_inst ( .DIN1(_46222), .DIN2(_46791), .Q(_46633) );
  nnd2s1 _47191_inst ( .DIN1(_46792), .DIN2(_46696), .Q(_46791) );
  hi1s1 _47192_inst ( .DIN(_46547), .Q(_46696) );
  nnd2s1 _47193_inst ( .DIN1(_46793), .DIN2(_46794), .Q(_46547) );
  nor2s1 _47194_inst ( .DIN1(_46795), .DIN2(_26575), .Q(_46794) );
  nor2s1 _47195_inst ( .DIN1(_26328), .DIN2(_46796), .Q(_46793) );
  nor2s1 _47196_inst ( .DIN1(_26249), .DIN2(_29221), .Q(_46792) );
  nnd2s1 _47197_inst ( .DIN1(_46797), .DIN2(_46785), .Q(_46222) );
  hi1s1 _47198_inst ( .DIN(_45211), .Q(_46785) );
  hi1s1 _47199_inst ( .DIN(_46715), .Q(_46788) );
  nor2s1 _47200_inst ( .DIN1(_46426), .DIN2(_46798), .Q(_46715) );
  and2s1 _47201_inst ( .DIN1(_27747), .DIN2(_46772), .Q(_46798) );
  nor2s1 _47202_inst ( .DIN1(_39516), .DIN2(_46753), .Q(_46426) );
  nnd2s1 _47203_inst ( .DIN1(_46799), .DIN2(_46800), .Q(_46778) );
  nnd2s1 _47204_inst ( .DIN1(_46801), .DIN2(_46802), .Q(_46799) );
  nor2s1 _47205_inst ( .DIN1(_46628), .DIN2(_46410), .Q(_46802) );
  hi1s1 _47206_inst ( .DIN(_46803), .Q(_46628) );
  nor2s1 _47207_inst ( .DIN1(_46306), .DIN2(_46704), .Q(_46801) );
  nnd2s1 _47208_inst ( .DIN1(_46627), .DIN2(_46804), .Q(_46704) );
  nnd2s1 _47209_inst ( .DIN1(_46440), .DIN2(_45194), .Q(_46804) );
  and2s1 _47210_inst ( .DIN1(_46805), .DIN2(_46806), .Q(_46627) );
  nnd2s1 _47211_inst ( .DIN1(_27747), .DIN2(_46701), .Q(_46806) );
  nnd2s1 _47212_inst ( .DIN1(_46692), .DIN2(_46441), .Q(_46805) );
  nnd2s1 _47213_inst ( .DIN1(_46423), .DIN2(_46527), .Q(_46306) );
  nnd2s1 _47214_inst ( .DIN1(_46739), .DIN2(_39523), .Q(_46527) );
  and2s1 _47215_inst ( .DIN1(_46807), .DIN2(_28218), .Q(_46739) );
  nor2s1 _47216_inst ( .DIN1(_2698), .DIN2(_46796), .Q(_46807) );
  nnd2s1 _47217_inst ( .DIN1(_45212), .DIN2(_46529), .Q(_46423) );
  and2s1 _47218_inst ( .DIN1(_46631), .DIN2(_46808), .Q(_46238) );
  nnd2s1 _47219_inst ( .DIN1(_46809), .DIN2(_46687), .Q(_46808) );
  nor2s1 _47220_inst ( .DIN1(_46258), .DIN2(_45547), .Q(_46809) );
  nnd2s1 _47221_inst ( .DIN1(_46810), .DIN2(_27747), .Q(_46631) );
  nor2s1 _47222_inst ( .DIN1(_26782), .DIN2(_46592), .Q(_46810) );
  nnd2s1 _47223_inst ( .DIN1(_46136), .DIN2(_46259), .Q(_46729) );
  nnd2s1 _47224_inst ( .DIN1(_46568), .DIN2(_46127), .Q(_46259) );
  hi1s1 _47225_inst ( .DIN(_46498), .Q(_46568) );
  nnd2s1 _47226_inst ( .DIN1(_46811), .DIN2(_46769), .Q(_46498) );
  nor2s1 _47227_inst ( .DIN1(_46812), .DIN2(_46813), .Q(_46811) );
  and2s1 _47228_inst ( .DIN1(_46814), .DIN2(_46815), .Q(_46136) );
  nor2s1 _47229_inst ( .DIN1(_46816), .DIN2(_46817), .Q(_46815) );
  nnd2s1 _47230_inst ( .DIN1(_46818), .DIN2(_46819), .Q(_46817) );
  nnd2s1 _47231_inst ( .DIN1(_46190), .DIN2(_46127), .Q(_46819) );
  nnd2s1 _47232_inst ( .DIN1(_46570), .DIN2(_46345), .Q(_46190) );
  nnd2s1 _47233_inst ( .DIN1(_46776), .DIN2(_46769), .Q(_46345) );
  nor2s1 _47234_inst ( .DIN1(_46534), .DIN2(_46210), .Q(_46570) );
  and2s1 _47235_inst ( .DIN1(_46771), .DIN2(_46750), .Q(_46210) );
  nor2s1 _47236_inst ( .DIN1(_46820), .DIN2(_46821), .Q(_46750) );
  hi1s1 _47237_inst ( .DIN(_46611), .Q(_46534) );
  nnd2s1 _47238_inst ( .DIN1(_46749), .DIN2(_46822), .Q(_46611) );
  or2s1 _47239_inst ( .DIN1(_46670), .DIN2(_26782), .Q(_46818) );
  nnd2s1 _47240_inst ( .DIN1(_46615), .DIN2(_46772), .Q(_46670) );
  nnd2s1 _47241_inst ( .DIN1(_46823), .DIN2(_46824), .Q(_46816) );
  nnd2s1 _47242_inst ( .DIN1(_46825), .DIN2(_46145), .Q(_46824) );
  nnd2s1 _47243_inst ( .DIN1(_46276), .DIN2(_46280), .Q(_46825) );
  nnd2s1 _47244_inst ( .DIN1(_27742), .DIN2(_46701), .Q(_46280) );
  nnd2s1 _47245_inst ( .DIN1(_45537), .DIN2(_46440), .Q(_46276) );
  nor2s1 _47246_inst ( .DIN1(_46601), .DIN2(_46255), .Q(_46823) );
  and2s1 _47247_inst ( .DIN1(_46118), .DIN2(_46720), .Q(_46255) );
  nnd2s1 _47248_inst ( .DIN1(_46826), .DIN2(_46827), .Q(_46720) );
  nnd2s1 _47249_inst ( .DIN1(_46726), .DIN2(_46440), .Q(_46827) );
  nnd2s1 _47250_inst ( .DIN1(_46687), .DIN2(_45537), .Q(_46826) );
  and2s1 _47251_inst ( .DIN1(_46615), .DIN2(_46209), .Q(_46601) );
  nor2s1 _47252_inst ( .DIN1(_46828), .DIN2(_46305), .Q(_46209) );
  nor2s1 _47253_inst ( .DIN1(_46829), .DIN2(_46830), .Q(_46814) );
  nnd2s1 _47254_inst ( .DIN1(_46287), .DIN2(_46831), .Q(_46830) );
  hi1s1 _47255_inst ( .DIN(_46336), .Q(_46831) );
  nnd2s1 _47256_inst ( .DIN1(_46832), .DIN2(_46833), .Q(_46336) );
  or2s1 _47257_inst ( .DIN1(_46257), .DIN2(_26782), .Q(_46833) );
  nnd2s1 _47258_inst ( .DIN1(_46834), .DIN2(_46694), .Q(_46257) );
  nor2s1 _47259_inst ( .DIN1(_46728), .DIN2(_29221), .Q(_46834) );
  nor2s1 _47260_inst ( .DIN1(_46835), .DIN2(_46836), .Q(_46832) );
  nor2s1 _47261_inst ( .DIN1(_46363), .DIN2(_46183), .Q(_46836) );
  nnd2s1 _47262_inst ( .DIN1(_46604), .DIN2(_46772), .Q(_46183) );
  hi1s1 _47263_inst ( .DIN(_46145), .Q(_46363) );
  nnd2s1 _47264_inst ( .DIN1(_26839), .DIN2(_26782), .Q(_46145) );
  hi1s1 _47265_inst ( .DIN(_46193), .Q(_46835) );
  nnd2s1 _47266_inst ( .DIN1(_46837), .DIN2(_46376), .Q(_46193) );
  nor2s1 _47267_inst ( .DIN1(_46305), .DIN2(_45550), .Q(_46837) );
  hi1s1 _47268_inst ( .DIN(_45198), .Q(_45550) );
  and2s1 _47269_inst ( .DIN1(_46838), .DIN2(_46839), .Q(_46287) );
  nor2s1 _47270_inst ( .DIN1(_46840), .DIN2(_46841), .Q(_46839) );
  nnd2s1 _47271_inst ( .DIN1(_46842), .DIN2(_46843), .Q(_46841) );
  nnd2s1 _47272_inst ( .DIN1(_46410), .DIN2(_46227), .Q(_46843) );
  nor2s1 _47273_inst ( .DIN1(_39516), .DIN2(_46592), .Q(_46410) );
  nnd2s1 _47274_inst ( .DIN1(_45208), .DIN2(_46844), .Q(_39516) );
  hi1s1 _47275_inst ( .DIN(_46239), .Q(_46842) );
  nnd2s1 _47276_inst ( .DIN1(_46501), .DIN2(_46845), .Q(_46239) );
  nnd2s1 _47277_inst ( .DIN1(_46594), .DIN2(_26840), .Q(_46845) );
  hi1s1 _47278_inst ( .DIN(_46361), .Q(_46594) );
  nnd2s1 _47279_inst ( .DIN1(_46846), .DIN2(_46717), .Q(_46361) );
  nor2s1 _47280_inst ( .DIN1(_28976), .DIN2(_46787), .Q(_46846) );
  hi1s1 _47281_inst ( .DIN(_46694), .Q(_46787) );
  nor2s1 _47282_inst ( .DIN1(_46847), .DIN2(_26468), .Q(_46694) );
  nnd2s1 _47283_inst ( .DIN1(_46614), .DIN2(_45197), .Q(_46501) );
  and2s1 _47284_inst ( .DIN1(_46687), .DIN2(_26840), .Q(_46614) );
  nnd2s1 _47285_inst ( .DIN1(_46848), .DIN2(_46849), .Q(_46840) );
  nnd2s1 _47286_inst ( .DIN1(_46850), .DIN2(_46127), .Q(_46849) );
  or2s1 _47287_inst ( .DIN1(_46198), .DIN2(_46470), .Q(_46850) );
  nnd2s1 _47288_inst ( .DIN1(_46360), .DIN2(_46152), .Q(_46470) );
  nnd2s1 _47289_inst ( .DIN1(_46741), .DIN2(_46771), .Q(_46152) );
  nnd2s1 _47290_inst ( .DIN1(_46851), .DIN2(_46163), .Q(_46198) );
  and2s1 _47291_inst ( .DIN1(_46332), .DIN2(_46299), .Q(_46163) );
  nnd2s1 _47292_inst ( .DIN1(_46738), .DIN2(_46769), .Q(_46299) );
  nor2s1 _47293_inst ( .DIN1(_46852), .DIN2(_46813), .Q(_46738) );
  nnd2s1 _47294_inst ( .DIN1(_46749), .DIN2(_46853), .Q(_46332) );
  nor2s1 _47295_inst ( .DIN1(_46854), .DIN2(_46813), .Q(_46749) );
  nor2s1 _47296_inst ( .DIN1(_46855), .DIN2(_46856), .Q(_46851) );
  and2s1 _47297_inst ( .DIN1(_46342), .DIN2(_46341), .Q(_46856) );
  hi1s1 _47298_inst ( .DIN(_46857), .Q(_46342) );
  hi1s1 _47299_inst ( .DIN(_46262), .Q(_46855) );
  nnd2s1 _47300_inst ( .DIN1(_46741), .DIN2(_46769), .Q(_46262) );
  and2s1 _47301_inst ( .DIN1(_46858), .DIN2(_26468), .Q(_46769) );
  nor2s1 _47302_inst ( .DIN1(_46859), .DIN2(_46860), .Q(_46741) );
  nor2s1 _47303_inst ( .DIN1(_46861), .DIN2(_46862), .Q(_46848) );
  nor2s1 _47304_inst ( .DIN1(_46863), .DIN2(_46305), .Q(_46862) );
  nor2s1 _47305_inst ( .DIN1(_46526), .DIN2(_46663), .Q(_46863) );
  nnd2s1 _47306_inst ( .DIN1(_46864), .DIN2(_46865), .Q(_46663) );
  nnd2s1 _47307_inst ( .DIN1(_46604), .DIN2(_46376), .Q(_46865) );
  nnd2s1 _47308_inst ( .DIN1(_45540), .DIN2(_46688), .Q(_46864) );
  nor2s1 _47309_inst ( .DIN1(_45211), .DIN2(_46368), .Q(_46526) );
  nnd2s1 _47310_inst ( .DIN1(_46866), .DIN2(_46822), .Q(_45211) );
  hi1s1 _47311_inst ( .DIN(_46249), .Q(_46861) );
  nnd2s1 _47312_inst ( .DIN1(_46867), .DIN2(_46692), .Q(_46249) );
  nor2s1 _47313_inst ( .DIN1(_46258), .DIN2(_46591), .Q(_46867) );
  hi1s1 _47314_inst ( .DIN(_45537), .Q(_46591) );
  nor2s1 _47315_inst ( .DIN1(_46868), .DIN2(_46869), .Q(_46838) );
  or2s1 _47316_inst ( .DIN1(_46530), .DIN2(_46334), .Q(_46869) );
  nnd2s1 _47317_inst ( .DIN1(_46870), .DIN2(_46871), .Q(_46334) );
  nnd2s1 _47318_inst ( .DIN1(_46872), .DIN2(_46687), .Q(_46871) );
  nor2s1 _47319_inst ( .DIN1(_46707), .DIN2(_26782), .Q(_46872) );
  nor2s1 _47320_inst ( .DIN1(_45540), .DIN2(_27742), .Q(_46707) );
  nor2s1 _47321_inst ( .DIN1(_46820), .DIN2(_46812), .Q(_27742) );
  nnd2s1 _47322_inst ( .DIN1(_46603), .DIN2(_46441), .Q(_46870) );
  nor2s1 _47323_inst ( .DIN1(_46860), .DIN2(_46821), .Q(_46441) );
  nor2s1 _47324_inst ( .DIN1(_46305), .DIN2(_46753), .Q(_46603) );
  nnd2s1 _47325_inst ( .DIN1(_46873), .DIN2(_46874), .Q(_46530) );
  nnd2s1 _47326_inst ( .DIN1(_46227), .DIN2(_46718), .Q(_46874) );
  nnd2s1 _47327_inst ( .DIN1(_46875), .DIN2(_46876), .Q(_46718) );
  nnd2s1 _47328_inst ( .DIN1(_46604), .DIN2(_46688), .Q(_46876) );
  hi1s1 _47329_inst ( .DIN(_46753), .Q(_46688) );
  nnd2s1 _47330_inst ( .DIN1(_46877), .DIN2(_46878), .Q(_46753) );
  nor2s1 _47331_inst ( .DIN1(_2699), .DIN2(_26363), .Q(_46877) );
  hi1s1 _47332_inst ( .DIN(_45205), .Q(_46604) );
  nnd2s1 _47333_inst ( .DIN1(_46866), .DIN2(_46853), .Q(_45205) );
  nnd2s1 _47334_inst ( .DIN1(_27743), .DIN2(_46687), .Q(_46875) );
  and2s1 _47335_inst ( .DIN1(_46879), .DIN2(_2684), .Q(_46687) );
  nor2s1 _47336_inst ( .DIN1(_46392), .DIN2(_46880), .Q(_46873) );
  nor2s1 _47337_inst ( .DIN1(_46699), .DIN2(_46305), .Q(_46880) );
  and2s1 _47338_inst ( .DIN1(_46881), .DIN2(_46882), .Q(_46699) );
  nnd2s1 _47339_inst ( .DIN1(_46883), .DIN2(_46772), .Q(_46882) );
  nor2s1 _47340_inst ( .DIN1(_46852), .DIN2(_45204), .Q(_46883) );
  nnd2s1 _47341_inst ( .DIN1(_46440), .DIN2(_45197), .Q(_46881) );
  hi1s1 _47342_inst ( .DIN(_45552), .Q(_45197) );
  nnd2s1 _47343_inst ( .DIN1(_46822), .DIN2(_46884), .Q(_45552) );
  hi1s1 _47344_inst ( .DIN(_46828), .Q(_46440) );
  and2s1 _47345_inst ( .DIN1(_46885), .DIN2(_45540), .Q(_46392) );
  and2s1 _47346_inst ( .DIN1(_46127), .DIN2(_46376), .Q(_46885) );
  nnd2s1 _47347_inst ( .DIN1(_46886), .DIN2(_46353), .Q(_46868) );
  and2s1 _47348_inst ( .DIN1(_46887), .DIN2(_46888), .Q(_46353) );
  nnd2s1 _47349_inst ( .DIN1(_46118), .DIN2(_46889), .Q(_46888) );
  nnd2s1 _47350_inst ( .DIN1(_46890), .DIN2(_46891), .Q(_46889) );
  nnd2s1 _47351_inst ( .DIN1(_46376), .DIN2(_45198), .Q(_46891) );
  nor2s1 _47352_inst ( .DIN1(_45204), .DIN2(_46812), .Q(_45198) );
  nor2s1 _47353_inst ( .DIN1(_46892), .DIN2(_46893), .Q(_46376) );
  nnd2s1 _47354_inst ( .DIN1(_39514), .DIN2(_46649), .Q(_46890) );
  hi1s1 _47355_inst ( .DIN(_46744), .Q(_46649) );
  nnd2s1 _47356_inst ( .DIN1(_46894), .DIN2(_46895), .Q(_46744) );
  nor2s1 _47357_inst ( .DIN1(_28976), .DIN2(_26225), .Q(_46894) );
  nnd2s1 _47358_inst ( .DIN1(_46495), .DIN2(_26840), .Q(_46887) );
  hi1s1 _47359_inst ( .DIN(_46231), .Q(_46495) );
  nnd2s1 _47360_inst ( .DIN1(_46716), .DIN2(_27740), .Q(_46231) );
  nor2s1 _47361_inst ( .DIN1(_46191), .DIN2(_46487), .Q(_46886) );
  nnd2s1 _47362_inst ( .DIN1(_46896), .DIN2(_46897), .Q(_46487) );
  nnd2s1 _47363_inst ( .DIN1(_46745), .DIN2(_46692), .Q(_46897) );
  nor2s1 _47364_inst ( .DIN1(_45541), .DIN2(_46305), .Q(_46745) );
  hi1s1 _47365_inst ( .DIN(_45194), .Q(_45541) );
  nor2s1 _47366_inst ( .DIN1(_45204), .DIN2(_46859), .Q(_45194) );
  nnd2s1 _47367_inst ( .DIN1(_46118), .DIN2(_46898), .Q(_46896) );
  nnd2s1 _47368_inst ( .DIN1(_46803), .DIN2(_46899), .Q(_46898) );
  nnd2s1 _47369_inst ( .DIN1(_46655), .DIN2(_39522), .Q(_46899) );
  hi1s1 _47370_inst ( .DIN(_45546), .Q(_39522) );
  nnd2s1 _47371_inst ( .DIN1(_45208), .DIN2(_46822), .Q(_45546) );
  nnd2s1 _47372_inst ( .DIN1(_46726), .DIN2(_46701), .Q(_46803) );
  nor2s1 _47373_inst ( .DIN1(_46860), .DIN2(_46812), .Q(_46726) );
  hi1s1 _47374_inst ( .DIN(_26782), .Q(_46118) );
  nnd2s1 _47375_inst ( .DIN1(_46900), .DIN2(_46901), .Q(_46191) );
  nnd2s1 _47376_inst ( .DIN1(_26840), .DIN2(_46902), .Q(_46901) );
  nnd2s1 _47377_inst ( .DIN1(_46157), .DIN2(_46248), .Q(_46902) );
  nnd2s1 _47378_inst ( .DIN1(_46655), .DIN2(_39523), .Q(_46248) );
  hi1s1 _47379_inst ( .DIN(_46580), .Q(_46157) );
  nnd2s1 _47380_inst ( .DIN1(_46362), .DIN2(_46903), .Q(_46580) );
  nnd2s1 _47381_inst ( .DIN1(_46529), .DIN2(_27740), .Q(_46903) );
  hi1s1 _47382_inst ( .DIN(_45551), .Q(_27740) );
  nnd2s1 _47383_inst ( .DIN1(_46866), .DIN2(_46844), .Q(_45551) );
  nnd2s1 _47384_inst ( .DIN1(_45196), .DIN2(_46716), .Q(_46362) );
  and2s1 _47385_inst ( .DIN1(_46904), .DIN2(_46905), .Q(_46716) );
  nor2s1 _47386_inst ( .DIN1(_2698), .DIN2(_28976), .Q(_46904) );
  nor2s1 _47387_inst ( .DIN1(_45204), .DIN2(_46821), .Q(_45196) );
  nnd2s1 _47388_inst ( .DIN1(_2718), .DIN2(_46906), .Q(_45204) );
  nnd2s1 _47389_inst ( .DIN1(_46525), .DIN2(_46127), .Q(_46900) );
  nor2s1 _47390_inst ( .DIN1(_46313), .DIN2(_46857), .Q(_46525) );
  nnd2s1 _47391_inst ( .DIN1(_46858), .DIN2(_2684), .Q(_46857) );
  and2s1 _47392_inst ( .DIN1(_46907), .DIN2(_46908), .Q(_46858) );
  nor2s1 _47393_inst ( .DIN1(_2699), .DIN2(_46909), .Q(_46908) );
  nor2s1 _47394_inst ( .DIN1(_2697), .DIN2(_26328), .Q(_46907) );
  nnd2s1 _47395_inst ( .DIN1(_46398), .DIN2(_46910), .Q(_46829) );
  nnd2s1 _47396_inst ( .DIN1(_46346), .DIN2(_26840), .Q(_46910) );
  and2s1 _47397_inst ( .DIN1(_46911), .DIN2(_46912), .Q(_46398) );
  nnd2s1 _47398_inst ( .DIN1(_26840), .DIN2(_46913), .Q(_46912) );
  nnd2s1 _47399_inst ( .DIN1(_46914), .DIN2(_46915), .Q(_46913) );
  nnd2s1 _47400_inst ( .DIN1(_27747), .DIN2(_46692), .Q(_46915) );
  nor2s1 _47401_inst ( .DIN1(_46852), .DIN2(_46820), .Q(_27747) );
  hi1s1 _47402_inst ( .DIN(_46706), .Q(_46914) );
  nnd2s1 _47403_inst ( .DIN1(_46916), .DIN2(_46917), .Q(_46706) );
  nnd2s1 _47404_inst ( .DIN1(_45540), .DIN2(_46692), .Q(_46917) );
  hi1s1 _47405_inst ( .DIN(_46592), .Q(_46692) );
  nnd2s1 _47406_inst ( .DIN1(_46918), .DIN2(_46878), .Q(_46592) );
  and2s1 _47407_inst ( .DIN1(_46919), .DIN2(_2684), .Q(_46878) );
  nor2s1 _47408_inst ( .DIN1(_37006), .DIN2(_26328), .Q(_46919) );
  nor2s1 _47409_inst ( .DIN1(_2697), .DIN2(_26225), .Q(_46918) );
  and2s1 _47410_inst ( .DIN1(_46822), .DIN2(_46920), .Q(_45540) );
  hi1s1 _47411_inst ( .DIN(_46852), .Q(_46822) );
  nnd2s1 _47412_inst ( .DIN1(_45537), .DIN2(_46701), .Q(_46916) );
  nor2s1 _47413_inst ( .DIN1(_46860), .DIN2(_46852), .Q(_45537) );
  nnd2s1 _47414_inst ( .DIN1(_26575), .DIN2(_26249), .Q(_46852) );
  nnd2s1 _47415_inst ( .DIN1(_46921), .DIN2(_2711), .Q(_46860) );
  nor2s1 _47416_inst ( .DIN1(_53521), .DIN2(_26692), .Q(_46921) );
  hi1s1 _47417_inst ( .DIN(_46305), .Q(_46112) );
  nnd2s1 _47418_inst ( .DIN1(_46127), .DIN2(_46800), .Q(_46305) );
  hi1s1 _47419_inst ( .DIN(______[21]), .Q(_46800) );
  or2s1 _47420_inst ( .DIN1(_46462), .DIN2(_26782), .Q(_46911) );
  nnd2s1 _47421_inst ( .DIN1(_27743), .DIN2(_46772), .Q(_46462) );
  hi1s1 _47422_inst ( .DIN(_46600), .Q(_46772) );
  nnd2s1 _47423_inst ( .DIN1(_46922), .DIN2(_46895), .Q(_46600) );
  hi1s1 _47424_inst ( .DIN(_46923), .Q(_46895) );
  nor2s1 _47425_inst ( .DIN1(_2699), .DIN2(_37006), .Q(_46922) );
  hi1s1 _47426_inst ( .DIN(_45532), .Q(_27743) );
  nnd2s1 _47427_inst ( .DIN1(_45208), .DIN2(_46853), .Q(_45532) );
  and2s1 _47428_inst ( .DIN1(_46924), .DIN2(_2711), .Q(_45208) );
  and2s1 _47429_inst ( .DIN1(_26692), .DIN2(_53521), .Q(_46924) );
  nnd2s1 _47430_inst ( .DIN1(_46925), .DIN2(_46926), .Q(____2___________[9])
         );
  nor2s1 _47431_inst ( .DIN1(_46927), .DIN2(_46928), .Q(_46926) );
  nnd2s1 _47432_inst ( .DIN1(_46929), .DIN2(_46930), .Q(_46928) );
  nor2s1 _47433_inst ( .DIN1(_46931), .DIN2(_46932), .Q(_46929) );
  nnd2s1 _47434_inst ( .DIN1(_46933), .DIN2(_46934), .Q(_46927) );
  nor2s1 _47435_inst ( .DIN1(_46935), .DIN2(_46936), .Q(_46934) );
  nor2s1 _47436_inst ( .DIN1(_46937), .DIN2(_46938), .Q(_46933) );
  nor2s1 _47437_inst ( .DIN1(_46939), .DIN2(_46940), .Q(_46925) );
  nnd2s1 _47438_inst ( .DIN1(_46941), .DIN2(_46942), .Q(_46940) );
  nor2s1 _47439_inst ( .DIN1(_46943), .DIN2(_46944), .Q(_46941) );
  nnd2s1 _47440_inst ( .DIN1(_46945), .DIN2(_46946), .Q(_46939) );
  nor2s1 _47441_inst ( .DIN1(_46947), .DIN2(_46948), .Q(_46945) );
  nnd2s1 _47442_inst ( .DIN1(_46949), .DIN2(_46950), .Q(____2___________[8])
         );
  nor2s1 _47443_inst ( .DIN1(_46951), .DIN2(_46952), .Q(_46950) );
  nnd2s1 _47444_inst ( .DIN1(_46953), .DIN2(_46954), .Q(_46952) );
  nnd2s1 _47445_inst ( .DIN1(_46955), .DIN2(_46956), .Q(_46954) );
  nor2s1 _47446_inst ( .DIN1(_46957), .DIN2(_46958), .Q(_46953) );
  nor2s1 _47447_inst ( .DIN1(_46959), .DIN2(_46960), .Q(_46958) );
  nor2s1 _47448_inst ( .DIN1(_46961), .DIN2(_46962), .Q(_46957) );
  nnd2s1 _47449_inst ( .DIN1(_46963), .DIN2(_46964), .Q(_46951) );
  nor2s1 _47450_inst ( .DIN1(_46965), .DIN2(_46966), .Q(_46964) );
  nor2s1 _47451_inst ( .DIN1(_46967), .DIN2(_46968), .Q(_46966) );
  nor2s1 _47452_inst ( .DIN1(_46969), .DIN2(_46970), .Q(_46967) );
  nor2s1 _47453_inst ( .DIN1(_46971), .DIN2(_46972), .Q(_46963) );
  nor2s1 _47454_inst ( .DIN1(_46973), .DIN2(_46974), .Q(_46972) );
  nor2s1 _47455_inst ( .DIN1(_26361), .DIN2(_46975), .Q(_46971) );
  nor2s1 _47456_inst ( .DIN1(_46976), .DIN2(_46977), .Q(_46949) );
  nnd2s1 _47457_inst ( .DIN1(_46978), .DIN2(_46979), .Q(_46977) );
  nor2s1 _47458_inst ( .DIN1(_46980), .DIN2(_46981), .Q(_46978) );
  nnd2s1 _47459_inst ( .DIN1(_46982), .DIN2(_46983), .Q(_46976) );
  nor2s1 _47460_inst ( .DIN1(_46984), .DIN2(_46985), .Q(_46983) );
  nor2s1 _47461_inst ( .DIN1(_46986), .DIN2(_46987), .Q(_46982) );
  nnd2s1 _47462_inst ( .DIN1(_46988), .DIN2(_46989), .Q(____2___________[7])
         );
  nor2s1 _47463_inst ( .DIN1(_46990), .DIN2(_46991), .Q(_46989) );
  nnd2s1 _47464_inst ( .DIN1(_46992), .DIN2(_46993), .Q(_46991) );
  nor2s1 _47465_inst ( .DIN1(_46994), .DIN2(_46995), .Q(_46993) );
  nor2s1 _47466_inst ( .DIN1(_46996), .DIN2(_46997), .Q(_46995) );
  nor2s1 _47467_inst ( .DIN1(_46968), .DIN2(_46998), .Q(_46994) );
  nor2s1 _47468_inst ( .DIN1(_46999), .DIN2(_47000), .Q(_46992) );
  nor2s1 _47469_inst ( .DIN1(_46973), .DIN2(_47001), .Q(_46999) );
  nnd2s1 _47470_inst ( .DIN1(_47002), .DIN2(_47003), .Q(_46990) );
  nor2s1 _47471_inst ( .DIN1(_47004), .DIN2(_47005), .Q(_47003) );
  nnd2s1 _47472_inst ( .DIN1(_47006), .DIN2(_47007), .Q(_47005) );
  nor2s1 _47473_inst ( .DIN1(_47008), .DIN2(_47009), .Q(_47002) );
  and2s1 _47474_inst ( .DIN1(_47010), .DIN2(_47011), .Q(_47009) );
  nor2s1 _47475_inst ( .DIN1(_47012), .DIN2(_47013), .Q(_46988) );
  nnd2s1 _47476_inst ( .DIN1(_47014), .DIN2(_47015), .Q(_47013) );
  nor2s1 _47477_inst ( .DIN1(_47016), .DIN2(_47017), .Q(_47015) );
  nor2s1 _47478_inst ( .DIN1(_47018), .DIN2(_47019), .Q(_47014) );
  nnd2s1 _47479_inst ( .DIN1(_47020), .DIN2(_47021), .Q(_47012) );
  nor2s1 _47480_inst ( .DIN1(_46932), .DIN2(_47022), .Q(_47021) );
  nnd2s1 _47481_inst ( .DIN1(_47023), .DIN2(_47024), .Q(_46932) );
  nnd2s1 _47482_inst ( .DIN1(_47025), .DIN2(_47026), .Q(_47024) );
  nnd2s1 _47483_inst ( .DIN1(_47027), .DIN2(_46956), .Q(_47023) );
  nor2s1 _47484_inst ( .DIN1(_47028), .DIN2(_47029), .Q(_47020) );
  nnd2s1 _47485_inst ( .DIN1(_47030), .DIN2(_47031), .Q(____2___________[6])
         );
  nor2s1 _47486_inst ( .DIN1(_47032), .DIN2(_47033), .Q(_47031) );
  nnd2s1 _47487_inst ( .DIN1(_47034), .DIN2(_47035), .Q(_47033) );
  nor2s1 _47488_inst ( .DIN1(_47036), .DIN2(_47037), .Q(_47035) );
  nor2s1 _47489_inst ( .DIN1(_47038), .DIN2(_47039), .Q(_47037) );
  nor2s1 _47490_inst ( .DIN1(_47040), .DIN2(_46975), .Q(_47036) );
  nor2s1 _47491_inst ( .DIN1(_47041), .DIN2(_47042), .Q(_47034) );
  nor2s1 _47492_inst ( .DIN1(_46996), .DIN2(_47043), .Q(_47042) );
  nor2s1 _47493_inst ( .DIN1(_47044), .DIN2(_47045), .Q(_47041) );
  nnd2s1 _47494_inst ( .DIN1(_47046), .DIN2(_47047), .Q(_47032) );
  nor2s1 _47495_inst ( .DIN1(_47048), .DIN2(_47049), .Q(_47047) );
  hi1s1 _47496_inst ( .DIN(_47050), .Q(_47049) );
  nor2s1 _47497_inst ( .DIN1(_47051), .DIN2(_47052), .Q(_47046) );
  nor2s1 _47498_inst ( .DIN1(_47053), .DIN2(_46973), .Q(_47052) );
  nor2s1 _47499_inst ( .DIN1(_47054), .DIN2(_47055), .Q(_47053) );
  hi1s1 _47500_inst ( .DIN(_47056), .Q(_47054) );
  nor2s1 _47501_inst ( .DIN1(_47057), .DIN2(_46968), .Q(_47051) );
  nor2s1 _47502_inst ( .DIN1(_47058), .DIN2(_47059), .Q(_47057) );
  nor2s1 _47503_inst ( .DIN1(_47060), .DIN2(_47061), .Q(_47030) );
  nnd2s1 _47504_inst ( .DIN1(_47062), .DIN2(_47063), .Q(_47061) );
  hi1s1 _47505_inst ( .DIN(_47064), .Q(_47063) );
  nor2s1 _47506_inst ( .DIN1(_47065), .DIN2(_47066), .Q(_47062) );
  nnd2s1 _47507_inst ( .DIN1(_47067), .DIN2(_47068), .Q(_47060) );
  nor2s1 _47508_inst ( .DIN1(_47069), .DIN2(_47070), .Q(_47068) );
  nor2s1 _47509_inst ( .DIN1(_47028), .DIN2(_47071), .Q(_47067) );
  nnd2s1 _47510_inst ( .DIN1(_47072), .DIN2(_47073), .Q(_47028) );
  nor2s1 _47511_inst ( .DIN1(_47074), .DIN2(_47075), .Q(_47073) );
  nnd2s1 _47512_inst ( .DIN1(_47076), .DIN2(_47077), .Q(_47075) );
  or2s1 _47513_inst ( .DIN1(_47078), .DIN2(_47079), .Q(_47077) );
  nnd2s1 _47514_inst ( .DIN1(_47080), .DIN2(_47081), .Q(_47076) );
  nnd2s1 _47515_inst ( .DIN1(_47082), .DIN2(_47083), .Q(_47074) );
  or2s1 _47516_inst ( .DIN1(_47084), .DIN2(_47040), .Q(_47082) );
  nor2s1 _47517_inst ( .DIN1(_47085), .DIN2(_47086), .Q(_47072) );
  or2s1 _47518_inst ( .DIN1(_46948), .DIN2(_47087), .Q(_47086) );
  nnd2s1 _47519_inst ( .DIN1(_47088), .DIN2(_47089), .Q(_46948) );
  nnd2s1 _47520_inst ( .DIN1(_47090), .DIN2(_47091), .Q(____2___________[5])
         );
  nor2s1 _47521_inst ( .DIN1(_47092), .DIN2(_47093), .Q(_47091) );
  nnd2s1 _47522_inst ( .DIN1(_47094), .DIN2(_47089), .Q(_47093) );
  nnd2s1 _47523_inst ( .DIN1(_47095), .DIN2(_47096), .Q(_47089) );
  nor2s1 _47524_inst ( .DIN1(_47097), .DIN2(_47098), .Q(_47094) );
  nor2s1 _47525_inst ( .DIN1(_47099), .DIN2(_47100), .Q(_47098) );
  nor2s1 _47526_inst ( .DIN1(_47079), .DIN2(_47101), .Q(_47097) );
  nnd2s1 _47527_inst ( .DIN1(_47102), .DIN2(_47103), .Q(_47092) );
  nor2s1 _47528_inst ( .DIN1(_47104), .DIN2(_47105), .Q(_47103) );
  nor2s1 _47529_inst ( .DIN1(_47106), .DIN2(_47107), .Q(_47102) );
  nor2s1 _47530_inst ( .DIN1(_46968), .DIN2(_47108), .Q(_47107) );
  nor2s1 _47531_inst ( .DIN1(_47109), .DIN2(_46996), .Q(_47106) );
  nor2s1 _47532_inst ( .DIN1(_47110), .DIN2(_47055), .Q(_47109) );
  nnd2s1 _47533_inst ( .DIN1(_47111), .DIN2(_47112), .Q(_47055) );
  nor2s1 _47534_inst ( .DIN1(_47113), .DIN2(_47114), .Q(_47111) );
  nor2s1 _47535_inst ( .DIN1(_47115), .DIN2(_47116), .Q(_47090) );
  nnd2s1 _47536_inst ( .DIN1(_47117), .DIN2(_47118), .Q(_47116) );
  hi1s1 _47537_inst ( .DIN(_47119), .Q(_47118) );
  nor2s1 _47538_inst ( .DIN1(_47120), .DIN2(_47121), .Q(_47117) );
  nnd2s1 _47539_inst ( .DIN1(_47122), .DIN2(_47123), .Q(_47115) );
  nor2s1 _47540_inst ( .DIN1(_47124), .DIN2(_47125), .Q(_47123) );
  nor2s1 _47541_inst ( .DIN1(_47017), .DIN2(_47126), .Q(_47122) );
  nnd2s1 _47542_inst ( .DIN1(_47127), .DIN2(_47128), .Q(____2___________[4])
         );
  nor2s1 _47543_inst ( .DIN1(_47129), .DIN2(_47130), .Q(_47128) );
  nnd2s1 _47544_inst ( .DIN1(_47131), .DIN2(_47132), .Q(_47130) );
  nnd2s1 _47545_inst ( .DIN1(_47133), .DIN2(_47134), .Q(_47132) );
  nnd2s1 _47546_inst ( .DIN1(_47135), .DIN2(_46956), .Q(_47131) );
  nnd2s1 _47547_inst ( .DIN1(_47136), .DIN2(_47137), .Q(_47129) );
  or2s1 _47548_inst ( .DIN1(_47138), .DIN2(_47079), .Q(_47137) );
  nor2s1 _47549_inst ( .DIN1(_47139), .DIN2(_47140), .Q(_47136) );
  nor2s1 _47550_inst ( .DIN1(_47141), .DIN2(_46973), .Q(_47140) );
  nor2s1 _47551_inst ( .DIN1(_47142), .DIN2(_47143), .Q(_47141) );
  nor2s1 _47552_inst ( .DIN1(_47144), .DIN2(_26361), .Q(_47139) );
  nor2s1 _47553_inst ( .DIN1(_47011), .DIN2(_47145), .Q(_47144) );
  nor2s1 _47554_inst ( .DIN1(_47146), .DIN2(_47147), .Q(_47127) );
  nnd2s1 _47555_inst ( .DIN1(_47148), .DIN2(_47149), .Q(_47147) );
  hi1s1 _47556_inst ( .DIN(_47150), .Q(_47148) );
  nnd2s1 _47557_inst ( .DIN1(_46979), .DIN2(_46946), .Q(_47146) );
  and2s1 _47558_inst ( .DIN1(_47151), .DIN2(_47152), .Q(_46946) );
  nor2s1 _47559_inst ( .DIN1(_47153), .DIN2(_47154), .Q(_47152) );
  nnd2s1 _47560_inst ( .DIN1(_47155), .DIN2(_47156), .Q(_47154) );
  nnd2s1 _47561_inst ( .DIN1(_47080), .DIN2(_47157), .Q(_47156) );
  nor2s1 _47562_inst ( .DIN1(_26361), .DIN2(_47158), .Q(_47153) );
  nor2s1 _47563_inst ( .DIN1(_47159), .DIN2(_47160), .Q(_47151) );
  and2s1 _47564_inst ( .DIN1(_47161), .DIN2(_47162), .Q(_46979) );
  nor2s1 _47565_inst ( .DIN1(_47163), .DIN2(_47164), .Q(_47162) );
  nnd2s1 _47566_inst ( .DIN1(_47165), .DIN2(_47166), .Q(_47164) );
  hi1s1 _47567_inst ( .DIN(_47167), .Q(_47166) );
  nor2s1 _47568_inst ( .DIN1(_47168), .DIN2(_47169), .Q(_47165) );
  nor2s1 _47569_inst ( .DIN1(_46996), .DIN2(_47056), .Q(_47168) );
  nnd2s1 _47570_inst ( .DIN1(_47170), .DIN2(_47171), .Q(_47163) );
  nor2s1 _47571_inst ( .DIN1(_47172), .DIN2(_47173), .Q(_47171) );
  nor2s1 _47572_inst ( .DIN1(_47174), .DIN2(_47175), .Q(_47170) );
  nor2s1 _47573_inst ( .DIN1(_47176), .DIN2(_47177), .Q(_47175) );
  hi1s1 _47574_inst ( .DIN(_47178), .Q(_47174) );
  nor2s1 _47575_inst ( .DIN1(_47179), .DIN2(_47180), .Q(_47161) );
  nnd2s1 _47576_inst ( .DIN1(_47181), .DIN2(_47182), .Q(_47180) );
  hi1s1 _47577_inst ( .DIN(_47069), .Q(_47182) );
  nor2s1 _47578_inst ( .DIN1(_47183), .DIN2(_47184), .Q(_47181) );
  nnd2s1 _47579_inst ( .DIN1(_47185), .DIN2(_47186), .Q(_47179) );
  hi1s1 _47580_inst ( .DIN(_47125), .Q(_47186) );
  nnd2s1 _47581_inst ( .DIN1(_47187), .DIN2(_47188), .Q(_47125) );
  nor2s1 _47582_inst ( .DIN1(_47189), .DIN2(_47190), .Q(_47187) );
  nor2s1 _47583_inst ( .DIN1(_46968), .DIN2(_47191), .Q(_47190) );
  nor2s1 _47584_inst ( .DIN1(_47176), .DIN2(_46998), .Q(_47189) );
  nor2s1 _47585_inst ( .DIN1(_47192), .DIN2(_47193), .Q(_47185) );
  nnd2s1 _47586_inst ( .DIN1(_47194), .DIN2(_47195), .Q(____2___________[3])
         );
  nor2s1 _47587_inst ( .DIN1(_47196), .DIN2(_47197), .Q(_47195) );
  nnd2s1 _47588_inst ( .DIN1(_47198), .DIN2(_47199), .Q(_47197) );
  nor2s1 _47589_inst ( .DIN1(_47200), .DIN2(_47201), .Q(_47198) );
  nor2s1 _47590_inst ( .DIN1(_46959), .DIN2(_47202), .Q(_47201) );
  nor2s1 _47591_inst ( .DIN1(_46961), .DIN2(_47108), .Q(_47200) );
  hi1s1 _47592_inst ( .DIN(_47203), .Q(_47108) );
  nnd2s1 _47593_inst ( .DIN1(_47204), .DIN2(_47205), .Q(_47196) );
  nor2s1 _47594_inst ( .DIN1(_47206), .DIN2(_47207), .Q(_47205) );
  nor2s1 _47595_inst ( .DIN1(_47208), .DIN2(_26361), .Q(_47207) );
  nor2s1 _47596_inst ( .DIN1(_46258), .DIN2(_47209), .Q(_47208) );
  hi1s1 _47597_inst ( .DIN(_47210), .Q(_47206) );
  nor2s1 _47598_inst ( .DIN1(_47211), .DIN2(_47212), .Q(_47204) );
  nor2s1 _47599_inst ( .DIN1(_47213), .DIN2(_47214), .Q(_47212) );
  nor2s1 _47600_inst ( .DIN1(_47215), .DIN2(_47099), .Q(_47211) );
  nor2s1 _47601_inst ( .DIN1(_46969), .DIN2(_47216), .Q(_47215) );
  nnd2s1 _47602_inst ( .DIN1(_47217), .DIN2(_47100), .Q(_47216) );
  nor2s1 _47603_inst ( .DIN1(_47218), .DIN2(_47219), .Q(_47194) );
  nnd2s1 _47604_inst ( .DIN1(_47220), .DIN2(_47149), .Q(_47219) );
  and2s1 _47605_inst ( .DIN1(_47221), .DIN2(_47222), .Q(_47149) );
  nor2s1 _47606_inst ( .DIN1(_47223), .DIN2(_47224), .Q(_47222) );
  nnd2s1 _47607_inst ( .DIN1(_47225), .DIN2(_47226), .Q(_47224) );
  nnd2s1 _47608_inst ( .DIN1(_47227), .DIN2(_26792), .Q(_47226) );
  nnd2s1 _47609_inst ( .DIN1(_47229), .DIN2(_47230), .Q(_47225) );
  nnd2s1 _47610_inst ( .DIN1(_47231), .DIN2(_47232), .Q(_47223) );
  nnd2s1 _47611_inst ( .DIN1(_47233), .DIN2(_47096), .Q(_47232) );
  nor2s1 _47612_inst ( .DIN1(_47234), .DIN2(_47235), .Q(_47231) );
  nor2s1 _47613_inst ( .DIN1(_47236), .DIN2(_47237), .Q(_47235) );
  nnd2s1 _47614_inst ( .DIN1(_47238), .DIN2(_47239), .Q(_47237) );
  hi1s1 _47615_inst ( .DIN(_47007), .Q(_47234) );
  nnd2s1 _47616_inst ( .DIN1(_47010), .DIN2(_47240), .Q(_47007) );
  nnd2s1 _47617_inst ( .DIN1(_47241), .DIN2(_47039), .Q(_47240) );
  nor2s1 _47618_inst ( .DIN1(_47242), .DIN2(_47243), .Q(_47241) );
  nor2s1 _47619_inst ( .DIN1(_47244), .DIN2(_47245), .Q(_47221) );
  or2s1 _47620_inst ( .DIN1(_47246), .DIN2(_47247), .Q(_47245) );
  nnd2s1 _47621_inst ( .DIN1(_47248), .DIN2(_47249), .Q(_47244) );
  nnd2s1 _47622_inst ( .DIN1(_47113), .DIN2(_46956), .Q(_47249) );
  nor2s1 _47623_inst ( .DIN1(_47065), .DIN2(_47250), .Q(_47220) );
  nnd2s1 _47624_inst ( .DIN1(_47251), .DIN2(_47252), .Q(_47065) );
  nor2s1 _47625_inst ( .DIN1(_47253), .DIN2(_47254), .Q(_47252) );
  nnd2s1 _47626_inst ( .DIN1(_47255), .DIN2(_47256), .Q(_47254) );
  hi1s1 _47627_inst ( .DIN(_47257), .Q(_47256) );
  nnd2s1 _47628_inst ( .DIN1(_47258), .DIN2(_47259), .Q(_47255) );
  nor2s1 _47629_inst ( .DIN1(_46959), .DIN2(_39742), .Q(_47258) );
  nor2s1 _47630_inst ( .DIN1(_47099), .DIN2(_46998), .Q(_47253) );
  nor2s1 _47631_inst ( .DIN1(_47260), .DIN2(_47261), .Q(_47251) );
  nnd2s1 _47632_inst ( .DIN1(_47262), .DIN2(_47263), .Q(_47261) );
  or2s1 _47633_inst ( .DIN1(_46997), .DIN2(_46973), .Q(_47263) );
  nnd2s1 _47634_inst ( .DIN1(_47264), .DIN2(_47134), .Q(_47262) );
  nnd2s1 _47635_inst ( .DIN1(_47265), .DIN2(_47266), .Q(_47218) );
  nor2s1 _47636_inst ( .DIN1(_46947), .DIN2(_47167), .Q(_47266) );
  nnd2s1 _47637_inst ( .DIN1(_47267), .DIN2(_47268), .Q(_47167) );
  nor2s1 _47638_inst ( .DIN1(_47269), .DIN2(_47270), .Q(_47268) );
  nnd2s1 _47639_inst ( .DIN1(_47271), .DIN2(_47272), .Q(_47270) );
  nnd2s1 _47640_inst ( .DIN1(_47273), .DIN2(_47096), .Q(_47271) );
  nor2s1 _47641_inst ( .DIN1(_26361), .DIN2(_47274), .Q(_47269) );
  nor2s1 _47642_inst ( .DIN1(_47275), .DIN2(_47276), .Q(_47267) );
  nnd2s1 _47643_inst ( .DIN1(_47277), .DIN2(_47278), .Q(_47276) );
  or2s1 _47644_inst ( .DIN1(_47279), .DIN2(_47213), .Q(_47278) );
  hi1s1 _47645_inst ( .DIN(_47280), .Q(_47277) );
  nnd2s1 _47646_inst ( .DIN1(_47281), .DIN2(_47282), .Q(_46947) );
  nnd2s1 _47647_inst ( .DIN1(_47230), .DIN2(_47283), .Q(_47282) );
  nnd2s1 _47648_inst ( .DIN1(_47284), .DIN2(_46962), .Q(_47283) );
  hi1s1 _47649_inst ( .DIN(_47169), .Q(_47281) );
  nnd2s1 _47650_inst ( .DIN1(_47285), .DIN2(_47286), .Q(_47169) );
  nnd2s1 _47651_inst ( .DIN1(_47287), .DIN2(_26792), .Q(_47286) );
  nnd2s1 _47652_inst ( .DIN1(_47288), .DIN2(_47289), .Q(_47285) );
  nor2s1 _47653_inst ( .DIN1(_47290), .DIN2(_46986), .Q(_47265) );
  nnd2s1 _47654_inst ( .DIN1(_47291), .DIN2(_47292), .Q(_46986) );
  nor2s1 _47655_inst ( .DIN1(_46935), .DIN2(_47293), .Q(_47292) );
  nor2s1 _47656_inst ( .DIN1(_47294), .DIN2(_47295), .Q(_47291) );
  nor2s1 _47657_inst ( .DIN1(_47296), .DIN2(_46959), .Q(_47295) );
  nor2s1 _47658_inst ( .DIN1(_47297), .DIN2(_47298), .Q(_47296) );
  hi1s1 _47659_inst ( .DIN(_47088), .Q(_47294) );
  nnd2s1 _47660_inst ( .DIN1(_47299), .DIN2(_47300), .Q(____2___________[2])
         );
  nor2s1 _47661_inst ( .DIN1(_47301), .DIN2(_47302), .Q(_47300) );
  nnd2s1 _47662_inst ( .DIN1(_47303), .DIN2(_47304), .Q(_47302) );
  nor2s1 _47663_inst ( .DIN1(_47305), .DIN2(_47306), .Q(_47303) );
  nor2s1 _47664_inst ( .DIN1(_47038), .DIN2(_47307), .Q(_47306) );
  nor2s1 _47665_inst ( .DIN1(_47308), .DIN2(_47044), .Q(_47305) );
  nnd2s1 _47666_inst ( .DIN1(_47309), .DIN2(_47310), .Q(_47301) );
  hi1s1 _47667_inst ( .DIN(_47104), .Q(_47310) );
  nor2s1 _47668_inst ( .DIN1(_46935), .DIN2(_47311), .Q(_47309) );
  hi1s1 _47669_inst ( .DIN(_47312), .Q(_46935) );
  nor2s1 _47670_inst ( .DIN1(_47313), .DIN2(_47314), .Q(_47299) );
  nnd2s1 _47671_inst ( .DIN1(_47315), .DIN2(_47316), .Q(_47314) );
  hi1s1 _47672_inst ( .DIN(_47317), .Q(_47316) );
  nor2s1 _47673_inst ( .DIN1(_47318), .DIN2(_47319), .Q(_47315) );
  nnd2s1 _47674_inst ( .DIN1(_47320), .DIN2(_47321), .Q(_47313) );
  hi1s1 _47675_inst ( .DIN(_47071), .Q(_47321) );
  nnd2s1 _47676_inst ( .DIN1(_47322), .DIN2(_47323), .Q(_47071) );
  nor2s1 _47677_inst ( .DIN1(_47324), .DIN2(_47325), .Q(_47323) );
  nor2s1 _47678_inst ( .DIN1(_47038), .DIN2(_46127), .Q(_47325) );
  nor2s1 _47679_inst ( .DIN1(_47326), .DIN2(_47017), .Q(_47322) );
  nor2s1 _47680_inst ( .DIN1(_46996), .DIN2(_47284), .Q(_47326) );
  nor2s1 _47681_inst ( .DIN1(_47327), .DIN2(_47260), .Q(_47320) );
  nnd2s1 _47682_inst ( .DIN1(_47328), .DIN2(_47329), .Q(_47260) );
  nnd2s1 _47683_inst ( .DIN1(_47330), .DIN2(_47331), .Q(_47329) );
  nor2s1 _47684_inst ( .DIN1(_37963), .DIN2(_47332), .Q(_47331) );
  nnd2s1 _47685_inst ( .DIN1(_40482), .DIN2(_47026), .Q(_47332) );
  nor2s1 _47686_inst ( .DIN1(_34215), .DIN2(_34484), .Q(_47330) );
  nor2s1 _47687_inst ( .DIN1(_47213), .DIN2(_47333), .Q(_47327) );
  nnd2s1 _47688_inst ( .DIN1(_47334), .DIN2(_47335), .Q(____2___________[1])
         );
  nor2s1 _47689_inst ( .DIN1(_47336), .DIN2(_47337), .Q(_47335) );
  nnd2s1 _47690_inst ( .DIN1(_47338), .DIN2(_47339), .Q(_47337) );
  nor2s1 _47691_inst ( .DIN1(_47340), .DIN2(_47341), .Q(_47339) );
  nor2s1 _47692_inst ( .DIN1(_46968), .DIN2(_47342), .Q(_47341) );
  nor2s1 _47693_inst ( .DIN1(_47038), .DIN2(_47343), .Q(_47340) );
  nor2s1 _47694_inst ( .DIN1(_47344), .DIN2(_47345), .Q(_47338) );
  nor2s1 _47695_inst ( .DIN1(_47040), .DIN2(_47346), .Q(_47345) );
  nor2s1 _47696_inst ( .DIN1(_46973), .DIN2(_47112), .Q(_47344) );
  nnd2s1 _47697_inst ( .DIN1(_47347), .DIN2(_47348), .Q(_47336) );
  nor2s1 _47698_inst ( .DIN1(_47349), .DIN2(_47350), .Q(_47348) );
  nnd2s1 _47699_inst ( .DIN1(_47351), .DIN2(_47352), .Q(_47350) );
  nnd2s1 _47700_inst ( .DIN1(_47353), .DIN2(_47354), .Q(_47351) );
  nnd2s1 _47701_inst ( .DIN1(_46960), .DIN2(_47355), .Q(_47354) );
  nor2s1 _47702_inst ( .DIN1(_46996), .DIN2(_47356), .Q(_47349) );
  nor2s1 _47703_inst ( .DIN1(_47357), .DIN2(_47358), .Q(_47347) );
  nor2s1 _47704_inst ( .DIN1(_46961), .DIN2(_47359), .Q(_47358) );
  nor2s1 _47705_inst ( .DIN1(_47079), .DIN2(_47308), .Q(_47357) );
  nor2s1 _47706_inst ( .DIN1(_47360), .DIN2(_47361), .Q(_47334) );
  nnd2s1 _47707_inst ( .DIN1(_47362), .DIN2(_47363), .Q(_47361) );
  nor2s1 _47708_inst ( .DIN1(_47319), .DIN2(_47364), .Q(_47363) );
  nnd2s1 _47709_inst ( .DIN1(_47365), .DIN2(_47366), .Q(_47319) );
  nor2s1 _47710_inst ( .DIN1(_47367), .DIN2(_47368), .Q(_47366) );
  nnd2s1 _47711_inst ( .DIN1(_47369), .DIN2(_47370), .Q(_47368) );
  nnd2s1 _47712_inst ( .DIN1(_47209), .DIN2(_47134), .Q(_47369) );
  nnd2s1 _47713_inst ( .DIN1(_47371), .DIN2(_47372), .Q(_47367) );
  nnd2s1 _47714_inst ( .DIN1(_47096), .DIN2(_47373), .Q(_47372) );
  nnd2s1 _47715_inst ( .DIN1(_47078), .DIN2(_47374), .Q(_47373) );
  nor2s1 _47716_inst ( .DIN1(_47375), .DIN2(_47376), .Q(_47078) );
  nor2s1 _47717_inst ( .DIN1(_47172), .DIN2(_47377), .Q(_47371) );
  nor2s1 _47718_inst ( .DIN1(_47378), .DIN2(_47379), .Q(_47365) );
  or2s1 _47719_inst ( .DIN1(_47380), .DIN2(_47381), .Q(_47379) );
  or2s1 _47720_inst ( .DIN1(_47382), .DIN2(_47126), .Q(_47378) );
  or2s1 _47721_inst ( .DIN1(_47383), .DIN2(_47384), .Q(_47126) );
  nor2s1 _47722_inst ( .DIN1(_47217), .DIN2(_46968), .Q(_47384) );
  nor2s1 _47723_inst ( .DIN1(_47385), .DIN2(_47386), .Q(_47362) );
  nnd2s1 _47724_inst ( .DIN1(_47387), .DIN2(_47388), .Q(_47360) );
  nor2s1 _47725_inst ( .DIN1(_47389), .DIN2(_47390), .Q(_47388) );
  nor2s1 _47726_inst ( .DIN1(_47017), .DIN2(_47391), .Q(_47387) );
  nnd2s1 _47727_inst ( .DIN1(_47392), .DIN2(_47393), .Q(_47017) );
  nor2s1 _47728_inst ( .DIN1(_47394), .DIN2(_47395), .Q(_47393) );
  nnd2s1 _47729_inst ( .DIN1(_47396), .DIN2(_47397), .Q(_47395) );
  nor2s1 _47730_inst ( .DIN1(_47398), .DIN2(_47399), .Q(_47392) );
  nnd2s1 _47731_inst ( .DIN1(_47400), .DIN2(_47401), .Q(_47399) );
  nnd2s1 _47732_inst ( .DIN1(_47142), .DIN2(_26792), .Q(_47400) );
  nnd2s1 _47733_inst ( .DIN1(_47402), .DIN2(_47403), .Q(____2___________[13])
         );
  nor2s1 _47734_inst ( .DIN1(_47404), .DIN2(_47405), .Q(_47403) );
  nnd2s1 _47735_inst ( .DIN1(_47406), .DIN2(_47407), .Q(_47405) );
  hi1s1 _47736_inst ( .DIN(_47159), .Q(_47407) );
  nnd2s1 _47737_inst ( .DIN1(_47408), .DIN2(_47409), .Q(_47159) );
  nor2s1 _47738_inst ( .DIN1(_47394), .DIN2(_47008), .Q(_47409) );
  hi1s1 _47739_inst ( .DIN(_47352), .Q(_47008) );
  and2s1 _47740_inst ( .DIN1(_47410), .DIN2(_47157), .Q(_47394) );
  nor2s1 _47741_inst ( .DIN1(_47411), .DIN2(_47087), .Q(_47408) );
  nnd2s1 _47742_inst ( .DIN1(_47412), .DIN2(_47304), .Q(_47087) );
  nnd2s1 _47743_inst ( .DIN1(_47413), .DIN2(_46956), .Q(_47304) );
  nor2s1 _47744_inst ( .DIN1(_47099), .DIN2(_47414), .Q(_47411) );
  nor2s1 _47745_inst ( .DIN1(_47415), .DIN2(_47280), .Q(_47406) );
  nnd2s1 _47746_inst ( .DIN1(_47416), .DIN2(_47417), .Q(_47404) );
  nor2s1 _47747_inst ( .DIN1(_47418), .DIN2(_47173), .Q(_47417) );
  hi1s1 _47748_inst ( .DIN(_47397), .Q(_47173) );
  nnd2s1 _47749_inst ( .DIN1(_47419), .DIN2(_47420), .Q(_47397) );
  nor2s1 _47750_inst ( .DIN1(_47099), .DIN2(_44202), .Q(_47419) );
  nor2s1 _47751_inst ( .DIN1(_47421), .DIN2(_47422), .Q(_47416) );
  nor2s1 _47752_inst ( .DIN1(_47079), .DIN2(_47202), .Q(_47422) );
  nor2s1 _47753_inst ( .DIN1(_47176), .DIN2(_47217), .Q(_47421) );
  nor2s1 _47754_inst ( .DIN1(_47423), .DIN2(_47424), .Q(_47402) );
  nnd2s1 _47755_inst ( .DIN1(_47425), .DIN2(_47426), .Q(_47424) );
  hi1s1 _47756_inst ( .DIN(_47427), .Q(_47426) );
  nor2s1 _47757_inst ( .DIN1(_47120), .DIN2(_47381), .Q(_47425) );
  or2s1 _47758_inst ( .DIN1(_47018), .DIN2(_47428), .Q(_47381) );
  and2s1 _47759_inst ( .DIN1(_47264), .DIN2(_47134), .Q(_47428) );
  nnd2s1 _47760_inst ( .DIN1(_47429), .DIN2(_47430), .Q(_47018) );
  nnd2s1 _47761_inst ( .DIN1(_47431), .DIN2(_46956), .Q(_47430) );
  nor2s1 _47762_inst ( .DIN1(_47432), .DIN2(_46938), .Q(_47429) );
  nor2s1 _47763_inst ( .DIN1(_47044), .DIN2(_47433), .Q(_46938) );
  hi1s1 _47764_inst ( .DIN(_47434), .Q(_47432) );
  nnd2s1 _47765_inst ( .DIN1(_47435), .DIN2(_47436), .Q(_47120) );
  nor2s1 _47766_inst ( .DIN1(_47437), .DIN2(_47438), .Q(_47436) );
  or2s1 _47767_inst ( .DIN1(_47257), .DIN2(_47172), .Q(_47438) );
  nor2s1 _47768_inst ( .DIN1(_47084), .DIN2(_46961), .Q(_47172) );
  nor2s1 _47769_inst ( .DIN1(_47250), .DIN2(_47439), .Q(_47435) );
  nnd2s1 _47770_inst ( .DIN1(_47440), .DIN2(_47441), .Q(_47439) );
  nnd2s1 _47771_inst ( .DIN1(_47442), .DIN2(_47157), .Q(_47441) );
  hi1s1 _47772_inst ( .DIN(_47443), .Q(_47440) );
  nnd2s1 _47773_inst ( .DIN1(_47444), .DIN2(_47445), .Q(_47423) );
  nor2s1 _47774_inst ( .DIN1(_47184), .DIN2(_46987), .Q(_47445) );
  nnd2s1 _47775_inst ( .DIN1(_47446), .DIN2(_47447), .Q(_46987) );
  nor2s1 _47776_inst ( .DIN1(_47448), .DIN2(_47449), .Q(_47447) );
  nnd2s1 _47777_inst ( .DIN1(_47450), .DIN2(_47451), .Q(_47449) );
  nor2s1 _47778_inst ( .DIN1(_46961), .DIN2(_47452), .Q(_47448) );
  nor2s1 _47779_inst ( .DIN1(_47453), .DIN2(_47142), .Q(_47452) );
  hi1s1 _47780_inst ( .DIN(_47454), .Q(_47142) );
  nor2s1 _47781_inst ( .DIN1(_47383), .DIN2(_47455), .Q(_47446) );
  or2s1 _47782_inst ( .DIN1(_47070), .DIN2(_47290), .Q(_47455) );
  nnd2s1 _47783_inst ( .DIN1(_47456), .DIN2(_47457), .Q(_47290) );
  nnd2s1 _47784_inst ( .DIN1(_47458), .DIN2(_47289), .Q(_47456) );
  nnd2s1 _47785_inst ( .DIN1(_47459), .DIN2(_47460), .Q(_47070) );
  nnd2s1 _47786_inst ( .DIN1(_46956), .DIN2(_47461), .Q(_47460) );
  nnd2s1 _47787_inst ( .DIN1(_47462), .DIN2(_47463), .Q(_47383) );
  nnd2s1 _47788_inst ( .DIN1(_47464), .DIN2(_46956), .Q(_47463) );
  nnd2s1 _47789_inst ( .DIN1(_47465), .DIN2(_47010), .Q(_47462) );
  nor2s1 _47790_inst ( .DIN1(_47466), .DIN2(_47066), .Q(_47444) );
  nnd2s1 _47791_inst ( .DIN1(_47467), .DIN2(_47468), .Q(_47066) );
  nor2s1 _47792_inst ( .DIN1(_47469), .DIN2(_47470), .Q(_47468) );
  nor2s1 _47793_inst ( .DIN1(_46996), .DIN2(_47279), .Q(_47470) );
  nor2s1 _47794_inst ( .DIN1(_47471), .DIN2(_47391), .Q(_47467) );
  nnd2s1 _47795_inst ( .DIN1(_47472), .DIN2(_47473), .Q(_47391) );
  nnd2s1 _47796_inst ( .DIN1(_47474), .DIN2(_47239), .Q(_47473) );
  nnd2s1 _47797_inst ( .DIN1(_47475), .DIN2(_47134), .Q(_47472) );
  nor2s1 _47798_inst ( .DIN1(_47040), .DIN2(_47476), .Q(_47471) );
  nnd2s1 _47799_inst ( .DIN1(_47477), .DIN2(_47478), .Q(____2___________[12])
         );
  nor2s1 _47800_inst ( .DIN1(_47479), .DIN2(_47480), .Q(_47478) );
  nnd2s1 _47801_inst ( .DIN1(_47481), .DIN2(_47482), .Q(_47480) );
  nor2s1 _47802_inst ( .DIN1(_47483), .DIN2(_47484), .Q(_47482) );
  nor2s1 _47803_inst ( .DIN1(_47040), .DIN2(_47039), .Q(_47484) );
  nor2s1 _47804_inst ( .DIN1(_46996), .DIN2(_47454), .Q(_47483) );
  nor2s1 _47805_inst ( .DIN1(_47485), .DIN2(_47486), .Q(_47481) );
  nor2s1 _47806_inst ( .DIN1(_47176), .DIN2(_47191), .Q(_47485) );
  nnd2s1 _47807_inst ( .DIN1(_47487), .DIN2(_47488), .Q(_47479) );
  nor2s1 _47808_inst ( .DIN1(_47489), .DIN2(_47490), .Q(_47488) );
  nor2s1 _47809_inst ( .DIN1(_47213), .DIN2(_47491), .Q(_47490) );
  nor2s1 _47810_inst ( .DIN1(_47229), .DIN2(_47288), .Q(_47491) );
  nor2s1 _47811_inst ( .DIN1(_47492), .DIN2(_47493), .Q(_47487) );
  nor2s1 _47812_inst ( .DIN1(_47308), .DIN2(_46959), .Q(_47493) );
  nor2s1 _47813_inst ( .DIN1(_47095), .DIN2(_47494), .Q(_47308) );
  nor2s1 _47814_inst ( .DIN1(_47495), .DIN2(_26361), .Q(_47492) );
  nor2s1 _47815_inst ( .DIN1(_47145), .DIN2(_47496), .Q(_47495) );
  nor2s1 _47816_inst ( .DIN1(_47497), .DIN2(_47498), .Q(_47477) );
  nnd2s1 _47817_inst ( .DIN1(_47499), .DIN2(_47500), .Q(_47498) );
  hi1s1 _47818_inst ( .DIN(_47501), .Q(_47500) );
  nor2s1 _47819_inst ( .DIN1(_47121), .DIN2(_47385), .Q(_47499) );
  nnd2s1 _47820_inst ( .DIN1(_47502), .DIN2(_47503), .Q(_47385) );
  nnd2s1 _47821_inst ( .DIN1(_46956), .DIN2(_47504), .Q(_47503) );
  nnd2s1 _47822_inst ( .DIN1(_47298), .DIN2(_47353), .Q(_47502) );
  nnd2s1 _47823_inst ( .DIN1(_47505), .DIN2(_47506), .Q(_47121) );
  nor2s1 _47824_inst ( .DIN1(_47507), .DIN2(_47508), .Q(_47506) );
  nnd2s1 _47825_inst ( .DIN1(_47509), .DIN2(_47510), .Q(_47508) );
  nnd2s1 _47826_inst ( .DIN1(_47134), .DIN2(_47511), .Q(_47509) );
  nnd2s1 _47827_inst ( .DIN1(_47512), .DIN2(_47513), .Q(_47511) );
  nnd2s1 _47828_inst ( .DIN1(_47450), .DIN2(_47272), .Q(_47507) );
  nor2s1 _47829_inst ( .DIN1(_47415), .DIN2(_47514), .Q(_47505) );
  nnd2s1 _47830_inst ( .DIN1(_47457), .DIN2(_47515), .Q(_47514) );
  nnd2s1 _47831_inst ( .DIN1(_47516), .DIN2(_47239), .Q(_47515) );
  nnd2s1 _47832_inst ( .DIN1(_47027), .DIN2(_47230), .Q(_47457) );
  nor2s1 _47833_inst ( .DIN1(_47038), .DIN2(_47517), .Q(_47415) );
  nnd2s1 _47834_inst ( .DIN1(_47518), .DIN2(_47519), .Q(_47497) );
  nor2s1 _47835_inst ( .DIN1(_47183), .DIN2(_47398), .Q(_47519) );
  nnd2s1 _47836_inst ( .DIN1(_47520), .DIN2(_47521), .Q(_47398) );
  nor2s1 _47837_inst ( .DIN1(_47522), .DIN2(_47523), .Q(_47521) );
  nor2s1 _47838_inst ( .DIN1(_46968), .DIN2(_47524), .Q(_47523) );
  nor2s1 _47839_inst ( .DIN1(_46961), .DIN2(_47525), .Q(_47522) );
  nor2s1 _47840_inst ( .DIN1(_47466), .DIN2(_47526), .Q(_47520) );
  nnd2s1 _47841_inst ( .DIN1(_47527), .DIN2(_47528), .Q(_47466) );
  nor2s1 _47842_inst ( .DIN1(_47529), .DIN2(_47530), .Q(_47528) );
  nor2s1 _47843_inst ( .DIN1(_46961), .DIN2(_47158), .Q(_47530) );
  nor2s1 _47844_inst ( .DIN1(_46959), .DIN2(_47531), .Q(_47529) );
  nor2s1 _47845_inst ( .DIN1(_47160), .DIN2(_47275), .Q(_47527) );
  nnd2s1 _47846_inst ( .DIN1(_47532), .DIN2(_47533), .Q(_47275) );
  nnd2s1 _47847_inst ( .DIN1(_47534), .DIN2(_47259), .Q(_47533) );
  hi1s1 _47848_inst ( .DIN(_47535), .Q(_47259) );
  nor2s1 _47849_inst ( .DIN1(_46968), .DIN2(_39745), .Q(_47534) );
  nnd2s1 _47850_inst ( .DIN1(_47536), .DIN2(_47239), .Q(_47532) );
  nnd2s1 _47851_inst ( .DIN1(_47537), .DIN2(_47538), .Q(_47160) );
  nnd2s1 _47852_inst ( .DIN1(_47539), .DIN2(_26792), .Q(_47538) );
  nor2s1 _47853_inst ( .DIN1(_47540), .DIN2(_47541), .Q(_47537) );
  nor2s1 _47854_inst ( .DIN1(_47099), .DIN2(_47542), .Q(_47541) );
  nor2s1 _47855_inst ( .DIN1(_47543), .DIN2(_47544), .Q(_47540) );
  nnd2s1 _47856_inst ( .DIN1(_47096), .DIN2(_38884), .Q(_47544) );
  nnd2s1 _47857_inst ( .DIN1(_35511), .DIN2(_47545), .Q(_47543) );
  nnd2s1 _47858_inst ( .DIN1(_47546), .DIN2(_47547), .Q(_47545) );
  nnd2s1 _47859_inst ( .DIN1(_37417), .DIN2(_40482), .Q(_47547) );
  nnd2s1 _47860_inst ( .DIN1(_43905), .DIN2(_40119), .Q(_47546) );
  nnd2s1 _47861_inst ( .DIN1(_47548), .DIN2(_47549), .Q(_47183) );
  nor2s1 _47862_inst ( .DIN1(_47004), .DIN2(_47550), .Q(_47549) );
  nor2s1 _47863_inst ( .DIN1(_47551), .DIN2(_47552), .Q(_47548) );
  and2s1 _47864_inst ( .DIN1(_47010), .DIN2(_47475), .Q(_47552) );
  nor2s1 _47865_inst ( .DIN1(_47044), .DIN2(_47553), .Q(_47551) );
  nor2s1 _47866_inst ( .DIN1(_47064), .DIN2(_47247), .Q(_47518) );
  nnd2s1 _47867_inst ( .DIN1(_47554), .DIN2(_47555), .Q(_47064) );
  nor2s1 _47868_inst ( .DIN1(_47556), .DIN2(_47557), .Q(_47555) );
  nnd2s1 _47869_inst ( .DIN1(_47558), .DIN2(_47559), .Q(_47557) );
  nnd2s1 _47870_inst ( .DIN1(_47143), .DIN2(_46956), .Q(_47559) );
  nnd2s1 _47871_inst ( .DIN1(_46970), .DIN2(_26792), .Q(_47558) );
  nnd2s1 _47872_inst ( .DIN1(_47560), .DIN2(_47561), .Q(_47556) );
  or2s1 _47873_inst ( .DIN1(_47342), .DIN2(_46968), .Q(_47561) );
  nor2s1 _47874_inst ( .DIN1(_47105), .DIN2(_47562), .Q(_47560) );
  nor2s1 _47875_inst ( .DIN1(_26361), .DIN2(_47563), .Q(_47562) );
  nor2s1 _47876_inst ( .DIN1(_47564), .DIN2(_47565), .Q(_47554) );
  nnd2s1 _47877_inst ( .DIN1(_47566), .DIN2(_47567), .Q(_47565) );
  hi1s1 _47878_inst ( .DIN(_47568), .Q(_47566) );
  nnd2s1 _47879_inst ( .DIN1(_47569), .DIN2(_47570), .Q(_47564) );
  hi1s1 _47880_inst ( .DIN(_47019), .Q(_47570) );
  nnd2s1 _47881_inst ( .DIN1(_47571), .DIN2(_47572), .Q(_47019) );
  nor2s1 _47882_inst ( .DIN1(_47573), .DIN2(_47574), .Q(_47572) );
  nnd2s1 _47883_inst ( .DIN1(_47575), .DIN2(_47576), .Q(_47574) );
  nnd2s1 _47884_inst ( .DIN1(_47577), .DIN2(_47081), .Q(_47576) );
  nnd2s1 _47885_inst ( .DIN1(_47135), .DIN2(_26792), .Q(_47575) );
  hi1s1 _47886_inst ( .DIN(_46962), .Q(_47135) );
  nnd2s1 _47887_inst ( .DIN1(_47178), .DIN2(_47312), .Q(_47573) );
  nnd2s1 _47888_inst ( .DIN1(_47010), .DIN2(_47578), .Q(_47312) );
  nor2s1 _47889_inst ( .DIN1(_47443), .DIN2(_47579), .Q(_47571) );
  nnd2s1 _47890_inst ( .DIN1(_46942), .DIN2(_47580), .Q(_47579) );
  nnd2s1 _47891_inst ( .DIN1(_47458), .DIN2(_47230), .Q(_47580) );
  hi1s1 _47892_inst ( .DIN(_47333), .Q(_47458) );
  nnd2s1 _47893_inst ( .DIN1(_47581), .DIN2(_47155), .Q(_47443) );
  nnd2s1 _47894_inst ( .DIN1(_47209), .DIN2(_26792), .Q(_47155) );
  hi1s1 _47895_inst ( .DIN(_47582), .Q(_47209) );
  nnd2s1 _47896_inst ( .DIN1(_47273), .DIN2(_47583), .Q(_47581) );
  nor2s1 _47897_inst ( .DIN1(_47584), .DIN2(_47585), .Q(_47569) );
  hi1s1 _47898_inst ( .DIN(_46930), .Q(_47585) );
  nor2s1 _47899_inst ( .DIN1(_47390), .DIN2(_47586), .Q(_46930) );
  nor2s1 _47900_inst ( .DIN1(_47587), .DIN2(_46961), .Q(_47586) );
  nnd2s1 _47901_inst ( .DIN1(_47588), .DIN2(_47589), .Q(_47390) );
  nnd2s1 _47902_inst ( .DIN1(_47590), .DIN2(_26792), .Q(_47589) );
  nnd2s1 _47903_inst ( .DIN1(_47591), .DIN2(_47592), .Q(_47590) );
  nor2s1 _47904_inst ( .DIN1(_47203), .DIN2(_47227), .Q(_47591) );
  hi1s1 _47905_inst ( .DIN(_46974), .Q(_47227) );
  nnd2s1 _47906_inst ( .DIN1(_47059), .DIN2(_47239), .Q(_47588) );
  nnd2s1 _47907_inst ( .DIN1(_47593), .DIN2(_47594), .Q(____2___________[11])
         );
  nor2s1 _47908_inst ( .DIN1(_47595), .DIN2(_47596), .Q(_47594) );
  nnd2s1 _47909_inst ( .DIN1(_47597), .DIN2(_47598), .Q(_47596) );
  nor2s1 _47910_inst ( .DIN1(_47599), .DIN2(_47600), .Q(_47598) );
  nor2s1 _47911_inst ( .DIN1(_46959), .DIN2(_47592), .Q(_47600) );
  hi1s1 _47912_inst ( .DIN(_47233), .Q(_47592) );
  nor2s1 _47913_inst ( .DIN1(_47601), .DIN2(_46996), .Q(_47599) );
  nor2s1 _47914_inst ( .DIN1(_47602), .DIN2(_47603), .Q(_47601) );
  nnd2s1 _47915_inst ( .DIN1(_47604), .DIN2(_47605), .Q(_47603) );
  nor2s1 _47916_inst ( .DIN1(_47437), .DIN2(_46943), .Q(_47597) );
  nnd2s1 _47917_inst ( .DIN1(_47606), .DIN2(_47607), .Q(_46943) );
  nor2s1 _47918_inst ( .DIN1(_47608), .DIN2(_47609), .Q(_47607) );
  nnd2s1 _47919_inst ( .DIN1(_47610), .DIN2(_47611), .Q(_47609) );
  nor2s1 _47920_inst ( .DIN1(_47257), .DIN2(_47469), .Q(_47611) );
  nor2s1 _47921_inst ( .DIN1(_26361), .DIN2(_47343), .Q(_47469) );
  nor2s1 _47922_inst ( .DIN1(_47355), .DIN2(_46961), .Q(_47257) );
  nor2s1 _47923_inst ( .DIN1(_47612), .DIN2(_47613), .Q(_47610) );
  nor2s1 _47924_inst ( .DIN1(_47176), .DIN2(_47614), .Q(_47613) );
  nor2s1 _47925_inst ( .DIN1(_47615), .DIN2(_47044), .Q(_47612) );
  nnd2s1 _47926_inst ( .DIN1(_47616), .DIN2(_47617), .Q(_47608) );
  nor2s1 _47927_inst ( .DIN1(_47048), .DIN2(_47618), .Q(_47617) );
  and2s1 _47928_inst ( .DIN1(_47504), .DIN2(_47289), .Q(_47048) );
  nor2s1 _47929_inst ( .DIN1(_47324), .DIN2(_47619), .Q(_47616) );
  nor2s1 _47930_inst ( .DIN1(_47620), .DIN2(_47621), .Q(_47606) );
  nnd2s1 _47931_inst ( .DIN1(_47622), .DIN2(_47623), .Q(_47621) );
  nor2s1 _47932_inst ( .DIN1(_47000), .DIN2(_47624), .Q(_47623) );
  nnd2s1 _47933_inst ( .DIN1(_47450), .DIN2(_47625), .Q(_47000) );
  nnd2s1 _47934_inst ( .DIN1(_47494), .DIN2(_47353), .Q(_47625) );
  nnd2s1 _47935_inst ( .DIN1(_47626), .DIN2(_47010), .Q(_47450) );
  nor2s1 _47936_inst ( .DIN1(_47389), .DIN2(_47124), .Q(_47622) );
  nnd2s1 _47937_inst ( .DIN1(_47627), .DIN2(_47199), .Q(_47124) );
  nnd2s1 _47938_inst ( .DIN1(_47475), .DIN2(_47026), .Q(_47199) );
  nor2s1 _47939_inst ( .DIN1(_47628), .DIN2(_47293), .Q(_47627) );
  hi1s1 _47940_inst ( .DIN(_47629), .Q(_47293) );
  nnd2s1 _47941_inst ( .DIN1(_47630), .DIN2(_47631), .Q(_47389) );
  nor2s1 _47942_inst ( .DIN1(_47632), .DIN2(_47633), .Q(_47631) );
  nnd2s1 _47943_inst ( .DIN1(_47510), .DIN2(_47459), .Q(_47633) );
  nnd2s1 _47944_inst ( .DIN1(_47634), .DIN2(_47635), .Q(_47459) );
  nor2s1 _47945_inst ( .DIN1(_46961), .DIN2(_47636), .Q(_47634) );
  nor2s1 _47946_inst ( .DIN1(_46973), .DIN2(_47279), .Q(_47632) );
  nor2s1 _47947_inst ( .DIN1(_47584), .DIN2(_47280), .Q(_47630) );
  nnd2s1 _47948_inst ( .DIN1(_47637), .DIN2(_47638), .Q(_47280) );
  nnd2s1 _47949_inst ( .DIN1(_47114), .DIN2(_47228), .Q(_47638) );
  nor2s1 _47950_inst ( .DIN1(_47639), .DIN2(_47640), .Q(_47114) );
  or2s1 _47951_inst ( .DIN1(_47641), .DIN2(_47642), .Q(_47639) );
  nnd2s1 _47952_inst ( .DIN1(_46956), .DIN2(_47110), .Q(_47637) );
  nor2s1 _47953_inst ( .DIN1(_47099), .DIN2(_47643), .Q(_47584) );
  nnd2s1 _47954_inst ( .DIN1(_47644), .DIN2(_47645), .Q(_47620) );
  nor2s1 _47955_inst ( .DIN1(_47646), .DIN2(_47647), .Q(_47645) );
  nor2s1 _47956_inst ( .DIN1(_46959), .DIN2(_47374), .Q(_47647) );
  hi1s1 _47957_inst ( .DIN(_47273), .Q(_47374) );
  nor2s1 _47958_inst ( .DIN1(_46973), .DIN2(_47333), .Q(_47646) );
  nor2s1 _47959_inst ( .DIN1(_47648), .DIN2(_47486), .Q(_47644) );
  nnd2s1 _47960_inst ( .DIN1(_47434), .DIN2(_47649), .Q(_47486) );
  hi1s1 _47961_inst ( .DIN(_47248), .Q(_47648) );
  nor2s1 _47962_inst ( .DIN1(_47418), .DIN2(_47650), .Q(_47248) );
  nor2s1 _47963_inst ( .DIN1(_47342), .DIN2(_47176), .Q(_47650) );
  nor2s1 _47964_inst ( .DIN1(_46973), .DIN2(_47359), .Q(_47437) );
  nnd2s1 _47965_inst ( .DIN1(_47651), .DIN2(_47652), .Q(_47595) );
  nor2s1 _47966_inst ( .DIN1(_47653), .DIN2(_47311), .Q(_47652) );
  and2s1 _47967_inst ( .DIN1(_47654), .DIN2(_47230), .Q(_47311) );
  nor2s1 _47968_inst ( .DIN1(_47655), .DIN2(_47656), .Q(_47651) );
  nor2s1 _47969_inst ( .DIN1(_47657), .DIN2(_26361), .Q(_47656) );
  nor2s1 _47970_inst ( .DIN1(_47243), .DIN2(_47658), .Q(_47657) );
  nor2s1 _47971_inst ( .DIN1(_47659), .DIN2(_46968), .Q(_47655) );
  nor2s1 _47972_inst ( .DIN1(_47203), .DIN2(_46970), .Q(_47659) );
  hi1s1 _47973_inst ( .DIN(_47660), .Q(_46970) );
  nor2s1 _47974_inst ( .DIN1(_47661), .DIN2(_47662), .Q(_47593) );
  nnd2s1 _47975_inst ( .DIN1(_47663), .DIN2(_47664), .Q(_47662) );
  hi1s1 _47976_inst ( .DIN(_47665), .Q(_47664) );
  nor2s1 _47977_inst ( .DIN1(_47364), .DIN2(_47501), .Q(_47663) );
  nnd2s1 _47978_inst ( .DIN1(_47666), .DIN2(_47667), .Q(_47501) );
  nnd2s1 _47979_inst ( .DIN1(_47080), .DIN2(_47239), .Q(_47667) );
  hi1s1 _47980_inst ( .DIN(_47217), .Q(_47080) );
  nnd2s1 _47981_inst ( .DIN1(_47668), .DIN2(_37701), .Q(_47217) );
  nor2s1 _47982_inst ( .DIN1(_37963), .DIN2(_47669), .Q(_47668) );
  nnd2s1 _47983_inst ( .DIN1(_47264), .DIN2(_47010), .Q(_47666) );
  nnd2s1 _47984_inst ( .DIN1(_47670), .DIN2(_47671), .Q(_47364) );
  nor2s1 _47985_inst ( .DIN1(_47004), .DIN2(_47672), .Q(_47671) );
  nor2s1 _47986_inst ( .DIN1(_47307), .DIN2(_47040), .Q(_47672) );
  hi1s1 _47987_inst ( .DIN(_47025), .Q(_47307) );
  nnd2s1 _47988_inst ( .DIN1(_47274), .DIN2(_46975), .Q(_47025) );
  nor2s1 _47989_inst ( .DIN1(_47284), .DIN2(_47213), .Q(_47004) );
  nor2s1 _47990_inst ( .DIN1(_47673), .DIN2(_47674), .Q(_47670) );
  nor2s1 _47991_inst ( .DIN1(_46959), .DIN2(_47587), .Q(_47674) );
  nor2s1 _47992_inst ( .DIN1(_47099), .DIN2(_47191), .Q(_47673) );
  nnd2s1 _47993_inst ( .DIN1(_47675), .DIN2(_47676), .Q(_47661) );
  nor2s1 _47994_inst ( .DIN1(_47677), .DIN2(_47678), .Q(_47676) );
  nor2s1 _47995_inst ( .DIN1(_47246), .DIN2(_47380), .Q(_47675) );
  nnd2s1 _47996_inst ( .DIN1(_47679), .DIN2(_47680), .Q(_47380) );
  nor2s1 _47997_inst ( .DIN1(_47681), .DIN2(_47682), .Q(_47680) );
  nnd2s1 _47998_inst ( .DIN1(_47683), .DIN2(_47684), .Q(_47682) );
  nnd2s1 _47999_inst ( .DIN1(_47134), .DIN2(_47685), .Q(_47684) );
  nnd2s1 _48000_inst ( .DIN1(_47039), .DIN2(_47512), .Q(_47685) );
  nnd2s1 _48001_inst ( .DIN1(_46969), .DIN2(_47157), .Q(_47683) );
  nnd2s1 _48002_inst ( .DIN1(_47451), .DIN2(_47050), .Q(_47681) );
  nor2s1 _48003_inst ( .DIN1(_47686), .DIN2(_47687), .Q(_47679) );
  or2s1 _48004_inst ( .DIN1(_47193), .DIN2(_47688), .Q(_47687) );
  nnd2s1 _48005_inst ( .DIN1(_47689), .DIN2(_47690), .Q(_47246) );
  nnd2s1 _48006_inst ( .DIN1(_47691), .DIN2(_47692), .Q(_47690) );
  nor2s1 _48007_inst ( .DIN1(_46959), .DIN2(_47693), .Q(_47692) );
  nnd2s1 _48008_inst ( .DIN1(_40119), .DIN2(_35511), .Q(_47693) );
  hi1s1 _48009_inst ( .DIN(_35507), .Q(_35511) );
  nor2s1 _48010_inst ( .DIN1(_39742), .DIN2(_47694), .Q(_47691) );
  nnd2s1 _48011_inst ( .DIN1(_47431), .DIN2(_47230), .Q(_47689) );
  nnd2s1 _48012_inst ( .DIN1(_47695), .DIN2(_47696), .Q(____2___________[10])
         );
  nor2s1 _48013_inst ( .DIN1(_47697), .DIN2(_47698), .Q(_47696) );
  nnd2s1 _48014_inst ( .DIN1(_47699), .DIN2(_47700), .Q(_47698) );
  nor2s1 _48015_inst ( .DIN1(_47701), .DIN2(_47702), .Q(_47700) );
  nor2s1 _48016_inst ( .DIN1(_47703), .DIN2(_47099), .Q(_47702) );
  nor2s1 _48017_inst ( .DIN1(_47704), .DIN2(_47705), .Q(_47703) );
  nnd2s1 _48018_inst ( .DIN1(_47706), .DIN2(_47660), .Q(_47705) );
  nor2s1 _48019_inst ( .DIN1(_39745), .DIN2(_47535), .Q(_47704) );
  nnd2s1 _48020_inst ( .DIN1(_47707), .DIN2(_37417), .Q(_47535) );
  nor2s1 _48021_inst ( .DIN1(_47708), .DIN2(_46973), .Q(_47701) );
  nor2s1 _48022_inst ( .DIN1(_47431), .DIN2(_47602), .Q(_47708) );
  nnd2s1 _48023_inst ( .DIN1(_47112), .DIN2(_46974), .Q(_47602) );
  nnd2s1 _48024_inst ( .DIN1(_47709), .DIN2(_47238), .Q(_46974) );
  hi1s1 _48025_inst ( .DIN(_47636), .Q(_47238) );
  nor2s1 _48026_inst ( .DIN1(_47710), .DIN2(_47192), .Q(_47699) );
  nnd2s1 _48027_inst ( .DIN1(_47711), .DIN2(_47712), .Q(_47192) );
  nor2s1 _48028_inst ( .DIN1(_47713), .DIN2(_47688), .Q(_47712) );
  nnd2s1 _48029_inst ( .DIN1(_47714), .DIN2(_47715), .Q(_47688) );
  nnd2s1 _48030_inst ( .DIN1(_47626), .DIN2(_47134), .Q(_47715) );
  and2s1 _48031_inst ( .DIN1(_47716), .DIN2(_47717), .Q(_47626) );
  nor2s1 _48032_inst ( .DIN1(_47718), .DIN2(_34484), .Q(_47716) );
  nnd2s1 _48033_inst ( .DIN1(_47719), .DIN2(_47157), .Q(_47714) );
  nor2s1 _48034_inst ( .DIN1(_47677), .DIN2(_47085), .Q(_47711) );
  nnd2s1 _48035_inst ( .DIN1(_47720), .DIN2(_47721), .Q(_47085) );
  or2s1 _48036_inst ( .DIN1(_47512), .DIN2(_47038), .Q(_47721) );
  nor2s1 _48037_inst ( .DIN1(_47722), .DIN2(_47723), .Q(_47720) );
  hi1s1 _48038_inst ( .DIN(_47724), .Q(_47723) );
  nnd2s1 _48039_inst ( .DIN1(_47725), .DIN2(_47726), .Q(_47677) );
  nnd2s1 _48040_inst ( .DIN1(_47727), .DIN2(_47081), .Q(_47726) );
  nnd2s1 _48041_inst ( .DIN1(_47728), .DIN2(_47353), .Q(_47725) );
  nor2s1 _48042_inst ( .DIN1(_47729), .DIN2(_47328), .Q(_47710) );
  nnd2s1 _48043_inst ( .DIN1(_47730), .DIN2(_47731), .Q(_47697) );
  nor2s1 _48044_inst ( .DIN1(_47618), .DIN2(_47732), .Q(_47731) );
  nor2s1 _48045_inst ( .DIN1(_47038), .DIN2(_47733), .Q(_47732) );
  nor2s1 _48046_inst ( .DIN1(_47133), .DIN2(_46258), .Q(_47733) );
  hi1s1 _48047_inst ( .DIN(_46975), .Q(_47133) );
  nnd2s1 _48048_inst ( .DIN1(_47734), .DIN2(_47735), .Q(_46975) );
  nor2s1 _48049_inst ( .DIN1(_34215), .DIN2(_47718), .Q(_47735) );
  nor2s1 _48050_inst ( .DIN1(_35368), .DIN2(_39745), .Q(_47734) );
  hi1s1 _48051_inst ( .DIN(_47401), .Q(_47618) );
  nnd2s1 _48052_inst ( .DIN1(_46956), .DIN2(_47229), .Q(_47401) );
  nor2s1 _48053_inst ( .DIN1(_47736), .DIN2(_47737), .Q(_47730) );
  nor2s1 _48054_inst ( .DIN1(_47738), .DIN2(_26361), .Q(_47737) );
  nor2s1 _48055_inst ( .DIN1(_47539), .DIN2(_47264), .Q(_47738) );
  and2s1 _48056_inst ( .DIN1(_47739), .DIN2(_47740), .Q(_47539) );
  nor2s1 _48057_inst ( .DIN1(_43602), .DIN2(_47741), .Q(_47739) );
  nor2s1 _48058_inst ( .DIN1(_47742), .DIN2(_47044), .Q(_47736) );
  nor2s1 _48059_inst ( .DIN1(_47233), .DIN2(_47743), .Q(_47742) );
  nor2s1 _48060_inst ( .DIN1(_47744), .DIN2(_47642), .Q(_47233) );
  nor2s1 _48061_inst ( .DIN1(_47745), .DIN2(_47746), .Q(_47695) );
  nnd2s1 _48062_inst ( .DIN1(_47747), .DIN2(_47748), .Q(_47746) );
  nor2s1 _48063_inst ( .DIN1(_47686), .DIN2(_47382), .Q(_47748) );
  nnd2s1 _48064_inst ( .DIN1(_47412), .DIN2(_47749), .Q(_47382) );
  nnd2s1 _48065_inst ( .DIN1(_47750), .DIN2(_47010), .Q(_47749) );
  and2s1 _48066_inst ( .DIN1(_47751), .DIN2(_47752), .Q(_47412) );
  nnd2s1 _48067_inst ( .DIN1(_47753), .DIN2(_33181), .Q(_47752) );
  nor2s1 _48068_inst ( .DIN1(_47099), .DIN2(_47754), .Q(_47753) );
  or2s1 _48069_inst ( .DIN1(_47513), .DIN2(_46961), .Q(_47751) );
  nnd2s1 _48070_inst ( .DIN1(_47755), .DIN2(_47756), .Q(_47686) );
  nnd2s1 _48071_inst ( .DIN1(_47442), .DIN2(_47239), .Q(_47756) );
  hi1s1 _48072_inst ( .DIN(_47177), .Q(_47442) );
  nnd2s1 _48073_inst ( .DIN1(_47757), .DIN2(_47157), .Q(_47755) );
  nor2s1 _48074_inst ( .DIN1(_47758), .DIN2(_47759), .Q(_47747) );
  nnd2s1 _48075_inst ( .DIN1(_47760), .DIN2(_47761), .Q(_47745) );
  nor2s1 _48076_inst ( .DIN1(_47526), .DIN2(_47568), .Q(_47761) );
  nnd2s1 _48077_inst ( .DIN1(_47762), .DIN2(_47763), .Q(_47568) );
  nnd2s1 _48078_inst ( .DIN1(_47287), .DIN2(_46956), .Q(_47763) );
  hi1s1 _48079_inst ( .DIN(_47359), .Q(_47287) );
  nnd2s1 _48080_inst ( .DIN1(_47764), .DIN2(_47765), .Q(_47359) );
  nor2s1 _48081_inst ( .DIN1(_26229), .DIN2(_47766), .Q(_47764) );
  nnd2s1 _48082_inst ( .DIN1(_47230), .DIN2(_47110), .Q(_47762) );
  nnd2s1 _48083_inst ( .DIN1(_47767), .DIN2(_47768), .Q(_47526) );
  hi1s1 _48084_inst ( .DIN(_47184), .Q(_47768) );
  nnd2s1 _48085_inst ( .DIN1(_47769), .DIN2(_47770), .Q(_47184) );
  nnd2s1 _48086_inst ( .DIN1(_47771), .DIN2(_47772), .Q(_47770) );
  nnd2s1 _48087_inst ( .DIN1(_47654), .DIN2(_46956), .Q(_47769) );
  and2s1 _48088_inst ( .DIN1(_47773), .DIN2(_37701), .Q(_47654) );
  nor2s1 _48089_inst ( .DIN1(_47774), .DIN2(_47694), .Q(_47773) );
  nor2s1 _48090_inst ( .DIN1(_46965), .DIN2(_47619), .Q(_47767) );
  hi1s1 _48091_inst ( .DIN(_47775), .Q(_47619) );
  nor2s1 _48092_inst ( .DIN1(_47119), .DIN2(_47150), .Q(_47760) );
  nnd2s1 _48093_inst ( .DIN1(_47776), .DIN2(_47777), .Q(_47150) );
  nor2s1 _48094_inst ( .DIN1(_47778), .DIN2(_47779), .Q(_47777) );
  nnd2s1 _48095_inst ( .DIN1(_47780), .DIN2(_47781), .Q(_47779) );
  nnd2s1 _48096_inst ( .DIN1(_47203), .DIN2(_47239), .Q(_47781) );
  nor2s1 _48097_inst ( .DIN1(_47642), .DIN2(_47636), .Q(_47203) );
  nnd2s1 _48098_inst ( .DIN1(_47453), .DIN2(_47157), .Q(_47780) );
  nnd2s1 _48099_inst ( .DIN1(_47434), .DIN2(_47050), .Q(_47778) );
  nnd2s1 _48100_inst ( .DIN1(_47027), .DIN2(_47289), .Q(_47050) );
  and2s1 _48101_inst ( .DIN1(_47782), .DIN2(_38714), .Q(_47027) );
  nor2s1 _48102_inst ( .DIN1(_31291), .DIN2(_47783), .Q(_47782) );
  nnd2s1 _48103_inst ( .DIN1(_47784), .DIN2(_47785), .Q(_47434) );
  nor2s1 _48104_inst ( .DIN1(_47099), .DIN2(_43602), .Q(_47785) );
  nor2s1 _48105_inst ( .DIN1(_47786), .DIN2(_47741), .Q(_47784) );
  nor2s1 _48106_inst ( .DIN1(_47787), .DIN2(_47788), .Q(_47776) );
  nnd2s1 _48107_inst ( .DIN1(_46942), .DIN2(_47789), .Q(_47788) );
  nnd2s1 _48108_inst ( .DIN1(_46955), .DIN2(_47230), .Q(_47789) );
  hi1s1 _48109_inst ( .DIN(_47043), .Q(_46955) );
  nnd2s1 _48110_inst ( .DIN1(_47790), .DIN2(_47791), .Q(_47787) );
  nnd2s1 _48111_inst ( .DIN1(_47375), .DIN2(_47583), .Q(_47791) );
  nnd2s1 _48112_inst ( .DIN1(_47096), .DIN2(_47494), .Q(_47790) );
  nnd2s1 _48113_inst ( .DIN1(_47792), .DIN2(_47793), .Q(_47119) );
  nor2s1 _48114_inst ( .DIN1(_47794), .DIN2(_47795), .Q(_47793) );
  nnd2s1 _48115_inst ( .DIN1(_47796), .DIN2(_47797), .Q(_47795) );
  nnd2s1 _48116_inst ( .DIN1(_46969), .DIN2(_47081), .Q(_47797) );
  hi1s1 _48117_inst ( .DIN(_47414), .Q(_46969) );
  nor2s1 _48118_inst ( .DIN1(_47798), .DIN2(_47799), .Q(_47796) );
  nor2s1 _48119_inst ( .DIN1(_47800), .DIN2(_47801), .Q(_47799) );
  nor2s1 _48120_inst ( .DIN1(_47802), .DIN2(_46996), .Q(_47798) );
  nor2s1 _48121_inst ( .DIN1(_47803), .DIN2(_47804), .Q(_47802) );
  nnd2s1 _48122_inst ( .DIN1(_47279), .DIN2(_47333), .Q(_47804) );
  nnd2s1 _48123_inst ( .DIN1(_47805), .DIN2(_47352), .Q(_47794) );
  nnd2s1 _48124_inst ( .DIN1(_47806), .DIN2(_47807), .Q(_47352) );
  nor2s1 _48125_inst ( .DIN1(_34215), .DIN2(_47808), .Q(_47807) );
  nnd2s1 _48126_inst ( .DIN1(_40732), .DIN2(_40482), .Q(_47808) );
  hi1s1 _48127_inst ( .DIN(_38163), .Q(_40482) );
  hi1s1 _48128_inst ( .DIN(_37963), .Q(_40732) );
  nor2s1 _48129_inst ( .DIN1(_47040), .DIN2(_34484), .Q(_47806) );
  nor2s1 _48130_inst ( .DIN1(_47418), .DIN2(_47550), .Q(_47805) );
  nor2s1 _48131_inst ( .DIN1(_46960), .DIN2(_46961), .Q(_47418) );
  nor2s1 _48132_inst ( .DIN1(_47809), .DIN2(_47810), .Q(_47792) );
  or2s1 _48133_inst ( .DIN1(_47247), .DIN2(_47678), .Q(_47810) );
  nnd2s1 _48134_inst ( .DIN1(_47811), .DIN2(_47812), .Q(_47678) );
  nnd2s1 _48135_inst ( .DIN1(_47376), .DIN2(_47583), .Q(_47812) );
  hi1s1 _48136_inst ( .DIN(_47553), .Q(_47376) );
  nnd2s1 _48137_inst ( .DIN1(_47298), .DIN2(_47096), .Q(_47811) );
  hi1s1 _48138_inst ( .DIN(_47045), .Q(_47298) );
  nnd2s1 _48139_inst ( .DIN1(_47813), .DIN2(_47814), .Q(_47247) );
  nnd2s1 _48140_inst ( .DIN1(_47461), .DIN2(_47230), .Q(_47814) );
  hi1s1 _48141_inst ( .DIN(_47605), .Q(_47461) );
  nor2s1 _48142_inst ( .DIN1(_46936), .DIN2(_47815), .Q(_47813) );
  nor2s1 _48143_inst ( .DIN1(_47040), .DIN2(_47343), .Q(_46936) );
  nnd2s1 _48144_inst ( .DIN1(_47816), .DIN2(_47817), .Q(_47343) );
  nor2s1 _48145_inst ( .DIN1(_47818), .DIN2(_47819), .Q(_47816) );
  nnd2s1 _48146_inst ( .DIN1(_47820), .DIN2(_47567), .Q(_47809) );
  and2s1 _48147_inst ( .DIN1(_47821), .DIN2(_47822), .Q(_47567) );
  nnd2s1 _48148_inst ( .DIN1(_47297), .DIN2(_47583), .Q(_47822) );
  nor2s1 _48149_inst ( .DIN1(_47823), .DIN2(_47824), .Q(_47821) );
  nor2s1 _48150_inst ( .DIN1(_47040), .DIN2(_47274), .Q(_47824) );
  nnd2s1 _48151_inst ( .DIN1(_47825), .DIN2(_43905), .Q(_47274) );
  nor2s1 _48152_inst ( .DIN1(_39742), .DIN2(_47800), .Q(_47825) );
  hi1s1 _48153_inst ( .DIN(_47451), .Q(_47823) );
  nnd2s1 _48154_inst ( .DIN1(_47011), .DIN2(_47228), .Q(_47451) );
  nor2s1 _48155_inst ( .DIN1(_47193), .DIN2(_47826), .Q(_47820) );
  or2s1 _48156_inst ( .DIN1(_47022), .DIN2(_47827), .Q(_47193) );
  and2s1 _48157_inst ( .DIN1(_47134), .DIN2(_47578), .Q(_47827) );
  nor2s1 _48158_inst ( .DIN1(_47828), .DIN2(_47669), .Q(_47578) );
  nnd2s1 _48159_inst ( .DIN1(_34490), .DIN2(_43900), .Q(_47828) );
  hi1s1 _48160_inst ( .DIN(_47829), .Q(_43900) );
  nnd2s1 _48161_inst ( .DIN1(_47830), .DIN2(_47831), .Q(_47022) );
  nnd2s1 _48162_inst ( .DIN1(_47832), .DIN2(_47833), .Q(_47831) );
  nor2s1 _48163_inst ( .DIN1(_46959), .DIN2(_47741), .Q(_47833) );
  nor2s1 _48164_inst ( .DIN1(_47834), .DIN2(_34485), .Q(_47832) );
  nor2s1 _48165_inst ( .DIN1(_47835), .DIN2(_47836), .Q(_47830) );
  nor2s1 _48166_inst ( .DIN1(_47837), .DIN2(_47838), .Q(_47836) );
  nnd2s1 _48167_inst ( .DIN1(_40867), .DIN2(_33181), .Q(_47838) );
  nnd2s1 _48168_inst ( .DIN1(_47740), .DIN2(_47010), .Q(_47837) );
  nor2s1 _48169_inst ( .DIN1(_46973), .DIN2(_47356), .Q(_47835) );
  nnd2s1 _48170_inst ( .DIN1(_47839), .DIN2(_47840), .Q(____2___________[0])
         );
  nor2s1 _48171_inst ( .DIN1(_47841), .DIN2(_47842), .Q(_47840) );
  nnd2s1 _48172_inst ( .DIN1(_47843), .DIN2(_47844), .Q(_47842) );
  nor2s1 _48173_inst ( .DIN1(_47845), .DIN2(_47846), .Q(_47844) );
  nor2s1 _48174_inst ( .DIN1(_47847), .DIN2(_46968), .Q(_47846) );
  nor2s1 _48175_inst ( .DIN1(_47848), .DIN2(_47849), .Q(_47847) );
  nnd2s1 _48176_inst ( .DIN1(_47850), .DIN2(_47851), .Q(_47849) );
  nnd2s1 _48177_inst ( .DIN1(_47852), .DIN2(_37961), .Q(_47851) );
  nor2s1 _48178_inst ( .DIN1(_43602), .DIN2(_47786), .Q(_47852) );
  nnd2s1 _48179_inst ( .DIN1(_47420), .DIN2(_37414), .Q(_47850) );
  nnd2s1 _48180_inst ( .DIN1(_47853), .DIN2(_47854), .Q(_47848) );
  nnd2s1 _48181_inst ( .DIN1(_47855), .DIN2(_47856), .Q(_47854) );
  hi1s1 _48182_inst ( .DIN(_47783), .Q(_47856) );
  nor2s1 _48183_inst ( .DIN1(_43906), .DIN2(_47857), .Q(_47855) );
  nor2s1 _48184_inst ( .DIN1(_47536), .DIN2(_47858), .Q(_47853) );
  hi1s1 _48185_inst ( .DIN(_47542), .Q(_47858) );
  nnd2s1 _48186_inst ( .DIN1(_47859), .DIN2(_47860), .Q(_47542) );
  and2s1 _48187_inst ( .DIN1(_47861), .DIN2(_47862), .Q(_47536) );
  nor2s1 _48188_inst ( .DIN1(_47863), .DIN2(_47040), .Q(_47845) );
  nor2s1 _48189_inst ( .DIN1(_47864), .DIN2(_47865), .Q(_47863) );
  nnd2s1 _48190_inst ( .DIN1(_47866), .DIN2(_47867), .Q(_47865) );
  nnd2s1 _48191_inst ( .DIN1(_47750), .DIN2(_52863), .Q(_47867) );
  hi1s1 _48192_inst ( .DIN(_47346), .Q(_47750) );
  hi1s1 _48193_inst ( .DIN(_47496), .Q(_47866) );
  nnd2s1 _48194_inst ( .DIN1(_47868), .DIN2(_47869), .Q(_47496) );
  nnd2s1 _48195_inst ( .DIN1(_47870), .DIN2(_40867), .Q(_47869) );
  nor2s1 _48196_inst ( .DIN1(_47871), .DIN2(_34485), .Q(_47870) );
  nnd2s1 _48197_inst ( .DIN1(_47872), .DIN2(_47873), .Q(_47864) );
  nnd2s1 _48198_inst ( .DIN1(_47772), .DIN2(_31809), .Q(_47873) );
  hi1s1 _48199_inst ( .DIN(_30174), .Q(_31809) );
  nor2s1 _48200_inst ( .DIN1(_47465), .DIN2(_47011), .Q(_47872) );
  nor2s1 _48201_inst ( .DIN1(_44202), .DIN2(_47754), .Q(_47011) );
  hi1s1 _48202_inst ( .DIN(_47563), .Q(_47465) );
  nnd2s1 _48203_inst ( .DIN1(_39740), .DIN2(_47420), .Q(_47563) );
  and2s1 _48204_inst ( .DIN1(_47874), .DIN2(_40867), .Q(_47420) );
  nor2s1 _48205_inst ( .DIN1(_46937), .DIN2(_47875), .Q(_47843) );
  nor2s1 _48206_inst ( .DIN1(_26361), .DIN2(_47513), .Q(_47875) );
  nnd2s1 _48207_inst ( .DIN1(_47876), .DIN2(_47877), .Q(_47513) );
  nor2s1 _48208_inst ( .DIN1(_31291), .DIN2(_45080), .Q(_47877) );
  nor2s1 _48209_inst ( .DIN1(_38162), .DIN2(_34485), .Q(_47876) );
  nor2s1 _48210_inst ( .DIN1(_46959), .DIN2(_47553), .Q(_46937) );
  nnd2s1 _48211_inst ( .DIN1(_47878), .DIN2(_37129), .Q(_47553) );
  nnd2s1 _48212_inst ( .DIN1(_47879), .DIN2(_47880), .Q(_47841) );
  nor2s1 _48213_inst ( .DIN1(_47881), .DIN2(_47882), .Q(_47880) );
  nor2s1 _48214_inst ( .DIN1(_47883), .DIN2(_47044), .Q(_47882) );
  nor2s1 _48215_inst ( .DIN1(_47884), .DIN2(_47728), .Q(_47883) );
  hi1s1 _48216_inst ( .DIN(_47531), .Q(_47728) );
  nnd2s1 _48217_inst ( .DIN1(_47885), .DIN2(_47886), .Q(_47531) );
  nor2s1 _48218_inst ( .DIN1(_33489), .DIN2(_43906), .Q(_47886) );
  nor2s1 _48219_inst ( .DIN1(_47887), .DIN2(_35993), .Q(_47885) );
  nor2s1 _48220_inst ( .DIN1(_43602), .DIN2(_47888), .Q(_47884) );
  nor2s1 _48221_inst ( .DIN1(_47176), .DIN2(_47889), .Q(_47881) );
  nor2s1 _48222_inst ( .DIN1(_47890), .DIN2(_47577), .Q(_47889) );
  nnd2s1 _48223_inst ( .DIN1(_47414), .DIN2(_47177), .Q(_47577) );
  nnd2s1 _48224_inst ( .DIN1(_47874), .DIN2(_47891), .Q(_47177) );
  nor2s1 _48225_inst ( .DIN1(_31291), .DIN2(_30174), .Q(_47891) );
  nor2s1 _48226_inst ( .DIN1(_47892), .DIN2(_35993), .Q(_47874) );
  nnd2s1 _48227_inst ( .DIN1(_47893), .DIN2(_33181), .Q(_47414) );
  hi1s1 _48228_inst ( .DIN(_34485), .Q(_33181) );
  nor2s1 _48229_inst ( .DIN1(_47754), .DIN2(_34485), .Q(_47890) );
  hi1s1 _48230_inst ( .DIN(_47081), .Q(_47176) );
  nor2s1 _48231_inst ( .DIN1(_47894), .DIN2(_47895), .Q(_47879) );
  nor2s1 _48232_inst ( .DIN1(_47896), .DIN2(_46996), .Q(_47895) );
  nor2s1 _48233_inst ( .DIN1(_47897), .DIN2(_47898), .Q(_47896) );
  nnd2s1 _48234_inst ( .DIN1(_47454), .DIN2(_47001), .Q(_47898) );
  nnd2s1 _48235_inst ( .DIN1(_47878), .DIN2(_37961), .Q(_47454) );
  hi1s1 _48236_inst ( .DIN(_47741), .Q(_37961) );
  nnd2s1 _48237_inst ( .DIN1(_47899), .DIN2(_2627), .Q(_47741) );
  nor2s1 _48238_inst ( .DIN1(_2628), .DIN2(_47900), .Q(_47899) );
  and2s1 _48239_inst ( .DIN1(_47862), .DIN2(_38853), .Q(_47878) );
  nor2s1 _48240_inst ( .DIN1(_34214), .DIN2(_33489), .Q(_47862) );
  nor2s1 _48241_inst ( .DIN1(_53348), .DIN2(_47356), .Q(_47897) );
  nnd2s1 _48242_inst ( .DIN1(_47859), .DIN2(_47740), .Q(_47356) );
  hi1s1 _48243_inst ( .DIN(_47871), .Q(_47740) );
  nor2s1 _48244_inst ( .DIN1(_44202), .DIN2(_43904), .Q(_47859) );
  nor2s1 _48245_inst ( .DIN1(_47901), .DIN2(_47099), .Q(_47894) );
  nor2s1 _48246_inst ( .DIN1(_47453), .DIN2(_47727), .Q(_47901) );
  hi1s1 _48247_inst ( .DIN(_47524), .Q(_47727) );
  nnd2s1 _48248_inst ( .DIN1(_47902), .DIN2(_47903), .Q(_47524) );
  nor2s1 _48249_inst ( .DIN1(_43906), .DIN2(_44202), .Q(_47902) );
  hi1s1 _48250_inst ( .DIN(_47525), .Q(_47453) );
  nnd2s1 _48251_inst ( .DIN1(_47904), .DIN2(_39740), .Q(_47525) );
  nor2s1 _48252_inst ( .DIN1(_31291), .DIN2(_47871), .Q(_47904) );
  nor2s1 _48253_inst ( .DIN1(_47905), .DIN2(_47906), .Q(_47839) );
  nnd2s1 _48254_inst ( .DIN1(_47907), .DIN2(_47908), .Q(_47906) );
  nor2s1 _48255_inst ( .DIN1(_47386), .DIN2(_47427), .Q(_47908) );
  nnd2s1 _48256_inst ( .DIN1(_47909), .DIN2(_47910), .Q(_47427) );
  nor2s1 _48257_inst ( .DIN1(_47911), .DIN2(_47912), .Q(_47910) );
  nnd2s1 _48258_inst ( .DIN1(_47913), .DIN2(_47178), .Q(_47912) );
  nnd2s1 _48259_inst ( .DIN1(_47914), .DIN2(_47771), .Q(_47178) );
  nor2s1 _48260_inst ( .DIN1(_39462), .DIN2(_47834), .Q(_47914) );
  nnd2s1 _48261_inst ( .DIN1(_47757), .DIN2(_47239), .Q(_47913) );
  hi1s1 _48262_inst ( .DIN(_46998), .Q(_47757) );
  nnd2s1 _48263_inst ( .DIN1(_39740), .DIN2(_47893), .Q(_46998) );
  nnd2s1 _48264_inst ( .DIN1(_47915), .DIN2(_47775), .Q(_47911) );
  nnd2s1 _48265_inst ( .DIN1(_47134), .DIN2(_47243), .Q(_47775) );
  and2s1 _48266_inst ( .DIN1(_47916), .DIN2(_47917), .Q(_47243) );
  nor2s1 _48267_inst ( .DIN1(_38163), .DIN2(_37413), .Q(_47917) );
  nor2s1 _48268_inst ( .DIN1(_34215), .DIN2(_47829), .Q(_47916) );
  nor2s1 _48269_inst ( .DIN1(_47722), .DIN2(_47104), .Q(_47915) );
  nor2s1 _48270_inst ( .DIN1(_47342), .DIN2(_47099), .Q(_47104) );
  nnd2s1 _48271_inst ( .DIN1(_47918), .DIN2(_47635), .Q(_47342) );
  nor2s1 _48272_inst ( .DIN1(_47919), .DIN2(_47920), .Q(_47918) );
  and2s1 _48273_inst ( .DIN1(_47921), .DIN2(_39740), .Q(_47722) );
  nor2s1 _48274_inst ( .DIN1(_47099), .DIN2(_47888), .Q(_47921) );
  nor2s1 _48275_inst ( .DIN1(_47922), .DIN2(_47923), .Q(_47909) );
  or2s1 _48276_inst ( .DIN1(_47029), .DIN2(_46980), .Q(_47923) );
  nnd2s1 _48277_inst ( .DIN1(_47924), .DIN2(_47925), .Q(_46980) );
  nor2s1 _48278_inst ( .DIN1(_47324), .DIN2(_47926), .Q(_47925) );
  nnd2s1 _48279_inst ( .DIN1(_47927), .DIN2(_47396), .Q(_47926) );
  nnd2s1 _48280_inst ( .DIN1(_47928), .DIN2(_47929), .Q(_47396) );
  nor2s1 _48281_inst ( .DIN1(_47099), .DIN2(_39462), .Q(_47929) );
  nor2s1 _48282_inst ( .DIN1(_47786), .DIN2(_34485), .Q(_47928) );
  hi1s1 _48283_inst ( .DIN(_47628), .Q(_47927) );
  nor2s1 _48284_inst ( .DIN1(_47930), .DIN2(_47328), .Q(_47628) );
  nnd2s1 _48285_inst ( .DIN1(_47931), .DIN2(_47932), .Q(_47328) );
  nor2s1 _48286_inst ( .DIN1(_46961), .DIN2(_37963), .Q(_47932) );
  nor2s1 _48287_inst ( .DIN1(_47800), .DIN2(_44319), .Q(_47931) );
  hi1s1 _48288_inst ( .DIN(_47933), .Q(_47800) );
  nor2s1 _48289_inst ( .DIN1(_47100), .DIN2(_46961), .Q(_47324) );
  nnd2s1 _48290_inst ( .DIN1(_47934), .DIN2(_47635), .Q(_47100) );
  nor2s1 _48291_inst ( .DIN1(_47826), .DIN2(_47935), .Q(_47924) );
  nnd2s1 _48292_inst ( .DIN1(_47936), .DIN2(_47937), .Q(_47935) );
  nnd2s1 _48293_inst ( .DIN1(_47375), .DIN2(_47353), .Q(_47937) );
  hi1s1 _48294_inst ( .DIN(_47615), .Q(_47375) );
  nnd2s1 _48295_inst ( .DIN1(_47938), .DIN2(_37129), .Q(_47615) );
  nor2s1 _48296_inst ( .DIN1(_47857), .DIN2(_47786), .Q(_47938) );
  nnd2s1 _48297_inst ( .DIN1(_47494), .DIN2(_47583), .Q(_47936) );
  hi1s1 _48298_inst ( .DIN(_47101), .Q(_47494) );
  nnd2s1 _48299_inst ( .DIN1(_47939), .DIN2(_47940), .Q(_47101) );
  nor2s1 _48300_inst ( .DIN1(_47829), .DIN2(_44319), .Q(_47939) );
  nnd2s1 _48301_inst ( .DIN1(_47941), .DIN2(_47370), .Q(_47826) );
  nnd2s1 _48302_inst ( .DIN1(_47143), .DIN2(_47228), .Q(_47370) );
  hi1s1 _48303_inst ( .DIN(_47604), .Q(_47143) );
  nnd2s1 _48304_inst ( .DIN1(_47942), .DIN2(_39740), .Q(_47604) );
  hi1s1 _48305_inst ( .DIN(_38713), .Q(_39740) );
  nor2s1 _48306_inst ( .DIN1(_43904), .DIN2(_47943), .Q(_47942) );
  nnd2s1 _48307_inst ( .DIN1(_47944), .DIN2(_47945), .Q(_43904) );
  or2s1 _48308_inst ( .DIN1(_47039), .DIN2(_47038), .Q(_47941) );
  hi1s1 _48309_inst ( .DIN(_47026), .Q(_47038) );
  nnd2s1 _48310_inst ( .DIN1(_47946), .DIN2(_37411), .Q(_47039) );
  hi1s1 _48311_inst ( .DIN(_47857), .Q(_37411) );
  nnd2s1 _48312_inst ( .DIN1(_47510), .DIN2(_47947), .Q(_47029) );
  nnd2s1 _48313_inst ( .DIN1(_47058), .DIN2(_47081), .Q(_47947) );
  nnd2s1 _48314_inst ( .DIN1(_47099), .DIN2(_46968), .Q(_47081) );
  hi1s1 _48315_inst ( .DIN(_47191), .Q(_47058) );
  nnd2s1 _48316_inst ( .DIN1(_47948), .DIN2(_37417), .Q(_47191) );
  hi1s1 _48317_inst ( .DIN(_47718), .Q(_37417) );
  nor2s1 _48318_inst ( .DIN1(_37413), .DIN2(_47669), .Q(_47948) );
  nnd2s1 _48319_inst ( .DIN1(_46258), .DIN2(_47134), .Q(_47510) );
  hi1s1 _48320_inst ( .DIN(_46127), .Q(_46258) );
  nnd2s1 _48321_inst ( .DIN1(_47949), .DIN2(_47707), .Q(_46127) );
  nor2s1 _48322_inst ( .DIN1(_38163), .DIN2(_35507), .Q(_47707) );
  nor2s1 _48323_inst ( .DIN1(_37963), .DIN2(_37413), .Q(_47949) );
  nnd2s1 _48324_inst ( .DIN1(_47950), .DIN2(_47951), .Q(_47922) );
  nnd2s1 _48325_inst ( .DIN1(_47803), .DIN2(_47230), .Q(_47951) );
  hi1s1 _48326_inst ( .DIN(_47284), .Q(_47803) );
  nnd2s1 _48327_inst ( .DIN1(_47952), .DIN2(_43905), .Q(_47284) );
  nor2s1 _48328_inst ( .DIN1(_44319), .DIN2(_47774), .Q(_47952) );
  nor2s1 _48329_inst ( .DIN1(_47953), .DIN2(_47954), .Q(_47950) );
  nor2s1 _48330_inst ( .DIN1(_46996), .DIN2(_46962), .Q(_47954) );
  nnd2s1 _48331_inst ( .DIN1(_47955), .DIN2(_47717), .Q(_46962) );
  nor2s1 _48332_inst ( .DIN1(_37413), .DIN2(_47718), .Q(_47955) );
  nor2s1 _48333_inst ( .DIN1(_26361), .DIN2(_47512), .Q(_47953) );
  nnd2s1 _48334_inst ( .DIN1(_47946), .DIN2(_37414), .Q(_47512) );
  hi1s1 _48335_inst ( .DIN(_44202), .Q(_37414) );
  and2s1 _48336_inst ( .DIN1(_47956), .DIN2(_37129), .Q(_47946) );
  nor2s1 _48337_inst ( .DIN1(_45080), .DIN2(_38162), .Q(_47956) );
  nnd2s1 _48338_inst ( .DIN1(_47957), .DIN2(_47958), .Q(_47386) );
  nor2s1 _48339_inst ( .DIN1(_47959), .DIN2(_47960), .Q(_47958) );
  nnd2s1 _48340_inst ( .DIN1(_47088), .DIN2(_47006), .Q(_47960) );
  hi1s1 _48341_inst ( .DIN(_47653), .Q(_47006) );
  nor2s1 _48342_inst ( .DIN1(_47801), .DIN2(_47774), .Q(_47653) );
  nnd2s1 _48343_inst ( .DIN1(_47961), .DIN2(_37701), .Q(_47801) );
  nor2s1 _48344_inst ( .DIN1(_37963), .DIN2(_26361), .Q(_47961) );
  nnd2s1 _48345_inst ( .DIN1(_47719), .DIN2(_47239), .Q(_47088) );
  and2s1 _48346_inst ( .DIN1(_47962), .DIN2(_47940), .Q(_47719) );
  nor2s1 _48347_inst ( .DIN1(_47718), .DIN2(_39742), .Q(_47962) );
  nor2s1 _48348_inst ( .DIN1(_47963), .DIN2(_46973), .Q(_47959) );
  nor2s1 _48349_inst ( .DIN1(_47464), .DIN2(_47229), .Q(_47963) );
  and2s1 _48350_inst ( .DIN1(_47964), .DIN2(_38884), .Q(_47229) );
  hi1s1 _48351_inst ( .DIN(_39742), .Q(_38884) );
  nnd2s1 _48352_inst ( .DIN1(_47965), .DIN2(_2571), .Q(_39742) );
  nor2s1 _48353_inst ( .DIN1(_47966), .DIN2(_26358), .Q(_47965) );
  nor2s1 _48354_inst ( .DIN1(_47669), .DIN2(_47718), .Q(_47964) );
  nnd2s1 _48355_inst ( .DIN1(_47944), .DIN2(_47967), .Q(_47718) );
  hi1s1 _48356_inst ( .DIN(_47214), .Q(_47464) );
  nnd2s1 _48357_inst ( .DIN1(_47968), .DIN2(_37418), .Q(_47214) );
  nor2s1 _48358_inst ( .DIN1(_47969), .DIN2(_47758), .Q(_47957) );
  nnd2s1 _48359_inst ( .DIN1(_47210), .DIN2(_47970), .Q(_47758) );
  nnd2s1 _48360_inst ( .DIN1(_47413), .DIN2(_47289), .Q(_47970) );
  and2s1 _48361_inst ( .DIN1(_47971), .DIN2(_47940), .Q(_47413) );
  nor2s1 _48362_inst ( .DIN1(_37413), .DIN2(_47829), .Q(_47971) );
  nnd2s1 _48363_inst ( .DIN1(_47410), .DIN2(_47239), .Q(_47210) );
  hi1s1 _48364_inst ( .DIN(_47099), .Q(_47239) );
  and2s1 _48365_inst ( .DIN1(_47972), .DIN2(_37418), .Q(_47410) );
  hi1s1 _48366_inst ( .DIN(_40731), .Q(_37418) );
  nor2s1 _48367_inst ( .DIN1(_47669), .DIN2(_34484), .Q(_47972) );
  nnd2s1 _48368_inst ( .DIN1(_35342), .DIN2(_40119), .Q(_47669) );
  hi1s1 _48369_inst ( .DIN(_35369), .Q(_40119) );
  hi1s1 _48370_inst ( .DIN(_34215), .Q(_35342) );
  nor2s1 _48371_inst ( .DIN1(_46996), .DIN2(_47333), .Q(_47969) );
  nnd2s1 _48372_inst ( .DIN1(_47968), .DIN2(_43905), .Q(_47333) );
  hi1s1 _48373_inst ( .DIN(_47694), .Q(_43905) );
  nor2s1 _48374_inst ( .DIN1(_44319), .DIN2(_47973), .Q(_47968) );
  nor2s1 _48375_inst ( .DIN1(_47665), .DIN2(_47759), .Q(_47907) );
  nnd2s1 _48376_inst ( .DIN1(_47974), .DIN2(_47975), .Q(_47759) );
  nnd2s1 _48377_inst ( .DIN1(_47010), .DIN2(_47976), .Q(_47975) );
  nnd2s1 _48378_inst ( .DIN1(_47582), .DIN2(_47084), .Q(_47976) );
  nnd2s1 _48379_inst ( .DIN1(_47977), .DIN2(_47860), .Q(_47084) );
  nor2s1 _48380_inst ( .DIN1(_31291), .DIN2(_43602), .Q(_47977) );
  nnd2s1 _48381_inst ( .DIN1(_47978), .DIN2(_40867), .Q(_47582) );
  nor2s1 _48382_inst ( .DIN1(_47857), .DIN2(_47943), .Q(_47978) );
  nnd2s1 _48383_inst ( .DIN1(_47273), .DIN2(_47353), .Q(_47974) );
  hi1s1 _48384_inst ( .DIN(_46959), .Q(_47353) );
  nor2s1 _48385_inst ( .DIN1(_47887), .DIN2(_47754), .Q(_47273) );
  or2s1 _48386_inst ( .DIN1(_47786), .DIN2(_43906), .Q(_47754) );
  nnd2s1 _48387_inst ( .DIN1(_47979), .DIN2(_47980), .Q(_47665) );
  nor2s1 _48388_inst ( .DIN1(_46965), .DIN2(_47713), .Q(_47980) );
  and2s1 _48389_inst ( .DIN1(_47242), .DIN2(_47134), .Q(_47713) );
  and2s1 _48390_inst ( .DIN1(_47981), .DIN2(_37701), .Q(_47242) );
  hi1s1 _48391_inst ( .DIN(_39745), .Q(_37701) );
  nor2s1 _48392_inst ( .DIN1(_47973), .DIN2(_40731), .Q(_47981) );
  nnd2s1 _48393_inst ( .DIN1(_47982), .DIN2(_47944), .Q(_40731) );
  nor2s1 _48394_inst ( .DIN1(_2628), .DIN2(_26340), .Q(_47982) );
  hi1s1 _48395_inst ( .DIN(_47717), .Q(_47973) );
  nor2s1 _48396_inst ( .DIN1(_35994), .DIN2(_35369), .Q(_47717) );
  and2s1 _48397_inst ( .DIN1(_47983), .DIN2(_47772), .Q(_46965) );
  nor2s1 _48398_inst ( .DIN1(_26361), .DIN2(_47857), .Q(_47983) );
  nor2s1 _48399_inst ( .DIN1(_47550), .DIN2(_47984), .Q(_47979) );
  nor2s1 _48400_inst ( .DIN1(_47138), .DIN2(_46959), .Q(_47984) );
  nor2s1 _48401_inst ( .DIN1(_47095), .DIN2(_47297), .Q(_47138) );
  hi1s1 _48402_inst ( .DIN(_47433), .Q(_47297) );
  nnd2s1 _48403_inst ( .DIN1(_47985), .DIN2(_40867), .Q(_47433) );
  hi1s1 _48404_inst ( .DIN(_47202), .Q(_47095) );
  nnd2s1 _48405_inst ( .DIN1(_47986), .DIN2(_47987), .Q(_47202) );
  nor2s1 _48406_inst ( .DIN1(_35507), .DIN2(_37413), .Q(_47987) );
  hi1s1 _48407_inst ( .DIN(_34490), .Q(_37413) );
  nnd2s1 _48408_inst ( .DIN1(_47988), .DIN2(_2598), .Q(_35507) );
  nor2s1 _48409_inst ( .DIN1(_2599), .DIN2(_26246), .Q(_47988) );
  nor2s1 _48410_inst ( .DIN1(_35369), .DIN2(_47694), .Q(_47986) );
  nnd2s1 _48411_inst ( .DIN1(_47989), .DIN2(_2637), .Q(_35369) );
  nor2s1 _48412_inst ( .DIN1(_46997), .DIN2(_46961), .Q(_47550) );
  nnd2s1 _48413_inst ( .DIN1(_47990), .DIN2(_40867), .Q(_46997) );
  nor2s1 _48414_inst ( .DIN1(_47783), .DIN2(_43602), .Q(_47990) );
  nnd2s1 _48415_inst ( .DIN1(_47991), .DIN2(_47992), .Q(_47905) );
  nor2s1 _48416_inst ( .DIN1(_46985), .DIN2(_47016), .Q(_47992) );
  nnd2s1 _48417_inst ( .DIN1(_47993), .DIN2(_47188), .Q(_47016) );
  nnd2s1 _48418_inst ( .DIN1(_47264), .DIN2(_47026), .Q(_47188) );
  nnd2s1 _48419_inst ( .DIN1(_47040), .DIN2(_26361), .Q(_47026) );
  and2s1 _48420_inst ( .DIN1(_47893), .DIN2(_38714), .Q(_47264) );
  hi1s1 _48421_inst ( .DIN(_43602), .Q(_38714) );
  nor2s1 _48422_inst ( .DIN1(_46931), .DIN2(_47994), .Q(_47993) );
  nor2s1 _48423_inst ( .DIN1(_47213), .DIN2(_47279), .Q(_47994) );
  nnd2s1 _48424_inst ( .DIN1(_47995), .DIN2(_34490), .Q(_47279) );
  nor2s1 _48425_inst ( .DIN1(_47966), .DIN2(_47996), .Q(_34490) );
  nor2s1 _48426_inst ( .DIN1(_47079), .DIN2(_47045), .Q(_46931) );
  nnd2s1 _48427_inst ( .DIN1(_47997), .DIN2(_33182), .Q(_47045) );
  nor2s1 _48428_inst ( .DIN1(_47829), .DIN2(_47774), .Q(_47997) );
  hi1s1 _48429_inst ( .DIN(_47940), .Q(_47774) );
  nnd2s1 _48430_inst ( .DIN1(_47998), .DIN2(_2628), .Q(_47829) );
  nor2s1 _48431_inst ( .DIN1(_47900), .DIN2(_26340), .Q(_47998) );
  hi1s1 _48432_inst ( .DIN(_47583), .Q(_47079) );
  nnd2s1 _48433_inst ( .DIN1(_46959), .DIN2(_47044), .Q(_47583) );
  nnd2s1 _48434_inst ( .DIN1(_47999), .DIN2(_48000), .Q(_46985) );
  or2s1 _48435_inst ( .DIN1(_47158), .DIN2(_47040), .Q(_48000) );
  nnd2s1 _48436_inst ( .DIN1(_48001), .DIN2(_47903), .Q(_47158) );
  nor2s1 _48437_inst ( .DIN1(_31291), .DIN2(_47887), .Q(_48001) );
  nor2s1 _48438_inst ( .DIN1(_47105), .DIN2(_47377), .Q(_47999) );
  hi1s1 _48439_inst ( .DIN(_47083), .Q(_47377) );
  nnd2s1 _48440_inst ( .DIN1(_47658), .DIN2(_47134), .Q(_47083) );
  hi1s1 _48441_inst ( .DIN(_47040), .Q(_47134) );
  hi1s1 _48442_inst ( .DIN(_47517), .Q(_47658) );
  nnd2s1 _48443_inst ( .DIN1(_33182), .DIN2(_47995), .Q(_47517) );
  and2s1 _48444_inst ( .DIN1(_48002), .DIN2(_38165), .Q(_47995) );
  hi1s1 _48445_inst ( .DIN(_35368), .Q(_38165) );
  nor2s1 _48446_inst ( .DIN1(_37963), .DIN2(_34215), .Q(_48002) );
  hi1s1 _48447_inst ( .DIN(_34484), .Q(_33182) );
  nnd2s1 _48448_inst ( .DIN1(_48003), .DIN2(_2575), .Q(_34484) );
  and2s1 _48449_inst ( .DIN1(_47431), .DIN2(_47289), .Q(_47105) );
  and2s1 _48450_inst ( .DIN1(_48004), .DIN2(_40867), .Q(_47431) );
  hi1s1 _48451_inst ( .DIN(_48005), .Q(_40867) );
  nor2s1 _48452_inst ( .DIN1(_47783), .DIN2(_34485), .Q(_48004) );
  nnd2s1 _48453_inst ( .DIN1(_48006), .DIN2(_2575), .Q(_34485) );
  nor2s1 _48454_inst ( .DIN1(_26229), .DIN2(_47996), .Q(_48006) );
  nor2s1 _48455_inst ( .DIN1(_47250), .DIN2(_47317), .Q(_47991) );
  nnd2s1 _48456_inst ( .DIN1(_48007), .DIN2(_48008), .Q(_47317) );
  nor2s1 _48457_inst ( .DIN1(_48009), .DIN2(_48010), .Q(_48008) );
  nnd2s1 _48458_inst ( .DIN1(_48011), .DIN2(_48012), .Q(_48010) );
  nnd2s1 _48459_inst ( .DIN1(_47096), .DIN2(_48013), .Q(_48012) );
  nnd2s1 _48460_inst ( .DIN1(_47587), .DIN2(_46960), .Q(_48013) );
  or2s1 _48461_inst ( .DIN1(_47236), .DIN2(_47819), .Q(_46960) );
  hi1s1 _48462_inst ( .DIN(_47743), .Q(_47587) );
  nor2s1 _48463_inst ( .DIN1(_47640), .DIN2(_48014), .Q(_47743) );
  nnd2s1 _48464_inst ( .DIN1(_47288), .DIN2(_46956), .Q(_48011) );
  hi1s1 _48465_inst ( .DIN(_46996), .Q(_46956) );
  hi1s1 _48466_inst ( .DIN(_47112), .Q(_47288) );
  nnd2s1 _48467_inst ( .DIN1(_48015), .DIN2(_48016), .Q(_47112) );
  nnd2s1 _48468_inst ( .DIN1(_47272), .DIN2(_47629), .Q(_48009) );
  nnd2s1 _48469_inst ( .DIN1(_47145), .DIN2(_47228), .Q(_47629) );
  hi1s1 _48470_inst ( .DIN(_47476), .Q(_47145) );
  nnd2s1 _48471_inst ( .DIN1(_48017), .DIN2(_47765), .Q(_47476) );
  hi1s1 _48472_inst ( .DIN(_48018), .Q(_47765) );
  nor2s1 _48473_inst ( .DIN1(_26398), .DIN2(_48019), .Q(_48017) );
  nnd2s1 _48474_inst ( .DIN1(_47474), .DIN2(_47157), .Q(_47272) );
  hi1s1 _48475_inst ( .DIN(_47614), .Q(_47474) );
  nnd2s1 _48476_inst ( .DIN1(_48020), .DIN2(_48021), .Q(_47614) );
  nor2s1 _48477_inst ( .DIN1(_26398), .DIN2(_48018), .Q(_48020) );
  nor2s1 _48478_inst ( .DIN1(_46984), .DIN2(_48022), .Q(_48007) );
  nnd2s1 _48479_inst ( .DIN1(_48023), .DIN2(_48024), .Q(_48022) );
  nnd2s1 _48480_inst ( .DIN1(_47475), .DIN2(_47010), .Q(_48024) );
  nor2s1 _48481_inst ( .DIN1(_47744), .DIN2(_47236), .Q(_47475) );
  hi1s1 _48482_inst ( .DIN(_47635), .Q(_47236) );
  nor2s1 _48483_inst ( .DIN1(_47766), .DIN2(_48025), .Q(_47635) );
  hi1s1 _48484_inst ( .DIN(_46944), .Q(_48023) );
  nnd2s1 _48485_inst ( .DIN1(_48026), .DIN2(_48027), .Q(_46944) );
  nor2s1 _48486_inst ( .DIN1(_48028), .DIN2(_48029), .Q(_48027) );
  nor2s1 _48487_inst ( .DIN1(_46961), .DIN2(_47660), .Q(_48029) );
  nnd2s1 _48488_inst ( .DIN1(_48030), .DIN2(_48031), .Q(_47660) );
  and2s1 _48489_inst ( .DIN1(_47110), .DIN2(_47230), .Q(_48028) );
  nor2s1 _48490_inst ( .DIN1(_48014), .DIN2(_48032), .Q(_47110) );
  nnd2s1 _48491_inst ( .DIN1(_47709), .DIN2(_48033), .Q(_48014) );
  nor2s1 _48492_inst ( .DIN1(_47966), .DIN2(_47766), .Q(_47709) );
  nnd2s1 _48493_inst ( .DIN1(_2598), .DIN2(_48034), .Q(_47766) );
  nor2s1 _48494_inst ( .DIN1(_47815), .DIN2(_48035), .Q(_48026) );
  nor2s1 _48495_inst ( .DIN1(_47213), .DIN2(_47605), .Q(_48035) );
  nnd2s1 _48496_inst ( .DIN1(_48036), .DIN2(_48037), .Q(_47605) );
  nor2s1 _48497_inst ( .DIN1(_2598), .DIN2(_48038), .Q(_48037) );
  nor2s1 _48498_inst ( .DIN1(_48025), .DIN2(_47636), .Q(_48036) );
  nnd2s1 _48499_inst ( .DIN1(_48039), .DIN2(_48040), .Q(_47636) );
  nor2s1 _48500_inst ( .DIN1(_2624), .DIN2(_48041), .Q(_48040) );
  nor2s1 _48501_inst ( .DIN1(_26417), .DIN2(_47641), .Q(_48039) );
  hi1s1 _48502_inst ( .DIN(_47289), .Q(_47213) );
  nnd2s1 _48503_inst ( .DIN1(_46973), .DIN2(_46996), .Q(_47289) );
  nnd2s1 _48504_inst ( .DIN1(_48042), .DIN2(_47228), .Q(_46996) );
  nor2s1 _48505_inst ( .DIN1(_47643), .DIN2(_46968), .Q(_47815) );
  nnd2s1 _48506_inst ( .DIN1(_48021), .DIN2(_48030), .Q(_47643) );
  hi1s1 _48507_inst ( .DIN(_47818), .Q(_48021) );
  nnd2s1 _48508_inst ( .DIN1(_48043), .DIN2(_26229), .Q(_47818) );
  nnd2s1 _48509_inst ( .DIN1(_47649), .DIN2(_48044), .Q(_46984) );
  or2s1 _48510_inst ( .DIN1(_47044), .DIN2(_47355), .Q(_48044) );
  nnd2s1 _48511_inst ( .DIN1(_48003), .DIN2(_48030), .Q(_47355) );
  nor2s1 _48512_inst ( .DIN1(_48018), .DIN2(_2598), .Q(_48030) );
  nnd2s1 _48513_inst ( .DIN1(_48045), .DIN2(_48016), .Q(_48018) );
  hi1s1 _48514_inst ( .DIN(_47920), .Q(_48016) );
  nor2s1 _48515_inst ( .DIN1(_2575), .DIN2(_47919), .Q(_48045) );
  nor2s1 _48516_inst ( .DIN1(_26229), .DIN2(_48038), .Q(_48003) );
  hi1s1 _48517_inst ( .DIN(_47096), .Q(_47044) );
  nor2s1 _48518_inst ( .DIN1(_48046), .DIN2(_46961), .Q(_47096) );
  nnd2s1 _48519_inst ( .DIN1(_47113), .DIN2(_47228), .Q(_47649) );
  nor2s1 _48520_inst ( .DIN1(_48047), .DIN2(_47642), .Q(_47113) );
  or2s1 _48521_inst ( .DIN1(_48032), .DIN2(_47920), .Q(_48047) );
  nnd2s1 _48522_inst ( .DIN1(_48048), .DIN2(_48049), .Q(_47250) );
  nor2s1 _48523_inst ( .DIN1(_47069), .DIN2(_48050), .Q(_48049) );
  nnd2s1 _48524_inst ( .DIN1(_46942), .DIN2(_47724), .Q(_48050) );
  nnd2s1 _48525_inst ( .DIN1(_47516), .DIN2(_47157), .Q(_47724) );
  and2s1 _48526_inst ( .DIN1(_48051), .DIN2(_48052), .Q(_47516) );
  nor2s1 _48527_inst ( .DIN1(_34215), .DIN2(_35368), .Q(_48052) );
  nnd2s1 _48528_inst ( .DIN1(_48053), .DIN2(_26246), .Q(_34215) );
  nor2s1 _48529_inst ( .DIN1(_44319), .DIN2(_47694), .Q(_48051) );
  nnd2s1 _48530_inst ( .DIN1(_48054), .DIN2(_47944), .Q(_47694) );
  and2s1 _48531_inst ( .DIN1(_2625), .DIN2(_2624), .Q(_47944) );
  nor2s1 _48532_inst ( .DIN1(_26340), .DIN2(_26273), .Q(_48054) );
  nnd2s1 _48533_inst ( .DIN1(_48055), .DIN2(_2571), .Q(_44319) );
  nor2s1 _48534_inst ( .DIN1(_26358), .DIN2(_48025), .Q(_48055) );
  and2s1 _48535_inst ( .DIN1(_48056), .DIN2(_48057), .Q(_46942) );
  nnd2s1 _48536_inst ( .DIN1(_47985), .DIN2(_48058), .Q(_48057) );
  nor2s1 _48537_inst ( .DIN1(_47099), .DIN2(_43906), .Q(_48058) );
  nnd2s1 _48538_inst ( .DIN1(_48059), .DIN2(_2625), .Q(_43906) );
  nor2s1 _48539_inst ( .DIN1(_2624), .DIN2(_48060), .Q(_48059) );
  nnd2s1 _48540_inst ( .DIN1(_48061), .DIN2(_47228), .Q(_47099) );
  hi1s1 _48541_inst ( .DIN(_48062), .Q(_48061) );
  nor2s1 _48542_inst ( .DIN1(_47857), .DIN2(_47783), .Q(_47985) );
  nnd2s1 _48543_inst ( .DIN1(_35510), .DIN2(_29039), .Q(_47783) );
  hi1s1 _48544_inst ( .DIN(_33489), .Q(_29039) );
  nnd2s1 _48545_inst ( .DIN1(_48063), .DIN2(_47772), .Q(_48056) );
  hi1s1 _48546_inst ( .DIN(_47888), .Q(_47772) );
  nnd2s1 _48547_inst ( .DIN1(_48064), .DIN2(_38166), .Q(_47888) );
  nor2s1 _48548_inst ( .DIN1(_45080), .DIN2(_39462), .Q(_48064) );
  nor2s1 _48549_inst ( .DIN1(_46959), .DIN2(_43602), .Q(_48063) );
  nnd2s1 _48550_inst ( .DIN1(_48031), .DIN2(_2575), .Q(_43602) );
  nnd2s1 _48551_inst ( .DIN1(_48046), .DIN2(_47228), .Q(_46959) );
  nor2s1 _48552_inst ( .DIN1(_26771), .DIN2(______[6]), .Q(_48046) );
  nnd2s1 _48553_inst ( .DIN1(_48065), .DIN2(_48066), .Q(_47069) );
  nnd2s1 _48554_inst ( .DIN1(_48067), .DIN2(_48068), .Q(_48066) );
  nor2s1 _48555_inst ( .DIN1(_48069), .DIN2(_37963), .Q(_48068) );
  nnd2s1 _48556_inst ( .DIN1(_48070), .DIN2(_48071), .Q(_37963) );
  nor2s1 _48557_inst ( .DIN1(_2628), .DIN2(_26417), .Q(_48070) );
  nor2s1 _48558_inst ( .DIN1(_47933), .DIN2(_47940), .Q(_48069) );
  nor2s1 _48559_inst ( .DIN1(_35994), .DIN2(_38163), .Q(_47940) );
  nnd2s1 _48560_inst ( .DIN1(_48072), .DIN2(_2637), .Q(_38163) );
  nor2s1 _48561_inst ( .DIN1(_26216), .DIN2(_26310), .Q(_48072) );
  nor2s1 _48562_inst ( .DIN1(_35994), .DIN2(_35368), .Q(_47933) );
  nnd2s1 _48563_inst ( .DIN1(_48073), .DIN2(_2643), .Q(_35368) );
  nor2s1 _48564_inst ( .DIN1(_2637), .DIN2(_26216), .Q(_48073) );
  nnd2s1 _48565_inst ( .DIN1(_48074), .DIN2(_2599), .Q(_35994) );
  nor2s1 _48566_inst ( .DIN1(_26246), .DIN2(_26398), .Q(_48074) );
  nor2s1 _48567_inst ( .DIN1(_47040), .DIN2(_39745), .Q(_48067) );
  nnd2s1 _48568_inst ( .DIN1(_48075), .DIN2(_48076), .Q(_39745) );
  nor2s1 _48569_inst ( .DIN1(_26229), .DIN2(_26358), .Q(_48076) );
  nor2s1 _48570_inst ( .DIN1(_26567), .DIN2(_26247), .Q(_48075) );
  nnd2s1 _48571_inst ( .DIN1(_48077), .DIN2(_47228), .Q(_47040) );
  nnd2s1 _48572_inst ( .DIN1(_28646), .DIN2(_26772), .Q(_48077) );
  nnd2s1 _48573_inst ( .DIN1(_48078), .DIN2(_48079), .Q(_48065) );
  and2s1 _48574_inst ( .DIN1(_47010), .DIN2(_37129), .Q(_48079) );
  nor2s1 _48575_inst ( .DIN1(_48060), .DIN2(_47900), .Q(_37129) );
  hi1s1 _48576_inst ( .DIN(_26361), .Q(_47010) );
  nor2s1 _48577_inst ( .DIN1(_44202), .DIN2(_47871), .Q(_48078) );
  nnd2s1 _48578_inst ( .DIN1(_38166), .DIN2(_28178), .Q(_47871) );
  hi1s1 _48579_inst ( .DIN(_38162), .Q(_38166) );
  nnd2s1 _48580_inst ( .DIN1(_48080), .DIN2(_48081), .Q(_44202) );
  nor2s1 _48581_inst ( .DIN1(_26358), .DIN2(_26247), .Q(_48080) );
  nor2s1 _48582_inst ( .DIN1(_46981), .DIN2(_47318), .Q(_48048) );
  nnd2s1 _48583_inst ( .DIN1(_48082), .DIN2(_48083), .Q(_47318) );
  nnd2s1 _48584_inst ( .DIN1(_47504), .DIN2(_47230), .Q(_48083) );
  hi1s1 _48585_inst ( .DIN(_46973), .Q(_47230) );
  nor2s1 _48586_inst ( .DIN1(_47642), .DIN2(_47819), .Q(_47504) );
  or2s1 _48587_inst ( .DIN1(_47919), .DIN2(_47641), .Q(_47819) );
  or2s1 _48588_inst ( .DIN1(_47900), .DIN2(_48041), .Q(_47919) );
  nnd2s1 _48589_inst ( .DIN1(_2624), .DIN2(_26417), .Q(_47900) );
  nnd2s1 _48590_inst ( .DIN1(_47817), .DIN2(_48031), .Q(_47642) );
  hi1s1 _48591_inst ( .DIN(_48019), .Q(_48031) );
  nor2s1 _48592_inst ( .DIN1(_2598), .DIN2(_2575), .Q(_47817) );
  hi1s1 _48593_inst ( .DIN(_47624), .Q(_48082) );
  nnd2s1 _48594_inst ( .DIN1(_48084), .DIN2(_48085), .Q(_47624) );
  nnd2s1 _48595_inst ( .DIN1(_48086), .DIN2(_47228), .Q(_48085) );
  nnd2s1 _48596_inst ( .DIN1(_47056), .DIN2(_47043), .Q(_48086) );
  nnd2s1 _48597_inst ( .DIN1(_47934), .DIN2(_48087), .Q(_47043) );
  nor2s1 _48598_inst ( .DIN1(_48019), .DIN2(_48088), .Q(_48087) );
  nnd2s1 _48599_inst ( .DIN1(_2598), .DIN2(_26567), .Q(_48088) );
  nor2s1 _48600_inst ( .DIN1(_47641), .DIN2(_47640), .Q(_47934) );
  nnd2s1 _48601_inst ( .DIN1(_48015), .DIN2(_48033), .Q(_47056) );
  hi1s1 _48602_inst ( .DIN(_47641), .Q(_48033) );
  nnd2s1 _48603_inst ( .DIN1(_48089), .DIN2(_48090), .Q(_47641) );
  nor2s1 _48604_inst ( .DIN1(_26665), .DIN2(_48091), .Q(_48090) );
  nnd2s1 _48605_inst ( .DIN1(_26246), .DIN2(_26216), .Q(_48091) );
  nor2s1 _48606_inst ( .DIN1(_26310), .DIN2(_26573), .Q(_48089) );
  and2s1 _48607_inst ( .DIN1(_48092), .DIN2(_48093), .Q(_48015) );
  nor2s1 _48608_inst ( .DIN1(_2575), .DIN2(_26398), .Q(_48093) );
  nor2s1 _48609_inst ( .DIN1(_48019), .DIN2(_48032), .Q(_48092) );
  nnd2s1 _48610_inst ( .DIN1(_48094), .DIN2(_48071), .Q(_48032) );
  nor2s1 _48611_inst ( .DIN1(_2628), .DIN2(_2625), .Q(_48094) );
  nnd2s1 _48612_inst ( .DIN1(_48043), .DIN2(_2576), .Q(_48019) );
  nnd2s1 _48613_inst ( .DIN1(_47059), .DIN2(_47157), .Q(_48084) );
  hi1s1 _48614_inst ( .DIN(_46968), .Q(_47157) );
  nnd2s1 _48615_inst ( .DIN1(_48062), .DIN2(_47228), .Q(_46968) );
  nnd2s1 _48616_inst ( .DIN1(______[6]), .DIN2(_26772), .Q(_48062) );
  hi1s1 _48617_inst ( .DIN(_47706), .Q(_47059) );
  nnd2s1 _48618_inst ( .DIN1(_48095), .DIN2(_48096), .Q(_47706) );
  nor2s1 _48619_inst ( .DIN1(_2598), .DIN2(_47966), .Q(_48096) );
  nnd2s1 _48620_inst ( .DIN1(_2576), .DIN2(_26567), .Q(_47966) );
  nor2s1 _48621_inst ( .DIN1(_48038), .DIN2(_47744), .Q(_48095) );
  or2s1 _48622_inst ( .DIN1(_47640), .DIN2(_47920), .Q(_47744) );
  nnd2s1 _48623_inst ( .DIN1(_48097), .DIN2(_48098), .Q(_47920) );
  nor2s1 _48624_inst ( .DIN1(_2590), .DIN2(_48099), .Q(_48098) );
  nnd2s1 _48625_inst ( .DIN1(_26573), .DIN2(_26310), .Q(_48099) );
  nor2s1 _48626_inst ( .DIN1(_26665), .DIN2(_26216), .Q(_48097) );
  nnd2s1 _48627_inst ( .DIN1(_48100), .DIN2(_48071), .Q(_47640) );
  nor2s1 _48628_inst ( .DIN1(_26273), .DIN2(_26417), .Q(_48100) );
  nnd2s1 _48629_inst ( .DIN1(_48101), .DIN2(_48102), .Q(_46981) );
  or2s1 _48630_inst ( .DIN1(_47001), .DIN2(_46973), .Q(_48102) );
  nnd2s1 _48631_inst ( .DIN1(_48103), .DIN2(_47228), .Q(_46973) );
  hi1s1 _48632_inst ( .DIN(_48042), .Q(_48103) );
  nnd2s1 _48633_inst ( .DIN1(______[6]), .DIN2(______[16]), .Q(_48042) );
  nnd2s1 _48634_inst ( .DIN1(_47861), .DIN2(_48104), .Q(_47001) );
  nor2s1 _48635_inst ( .DIN1(_33489), .DIN2(_35993), .Q(_48104) );
  nnd2s1 _48636_inst ( .DIN1(_47989), .DIN2(_26573), .Q(_33489) );
  nor2s1 _48637_inst ( .DIN1(_2643), .DIN2(_2642), .Q(_47989) );
  nor2s1 _48638_inst ( .DIN1(_48005), .DIN2(_38713), .Q(_47861) );
  nnd2s1 _48639_inst ( .DIN1(_48081), .DIN2(_48105), .Q(_38713) );
  nnd2s1 _48640_inst ( .DIN1(_48106), .DIN2(_48071), .Q(_48005) );
  nor2s1 _48641_inst ( .DIN1(_26340), .DIN2(_2624), .Q(_48071) );
  nor2s1 _48642_inst ( .DIN1(_2625), .DIN2(_26273), .Q(_48106) );
  nor2s1 _48643_inst ( .DIN1(_47489), .DIN2(_48107), .Q(_48101) );
  nor2s1 _48644_inst ( .DIN1(_48108), .DIN2(_26361), .Q(_48107) );
  and2s1 _48645_inst ( .DIN1(_47868), .DIN2(_47346), .Q(_48108) );
  nnd2s1 _48646_inst ( .DIN1(_48109), .DIN2(_38853), .Q(_47346) );
  hi1s1 _48647_inst ( .DIN(_47887), .Q(_38853) );
  nnd2s1 _48648_inst ( .DIN1(_48043), .DIN2(_48110), .Q(_47887) );
  nor2s1 _48649_inst ( .DIN1(_26247), .DIN2(_53516), .Q(_48043) );
  nor2s1 _48650_inst ( .DIN1(_31291), .DIN2(_47786), .Q(_48109) );
  nnd2s1 _48651_inst ( .DIN1(_35370), .DIN2(_35510), .Q(_47786) );
  hi1s1 _48652_inst ( .DIN(_45080), .Q(_35510) );
  nnd2s1 _48653_inst ( .DIN1(_48053), .DIN2(_2590), .Q(_45080) );
  nor2s1 _48654_inst ( .DIN1(_2599), .DIN2(_2598), .Q(_48053) );
  nnd2s1 _48655_inst ( .DIN1(_48111), .DIN2(_47860), .Q(_47868) );
  hi1s1 _48656_inst ( .DIN(_47834), .Q(_47860) );
  nnd2s1 _48657_inst ( .DIN1(_35370), .DIN2(_28178), .Q(_47834) );
  hi1s1 _48658_inst ( .DIN(_34214), .Q(_28178) );
  nnd2s1 _48659_inst ( .DIN1(_48112), .DIN2(_2599), .Q(_34214) );
  nor2s1 _48660_inst ( .DIN1(_2598), .DIN2(_26246), .Q(_48112) );
  hi1s1 _48661_inst ( .DIN(_47892), .Q(_35370) );
  nnd2s1 _48662_inst ( .DIN1(_48113), .DIN2(_2637), .Q(_47892) );
  nor2s1 _48663_inst ( .DIN1(_2643), .DIN2(_26216), .Q(_48113) );
  nor2s1 _48664_inst ( .DIN1(_31291), .DIN2(_47857), .Q(_48111) );
  nnd2s1 _48665_inst ( .DIN1(_48081), .DIN2(_48034), .Q(_47857) );
  hi1s1 _48666_inst ( .DIN(_48038), .Q(_48034) );
  nnd2s1 _48667_inst ( .DIN1(_53516), .DIN2(_26247), .Q(_48038) );
  nor2s1 _48668_inst ( .DIN1(_2576), .DIN2(_2575), .Q(_48081) );
  nnd2s1 _48669_inst ( .DIN1(_48114), .DIN2(_47967), .Q(_31291) );
  hi1s1 _48670_inst ( .DIN(_48041), .Q(_47967) );
  nnd2s1 _48671_inst ( .DIN1(_26273), .DIN2(_26340), .Q(_48041) );
  and2s1 _48672_inst ( .DIN1(_47771), .DIN2(_47893), .Q(_47489) );
  nor2s1 _48673_inst ( .DIN1(_47943), .DIN2(_39462), .Q(_47893) );
  nnd2s1 _48674_inst ( .DIN1(_48114), .DIN2(_47945), .Q(_39462) );
  hi1s1 _48675_inst ( .DIN(_48060), .Q(_47945) );
  nnd2s1 _48676_inst ( .DIN1(_2628), .DIN2(_26340), .Q(_48060) );
  nor2s1 _48677_inst ( .DIN1(_2625), .DIN2(_2624), .Q(_48114) );
  hi1s1 _48678_inst ( .DIN(_47903), .Q(_47943) );
  nor2s1 _48679_inst ( .DIN1(_35993), .DIN2(_38162), .Q(_47903) );
  nnd2s1 _48680_inst ( .DIN1(_48115), .DIN2(_2643), .Q(_38162) );
  nor2s1 _48681_inst ( .DIN1(_2642), .DIN2(_2637), .Q(_48115) );
  nnd2s1 _48682_inst ( .DIN1(_48116), .DIN2(_2598), .Q(_35993) );
  nor2s1 _48683_inst ( .DIN1(_2599), .DIN2(_2590), .Q(_48116) );
  nor2s1 _48684_inst ( .DIN1(_30174), .DIN2(_26361), .Q(_47771) );
  nor2s1 _48685_inst ( .DIN1(______[6]), .DIN2(______[16]), .Q(_48117) );
  nnd2s1 _48686_inst ( .DIN1(_48110), .DIN2(_48105), .Q(_30174) );
  hi1s1 _48687_inst ( .DIN(_47996), .Q(_48105) );
  nnd2s1 _48688_inst ( .DIN1(_26247), .DIN2(_26358), .Q(_47996) );
  hi1s1 _48689_inst ( .DIN(_48025), .Q(_48110) );
  nnd2s1 _48690_inst ( .DIN1(_2575), .DIN2(_26229), .Q(_48025) );
  nnd2s1 _48691_inst ( .DIN1(_48118), .DIN2(_48119), .Q(____1___________[9])
         );
  nor2s1 _48692_inst ( .DIN1(_48120), .DIN2(_48121), .Q(_48119) );
  nnd2s1 _48693_inst ( .DIN1(_48122), .DIN2(_48123), .Q(_48121) );
  nnd2s1 _48694_inst ( .DIN1(_26768), .DIN2(_48124), .Q(_48123) );
  nnd2s1 _48695_inst ( .DIN1(_48125), .DIN2(_48126), .Q(_48124) );
  nor2s1 _48696_inst ( .DIN1(_48127), .DIN2(_48128), .Q(_48125) );
  nnd2s1 _48697_inst ( .DIN1(_48129), .DIN2(_48130), .Q(_48122) );
  nnd2s1 _48698_inst ( .DIN1(_48131), .DIN2(_48132), .Q(_48129) );
  nor2s1 _48699_inst ( .DIN1(_48133), .DIN2(_48134), .Q(_48131) );
  nnd2s1 _48700_inst ( .DIN1(_48135), .DIN2(_48136), .Q(_48120) );
  nnd2s1 _48701_inst ( .DIN1(_48137), .DIN2(_48138), .Q(_48136) );
  nnd2s1 _48702_inst ( .DIN1(_48139), .DIN2(_48140), .Q(_48138) );
  and2s1 _48703_inst ( .DIN1(_48141), .DIN2(_48142), .Q(_48135) );
  nor2s1 _48704_inst ( .DIN1(_48143), .DIN2(_48144), .Q(_48118) );
  or2s1 _48705_inst ( .DIN1(_48145), .DIN2(_48146), .Q(_48144) );
  nnd2s1 _48706_inst ( .DIN1(_48147), .DIN2(_48148), .Q(_48143) );
  nor2s1 _48707_inst ( .DIN1(_48149), .DIN2(_48150), .Q(_48147) );
  nnd2s1 _48708_inst ( .DIN1(_48151), .DIN2(_48152), .Q(____1___________[8])
         );
  nor2s1 _48709_inst ( .DIN1(_48153), .DIN2(_48154), .Q(_48152) );
  or2s1 _48710_inst ( .DIN1(_48155), .DIN2(_48150), .Q(_48154) );
  nnd2s1 _48711_inst ( .DIN1(_48156), .DIN2(_48157), .Q(_48150) );
  nor2s1 _48712_inst ( .DIN1(_48158), .DIN2(_48159), .Q(_48157) );
  nnd2s1 _48713_inst ( .DIN1(_48160), .DIN2(_48161), .Q(_48159) );
  nnd2s1 _48714_inst ( .DIN1(_48162), .DIN2(_48130), .Q(_48161) );
  nnd2s1 _48715_inst ( .DIN1(_48163), .DIN2(_48164), .Q(_48162) );
  and2s1 _48716_inst ( .DIN1(_48165), .DIN2(_48166), .Q(_48163) );
  nnd2s1 _48717_inst ( .DIN1(_48137), .DIN2(_48167), .Q(_48160) );
  nor2s1 _48718_inst ( .DIN1(_48168), .DIN2(_48169), .Q(_48156) );
  nnd2s1 _48719_inst ( .DIN1(_48170), .DIN2(_48171), .Q(_48153) );
  nnd2s1 _48720_inst ( .DIN1(_48172), .DIN2(_48173), .Q(_48171) );
  nnd2s1 _48721_inst ( .DIN1(_48174), .DIN2(_48175), .Q(_48172) );
  nor2s1 _48722_inst ( .DIN1(_48176), .DIN2(_48177), .Q(_48170) );
  nor2s1 _48723_inst ( .DIN1(_48178), .DIN2(_26783), .Q(_48177) );
  nor2s1 _48724_inst ( .DIN1(_48180), .DIN2(_48181), .Q(_48178) );
  nnd2s1 _48725_inst ( .DIN1(_48182), .DIN2(_48183), .Q(_48181) );
  nor2s1 _48726_inst ( .DIN1(_48134), .DIN2(_48184), .Q(_48183) );
  nor2s1 _48727_inst ( .DIN1(_48185), .DIN2(_48186), .Q(_48182) );
  nnd2s1 _48728_inst ( .DIN1(_48187), .DIN2(_48188), .Q(_48180) );
  nor2s1 _48729_inst ( .DIN1(_48189), .DIN2(_48190), .Q(_48188) );
  and2s1 _48730_inst ( .DIN1(_48191), .DIN2(_48192), .Q(_48187) );
  nor2s1 _48731_inst ( .DIN1(_48193), .DIN2(_48194), .Q(_48151) );
  nnd2s1 _48732_inst ( .DIN1(_48195), .DIN2(_48196), .Q(_48194) );
  nnd2s1 _48733_inst ( .DIN1(_48197), .DIN2(_48198), .Q(_48193) );
  hi1s1 _48734_inst ( .DIN(_48199), .Q(_48198) );
  nor2s1 _48735_inst ( .DIN1(_48200), .DIN2(_48201), .Q(_48197) );
  nnd2s1 _48736_inst ( .DIN1(_48202), .DIN2(_48203), .Q(____1___________[7])
         );
  nor2s1 _48737_inst ( .DIN1(_48204), .DIN2(_48205), .Q(_48203) );
  nnd2s1 _48738_inst ( .DIN1(_48206), .DIN2(_48207), .Q(_48205) );
  nor2s1 _48739_inst ( .DIN1(_48208), .DIN2(_48145), .Q(_48206) );
  nnd2s1 _48740_inst ( .DIN1(_48209), .DIN2(_48210), .Q(_48145) );
  nor2s1 _48741_inst ( .DIN1(_48211), .DIN2(_48212), .Q(_48210) );
  nnd2s1 _48742_inst ( .DIN1(_48213), .DIN2(_48214), .Q(_48212) );
  nnd2s1 _48743_inst ( .DIN1(_48215), .DIN2(_26769), .Q(_48214) );
  nor2s1 _48744_inst ( .DIN1(_48216), .DIN2(_48217), .Q(_48213) );
  nor2s1 _48745_inst ( .DIN1(_26844), .DIN2(_48219), .Q(_48217) );
  nor2s1 _48746_inst ( .DIN1(_48220), .DIN2(_48221), .Q(_48216) );
  nor2s1 _48747_inst ( .DIN1(_48222), .DIN2(_48223), .Q(_48221) );
  or2s1 _48748_inst ( .DIN1(_48224), .DIN2(_48225), .Q(_48223) );
  nnd2s1 _48749_inst ( .DIN1(_48226), .DIN2(_48175), .Q(_48222) );
  nnd2s1 _48750_inst ( .DIN1(_48227), .DIN2(_48228), .Q(_48211) );
  and2s1 _48751_inst ( .DIN1(_48229), .DIN2(_48230), .Q(_48228) );
  and2s1 _48752_inst ( .DIN1(_48231), .DIN2(_48232), .Q(_48227) );
  nor2s1 _48753_inst ( .DIN1(_48233), .DIN2(_48234), .Q(_48209) );
  nnd2s1 _48754_inst ( .DIN1(_48235), .DIN2(_48236), .Q(_48234) );
  nor2s1 _48755_inst ( .DIN1(_48237), .DIN2(_48238), .Q(_48235) );
  nnd2s1 _48756_inst ( .DIN1(_48239), .DIN2(_48240), .Q(_48233) );
  nor2s1 _48757_inst ( .DIN1(_48241), .DIN2(_48242), .Q(_48240) );
  nor2s1 _48758_inst ( .DIN1(_48243), .DIN2(_48244), .Q(_48239) );
  nor2s1 _48759_inst ( .DIN1(_48220), .DIN2(_48245), .Q(_48208) );
  nnd2s1 _48760_inst ( .DIN1(_48246), .DIN2(_48247), .Q(_48204) );
  nnd2s1 _48761_inst ( .DIN1(_26769), .DIN2(_48248), .Q(_48247) );
  nnd2s1 _48762_inst ( .DIN1(_48249), .DIN2(_48250), .Q(_48248) );
  nor2s1 _48763_inst ( .DIN1(_48251), .DIN2(_48252), .Q(_48250) );
  nnd2s1 _48764_inst ( .DIN1(_48253), .DIN2(_48254), .Q(_48252) );
  nor2s1 _48765_inst ( .DIN1(_48255), .DIN2(_48256), .Q(_48249) );
  nnd2s1 _48766_inst ( .DIN1(_48257), .DIN2(_48258), .Q(_48256) );
  hi1s1 _48767_inst ( .DIN(_48259), .Q(_48257) );
  nor2s1 _48768_inst ( .DIN1(_48260), .DIN2(_48261), .Q(_48246) );
  nor2s1 _48769_inst ( .DIN1(_48262), .DIN2(_26843), .Q(_48261) );
  nor2s1 _48770_inst ( .DIN1(_48263), .DIN2(_48264), .Q(_48262) );
  nnd2s1 _48771_inst ( .DIN1(_48265), .DIN2(_48165), .Q(_48264) );
  hi1s1 _48772_inst ( .DIN(_48266), .Q(_48260) );
  nor2s1 _48773_inst ( .DIN1(_48267), .DIN2(_48268), .Q(_48202) );
  or2s1 _48774_inst ( .DIN1(_48269), .DIN2(_48270), .Q(_48268) );
  nnd2s1 _48775_inst ( .DIN1(_48271), .DIN2(_48272), .Q(_48267) );
  nor2s1 _48776_inst ( .DIN1(_48273), .DIN2(_48274), .Q(_48271) );
  nnd2s1 _48777_inst ( .DIN1(_48275), .DIN2(_48276), .Q(____1___________[6])
         );
  nor2s1 _48778_inst ( .DIN1(_48277), .DIN2(_48278), .Q(_48276) );
  nnd2s1 _48779_inst ( .DIN1(_48279), .DIN2(_48280), .Q(_48278) );
  nor2s1 _48780_inst ( .DIN1(_48281), .DIN2(_48282), .Q(_48279) );
  nor2s1 _48781_inst ( .DIN1(_48220), .DIN2(_48283), .Q(_48282) );
  nor2s1 _48782_inst ( .DIN1(_48284), .DIN2(_39097), .Q(_48281) );
  nnd2s1 _48783_inst ( .DIN1(_48285), .DIN2(_48286), .Q(_48277) );
  nnd2s1 _48784_inst ( .DIN1(_26768), .DIN2(_48287), .Q(_48286) );
  nnd2s1 _48785_inst ( .DIN1(_48288), .DIN2(_48289), .Q(_48287) );
  nor2s1 _48786_inst ( .DIN1(_48290), .DIN2(_48291), .Q(_48289) );
  nor2s1 _48787_inst ( .DIN1(_48259), .DIN2(_48292), .Q(_48288) );
  nor2s1 _48788_inst ( .DIN1(_48293), .DIN2(_48294), .Q(_48285) );
  nor2s1 _48789_inst ( .DIN1(_48295), .DIN2(_26843), .Q(_48294) );
  nor2s1 _48790_inst ( .DIN1(_48296), .DIN2(_48297), .Q(_48295) );
  or2s1 _48791_inst ( .DIN1(_48186), .DIN2(_48184), .Q(_48297) );
  nnd2s1 _48792_inst ( .DIN1(_48140), .DIN2(_48298), .Q(_48296) );
  nor2s1 _48793_inst ( .DIN1(_48299), .DIN2(_48300), .Q(_48275) );
  nnd2s1 _48794_inst ( .DIN1(_48301), .DIN2(_48302), .Q(_48300) );
  nor2s1 _48795_inst ( .DIN1(_48303), .DIN2(_48304), .Q(_48301) );
  nnd2s1 _48796_inst ( .DIN1(_48305), .DIN2(_48306), .Q(_48299) );
  nor2s1 _48797_inst ( .DIN1(_48199), .DIN2(_48307), .Q(_48305) );
  nnd2s1 _48798_inst ( .DIN1(_48308), .DIN2(_48309), .Q(_48199) );
  nor2s1 _48799_inst ( .DIN1(_48310), .DIN2(_48311), .Q(_48309) );
  nor2s1 _48800_inst ( .DIN1(_34671), .DIN2(_48312), .Q(_48311) );
  nor2s1 _48801_inst ( .DIN1(_48313), .DIN2(_26844), .Q(_48310) );
  nor2s1 _48802_inst ( .DIN1(_48314), .DIN2(_48315), .Q(_48313) );
  nor2s1 _48803_inst ( .DIN1(_48316), .DIN2(_48317), .Q(_48314) );
  nor2s1 _48804_inst ( .DIN1(_48318), .DIN2(_48319), .Q(_48308) );
  nor2s1 _48805_inst ( .DIN1(_48220), .DIN2(_48320), .Q(_48318) );
  nnd2s1 _48806_inst ( .DIN1(_48321), .DIN2(_48322), .Q(____1___________[5])
         );
  nor2s1 _48807_inst ( .DIN1(_48323), .DIN2(_48324), .Q(_48322) );
  nnd2s1 _48808_inst ( .DIN1(_48148), .DIN2(_48325), .Q(_48324) );
  hi1s1 _48809_inst ( .DIN(_48241), .Q(_48325) );
  nnd2s1 _48810_inst ( .DIN1(_48326), .DIN2(_48327), .Q(_48241) );
  nor2s1 _48811_inst ( .DIN1(_48328), .DIN2(_48329), .Q(_48327) );
  or2s1 _48812_inst ( .DIN1(_48330), .DIN2(_48293), .Q(_48329) );
  hi1s1 _48813_inst ( .DIN(_48331), .Q(_48293) );
  nor2s1 _48814_inst ( .DIN1(_48332), .DIN2(_48333), .Q(_48328) );
  nor2s1 _48815_inst ( .DIN1(_48334), .DIN2(_48335), .Q(_48333) );
  nor2s1 _48816_inst ( .DIN1(_48336), .DIN2(_48337), .Q(_48326) );
  nnd2s1 _48817_inst ( .DIN1(_48338), .DIN2(_48339), .Q(_48337) );
  and2s1 _48818_inst ( .DIN1(_48340), .DIN2(_48341), .Q(_48148) );
  nor2s1 _48819_inst ( .DIN1(_48342), .DIN2(_48343), .Q(_48341) );
  nnd2s1 _48820_inst ( .DIN1(_48344), .DIN2(_48345), .Q(_48343) );
  nnd2s1 _48821_inst ( .DIN1(_48346), .DIN2(_48173), .Q(_48345) );
  nnd2s1 _48822_inst ( .DIN1(_48174), .DIN2(_48347), .Q(_48346) );
  nnd2s1 _48823_inst ( .DIN1(_48348), .DIN2(_48130), .Q(_48344) );
  nnd2s1 _48824_inst ( .DIN1(_48349), .DIN2(_48253), .Q(_48348) );
  hi1s1 _48825_inst ( .DIN(_48350), .Q(_48253) );
  nor2s1 _48826_inst ( .DIN1(_48351), .DIN2(_48352), .Q(_48340) );
  nnd2s1 _48827_inst ( .DIN1(_48353), .DIN2(_48354), .Q(_48323) );
  nnd2s1 _48828_inst ( .DIN1(_26769), .DIN2(_48355), .Q(_48354) );
  nnd2s1 _48829_inst ( .DIN1(_48356), .DIN2(_48357), .Q(_48355) );
  nor2s1 _48830_inst ( .DIN1(_48358), .DIN2(_48359), .Q(_48357) );
  nnd2s1 _48831_inst ( .DIN1(_48360), .DIN2(_48265), .Q(_48359) );
  hi1s1 _48832_inst ( .DIN(_48245), .Q(_48358) );
  nor2s1 _48833_inst ( .DIN1(_48361), .DIN2(_48362), .Q(_48356) );
  nor2s1 _48834_inst ( .DIN1(_48363), .DIN2(_48364), .Q(_48353) );
  nor2s1 _48835_inst ( .DIN1(_48365), .DIN2(_26844), .Q(_48364) );
  nor2s1 _48836_inst ( .DIN1(_48185), .DIN2(_48366), .Q(_48365) );
  nnd2s1 _48837_inst ( .DIN1(_48367), .DIN2(_48368), .Q(_48366) );
  nnd2s1 _48838_inst ( .DIN1(_48369), .DIN2(_48370), .Q(_48185) );
  nor2s1 _48839_inst ( .DIN1(_48332), .DIN2(_48371), .Q(_48363) );
  nor2s1 _48840_inst ( .DIN1(_48251), .DIN2(_48372), .Q(_48371) );
  nor2s1 _48841_inst ( .DIN1(_48373), .DIN2(_48374), .Q(_48321) );
  or2s1 _48842_inst ( .DIN1(_48375), .DIN2(_48376), .Q(_48374) );
  nnd2s1 _48843_inst ( .DIN1(_48377), .DIN2(_48272), .Q(_48373) );
  and2s1 _48844_inst ( .DIN1(_48378), .DIN2(_48379), .Q(_48272) );
  nnd2s1 _48845_inst ( .DIN1(_48380), .DIN2(_26768), .Q(_48379) );
  nor2s1 _48846_inst ( .DIN1(_48381), .DIN2(_48382), .Q(_48378) );
  nor2s1 _48847_inst ( .DIN1(_26843), .DIN2(_48383), .Q(_48382) );
  nnd2s1 _48848_inst ( .DIN1(_48384), .DIN2(_48385), .Q(____1___________[4])
         );
  nor2s1 _48849_inst ( .DIN1(_48386), .DIN2(_48387), .Q(_48385) );
  nnd2s1 _48850_inst ( .DIN1(_48388), .DIN2(_48389), .Q(_48387) );
  hi1s1 _48851_inst ( .DIN(_48242), .Q(_48389) );
  nnd2s1 _48852_inst ( .DIN1(_48390), .DIN2(_48391), .Q(_48242) );
  nnd2s1 _48853_inst ( .DIN1(_48392), .DIN2(_47729), .Q(_48391) );
  nnd2s1 _48854_inst ( .DIN1(_48315), .DIN2(_48173), .Q(_48390) );
  nor2s1 _48855_inst ( .DIN1(_48393), .DIN2(_48394), .Q(_48388) );
  nor2s1 _48856_inst ( .DIN1(_48395), .DIN2(_26783), .Q(_48393) );
  nor2s1 _48857_inst ( .DIN1(_48396), .DIN2(_48397), .Q(_48395) );
  nnd2s1 _48858_inst ( .DIN1(_48398), .DIN2(_48399), .Q(_48397) );
  nnd2s1 _48859_inst ( .DIN1(_48400), .DIN2(_48401), .Q(_48398) );
  nnd2s1 _48860_inst ( .DIN1(_48402), .DIN2(_48403), .Q(_48396) );
  nnd2s1 _48861_inst ( .DIN1(_48404), .DIN2(_48405), .Q(_48386) );
  nor2s1 _48862_inst ( .DIN1(_48406), .DIN2(_48407), .Q(_48405) );
  hi1s1 _48863_inst ( .DIN(_48408), .Q(_48406) );
  nor2s1 _48864_inst ( .DIN1(_48409), .DIN2(_48410), .Q(_48404) );
  nor2s1 _48865_inst ( .DIN1(_48411), .DIN2(_26844), .Q(_48410) );
  nor2s1 _48866_inst ( .DIN1(_48412), .DIN2(_48413), .Q(_48411) );
  nnd2s1 _48867_inst ( .DIN1(_48414), .DIN2(_48415), .Q(_48413) );
  nor2s1 _48868_inst ( .DIN1(_48416), .DIN2(_48417), .Q(_48384) );
  nnd2s1 _48869_inst ( .DIN1(_48418), .DIN2(_48419), .Q(_48417) );
  hi1s1 _48870_inst ( .DIN(_48420), .Q(_48419) );
  nor2s1 _48871_inst ( .DIN1(_48421), .DIN2(_48422), .Q(_48418) );
  nnd2s1 _48872_inst ( .DIN1(_48423), .DIN2(_48424), .Q(_48416) );
  nor2s1 _48873_inst ( .DIN1(_48351), .DIN2(_48200), .Q(_48424) );
  nnd2s1 _48874_inst ( .DIN1(_48142), .DIN2(_48425), .Q(_48200) );
  nnd2s1 _48875_inst ( .DIN1(_48426), .DIN2(_48427), .Q(_48351) );
  nnd2s1 _48876_inst ( .DIN1(_48255), .DIN2(_48173), .Q(_48427) );
  nor2s1 _48877_inst ( .DIN1(_48303), .DIN2(_48428), .Q(_48423) );
  nnd2s1 _48878_inst ( .DIN1(_48429), .DIN2(_48430), .Q(_48303) );
  nor2s1 _48879_inst ( .DIN1(_48431), .DIN2(_48432), .Q(_48430) );
  nnd2s1 _48880_inst ( .DIN1(_48433), .DIN2(_48434), .Q(_48432) );
  or2s1 _48881_inst ( .DIN1(_48370), .DIN2(_26806), .Q(_48434) );
  or2s1 _48882_inst ( .DIN1(_26783), .DIN2(_48435), .Q(_48433) );
  nnd2s1 _48883_inst ( .DIN1(_48436), .DIN2(_48437), .Q(_48431) );
  nnd2s1 _48884_inst ( .DIN1(_48137), .DIN2(_48438), .Q(_48437) );
  or2s1 _48885_inst ( .DIN1(_48167), .DIN2(_48439), .Q(_48438) );
  nnd2s1 _48886_inst ( .DIN1(_48440), .DIN2(_48441), .Q(_48167) );
  nnd2s1 _48887_inst ( .DIN1(_34673), .DIN2(_48442), .Q(_48441) );
  and2s1 _48888_inst ( .DIN1(_48443), .DIN2(_48232), .Q(_48436) );
  nor2s1 _48889_inst ( .DIN1(_48444), .DIN2(_48445), .Q(_48429) );
  or2s1 _48890_inst ( .DIN1(_48446), .DIN2(_48447), .Q(_48445) );
  or2s1 _48891_inst ( .DIN1(_48448), .DIN2(_48342), .Q(_48444) );
  nnd2s1 _48892_inst ( .DIN1(_48449), .DIN2(_48450), .Q(_48342) );
  nnd2s1 _48893_inst ( .DIN1(_48451), .DIN2(_48452), .Q(_48450) );
  nor2s1 _48894_inst ( .DIN1(_38283), .DIN2(_37533), .Q(_48451) );
  nnd2s1 _48895_inst ( .DIN1(_48453), .DIN2(_48137), .Q(_48449) );
  nnd2s1 _48896_inst ( .DIN1(_48454), .DIN2(_48455), .Q(____1___________[3])
         );
  nor2s1 _48897_inst ( .DIN1(_48456), .DIN2(_48457), .Q(_48455) );
  nnd2s1 _48898_inst ( .DIN1(_48458), .DIN2(_48426), .Q(_48457) );
  nnd2s1 _48899_inst ( .DIN1(_48459), .DIN2(_48130), .Q(_48426) );
  nor2s1 _48900_inst ( .DIN1(_48460), .DIN2(_48461), .Q(_48458) );
  nor2s1 _48901_inst ( .DIN1(_48462), .DIN2(_26783), .Q(_48461) );
  nor2s1 _48902_inst ( .DIN1(_48463), .DIN2(_48255), .Q(_48462) );
  nor2s1 _48903_inst ( .DIN1(_48464), .DIN2(_26843), .Q(_48460) );
  nor2s1 _48904_inst ( .DIN1(_48465), .DIN2(_48466), .Q(_48464) );
  nnd2s1 _48905_inst ( .DIN1(_48467), .DIN2(_48468), .Q(_48456) );
  nor2s1 _48906_inst ( .DIN1(_48469), .DIN2(_48470), .Q(_48467) );
  nor2s1 _48907_inst ( .DIN1(_48471), .DIN2(_48472), .Q(_48454) );
  or2s1 _48908_inst ( .DIN1(_48473), .DIN2(_48474), .Q(_48472) );
  nnd2s1 _48909_inst ( .DIN1(_48475), .DIN2(_48195), .Q(_48471) );
  and2s1 _48910_inst ( .DIN1(_48476), .DIN2(_48477), .Q(_48195) );
  nor2s1 _48911_inst ( .DIN1(_48478), .DIN2(_48479), .Q(_48477) );
  nnd2s1 _48912_inst ( .DIN1(_48480), .DIN2(_48481), .Q(_48479) );
  nnd2s1 _48913_inst ( .DIN1(_26768), .DIN2(_48482), .Q(_48481) );
  nnd2s1 _48914_inst ( .DIN1(_48483), .DIN2(_48126), .Q(_48482) );
  nor2s1 _48915_inst ( .DIN1(_48484), .DIN2(_48361), .Q(_48483) );
  nnd2s1 _48916_inst ( .DIN1(_48485), .DIN2(_48130), .Q(_48480) );
  nnd2s1 _48917_inst ( .DIN1(_48486), .DIN2(_48487), .Q(_48478) );
  nnd2s1 _48918_inst ( .DIN1(_48137), .DIN2(_48488), .Q(_48486) );
  nnd2s1 _48919_inst ( .DIN1(_48489), .DIN2(_48490), .Q(_48488) );
  nor2s1 _48920_inst ( .DIN1(_48491), .DIN2(_48350), .Q(_48489) );
  nor2s1 _48921_inst ( .DIN1(_48492), .DIN2(_48493), .Q(_48476) );
  nnd2s1 _48922_inst ( .DIN1(_48280), .DIN2(_48494), .Q(_48493) );
  hi1s1 _48923_inst ( .DIN(_48495), .Q(_48494) );
  and2s1 _48924_inst ( .DIN1(_48496), .DIN2(_48497), .Q(_48280) );
  nnd2s1 _48925_inst ( .DIN1(_48498), .DIN2(_48499), .Q(_48497) );
  nor2s1 _48926_inst ( .DIN1(_48332), .DIN2(_37555), .Q(_48498) );
  nnd2s1 _48927_inst ( .DIN1(_48500), .DIN2(_48501), .Q(_48492) );
  nnd2s1 _48928_inst ( .DIN1(_48392), .DIN2(_47930), .Q(_48501) );
  hi1s1 _48929_inst ( .DIN(_48502), .Q(_48392) );
  hi1s1 _48930_inst ( .DIN(_48503), .Q(_48500) );
  nor2s1 _48931_inst ( .DIN1(_48243), .DIN2(_48146), .Q(_48475) );
  nnd2s1 _48932_inst ( .DIN1(_48504), .DIN2(_48505), .Q(_48146) );
  nnd2s1 _48933_inst ( .DIN1(_48506), .DIN2(_48130), .Q(_48505) );
  nor2s1 _48934_inst ( .DIN1(_48507), .DIN2(_48508), .Q(_48504) );
  and2s1 _48935_inst ( .DIN1(_48292), .DIN2(_48137), .Q(_48508) );
  nnd2s1 _48936_inst ( .DIN1(_48360), .DIN2(_48509), .Q(_48292) );
  nnd2s1 _48937_inst ( .DIN1(_34677), .DIN2(_48499), .Q(_48509) );
  nnd2s1 _48938_inst ( .DIN1(_48510), .DIN2(_48511), .Q(_48243) );
  or2s1 _48939_inst ( .DIN1(_34671), .DIN2(_48284), .Q(_48511) );
  nor2s1 _48940_inst ( .DIN1(_48409), .DIN2(_48512), .Q(_48510) );
  nor2s1 _48941_inst ( .DIN1(_48513), .DIN2(_26844), .Q(_48512) );
  nor2s1 _48942_inst ( .DIN1(_48514), .DIN2(_48515), .Q(_48513) );
  nor2s1 _48943_inst ( .DIN1(_48284), .DIN2(_33614), .Q(_48409) );
  nnd2s1 _48944_inst ( .DIN1(_48516), .DIN2(_48517), .Q(____1___________[2])
         );
  nor2s1 _48945_inst ( .DIN1(_48518), .DIN2(_48519), .Q(_48517) );
  nnd2s1 _48946_inst ( .DIN1(_48520), .DIN2(_48196), .Q(_48519) );
  and2s1 _48947_inst ( .DIN1(_48521), .DIN2(_48522), .Q(_48196) );
  nor2s1 _48948_inst ( .DIN1(_48523), .DIN2(_48524), .Q(_48522) );
  nnd2s1 _48949_inst ( .DIN1(_48525), .DIN2(_48232), .Q(_48524) );
  nnd2s1 _48950_inst ( .DIN1(_48137), .DIN2(_48255), .Q(_48525) );
  nnd2s1 _48951_inst ( .DIN1(_48408), .DIN2(_48266), .Q(_48523) );
  nnd2s1 _48952_inst ( .DIN1(_48137), .DIN2(_48526), .Q(_48408) );
  nnd2s1 _48953_inst ( .DIN1(_48245), .DIN2(_48527), .Q(_48526) );
  nor2s1 _48954_inst ( .DIN1(_48528), .DIN2(_48529), .Q(_48521) );
  nnd2s1 _48955_inst ( .DIN1(_48530), .DIN2(_48531), .Q(_48529) );
  nnd2s1 _48956_inst ( .DIN1(_48532), .DIN2(_48173), .Q(_48531) );
  nnd2s1 _48957_inst ( .DIN1(_48533), .DIN2(_26769), .Q(_48530) );
  nor2s1 _48958_inst ( .DIN1(_48534), .DIN2(_48244), .Q(_48520) );
  nnd2s1 _48959_inst ( .DIN1(_48535), .DIN2(_48536), .Q(_48244) );
  and2s1 _48960_inst ( .DIN1(_48496), .DIN2(_48468), .Q(_48536) );
  nnd2s1 _48961_inst ( .DIN1(_48537), .DIN2(_48538), .Q(_48496) );
  nnd2s1 _48962_inst ( .DIN1(_48539), .DIN2(_48540), .Q(_48538) );
  nnd2s1 _48963_inst ( .DIN1(_36977), .DIN2(_48137), .Q(_48540) );
  nnd2s1 _48964_inst ( .DIN1(_48541), .DIN2(_26768), .Q(_48539) );
  nor2s1 _48965_inst ( .DIN1(_48542), .DIN2(_48543), .Q(_48535) );
  nor2s1 _48966_inst ( .DIN1(_48332), .DIN2(_48544), .Q(_48543) );
  nor2s1 _48967_inst ( .DIN1(_48412), .DIN2(_48545), .Q(_48544) );
  nor2s1 _48968_inst ( .DIN1(_48546), .DIN2(_48547), .Q(_48542) );
  nnd2s1 _48969_inst ( .DIN1(_26769), .DIN2(_48548), .Q(_48547) );
  nor2s1 _48970_inst ( .DIN1(_48549), .DIN2(_26783), .Q(_48534) );
  nor2s1 _48971_inst ( .DIN1(_48550), .DIN2(_48551), .Q(_48549) );
  nnd2s1 _48972_inst ( .DIN1(_48139), .DIN2(_48166), .Q(_48551) );
  nnd2s1 _48973_inst ( .DIN1(_48552), .DIN2(_48347), .Q(_48550) );
  nor2s1 _48974_inst ( .DIN1(_48553), .DIN2(_48459), .Q(_48552) );
  hi1s1 _48975_inst ( .DIN(_48554), .Q(_48459) );
  nnd2s1 _48976_inst ( .DIN1(_48555), .DIN2(_48556), .Q(_48518) );
  nnd2s1 _48977_inst ( .DIN1(_48557), .DIN2(_48130), .Q(_48556) );
  nnd2s1 _48978_inst ( .DIN1(_48558), .DIN2(_48367), .Q(_48557) );
  and2s1 _48979_inst ( .DIN1(_48414), .DIN2(_48265), .Q(_48558) );
  nor2s1 _48980_inst ( .DIN1(_48559), .DIN2(_48560), .Q(_48555) );
  nor2s1 _48981_inst ( .DIN1(_48561), .DIN2(_26843), .Q(_48560) );
  nor2s1 _48982_inst ( .DIN1(_48251), .DIN2(_48562), .Q(_48561) );
  hi1s1 _48983_inst ( .DIN(_48563), .Q(_48251) );
  hi1s1 _48984_inst ( .DIN(_48564), .Q(_48559) );
  nor2s1 _48985_inst ( .DIN1(_48565), .DIN2(_48566), .Q(_48516) );
  nnd2s1 _48986_inst ( .DIN1(_48567), .DIN2(_48568), .Q(_48566) );
  hi1s1 _48987_inst ( .DIN(_48569), .Q(_48567) );
  nnd2s1 _48988_inst ( .DIN1(_48570), .DIN2(_48571), .Q(_48565) );
  hi1s1 _48989_inst ( .DIN(_48421), .Q(_48571) );
  nnd2s1 _48990_inst ( .DIN1(_48572), .DIN2(_48573), .Q(_48421) );
  or2s1 _48991_inst ( .DIN1(_48174), .DIN2(_26783), .Q(_48573) );
  nor2s1 _48992_inst ( .DIN1(_48574), .DIN2(_48575), .Q(_48572) );
  nor2s1 _48993_inst ( .DIN1(_26843), .DIN2(_48576), .Q(_48575) );
  nor2s1 _48994_inst ( .DIN1(_48220), .DIN2(_48577), .Q(_48574) );
  nor2s1 _48995_inst ( .DIN1(_48270), .DIN2(_48376), .Q(_48570) );
  nnd2s1 _48996_inst ( .DIN1(_48578), .DIN2(_48579), .Q(_48376) );
  nor2s1 _48997_inst ( .DIN1(_48580), .DIN2(_48581), .Q(_48579) );
  nnd2s1 _48998_inst ( .DIN1(_48582), .DIN2(_48583), .Q(_48581) );
  and2s1 _48999_inst ( .DIN1(_48584), .DIN2(_48585), .Q(_48583) );
  nor2s1 _49000_inst ( .DIN1(_48507), .DIN2(_48586), .Q(_48582) );
  nor2s1 _49001_inst ( .DIN1(_48587), .DIN2(_48312), .Q(_48586) );
  nor2s1 _49002_inst ( .DIN1(_48588), .DIN2(_48589), .Q(_48587) );
  nnd2s1 _49003_inst ( .DIN1(_48590), .DIN2(_48591), .Q(_48580) );
  nor2s1 _49004_inst ( .DIN1(_48592), .DIN2(_48593), .Q(_48591) );
  hi1s1 _49005_inst ( .DIN(_48594), .Q(_48593) );
  nor2s1 _49006_inst ( .DIN1(_48595), .DIN2(_48596), .Q(_48590) );
  hi1s1 _49007_inst ( .DIN(_48597), .Q(_48595) );
  nor2s1 _49008_inst ( .DIN1(_48598), .DIN2(_48599), .Q(_48578) );
  nnd2s1 _49009_inst ( .DIN1(_48600), .DIN2(_48601), .Q(_48599) );
  nor2s1 _49010_inst ( .DIN1(_48201), .DIN2(_48428), .Q(_48600) );
  nnd2s1 _49011_inst ( .DIN1(_48602), .DIN2(_48603), .Q(_48428) );
  nor2s1 _49012_inst ( .DIN1(_48604), .DIN2(_48605), .Q(_48602) );
  nor2s1 _49013_inst ( .DIN1(_48332), .DIN2(_48606), .Q(_48605) );
  nor2s1 _49014_inst ( .DIN1(_26783), .DIN2(_48165), .Q(_48604) );
  nnd2s1 _49015_inst ( .DIN1(_48607), .DIN2(_48608), .Q(_48201) );
  nnd2s1 _49016_inst ( .DIN1(_48128), .DIN2(_48137), .Q(_48608) );
  nnd2s1 _49017_inst ( .DIN1(_48465), .DIN2(_48173), .Q(_48607) );
  nnd2s1 _49018_inst ( .DIN1(_48609), .DIN2(_48610), .Q(_48598) );
  nor2s1 _49019_inst ( .DIN1(_48611), .DIN2(_48612), .Q(_48610) );
  nor2s1 _49020_inst ( .DIN1(_48613), .DIN2(_26843), .Q(_48612) );
  nor2s1 _49021_inst ( .DIN1(_48614), .DIN2(_48615), .Q(_48613) );
  nnd2s1 _49022_inst ( .DIN1(_48435), .DIN2(_48616), .Q(_48615) );
  nor2s1 _49023_inst ( .DIN1(_48133), .DIN2(_46961), .Q(_48435) );
  hi1s1 _49024_inst ( .DIN(_48192), .Q(_48133) );
  nnd2s1 _49025_inst ( .DIN1(_48617), .DIN2(_48258), .Q(_48614) );
  nnd2s1 _49026_inst ( .DIN1(_48618), .DIN2(_48400), .Q(_48258) );
  nor2s1 _49027_inst ( .DIN1(_48619), .DIN2(_48620), .Q(_48617) );
  nor2s1 _49028_inst ( .DIN1(_48621), .DIN2(_26783), .Q(_48611) );
  nor2s1 _49029_inst ( .DIN1(_48622), .DIN2(_48623), .Q(_48621) );
  nnd2s1 _49030_inst ( .DIN1(_48415), .DIN2(_48624), .Q(_48623) );
  hi1s1 _49031_inst ( .DIN(_48625), .Q(_48622) );
  nor2s1 _49032_inst ( .DIN1(_48626), .DIN2(_48503), .Q(_48609) );
  nnd2s1 _49033_inst ( .DIN1(_48627), .DIN2(_48628), .Q(_48503) );
  nnd2s1 _49034_inst ( .DIN1(_48380), .DIN2(_48137), .Q(_48628) );
  hi1s1 _49035_inst ( .DIN(_48629), .Q(_48380) );
  nor2s1 _49036_inst ( .DIN1(_48220), .DIN2(_48630), .Q(_48626) );
  or2s1 _49037_inst ( .DIN1(_48631), .DIN2(_48307), .Q(_48270) );
  nnd2s1 _49038_inst ( .DIN1(_48632), .DIN2(_48633), .Q(_48307) );
  nnd2s1 _49039_inst ( .DIN1(_48634), .DIN2(_48130), .Q(_48633) );
  nnd2s1 _49040_inst ( .DIN1(_48189), .DIN2(_48137), .Q(_48632) );
  or2s1 _49041_inst ( .DIN1(_48635), .DIN2(_48636), .Q(_48631) );
  nor2s1 _49042_inst ( .DIN1(_48332), .DIN2(_48140), .Q(_48636) );
  nor2s1 _49043_inst ( .DIN1(_48637), .DIN2(_26843), .Q(_48635) );
  nor2s1 _49044_inst ( .DIN1(_48439), .DIN2(_48638), .Q(_48637) );
  hi1s1 _49045_inst ( .DIN(_48639), .Q(_48439) );
  nnd2s1 _49046_inst ( .DIN1(_48640), .DIN2(_48641), .Q(____1___________[1])
         );
  nor2s1 _49047_inst ( .DIN1(_48642), .DIN2(_48643), .Q(_48641) );
  nnd2s1 _49048_inst ( .DIN1(_48644), .DIN2(_48339), .Q(_48643) );
  and2s1 _49049_inst ( .DIN1(_48645), .DIN2(_48646), .Q(_48339) );
  nnd2s1 _49050_inst ( .DIN1(_48647), .DIN2(_48173), .Q(_48646) );
  nnd2s1 _49051_inst ( .DIN1(_48648), .DIN2(_48649), .Q(_48647) );
  nnd2s1 _49052_inst ( .DIN1(_48650), .DIN2(_48137), .Q(_48645) );
  hi1s1 _49053_inst ( .DIN(_48168), .Q(_48644) );
  nnd2s1 _49054_inst ( .DIN1(_48651), .DIN2(_48652), .Q(_48168) );
  or2s1 _49055_inst ( .DIN1(_48367), .DIN2(_26806), .Q(_48652) );
  nnd2s1 _49056_inst ( .DIN1(_48653), .DIN2(_48654), .Q(_48642) );
  nnd2s1 _49057_inst ( .DIN1(_26768), .DIN2(_48655), .Q(_48654) );
  nnd2s1 _49058_inst ( .DIN1(_48656), .DIN2(_48657), .Q(_48655) );
  hi1s1 _49059_inst ( .DIN(_48658), .Q(_48657) );
  nor2s1 _49060_inst ( .DIN1(_48532), .DIN2(_48659), .Q(_48656) );
  and2s1 _49061_inst ( .DIN1(_36977), .DIN2(_48537), .Q(_48659) );
  nor2s1 _49062_inst ( .DIN1(_48660), .DIN2(_48661), .Q(_48653) );
  nor2s1 _49063_inst ( .DIN1(_48662), .DIN2(_26844), .Q(_48661) );
  and2s1 _49064_inst ( .DIN1(_48132), .DIN2(_48663), .Q(_48662) );
  nor2s1 _49065_inst ( .DIN1(_48362), .DIN2(_48664), .Q(_48132) );
  hi1s1 _49066_inst ( .DIN(_48490), .Q(_48362) );
  nor2s1 _49067_inst ( .DIN1(_48665), .DIN2(_48666), .Q(_48640) );
  nnd2s1 _49068_inst ( .DIN1(_48667), .DIN2(_48668), .Q(_48666) );
  hi1s1 _49069_inst ( .DIN(_48669), .Q(_48668) );
  nnd2s1 _49070_inst ( .DIN1(_48670), .DIN2(_48671), .Q(_48665) );
  hi1s1 _49071_inst ( .DIN(_48672), .Q(_48671) );
  nor2s1 _49072_inst ( .DIN1(_48273), .DIN2(_48474), .Q(_48670) );
  nnd2s1 _49073_inst ( .DIN1(_48673), .DIN2(_48674), .Q(_48474) );
  nor2s1 _49074_inst ( .DIN1(_48675), .DIN2(_48676), .Q(_48674) );
  nnd2s1 _49075_inst ( .DIN1(_48677), .DIN2(_48678), .Q(_48676) );
  nnd2s1 _49076_inst ( .DIN1(_48679), .DIN2(_48173), .Q(_48678) );
  nnd2s1 _49077_inst ( .DIN1(_48245), .DIN2(_48283), .Q(_48679) );
  or2s1 _49078_inst ( .DIN1(_35696), .DIN2(_48680), .Q(_48677) );
  nnd2s1 _49079_inst ( .DIN1(_48564), .DIN2(_48597), .Q(_48675) );
  nnd2s1 _49080_inst ( .DIN1(_26769), .DIN2(_48681), .Q(_48597) );
  nnd2s1 _49081_inst ( .DIN1(_48254), .DIN2(_48226), .Q(_48681) );
  nnd2s1 _49082_inst ( .DIN1(_48291), .DIN2(_48130), .Q(_48564) );
  nor2s1 _49083_inst ( .DIN1(_48682), .DIN2(_48683), .Q(_48673) );
  nnd2s1 _49084_inst ( .DIN1(_48603), .DIN2(_48684), .Q(_48683) );
  or2s1 _49085_inst ( .DIN1(_48383), .DIN2(_26783), .Q(_48684) );
  nnd2s1 _49086_inst ( .DIN1(_48137), .DIN2(_48224), .Q(_48603) );
  nnd2s1 _49087_inst ( .DIN1(_48487), .DIN2(_48685), .Q(_48273) );
  or2s1 _49088_inst ( .DIN1(_48686), .DIN2(_26844), .Q(_48685) );
  nnd2s1 _49089_inst ( .DIN1(_48687), .DIN2(_48688), .Q(____1___________[11])
         );
  nor2s1 _49090_inst ( .DIN1(_48689), .DIN2(_48690), .Q(_48688) );
  nnd2s1 _49091_inst ( .DIN1(_48691), .DIN2(_48338), .Q(_48690) );
  and2s1 _49092_inst ( .DIN1(_48692), .DIN2(_48693), .Q(_48338) );
  nnd2s1 _49093_inst ( .DIN1(_48491), .DIN2(_26769), .Q(_48693) );
  nnd2s1 _49094_inst ( .DIN1(_48190), .DIN2(_48137), .Q(_48692) );
  nor2s1 _49095_inst ( .DIN1(_48694), .DIN2(_48695), .Q(_48691) );
  nor2s1 _49096_inst ( .DIN1(_47729), .DIN2(_48502), .Q(_48695) );
  hi1s1 _49097_inst ( .DIN(_47930), .Q(_47729) );
  nor2s1 _49098_inst ( .DIN1(_35781), .DIN2(_48680), .Q(_48694) );
  hi1s1 _49099_inst ( .DIN(_34673), .Q(_35781) );
  nnd2s1 _49100_inst ( .DIN1(_48696), .DIN2(_48697), .Q(_48689) );
  nnd2s1 _49101_inst ( .DIN1(_48137), .DIN2(_48698), .Q(_48697) );
  nnd2s1 _49102_inst ( .DIN1(_48699), .DIN2(_48139), .Q(_48698) );
  nor2s1 _49103_inst ( .DIN1(_48545), .DIN2(_48634), .Q(_48699) );
  hi1s1 _49104_inst ( .DIN(_48126), .Q(_48634) );
  nnd2s1 _49105_inst ( .DIN1(_48700), .DIN2(_34678), .Q(_48126) );
  nor2s1 _49106_inst ( .DIN1(_48596), .DIN2(_48701), .Q(_48696) );
  nor2s1 _49107_inst ( .DIN1(_48702), .DIN2(_26783), .Q(_48701) );
  nor2s1 _49108_inst ( .DIN1(_48703), .DIN2(_48263), .Q(_48702) );
  nnd2s1 _49109_inst ( .DIN1(_48349), .DIN2(_48606), .Q(_48263) );
  hi1s1 _49110_inst ( .DIN(_48134), .Q(_48606) );
  hi1s1 _49111_inst ( .DIN(_48704), .Q(_48703) );
  and2s1 _49112_inst ( .DIN1(_26768), .DIN2(_48705), .Q(_48596) );
  nnd2s1 _49113_inst ( .DIN1(_48191), .DIN2(_48706), .Q(_48705) );
  nor2s1 _49114_inst ( .DIN1(_48707), .DIN2(_48708), .Q(_48687) );
  nnd2s1 _49115_inst ( .DIN1(_48709), .DIN2(_48710), .Q(_48708) );
  nor2s1 _49116_inst ( .DIN1(_48569), .DIN2(_48672), .Q(_48709) );
  nnd2s1 _49117_inst ( .DIN1(_48711), .DIN2(_48712), .Q(_48672) );
  nor2s1 _49118_inst ( .DIN1(_48713), .DIN2(_48714), .Q(_48712) );
  nor2s1 _49119_inst ( .DIN1(_48715), .DIN2(_26843), .Q(_48714) );
  nor2s1 _49120_inst ( .DIN1(_48716), .DIN2(_48717), .Q(_48715) );
  nnd2s1 _49121_inst ( .DIN1(_47228), .DIN2(_48629), .Q(_48717) );
  hi1s1 _49122_inst ( .DIN(_48232), .Q(_48713) );
  nnd2s1 _49123_inst ( .DIN1(_48718), .DIN2(_48618), .Q(_48232) );
  nor2s1 _49124_inst ( .DIN1(_48332), .DIN2(_48719), .Q(_48718) );
  nor2s1 _49125_inst ( .DIN1(_48720), .DIN2(_48375), .Q(_48711) );
  nnd2s1 _49126_inst ( .DIN1(_48721), .DIN2(_48722), .Q(_48375) );
  nnd2s1 _49127_inst ( .DIN1(_48723), .DIN2(_48499), .Q(_48722) );
  nor2s1 _49128_inst ( .DIN1(_37555), .DIN2(_26844), .Q(_48723) );
  nnd2s1 _49129_inst ( .DIN1(_48485), .DIN2(_26768), .Q(_48721) );
  hi1s1 _49130_inst ( .DIN(_48140), .Q(_48485) );
  nnd2s1 _49131_inst ( .DIN1(_48589), .DIN2(_48499), .Q(_48140) );
  hi1s1 _49132_inst ( .DIN(_48546), .Q(_48499) );
  nor2s1 _49133_inst ( .DIN1(_48332), .DIN2(_48165), .Q(_48720) );
  or2s1 _49134_inst ( .DIN1(_48719), .DIN2(_48724), .Q(_48165) );
  nnd2s1 _49135_inst ( .DIN1(_48443), .DIN2(_48725), .Q(_48569) );
  or2s1 _49136_inst ( .DIN1(_39095), .DIN2(_48312), .Q(_48725) );
  nnd2s1 _49137_inst ( .DIN1(_48726), .DIN2(_48137), .Q(_48312) );
  nnd2s1 _49138_inst ( .DIN1(_48727), .DIN2(_48728), .Q(_48443) );
  nor2s1 _49139_inst ( .DIN1(_37550), .DIN2(_26783), .Q(_48728) );
  nnd2s1 _49140_inst ( .DIN1(_48729), .DIN2(_48730), .Q(_48707) );
  hi1s1 _49141_inst ( .DIN(_48422), .Q(_48730) );
  nnd2s1 _49142_inst ( .DIN1(_48731), .DIN2(_48732), .Q(_48422) );
  nor2s1 _49143_inst ( .DIN1(_48733), .DIN2(_48734), .Q(_48732) );
  nnd2s1 _49144_inst ( .DIN1(_48487), .DIN2(_48266), .Q(_48734) );
  nnd2s1 _49145_inst ( .DIN1(_48735), .DIN2(_35706), .Q(_48266) );
  nor2s1 _49146_inst ( .DIN1(_26843), .DIN2(_48546), .Q(_48735) );
  nnd2s1 _49147_inst ( .DIN1(_48619), .DIN2(_26769), .Q(_48487) );
  nor2s1 _49148_inst ( .DIN1(_48736), .DIN2(_26783), .Q(_48733) );
  and2s1 _49149_inst ( .DIN1(_48648), .DIN2(_48320), .Q(_48736) );
  nor2s1 _49150_inst ( .DIN1(_48737), .DIN2(_48738), .Q(_48731) );
  nor2s1 _49151_inst ( .DIN1(_48739), .DIN2(_26843), .Q(_48738) );
  nor2s1 _49152_inst ( .DIN1(_48740), .DIN2(_48741), .Q(_48739) );
  nnd2s1 _49153_inst ( .DIN1(_48367), .DIN2(_48630), .Q(_48741) );
  nnd2s1 _49154_inst ( .DIN1(_48742), .DIN2(_48649), .Q(_48740) );
  hi1s1 _49155_inst ( .DIN(_48650), .Q(_48742) );
  nor2s1 _49156_inst ( .DIN1(_48332), .DIN2(_48743), .Q(_48737) );
  nor2s1 _49157_inst ( .DIN1(_48334), .DIN2(_48350), .Q(_48743) );
  hi1s1 _49158_inst ( .DIN(_48744), .Q(_48334) );
  nor2s1 _49159_inst ( .DIN1(_48237), .DIN2(_48274), .Q(_48729) );
  nnd2s1 _49160_inst ( .DIN1(_48745), .DIN2(_48746), .Q(_48274) );
  nnd2s1 _49161_inst ( .DIN1(_48184), .DIN2(_26768), .Q(_48746) );
  nnd2s1 _49162_inst ( .DIN1(_48747), .DIN2(_48748), .Q(_48237) );
  or2s1 _49163_inst ( .DIN1(_48414), .DIN2(_26783), .Q(_48748) );
  nnd2s1 _49164_inst ( .DIN1(_48372), .DIN2(_48137), .Q(_48747) );
  nnd2s1 _49165_inst ( .DIN1(_48749), .DIN2(_48750), .Q(____1___________[10])
         );
  nor2s1 _49166_inst ( .DIN1(_48751), .DIN2(_48752), .Q(_48750) );
  nnd2s1 _49167_inst ( .DIN1(_48753), .DIN2(_48754), .Q(_48752) );
  hi1s1 _49168_inst ( .DIN(_48755), .Q(_48754) );
  nor2s1 _49169_inst ( .DIN1(_48495), .DIN2(_48319), .Q(_48753) );
  nnd2s1 _49170_inst ( .DIN1(_48756), .DIN2(_48229), .Q(_48319) );
  hi1s1 _49171_inst ( .DIN(_48660), .Q(_48229) );
  nor2s1 _49172_inst ( .DIN1(_48415), .DIN2(_48332), .Q(_48660) );
  nnd2s1 _49173_inst ( .DIN1(_48757), .DIN2(_48758), .Q(_48415) );
  nor2s1 _49174_inst ( .DIN1(_48759), .DIN2(_48760), .Q(_48758) );
  nor2s1 _49175_inst ( .DIN1(_48724), .DIN2(_48761), .Q(_48757) );
  nnd2s1 _49176_inst ( .DIN1(_26768), .DIN2(_48762), .Q(_48756) );
  nnd2s1 _49177_inst ( .DIN1(_48630), .DIN2(_48368), .Q(_48762) );
  nnd2s1 _49178_inst ( .DIN1(_48763), .DIN2(_48764), .Q(_48495) );
  nnd2s1 _49179_inst ( .DIN1(_46961), .DIN2(_48173), .Q(_48764) );
  nnd2s1 _49180_inst ( .DIN1(_48765), .DIN2(_39091), .Q(_47228) );
  nnd2s1 _49181_inst ( .DIN1(_48650), .DIN2(_26769), .Q(_48763) );
  nnd2s1 _49182_inst ( .DIN1(_48766), .DIN2(_48767), .Q(_48751) );
  nor2s1 _49183_inst ( .DIN1(_48768), .DIN2(_48769), .Q(_48767) );
  nor2s1 _49184_inst ( .DIN1(_48332), .DIN2(_48369), .Q(_48769) );
  hi1s1 _49185_inst ( .DIN(_48412), .Q(_48369) );
  hi1s1 _49186_inst ( .DIN(_48142), .Q(_48768) );
  nnd2s1 _49187_inst ( .DIN1(_48290), .DIN2(_48173), .Q(_48142) );
  hi1s1 _49188_inst ( .DIN(_48624), .Q(_48290) );
  nor2s1 _49189_inst ( .DIN1(_48770), .DIN2(_48771), .Q(_48766) );
  nor2s1 _49190_inst ( .DIN1(_26844), .DIN2(_48704), .Q(_48771) );
  nor2s1 _49191_inst ( .DIN1(_48220), .DIN2(_48298), .Q(_48770) );
  nor2s1 _49192_inst ( .DIN1(_48772), .DIN2(_48773), .Q(_48749) );
  nnd2s1 _49193_inst ( .DIN1(_48774), .DIN2(_48710), .Q(_48773) );
  and2s1 _49194_inst ( .DIN1(_48775), .DIN2(_48776), .Q(_48710) );
  nor2s1 _49195_inst ( .DIN1(_48777), .DIN2(_48778), .Q(_48776) );
  nnd2s1 _49196_inst ( .DIN1(_48779), .DIN2(_48780), .Q(_48778) );
  nnd2s1 _49197_inst ( .DIN1(_48137), .DIN2(_48781), .Q(_48780) );
  nnd2s1 _49198_inst ( .DIN1(_48782), .DIN2(_48783), .Q(_48781) );
  nor2s1 _49199_inst ( .DIN1(_48532), .DIN2(_48127), .Q(_48783) );
  hi1s1 _49200_inst ( .DIN(_48360), .Q(_48532) );
  nor2s1 _49201_inst ( .DIN1(_48186), .DIN2(_48506), .Q(_48782) );
  nnd2s1 _49202_inst ( .DIN1(_48399), .DIN2(_48784), .Q(_48186) );
  nor2s1 _49203_inst ( .DIN1(_48785), .DIN2(_48786), .Q(_48779) );
  nor2s1 _49204_inst ( .DIN1(_48787), .DIN2(_26783), .Q(_48786) );
  nor2s1 _49205_inst ( .DIN1(_48788), .DIN2(_48789), .Q(_48787) );
  nnd2s1 _49206_inst ( .DIN1(_48639), .DIN2(_48686), .Q(_48789) );
  nor2s1 _49207_inst ( .DIN1(_48790), .DIN2(_48791), .Q(_48785) );
  nnd2s1 _49208_inst ( .DIN1(_33611), .DIN2(_48541), .Q(_48791) );
  nnd2s1 _49209_inst ( .DIN1(_48792), .DIN2(_48425), .Q(_48777) );
  nnd2s1 _49210_inst ( .DIN1(_48638), .DIN2(_48130), .Q(_48425) );
  nor2s1 _49211_inst ( .DIN1(_48592), .DIN2(_48330), .Q(_48792) );
  nor2s1 _49212_inst ( .DIN1(_48793), .DIN2(_48794), .Q(_48775) );
  nnd2s1 _49213_inst ( .DIN1(_48795), .DIN2(_48568), .Q(_48794) );
  and2s1 _49214_inst ( .DIN1(_48796), .DIN2(_48797), .Q(_48568) );
  nnd2s1 _49215_inst ( .DIN1(_48137), .DIN2(_48798), .Q(_48797) );
  nnd2s1 _49216_inst ( .DIN1(_48283), .DIN2(_48799), .Q(_48798) );
  nnd2s1 _49217_inst ( .DIN1(_48620), .DIN2(_26768), .Q(_48796) );
  nor2s1 _49218_inst ( .DIN1(_48155), .DIN2(_48447), .Q(_48795) );
  nnd2s1 _49219_inst ( .DIN1(_48800), .DIN2(_48801), .Q(_48447) );
  nor2s1 _49220_inst ( .DIN1(_48802), .DIN2(_48803), .Q(_48801) );
  nnd2s1 _49221_inst ( .DIN1(_48468), .DIN2(_48231), .Q(_48803) );
  nnd2s1 _49222_inst ( .DIN1(_48804), .DIN2(_48137), .Q(_48468) );
  nor2s1 _49223_inst ( .DIN1(_48805), .DIN2(_38460), .Q(_48804) );
  nor2s1 _49224_inst ( .DIN1(_48806), .DIN2(_48807), .Q(_48805) );
  nor2s1 _49225_inst ( .DIN1(_42270), .DIN2(_39092), .Q(_48807) );
  nor2s1 _49226_inst ( .DIN1(_37533), .DIN2(_38279), .Q(_48806) );
  nor2s1 _49227_inst ( .DIN1(_26783), .DIN2(_48226), .Q(_48802) );
  nor2s1 _49228_inst ( .DIN1(_48169), .DIN2(_48808), .Q(_48800) );
  nnd2s1 _49229_inst ( .DIN1(_48809), .DIN2(_48810), .Q(_48808) );
  nnd2s1 _49230_inst ( .DIN1(_48463), .DIN2(_48137), .Q(_48810) );
  hi1s1 _49231_inst ( .DIN(_48811), .Q(_48809) );
  nnd2s1 _49232_inst ( .DIN1(_48812), .DIN2(_48813), .Q(_48169) );
  nnd2s1 _49233_inst ( .DIN1(_26769), .DIN2(_48814), .Q(_48813) );
  nnd2s1 _49234_inst ( .DIN1(_48815), .DIN2(_48219), .Q(_48814) );
  nnd2s1 _49235_inst ( .DIN1(_48361), .DIN2(_48137), .Q(_48812) );
  nnd2s1 _49236_inst ( .DIN1(_48816), .DIN2(_48817), .Q(_48155) );
  nnd2s1 _49237_inst ( .DIN1(_48818), .DIN2(_48137), .Q(_48817) );
  nnd2s1 _49238_inst ( .DIN1(_26768), .DIN2(_48224), .Q(_48816) );
  nnd2s1 _49239_inst ( .DIN1(_48819), .DIN2(_48820), .Q(_48793) );
  hi1s1 _49240_inst ( .DIN(_48821), .Q(_48820) );
  nor2s1 _49241_inst ( .DIN1(_48822), .DIN2(_48238), .Q(_48819) );
  nnd2s1 _49242_inst ( .DIN1(_48823), .DIN2(_48824), .Q(_48238) );
  nnd2s1 _49243_inst ( .DIN1(_48484), .DIN2(_26769), .Q(_48824) );
  nor2s1 _49244_inst ( .DIN1(_48825), .DIN2(_48826), .Q(_48823) );
  nor2s1 _49245_inst ( .DIN1(_48827), .DIN2(_48828), .Q(_48826) );
  nnd2s1 _49246_inst ( .DIN1(_34673), .DIN2(_35997), .Q(_48828) );
  hi1s1 _49247_inst ( .DIN(_38261), .Q(_35997) );
  hi1s1 _49248_inst ( .DIN(_48829), .Q(_48825) );
  nor2s1 _49249_inst ( .DIN1(_48830), .DIN2(_48332), .Q(_48822) );
  nor2s1 _49250_inst ( .DIN1(_48831), .DIN2(_48832), .Q(_48830) );
  or2s1 _49251_inst ( .DIN1(_48259), .DIN2(_48128), .Q(_48832) );
  nnd2s1 _49252_inst ( .DIN1(_48166), .DIN2(_48554), .Q(_48831) );
  nor2s1 _49253_inst ( .DIN1(_48473), .DIN2(_48669), .Q(_48774) );
  nnd2s1 _49254_inst ( .DIN1(_48833), .DIN2(_48601), .Q(_48669) );
  and2s1 _49255_inst ( .DIN1(_48502), .DIN2(_48230), .Q(_48601) );
  nnd2s1 _49256_inst ( .DIN1(_48834), .DIN2(_48400), .Q(_48230) );
  hi1s1 _49257_inst ( .DIN(_48317), .Q(_48400) );
  nor2s1 _49258_inst ( .DIN1(_48332), .DIN2(_48316), .Q(_48834) );
  nnd2s1 _49259_inst ( .DIN1(_48835), .DIN2(_48836), .Q(_48502) );
  nor2s1 _49260_inst ( .DIN1(_48332), .DIN2(_36022), .Q(_48836) );
  nor2s1 _49261_inst ( .DIN1(_34827), .DIN2(_33614), .Q(_48835) );
  nor2s1 _49262_inst ( .DIN1(_48837), .DIN2(_48838), .Q(_48833) );
  nor2s1 _49263_inst ( .DIN1(_26783), .DIN2(_48174), .Q(_48838) );
  nor2s1 _49264_inst ( .DIN1(_48839), .DIN2(_26844), .Q(_48837) );
  nnd2s1 _49265_inst ( .DIN1(_48840), .DIN2(_48377), .Q(_48473) );
  and2s1 _49266_inst ( .DIN1(_48841), .DIN2(_48842), .Q(_48377) );
  nnd2s1 _49267_inst ( .DIN1(_48716), .DIN2(_26768), .Q(_48842) );
  hi1s1 _49268_inst ( .DIN(_48175), .Q(_48716) );
  nor2s1 _49269_inst ( .DIN1(_48843), .DIN2(_48394), .Q(_48841) );
  nor2s1 _49270_inst ( .DIN1(_48220), .DIN2(_48139), .Q(_48394) );
  nor2s1 _49271_inst ( .DIN1(_48844), .DIN2(_26844), .Q(_48843) );
  nor2s1 _49272_inst ( .DIN1(_48553), .DIN2(_48184), .Q(_48844) );
  hi1s1 _49273_inst ( .DIN(_48577), .Q(_48184) );
  hi1s1 _49274_inst ( .DIN(_48320), .Q(_48553) );
  nor2s1 _49275_inst ( .DIN1(_48381), .DIN2(_48845), .Q(_48840) );
  nor2s1 _49276_inst ( .DIN1(_48846), .DIN2(_48332), .Q(_48845) );
  nor2s1 _49277_inst ( .DIN1(_48847), .DIN2(_48848), .Q(_48846) );
  nnd2s1 _49278_inst ( .DIN1(_48563), .DIN2(_48414), .Q(_48848) );
  nnd2s1 _49279_inst ( .DIN1(_48849), .DIN2(_39096), .Q(_48563) );
  nnd2s1 _49280_inst ( .DIN1(_48850), .DIN2(_48851), .Q(_48847) );
  nnd2s1 _49281_inst ( .DIN1(_48852), .DIN2(_27082), .Q(_48851) );
  nnd2s1 _49282_inst ( .DIN1(_48853), .DIN2(_48854), .Q(_48852) );
  nor2s1 _49283_inst ( .DIN1(_48619), .DIN2(_48855), .Q(_48854) );
  nnd2s1 _49284_inst ( .DIN1(_48815), .DIN2(_48349), .Q(_48855) );
  hi1s1 _49285_inst ( .DIN(_48533), .Q(_48349) );
  and2s1 _49286_inst ( .DIN1(_48856), .DIN2(_34678), .Q(_48619) );
  nor2s1 _49287_inst ( .DIN1(_34828), .DIN2(_41220), .Q(_48856) );
  nor2s1 _49288_inst ( .DIN1(_48620), .DIN2(_48788), .Q(_48853) );
  nnd2s1 _49289_inst ( .DIN1(_48383), .DIN2(_48857), .Q(_48788) );
  nnd2s1 _49290_inst ( .DIN1(_48588), .DIN2(_48726), .Q(_48857) );
  nnd2s1 _49291_inst ( .DIN1(_48765), .DIN2(_35700), .Q(_48383) );
  hi1s1 _49292_inst ( .DIN(_39095), .Q(_35700) );
  nnd2s1 _49293_inst ( .DIN1(______[24]), .DIN2(_48858), .Q(_48850) );
  nnd2s1 _49294_inst ( .DIN1(_48625), .DIN2(_48629), .Q(_48858) );
  nnd2s1 _49295_inst ( .DIN1(_34678), .DIN2(_48726), .Q(_48629) );
  and2s1 _49296_inst ( .DIN1(_48859), .DIN2(_34673), .Q(_48381) );
  nor2s1 _49297_inst ( .DIN1(_48220), .DIN2(_48860), .Q(_48859) );
  nnd2s1 _49298_inst ( .DIN1(_48861), .DIN2(_48862), .Q(_48772) );
  hi1s1 _49299_inst ( .DIN(_48863), .Q(_48862) );
  nor2s1 _49300_inst ( .DIN1(_48446), .DIN2(_48864), .Q(_48861) );
  hi1s1 _49301_inst ( .DIN(_48306), .Q(_48864) );
  nor2s1 _49302_inst ( .DIN1(_48528), .DIN2(_48865), .Q(_48306) );
  nor2s1 _49303_inst ( .DIN1(_48367), .DIN2(_26783), .Q(_48865) );
  nnd2s1 _49304_inst ( .DIN1(_48866), .DIN2(_48867), .Q(_48367) );
  nor2s1 _49305_inst ( .DIN1(_48868), .DIN2(_48316), .Q(_48866) );
  nnd2s1 _49306_inst ( .DIN1(_48869), .DIN2(_48870), .Q(_48528) );
  nnd2s1 _49307_inst ( .DIN1(_48664), .DIN2(_48130), .Q(_48870) );
  nor2s1 _49308_inst ( .DIN1(_48871), .DIN2(_48872), .Q(_48869) );
  nor2s1 _49309_inst ( .DIN1(_26844), .DIN2(_48648), .Q(_48872) );
  nnd2s1 _49310_inst ( .DIN1(_48873), .DIN2(_48401), .Q(_48648) );
  nor2s1 _49311_inst ( .DIN1(_48874), .DIN2(_48875), .Q(_48873) );
  nor2s1 _49312_inst ( .DIN1(_26783), .DIN2(_48649), .Q(_48871) );
  nnd2s1 _49313_inst ( .DIN1(_48876), .DIN2(_48867), .Q(_48649) );
  nor2s1 _49314_inst ( .DIN1(_48877), .DIN2(_48759), .Q(_48867) );
  nor2s1 _49315_inst ( .DIN1(_48868), .DIN2(_48724), .Q(_48876) );
  nnd2s1 _49316_inst ( .DIN1(_48878), .DIN2(_48879), .Q(_48446) );
  nor2s1 _49317_inst ( .DIN1(_48880), .DIN2(_48881), .Q(_48879) );
  nnd2s1 _49318_inst ( .DIN1(_48882), .DIN2(_48594), .Q(_48881) );
  hi1s1 _49319_inst ( .DIN(_48651), .Q(_48880) );
  nnd2s1 _49320_inst ( .DIN1(_48883), .DIN2(_48618), .Q(_48651) );
  nor2s1 _49321_inst ( .DIN1(_48332), .DIN2(_48317), .Q(_48883) );
  nor2s1 _49322_inst ( .DIN1(_48884), .DIN2(_48269), .Q(_48878) );
  nor2s1 _49323_inst ( .DIN1(_48220), .DIN2(_48885), .Q(_48884) );
  nnd2s1 _49324_inst ( .DIN1(_48886), .DIN2(_48887), .Q(____1___________[0])
         );
  nor2s1 _49325_inst ( .DIN1(_48888), .DIN2(_48889), .Q(_48887) );
  nnd2s1 _49326_inst ( .DIN1(_48890), .DIN2(_48891), .Q(_48889) );
  nnd2s1 _49327_inst ( .DIN1(_26769), .DIN2(_48892), .Q(_48891) );
  nnd2s1 _49328_inst ( .DIN1(_48893), .DIN2(_48894), .Q(_48892) );
  nor2s1 _49329_inst ( .DIN1(_48895), .DIN2(_48896), .Q(_48894) );
  nnd2s1 _49330_inst ( .DIN1(_48897), .DIN2(_48898), .Q(_48896) );
  nnd2s1 _49331_inst ( .DIN1(_48899), .DIN2(_36583), .Q(_48898) );
  nor2s1 _49332_inst ( .DIN1(_26331), .DIN2(_48860), .Q(_48899) );
  hi1s1 _49333_inst ( .DIN(_48442), .Q(_48860) );
  nnd2s1 _49334_inst ( .DIN1(_48537), .DIN2(_48900), .Q(_48897) );
  nnd2s1 _49335_inst ( .DIN1(_38279), .DIN2(_48901), .Q(_48900) );
  nnd2s1 _49336_inst ( .DIN1(_36977), .DIN2(_53517), .Q(_48901) );
  nor2s1 _49337_inst ( .DIN1(_31103), .DIN2(_37533), .Q(_48537) );
  nnd2s1 _49338_inst ( .DIN1(_48902), .DIN2(_48903), .Q(_48895) );
  nnd2s1 _49339_inst ( .DIN1(_48904), .DIN2(_48905), .Q(_48903) );
  nor2s1 _49340_inst ( .DIN1(_32015), .DIN2(_26481), .Q(_48905) );
  nor2s1 _49341_inst ( .DIN1(_48664), .DIN2(_48491), .Q(_48902) );
  hi1s1 _49342_inst ( .DIN(_48885), .Q(_48491) );
  nnd2s1 _49343_inst ( .DIN1(_48906), .DIN2(_36977), .Q(_48885) );
  nor2s1 _49344_inst ( .DIN1(_31103), .DIN2(_37557), .Q(_48906) );
  and2s1 _49345_inst ( .DIN1(_48401), .DIN2(_48907), .Q(_48664) );
  nnd2s1 _49346_inst ( .DIN1(_48908), .DIN2(_48909), .Q(_48907) );
  nnd2s1 _49347_inst ( .DIN1(_48910), .DIN2(_48911), .Q(_48909) );
  nor2s1 _49348_inst ( .DIN1(_48912), .DIN2(_48913), .Q(_48910) );
  or2s1 _49349_inst ( .DIN1(_48761), .DIN2(_48874), .Q(_48908) );
  nor2s1 _49350_inst ( .DIN1(_48914), .DIN2(_48915), .Q(_48893) );
  nnd2s1 _49351_inst ( .DIN1(_48916), .DIN2(_48839), .Q(_48915) );
  nor2s1 _49352_inst ( .DIN1(_48134), .DIN2(_48315), .Q(_48839) );
  hi1s1 _49353_inst ( .DIN(_48706), .Q(_48315) );
  nnd2s1 _49354_inst ( .DIN1(_48917), .DIN2(_48401), .Q(_48706) );
  hi1s1 _49355_inst ( .DIN(_48316), .Q(_48401) );
  nor2s1 _49356_inst ( .DIN1(_48875), .DIN2(_48918), .Q(_48917) );
  nor2s1 _49357_inst ( .DIN1(_48919), .DIN2(_48316), .Q(_48134) );
  hi1s1 _49358_inst ( .DIN(_48920), .Q(_48916) );
  nnd2s1 _49359_inst ( .DIN1(_48663), .DIN2(_48616), .Q(_48914) );
  and2s1 _49360_inst ( .DIN1(_48921), .DIN2(_48815), .Q(_48616) );
  nnd2s1 _49361_inst ( .DIN1(_48922), .DIN2(_36977), .Q(_48815) );
  nor2s1 _49362_inst ( .DIN1(_32015), .DIN2(_37557), .Q(_48922) );
  nor2s1 _49363_inst ( .DIN1(_48923), .DIN2(_48515), .Q(_48921) );
  nor2s1 _49364_inst ( .DIN1(_34672), .DIN2(_48924), .Q(_48515) );
  nor2s1 _49365_inst ( .DIN1(_48255), .DIN2(_48412), .Q(_48663) );
  nor2s1 _49366_inst ( .DIN1(_48919), .DIN2(_48724), .Q(_48412) );
  nnd2s1 _49367_inst ( .DIN1(_48704), .DIN2(_48298), .Q(_48255) );
  nnd2s1 _49368_inst ( .DIN1(_48925), .DIN2(_48926), .Q(_48298) );
  nor2s1 _49369_inst ( .DIN1(_48875), .DIN2(_48927), .Q(_48925) );
  nnd2s1 _49370_inst ( .DIN1(_48928), .DIN2(_48929), .Q(_48704) );
  nor2s1 _49371_inst ( .DIN1(_48930), .DIN2(_48913), .Q(_48928) );
  nor2s1 _49372_inst ( .DIN1(_48931), .DIN2(_48932), .Q(_48890) );
  nor2s1 _49373_inst ( .DIN1(_48220), .DIN2(_48933), .Q(_48932) );
  nor2s1 _49374_inst ( .DIN1(_48934), .DIN2(_48935), .Q(_48933) );
  nnd2s1 _49375_inst ( .DIN1(_48936), .DIN2(_48360), .Q(_48935) );
  nnd2s1 _49376_inst ( .DIN1(_48727), .DIN2(_34678), .Q(_48360) );
  nnd2s1 _49377_inst ( .DIN1(_48937), .DIN2(_36586), .Q(_48936) );
  nnd2s1 _49378_inst ( .DIN1(_48938), .DIN2(_48226), .Q(_48934) );
  nnd2s1 _49379_inst ( .DIN1(_48939), .DIN2(_34399), .Q(_48226) );
  nor2s1 _49380_inst ( .DIN1(_48940), .DIN2(_48453), .Q(_48938) );
  and2s1 _49381_inst ( .DIN1(_48941), .DIN2(_36583), .Q(_48453) );
  hi1s1 _49382_inst ( .DIN(_48219), .Q(_48940) );
  nnd2s1 _49383_inst ( .DIN1(_48942), .DIN2(_35755), .Q(_48219) );
  nor2s1 _49384_inst ( .DIN1(_48332), .DIN2(_48943), .Q(_48931) );
  nor2s1 _49385_inst ( .DIN1(_48335), .DIN2(_48259), .Q(_48943) );
  nnd2s1 _49386_inst ( .DIN1(_48490), .DIN2(_48164), .Q(_48259) );
  nnd2s1 _49387_inst ( .DIN1(_34399), .DIN2(_48442), .Q(_48164) );
  nnd2s1 _49388_inst ( .DIN1(_48941), .DIN2(_48944), .Q(_48490) );
  nor2s1 _49389_inst ( .DIN1(_38460), .DIN2(_42209), .Q(_48941) );
  hi1s1 _49390_inst ( .DIN(_48399), .Q(_48335) );
  nnd2s1 _49391_inst ( .DIN1(_48945), .DIN2(_38071), .Q(_48399) );
  hi1s1 _49392_inst ( .DIN(_48946), .Q(_38071) );
  nor2s1 _49393_inst ( .DIN1(_32015), .DIN2(_36611), .Q(_48945) );
  nnd2s1 _49394_inst ( .DIN1(_48947), .DIN2(_48948), .Q(_48888) );
  nor2s1 _49395_inst ( .DIN1(_48176), .DIN2(_48949), .Q(_48948) );
  nor2s1 _49396_inst ( .DIN1(_48680), .DIN2(_48950), .Q(_48949) );
  nnd2s1 _49397_inst ( .DIN1(_36586), .DIN2(_53108), .Q(_48950) );
  hi1s1 _49398_inst ( .DIN(_37533), .Q(_36586) );
  hi1s1 _49399_inst ( .DIN(_48882), .Q(_48176) );
  nnd2s1 _49400_inst ( .DIN1(_48514), .DIN2(_26769), .Q(_48882) );
  and2s1 _49401_inst ( .DIN1(_48951), .DIN2(_34673), .Q(_48514) );
  nor2s1 _49402_inst ( .DIN1(_48952), .DIN2(_48953), .Q(_48947) );
  nor2s1 _49403_inst ( .DIN1(_48954), .DIN2(_26843), .Q(_48953) );
  nor2s1 _49404_inst ( .DIN1(_48955), .DIN2(_48658), .Q(_48954) );
  nnd2s1 _49405_inst ( .DIN1(_48956), .DIN2(_48957), .Q(_48658) );
  nor2s1 _49406_inst ( .DIN1(_48350), .DIN2(_48361), .Q(_48957) );
  and2s1 _49407_inst ( .DIN1(_48958), .DIN2(_48589), .Q(_48361) );
  nor2s1 _49408_inst ( .DIN1(_34827), .DIN2(_41221), .Q(_48958) );
  nor2s1 _49409_inst ( .DIN1(_48959), .DIN2(_48874), .Q(_48350) );
  nor2s1 _49410_inst ( .DIN1(_48225), .DIN2(_48466), .Q(_48956) );
  nnd2s1 _49411_inst ( .DIN1(_48744), .DIN2(_48624), .Q(_48466) );
  nnd2s1 _49412_inst ( .DIN1(_48960), .DIN2(_48926), .Q(_48624) );
  nor2s1 _49413_inst ( .DIN1(_48761), .DIN2(_48961), .Q(_48960) );
  nnd2s1 _49414_inst ( .DIN1(_48962), .DIN2(_48963), .Q(_48744) );
  nor2s1 _49415_inst ( .DIN1(_48759), .DIN2(_48927), .Q(_48962) );
  nnd2s1 _49416_inst ( .DIN1(_48320), .DIN2(_48630), .Q(_48225) );
  or2s1 _49417_inst ( .DIN1(_48317), .DIN2(_48961), .Q(_48630) );
  nnd2s1 _49418_inst ( .DIN1(_48964), .DIN2(_48965), .Q(_48317) );
  nor2s1 _49419_inst ( .DIN1(_48877), .DIN2(_48966), .Q(_48965) );
  nnd2s1 _49420_inst ( .DIN1(_26430), .DIN2(_26278), .Q(_48966) );
  nor2s1 _49421_inst ( .DIN1(_48759), .DIN2(_26633), .Q(_48964) );
  nnd2s1 _49422_inst ( .DIN1(_48967), .DIN2(_48618), .Q(_48320) );
  hi1s1 _49423_inst ( .DIN(_48927), .Q(_48618) );
  nor2s1 _49424_inst ( .DIN1(_48874), .DIN2(_48761), .Q(_48967) );
  nor2s1 _49425_inst ( .DIN1(_48924), .DIN2(_34396), .Q(_48955) );
  nor2s1 _49426_inst ( .DIN1(_48968), .DIN2(_39092), .Q(_48952) );
  nor2s1 _49427_inst ( .DIN1(_48969), .DIN2(_48970), .Q(_48968) );
  nor2s1 _49428_inst ( .DIN1(_42270), .DIN2(_48790), .Q(_48970) );
  nor2s1 _49429_inst ( .DIN1(_38283), .DIN2(_48827), .Q(_48969) );
  nor2s1 _49430_inst ( .DIN1(_48971), .DIN2(_48972), .Q(_48886) );
  nnd2s1 _49431_inst ( .DIN1(_48973), .DIN2(_48667), .Q(_48972) );
  and2s1 _49432_inst ( .DIN1(_48974), .DIN2(_48975), .Q(_48667) );
  nor2s1 _49433_inst ( .DIN1(_48976), .DIN2(_48977), .Q(_48975) );
  nnd2s1 _49434_inst ( .DIN1(_48978), .DIN2(_48979), .Q(_48977) );
  nnd2s1 _49435_inst ( .DIN1(_48980), .DIN2(_48173), .Q(_48979) );
  nnd2s1 _49436_inst ( .DIN1(_48981), .DIN2(_48577), .Q(_48980) );
  nnd2s1 _49437_inst ( .DIN1(_48588), .DIN2(_48982), .Q(_48577) );
  hi1s1 _49438_inst ( .DIN(_39097), .Q(_48588) );
  nnd2s1 _49439_inst ( .DIN1(_48983), .DIN2(_48984), .Q(_39097) );
  nor2s1 _49440_inst ( .DIN1(_48215), .DIN2(_48463), .Q(_48981) );
  hi1s1 _49441_inst ( .DIN(_48347), .Q(_48463) );
  nnd2s1 _49442_inst ( .DIN1(_48985), .DIN2(_39096), .Q(_48347) );
  nor2s1 _49443_inst ( .DIN1(_32015), .DIN2(_42270), .Q(_48985) );
  hi1s1 _49444_inst ( .DIN(_48799), .Q(_48215) );
  nnd2s1 _49445_inst ( .DIN1(_48986), .DIN2(_34678), .Q(_48799) );
  nor2s1 _49446_inst ( .DIN1(_38284), .DIN2(_34827), .Q(_48986) );
  nnd2s1 _49447_inst ( .DIN1(_26768), .DIN2(_48506), .Q(_48978) );
  nnd2s1 _49448_inst ( .DIN1(_48265), .DIN2(_48370), .Q(_48506) );
  nnd2s1 _49449_inst ( .DIN1(_48987), .DIN2(_39078), .Q(_48370) );
  nnd2s1 _49450_inst ( .DIN1(_48988), .DIN2(_38072), .Q(_48265) );
  nor2s1 _49451_inst ( .DIN1(_38460), .DIN2(_37557), .Q(_48988) );
  nnd2s1 _49452_inst ( .DIN1(_48989), .DIN2(_48585), .Q(_48976) );
  nnd2s1 _49453_inst ( .DIN1(_48990), .DIN2(_34677), .Q(_48585) );
  nor2s1 _49454_inst ( .DIN1(_48332), .DIN2(_48546), .Q(_48990) );
  nnd2s1 _49455_inst ( .DIN1(_48137), .DIN2(_48991), .Q(_48989) );
  nnd2s1 _49456_inst ( .DIN1(_48992), .DIN2(_48414), .Q(_48991) );
  nnd2s1 _49457_inst ( .DIN1(_48939), .DIN2(_36583), .Q(_48414) );
  nor2s1 _49458_inst ( .DIN1(_38460), .DIN2(_48946), .Q(_48939) );
  nor2s1 _49459_inst ( .DIN1(_48304), .DIN2(_48993), .Q(_48974) );
  nnd2s1 _49460_inst ( .DIN1(_48207), .DIN2(_48236), .Q(_48993) );
  and2s1 _49461_inst ( .DIN1(_48994), .DIN2(_48995), .Q(_48236) );
  nnd2s1 _49462_inst ( .DIN1(_48996), .DIN2(_48997), .Q(_48995) );
  nor2s1 _49463_inst ( .DIN1(_48332), .DIN2(_38460), .Q(_48997) );
  nor2s1 _49464_inst ( .DIN1(_42209), .DIN2(_36611), .Q(_48996) );
  nnd2s1 _49465_inst ( .DIN1(_48727), .DIN2(_48998), .Q(_48994) );
  nor2s1 _49466_inst ( .DIN1(_37550), .DIN2(_26843), .Q(_48998) );
  nor2s1 _49467_inst ( .DIN1(_41221), .DIN2(_34828), .Q(_48727) );
  and2s1 _49468_inst ( .DIN1(_48999), .DIN2(_49000), .Q(_48207) );
  nnd2s1 _49469_inst ( .DIN1(_48128), .DIN2(_48130), .Q(_49000) );
  nor2s1 _49470_inst ( .DIN1(_33613), .DIN2(_48546), .Q(_48128) );
  hi1s1 _49471_inst ( .DIN(_34678), .Q(_33613) );
  nor2s1 _49472_inst ( .DIN1(_49001), .DIN2(_48912), .Q(_34678) );
  nnd2s1 _49473_inst ( .DIN1(_26324), .DIN2(_38028), .Q(_49001) );
  nnd2s1 _49474_inst ( .DIN1(_48127), .DIN2(_48173), .Q(_48999) );
  hi1s1 _49475_inst ( .DIN(_48527), .Q(_48127) );
  nnd2s1 _49476_inst ( .DIN1(_49002), .DIN2(_38486), .Q(_48527) );
  nor2s1 _49477_inst ( .DIN1(_36022), .DIN2(_37555), .Q(_49002) );
  nnd2s1 _49478_inst ( .DIN1(_49003), .DIN2(_49004), .Q(_48304) );
  nnd2s1 _49479_inst ( .DIN1(_48484), .DIN2(_48173), .Q(_49004) );
  hi1s1 _49480_inst ( .DIN(_48576), .Q(_48484) );
  nnd2s1 _49481_inst ( .DIN1(_49005), .DIN2(_34669), .Q(_48576) );
  nor2s1 _49482_inst ( .DIN1(_39417), .DIN2(_41221), .Q(_49005) );
  nnd2s1 _49483_inst ( .DIN1(_49006), .DIN2(_2472), .Q(_41221) );
  nor2s1 _49484_inst ( .DIN1(_2473), .DIN2(_49007), .Q(_49006) );
  nor2s1 _49485_inst ( .DIN1(_48592), .DIN2(_49008), .Q(_49003) );
  nor2s1 _49486_inst ( .DIN1(_49009), .DIN2(_26783), .Q(_49008) );
  nor2s1 _49487_inst ( .DIN1(_48620), .DIN2(_49010), .Q(_49009) );
  hi1s1 _49488_inst ( .DIN(_48139), .Q(_49010) );
  nnd2s1 _49489_inst ( .DIN1(_36587), .DIN2(_48442), .Q(_48139) );
  hi1s1 _49490_inst ( .DIN(_39092), .Q(_36587) );
  and2s1 _49491_inst ( .DIN1(_48982), .DIN2(_39091), .Q(_48620) );
  hi1s1 _49492_inst ( .DIN(_37550), .Q(_39091) );
  nnd2s1 _49493_inst ( .DIN1(_49011), .DIN2(_49012), .Q(_37550) );
  nor2s1 _49494_inst ( .DIN1(_2429), .DIN2(_49013), .Q(_49011) );
  and2s1 _49495_inst ( .DIN1(_49014), .DIN2(_48726), .Q(_48592) );
  nor2s1 _49496_inst ( .DIN1(_48220), .DIN2(_33614), .Q(_49014) );
  nor2s1 _49497_inst ( .DIN1(_48420), .DIN2(_48682), .Q(_48973) );
  nnd2s1 _49498_inst ( .DIN1(_49015), .DIN2(_49016), .Q(_48682) );
  nor2s1 _49499_inst ( .DIN1(_49017), .DIN2(_49018), .Q(_49016) );
  nnd2s1 _49500_inst ( .DIN1(_48231), .DIN2(_48829), .Q(_49018) );
  nnd2s1 _49501_inst ( .DIN1(_49019), .DIN2(_48442), .Q(_48829) );
  nor2s1 _49502_inst ( .DIN1(_26783), .DIN2(_37533), .Q(_49019) );
  nnd2s1 _49503_inst ( .DIN1(_48137), .DIN2(_48923), .Q(_48231) );
  and2s1 _49504_inst ( .DIN1(_49020), .DIN2(_35617), .Q(_48923) );
  nor2s1 _49505_inst ( .DIN1(_38283), .DIN2(_35784), .Q(_49020) );
  nnd2s1 _49506_inst ( .DIN1(_48983), .DIN2(_38028), .Q(_35784) );
  nnd2s1 _49507_inst ( .DIN1(_48331), .DIN2(_48594), .Q(_49017) );
  nnd2s1 _49508_inst ( .DIN1(_49021), .DIN2(_48452), .Q(_48594) );
  hi1s1 _49509_inst ( .DIN(_48790), .Q(_48452) );
  nnd2s1 _49510_inst ( .DIN1(_35617), .DIN2(_26768), .Q(_48790) );
  nor2s1 _49511_inst ( .DIN1(_42270), .DIN2(_34396), .Q(_49021) );
  hi1s1 _49512_inst ( .DIN(_39078), .Q(_34396) );
  nor2s1 _49513_inst ( .DIN1(_48874), .DIN2(_26324), .Q(_39078) );
  nnd2s1 _49514_inst ( .DIN1(_49012), .DIN2(_49022), .Q(_48874) );
  nnd2s1 _49515_inst ( .DIN1(_48137), .DIN2(_49023), .Q(_48331) );
  nnd2s1 _49516_inst ( .DIN1(_48191), .DIN2(_48625), .Q(_49023) );
  nnd2s1 _49517_inst ( .DIN1(_49024), .DIN2(_48944), .Q(_48625) );
  hi1s1 _49518_inst ( .DIN(_35758), .Q(_48944) );
  nnd2s1 _49519_inst ( .DIN1(_49025), .DIN2(_49012), .Q(_35758) );
  nor2s1 _49520_inst ( .DIN1(_2429), .DIN2(_48759), .Q(_49025) );
  nor2s1 _49521_inst ( .DIN1(_32015), .DIN2(_48946), .Q(_49024) );
  nnd2s1 _49522_inst ( .DIN1(_49026), .DIN2(_49027), .Q(_48946) );
  nnd2s1 _49523_inst ( .DIN1(_48765), .DIN2(_34669), .Q(_48191) );
  nor2s1 _49524_inst ( .DIN1(_38284), .DIN2(_39417), .Q(_48765) );
  nor2s1 _49525_inst ( .DIN1(_48352), .DIN2(_49028), .Q(_49015) );
  nnd2s1 _49526_inst ( .DIN1(_49029), .DIN2(_49030), .Q(_49028) );
  nnd2s1 _49527_inst ( .DIN1(_49031), .DIN2(_48130), .Q(_49030) );
  nnd2s1 _49528_inst ( .DIN1(_48166), .DIN2(_48192), .Q(_49031) );
  nnd2s1 _49529_inst ( .DIN1(_49032), .DIN2(_35755), .Q(_48192) );
  hi1s1 _49530_inst ( .DIN(_35785), .Q(_35755) );
  nnd2s1 _49531_inst ( .DIN1(_49033), .DIN2(_36583), .Q(_48166) );
  hi1s1 _49532_inst ( .DIN(_37557), .Q(_36583) );
  nor2s1 _49533_inst ( .DIN1(_32015), .DIN2(_38261), .Q(_49033) );
  nnd2s1 _49534_inst ( .DIN1(_48218), .DIN2(_48920), .Q(_49029) );
  nnd2s1 _49535_inst ( .DIN1(_48440), .DIN2(_49034), .Q(_48920) );
  nnd2s1 _49536_inst ( .DIN1(_49032), .DIN2(_34673), .Q(_49034) );
  nor2s1 _49537_inst ( .DIN1(_49013), .DIN2(_48877), .Q(_34673) );
  nor2s1 _49538_inst ( .DIN1(_31103), .DIN2(_38261), .Q(_49032) );
  nnd2s1 _49539_inst ( .DIN1(_48951), .DIN2(_33611), .Q(_48440) );
  nor2s1 _49540_inst ( .DIN1(_32015), .DIN2(_38283), .Q(_48951) );
  nnd2s1 _49541_inst ( .DIN1(_49035), .DIN2(_49036), .Q(_48352) );
  nor2s1 _49542_inst ( .DIN1(_48407), .DIN2(_49037), .Q(_49036) );
  nor2s1 _49543_inst ( .DIN1(_48220), .DIN2(_48639), .Q(_49037) );
  nnd2s1 _49544_inst ( .DIN1(_49038), .DIN2(_37556), .Q(_48639) );
  nor2s1 _49545_inst ( .DIN1(_32015), .DIN2(_36021), .Q(_49038) );
  and2s1 _49546_inst ( .DIN1(_48904), .DIN2(_49039), .Q(_48407) );
  nor2s1 _49547_inst ( .DIN1(_32015), .DIN2(_26844), .Q(_49039) );
  nor2s1 _49548_inst ( .DIN1(_38261), .DIN2(_35695), .Q(_48904) );
  nor2s1 _49549_inst ( .DIN1(_48821), .DIN2(_48811), .Q(_49035) );
  nnd2s1 _49550_inst ( .DIN1(_49040), .DIN2(_49041), .Q(_48811) );
  nnd2s1 _49551_inst ( .DIN1(_49042), .DIN2(_27937), .Q(_49041) );
  nor2s1 _49552_inst ( .DIN1(_48827), .DIN2(_42270), .Q(_49042) );
  hi1s1 _49553_inst ( .DIN(_49043), .Q(_48827) );
  nnd2s1 _49554_inst ( .DIN1(_49044), .DIN2(_35706), .Q(_49040) );
  nor2s1 _49555_inst ( .DIN1(_26783), .DIN2(_48546), .Q(_49044) );
  nnd2s1 _49556_inst ( .DIN1(_38031), .DIN2(_38486), .Q(_48546) );
  hi1s1 _49557_inst ( .DIN(_41220), .Q(_38031) );
  nnd2s1 _49558_inst ( .DIN1(_49045), .DIN2(_49046), .Q(_48821) );
  nnd2s1 _49559_inst ( .DIN1(_49047), .DIN2(_49048), .Q(_49046) );
  nor2s1 _49560_inst ( .DIN1(_26783), .DIN2(_38283), .Q(_49048) );
  nor2s1 _49561_inst ( .DIN1(_31103), .DIN2(_39092), .Q(_49047) );
  nnd2s1 _49562_inst ( .DIN1(_49049), .DIN2(_49050), .Q(_39092) );
  nor2s1 _49563_inst ( .DIN1(_2429), .DIN2(_49051), .Q(_49049) );
  nnd2s1 _49564_inst ( .DIN1(_49052), .DIN2(_49043), .Q(_49045) );
  nor2s1 _49565_inst ( .DIN1(_31103), .DIN2(_26844), .Q(_49043) );
  nor2s1 _49566_inst ( .DIN1(_49053), .DIN2(_37533), .Q(_49052) );
  nnd2s1 _49567_inst ( .DIN1(_38027), .DIN2(_49022), .Q(_37533) );
  nor2s1 _49568_inst ( .DIN1(_38072), .DIN2(_48541), .Q(_49053) );
  hi1s1 _49569_inst ( .DIN(_42209), .Q(_48541) );
  hi1s1 _49570_inst ( .DIN(_38279), .Q(_38072) );
  nnd2s1 _49571_inst ( .DIN1(_49054), .DIN2(_49055), .Q(_38279) );
  nnd2s1 _49572_inst ( .DIN1(_49056), .DIN2(_49057), .Q(_48420) );
  nor2s1 _49573_inst ( .DIN1(_49058), .DIN2(_48158), .Q(_49057) );
  nor2s1 _49574_inst ( .DIN1(_26783), .DIN2(_48283), .Q(_48158) );
  nnd2s1 _49575_inst ( .DIN1(_48982), .DIN2(_48589), .Q(_48283) );
  nor2s1 _49576_inst ( .DIN1(_48332), .DIN2(_49059), .Q(_49058) );
  nor2s1 _49577_inst ( .DIN1(_48545), .DIN2(_48533), .Q(_49059) );
  nor2s1 _49578_inst ( .DIN1(_48719), .DIN2(_48316), .Q(_48533) );
  nnd2s1 _49579_inst ( .DIN1(_49026), .DIN2(_49055), .Q(_48316) );
  nor2s1 _49580_inst ( .DIN1(_53518), .DIN2(_26580), .Q(_49026) );
  or2s1 _49581_inst ( .DIN1(_48761), .DIN2(_48918), .Q(_48719) );
  nnd2s1 _49582_inst ( .DIN1(_49060), .DIN2(_49061), .Q(_48761) );
  nor2s1 _49583_inst ( .DIN1(_53520), .DIN2(_2429), .Q(_49061) );
  nor2s1 _49584_inst ( .DIN1(_2320), .DIN2(_26633), .Q(_49060) );
  hi1s1 _49585_inst ( .DIN(_48368), .Q(_48545) );
  nnd2s1 _49586_inst ( .DIN1(_49062), .DIN2(_48926), .Q(_48368) );
  nor2s1 _49587_inst ( .DIN1(_49051), .DIN2(_48912), .Q(_48926) );
  nor2s1 _49588_inst ( .DIN1(_48875), .DIN2(_48961), .Q(_49062) );
  nor2s1 _49589_inst ( .DIN1(_48336), .DIN2(_48863), .Q(_49056) );
  nnd2s1 _49590_inst ( .DIN1(_48584), .DIN2(_49063), .Q(_48863) );
  nnd2s1 _49591_inst ( .DIN1(_48291), .DIN2(_48137), .Q(_49063) );
  and2s1 _49592_inst ( .DIN1(_49064), .DIN2(_34669), .Q(_48291) );
  hi1s1 _49593_inst ( .DIN(_33614), .Q(_34669) );
  nnd2s1 _49594_inst ( .DIN1(_49065), .DIN2(_49066), .Q(_33614) );
  hi1s1 _49595_inst ( .DIN(_48469), .Q(_48584) );
  nor2s1 _49596_inst ( .DIN1(_39095), .DIN2(_48284), .Q(_48469) );
  nnd2s1 _49597_inst ( .DIN1(_48726), .DIN2(_26769), .Q(_48284) );
  nor2s1 _49598_inst ( .DIN1(_34828), .DIN2(_38284), .Q(_48726) );
  nnd2s1 _49599_inst ( .DIN1(_49067), .DIN2(_49068), .Q(_38284) );
  nnd2s1 _49600_inst ( .DIN1(_48983), .DIN2(_49022), .Q(_39095) );
  nnd2s1 _49601_inst ( .DIN1(_49069), .DIN2(_49070), .Q(_48336) );
  or2s1 _49602_inst ( .DIN1(_48784), .DIN2(_26806), .Q(_49070) );
  nnd2s1 _49603_inst ( .DIN1(_49071), .DIN2(_34676), .Q(_48784) );
  nor2s1 _49604_inst ( .DIN1(_38283), .DIN2(_31103), .Q(_49071) );
  nnd2s1 _49605_inst ( .DIN1(_48189), .DIN2(_26768), .Q(_49069) );
  and2s1 _49606_inst ( .DIN1(_49064), .DIN2(_34677), .Q(_48189) );
  hi1s1 _49607_inst ( .DIN(_35757), .Q(_34677) );
  nnd2s1 _49608_inst ( .DIN1(_49066), .DIN2(_49022), .Q(_35757) );
  hi1s1 _49609_inst ( .DIN(_49051), .Q(_49022) );
  nor2s1 _49610_inst ( .DIN1(_36022), .DIN2(_34828), .Q(_49064) );
  nnd2s1 _49611_inst ( .DIN1(_49072), .DIN2(_2395), .Q(_34828) );
  nor2s1 _49612_inst ( .DIN1(_2320), .DIN2(_26278), .Q(_49072) );
  nnd2s1 _49613_inst ( .DIN1(_49073), .DIN2(_48302), .Q(_48971) );
  and2s1 _49614_inst ( .DIN1(_49074), .DIN2(_49075), .Q(_48302) );
  nor2s1 _49615_inst ( .DIN1(_48330), .DIN2(_49076), .Q(_49075) );
  nnd2s1 _49616_inst ( .DIN1(_48745), .DIN2(_48141), .Q(_49076) );
  nnd2s1 _49617_inst ( .DIN1(_26769), .DIN2(_49077), .Q(_48141) );
  nnd2s1 _49618_inst ( .DIN1(_49078), .DIN2(_48245), .Q(_49077) );
  nnd2s1 _49619_inst ( .DIN1(_49079), .DIN2(_38486), .Q(_48245) );
  hi1s1 _49620_inst ( .DIN(_34827), .Q(_38486) );
  nnd2s1 _49621_inst ( .DIN1(_49080), .DIN2(_53520), .Q(_34827) );
  nor2s1 _49622_inst ( .DIN1(_2395), .DIN2(_2320), .Q(_49080) );
  nor2s1 _49623_inst ( .DIN1(_37555), .DIN2(_38280), .Q(_49079) );
  nor2s1 _49624_inst ( .DIN1(_48650), .DIN2(_48638), .Q(_49078) );
  and2s1 _49625_inst ( .DIN1(_48700), .DIN2(_48548), .Q(_48638) );
  hi1s1 _49626_inst ( .DIN(_37555), .Q(_48548) );
  nnd2s1 _49627_inst ( .DIN1(_48983), .DIN2(_49065), .Q(_37555) );
  nor2s1 _49628_inst ( .DIN1(_48760), .DIN2(_26324), .Q(_48983) );
  nor2s1 _49629_inst ( .DIN1(_39417), .DIN2(_36022), .Q(_48700) );
  nnd2s1 _49630_inst ( .DIN1(_49081), .DIN2(_49082), .Q(_36022) );
  nor2s1 _49631_inst ( .DIN1(_2473), .DIN2(_2472), .Q(_49081) );
  nor2s1 _49632_inst ( .DIN1(_48918), .DIN2(_48959), .Q(_48650) );
  hi1s1 _49633_inst ( .DIN(_48929), .Q(_48959) );
  nor2s1 _49634_inst ( .DIN1(_48724), .DIN2(_48875), .Q(_48929) );
  nnd2s1 _49635_inst ( .DIN1(_49067), .DIN2(_49054), .Q(_48724) );
  nor2s1 _49636_inst ( .DIN1(_2472), .DIN2(_26303), .Q(_49067) );
  nnd2s1 _49637_inst ( .DIN1(_48984), .DIN2(_49083), .Q(_48918) );
  hi1s1 _49638_inst ( .DIN(_48470), .Q(_48745) );
  nor2s1 _49639_inst ( .DIN1(_48174), .DIN2(_26844), .Q(_48470) );
  or2s1 _49640_inst ( .DIN1(_48919), .DIN2(_48927), .Q(_48174) );
  nnd2s1 _49641_inst ( .DIN1(_49027), .DIN2(_49068), .Q(_48927) );
  nnd2s1 _49642_inst ( .DIN1(_48963), .DIN2(_49065), .Q(_48919) );
  nor2s1 _49643_inst ( .DIN1(_48680), .DIN2(_37557), .Q(_48330) );
  nnd2s1 _49644_inst ( .DIN1(_49084), .DIN2(_48984), .Q(_37557) );
  nor2s1 _49645_inst ( .DIN1(_26324), .DIN2(_48930), .Q(_49084) );
  hi1s1 _49646_inst ( .DIN(_49012), .Q(_48930) );
  nnd2s1 _49647_inst ( .DIN1(_48442), .DIN2(_48137), .Q(_48680) );
  nor2s1 _49648_inst ( .DIN1(_36021), .DIN2(_38460), .Q(_48442) );
  nor2s1 _49649_inst ( .DIN1(_48755), .DIN2(_49085), .Q(_49074) );
  nnd2s1 _49650_inst ( .DIN1(_49086), .DIN2(_49087), .Q(_49085) );
  nnd2s1 _49651_inst ( .DIN1(_26768), .DIN2(_49088), .Q(_49087) );
  nnd2s1 _49652_inst ( .DIN1(_48554), .DIN2(_48175), .Q(_49088) );
  nnd2s1 _49653_inst ( .DIN1(_49089), .DIN2(_48963), .Q(_48175) );
  nor2s1 _49654_inst ( .DIN1(_48875), .DIN2(_48760), .Q(_48963) );
  hi1s1 _49655_inst ( .DIN(_48911), .Q(_48875) );
  nor2s1 _49656_inst ( .DIN1(_48868), .DIN2(_2429), .Q(_48911) );
  nnd2s1 _49657_inst ( .DIN1(_49090), .DIN2(_2320), .Q(_48868) );
  nor2s1 _49658_inst ( .DIN1(_48759), .DIN2(_48961), .Q(_49089) );
  nnd2s1 _49659_inst ( .DIN1(_49091), .DIN2(_49054), .Q(_48961) );
  nnd2s1 _49660_inst ( .DIN1(_48987), .DIN2(_39096), .Q(_48554) );
  hi1s1 _49661_inst ( .DIN(_34672), .Q(_39096) );
  nnd2s1 _49662_inst ( .DIN1(_49092), .DIN2(_49050), .Q(_34672) );
  hi1s1 _49663_inst ( .DIN(_48760), .Q(_49050) );
  nnd2s1 _49664_inst ( .DIN1(_2439), .DIN2(_26714), .Q(_48760) );
  nor2s1 _49665_inst ( .DIN1(_2429), .DIN2(_48913), .Q(_49092) );
  nor2s1 _49666_inst ( .DIN1(_36021), .DIN2(_31103), .Q(_48987) );
  nnd2s1 _49667_inst ( .DIN1(_48224), .DIN2(_48173), .Q(_49086) );
  nnd2s1 _49668_inst ( .DIN1(_49093), .DIN2(_49094), .Q(_48224) );
  nnd2s1 _49669_inst ( .DIN1(_48849), .DIN2(_34676), .Q(_49094) );
  nor2s1 _49670_inst ( .DIN1(_48877), .DIN2(_49051), .Q(_34676) );
  nnd2s1 _49671_inst ( .DIN1(_2440), .DIN2(_26725), .Q(_49051) );
  or2s1 _49672_inst ( .DIN1(_35785), .DIN2(_48924), .Q(_49093) );
  nnd2s1 _49673_inst ( .DIN1(_36977), .DIN2(_35617), .Q(_48924) );
  hi1s1 _49674_inst ( .DIN(_38460), .Q(_35617) );
  hi1s1 _49675_inst ( .DIN(_42270), .Q(_36977) );
  nnd2s1 _49676_inst ( .DIN1(_49068), .DIN2(_49055), .Q(_42270) );
  nnd2s1 _49677_inst ( .DIN1(_49095), .DIN2(_49012), .Q(_35785) );
  nor2s1 _49678_inst ( .DIN1(_26324), .DIN2(_48759), .Q(_49095) );
  nnd2s1 _49679_inst ( .DIN1(_49096), .DIN2(_49097), .Q(_48755) );
  nnd2s1 _49680_inst ( .DIN1(_48372), .DIN2(_48130), .Q(_49097) );
  hi1s1 _49681_inst ( .DIN(_48403), .Q(_48372) );
  nnd2s1 _49682_inst ( .DIN1(_48937), .DIN2(_37556), .Q(_48403) );
  hi1s1 _49683_inst ( .DIN(_35695), .Q(_37556) );
  nnd2s1 _49684_inst ( .DIN1(_38027), .DIN2(_48984), .Q(_35695) );
  hi1s1 _49685_inst ( .DIN(_48913), .Q(_48984) );
  nor2s1 _49686_inst ( .DIN1(_38283), .DIN2(_38460), .Q(_48937) );
  nnd2s1 _49687_inst ( .DIN1(_49098), .DIN2(_2473), .Q(_38283) );
  nor2s1 _49688_inst ( .DIN1(_2472), .DIN2(_49007), .Q(_49098) );
  nnd2s1 _49689_inst ( .DIN1(_48190), .DIN2(_48173), .Q(_49096) );
  hi1s1 _49690_inst ( .DIN(_48402), .Q(_48190) );
  nnd2s1 _49691_inst ( .DIN1(_48942), .DIN2(_34399), .Q(_48402) );
  hi1s1 _49692_inst ( .DIN(_35696), .Q(_34399) );
  nnd2s1 _49693_inst ( .DIN1(_49099), .DIN2(_49065), .Q(_35696) );
  nor2s1 _49694_inst ( .DIN1(_2429), .DIN2(_48912), .Q(_49099) );
  nor2s1 _49695_inst ( .DIN1(_38460), .DIN2(_38261), .Q(_48942) );
  nnd2s1 _49696_inst ( .DIN1(_49100), .DIN2(_49027), .Q(_38261) );
  nnd2s1 _49697_inst ( .DIN1(_49090), .DIN2(_26430), .Q(_38460) );
  nor2s1 _49698_inst ( .DIN1(_53520), .DIN2(_2395), .Q(_49090) );
  nor2s1 _49699_inst ( .DIN1(_48269), .DIN2(_48448), .Q(_49073) );
  or2s1 _49700_inst ( .DIN1(_48507), .DIN2(_48149), .Q(_48448) );
  nor2s1 _49701_inst ( .DIN1(_48254), .DIN2(_48220), .Q(_48149) );
  hi1s1 _49702_inst ( .DIN(_48173), .Q(_48220) );
  nnd2s1 _49703_inst ( .DIN1(_26843), .DIN2(_26783), .Q(_48173) );
  hi1s1 _49704_inst ( .DIN(_48818), .Q(_48254) );
  nor2s1 _49705_inst ( .DIN1(_49101), .DIN2(_31103), .Q(_48818) );
  nnd2s1 _49706_inst ( .DIN1(_49102), .DIN2(_2395), .Q(_31103) );
  nor2s1 _49707_inst ( .DIN1(_53520), .DIN2(_26430), .Q(_49102) );
  or2s1 _49708_inst ( .DIN1(_36611), .DIN2(_36021), .Q(_49101) );
  nnd2s1 _49709_inst ( .DIN1(_49100), .DIN2(_49055), .Q(_36021) );
  nor2s1 _49710_inst ( .DIN1(_26642), .DIN2(_2474), .Q(_49055) );
  nor2s1 _49711_inst ( .DIN1(_53518), .DIN2(_2473), .Q(_49100) );
  hi1s1 _49712_inst ( .DIN(_33611), .Q(_36611) );
  nor2s1 _49713_inst ( .DIN1(_48913), .DIN2(_48877), .Q(_33611) );
  nnd2s1 _49714_inst ( .DIN1(_2429), .DIN2(_49083), .Q(_48877) );
  nnd2s1 _49715_inst ( .DIN1(_2432), .DIN2(_26316), .Q(_48913) );
  nor2s1 _49716_inst ( .DIN1(_48686), .DIN2(_48332), .Q(_48507) );
  nnd2s1 _49717_inst ( .DIN1(_48849), .DIN2(_27937), .Q(_48686) );
  hi1s1 _49718_inst ( .DIN(_35694), .Q(_27937) );
  nnd2s1 _49719_inst ( .DIN1(_38028), .DIN2(_49066), .Q(_35694) );
  and2s1 _49720_inst ( .DIN1(_49083), .DIN2(_26324), .Q(_49066) );
  nor2s1 _49721_inst ( .DIN1(_26714), .DIN2(_2439), .Q(_49083) );
  hi1s1 _49722_inst ( .DIN(_48759), .Q(_38028) );
  nnd2s1 _49723_inst ( .DIN1(_26316), .DIN2(_26725), .Q(_48759) );
  nor2s1 _49724_inst ( .DIN1(_32015), .DIN2(_42209), .Q(_48849) );
  nnd2s1 _49725_inst ( .DIN1(_49103), .DIN2(_2472), .Q(_42209) );
  nor2s1 _49726_inst ( .DIN1(_49007), .DIN2(_26580), .Q(_49103) );
  hi1s1 _49727_inst ( .DIN(_49082), .Q(_49007) );
  nor2s1 _49728_inst ( .DIN1(_26303), .DIN2(_53518), .Q(_49082) );
  nnd2s1 _49729_inst ( .DIN1(_49104), .DIN2(_2320), .Q(_32015) );
  nor2s1 _49730_inst ( .DIN1(_2395), .DIN2(_26278), .Q(_49104) );
  nnd2s1 _49731_inst ( .DIN1(_48627), .DIN2(_49105), .Q(_48269) );
  nnd2s1 _49732_inst ( .DIN1(_48465), .DIN2(_48137), .Q(_49105) );
  and2s1 _49733_inst ( .DIN1(_48982), .DIN2(_35706), .Q(_48465) );
  hi1s1 _49734_inst ( .DIN(_37551), .Q(_35706) );
  nnd2s1 _49735_inst ( .DIN1(_49106), .DIN2(_49012), .Q(_37551) );
  nor2s1 _49736_inst ( .DIN1(_53519), .DIN2(_2439), .Q(_49012) );
  nor2s1 _49737_inst ( .DIN1(_26324), .DIN2(_49013), .Q(_49106) );
  nor2s1 _49738_inst ( .DIN1(_41220), .DIN2(_39417), .Q(_48982) );
  nnd2s1 _49739_inst ( .DIN1(_49054), .DIN2(_49027), .Q(_41220) );
  nor2s1 _49740_inst ( .DIN1(_2474), .DIN2(_2472), .Q(_49027) );
  and2s1 _49741_inst ( .DIN1(_53518), .DIN2(_26580), .Q(_49054) );
  nnd2s1 _49742_inst ( .DIN1(_48562), .DIN2(_26769), .Q(_48627) );
  hi1s1 _49743_inst ( .DIN(_48992), .Q(_48562) );
  nnd2s1 _49744_inst ( .DIN1(_49107), .DIN2(_48589), .Q(_48992) );
  hi1s1 _49745_inst ( .DIN(_34671), .Q(_48589) );
  nnd2s1 _49746_inst ( .DIN1(_38027), .DIN2(_49065), .Q(_34671) );
  hi1s1 _49747_inst ( .DIN(_49013), .Q(_49065) );
  nnd2s1 _49748_inst ( .DIN1(_2432), .DIN2(_2440), .Q(_49013) );
  nor2s1 _49749_inst ( .DIN1(_48912), .DIN2(_26324), .Q(_38027) );
  nnd2s1 _49750_inst ( .DIN1(_2439), .DIN2(_53519), .Q(_48912) );
  nor2s1 _49751_inst ( .DIN1(_39417), .DIN2(_38280), .Q(_49107) );
  nnd2s1 _49752_inst ( .DIN1(_49091), .DIN2(_49068), .Q(_38280) );
  and2s1 _49753_inst ( .DIN1(_53518), .DIN2(_2473), .Q(_49068) );
  nor2s1 _49754_inst ( .DIN1(_26303), .DIN2(_26642), .Q(_49091) );
  nnd2s1 _49755_inst ( .DIN1(_49108), .DIN2(_2395), .Q(_39417) );
  nor2s1 _49756_inst ( .DIN1(_26278), .DIN2(_26430), .Q(_49108) );
  nnd2s1 _49757_inst ( .DIN1(_49109), .DIN2(_49110), .Q(____0___________[9])
         );
  nor2s1 _49758_inst ( .DIN1(_49111), .DIN2(_49112), .Q(_49110) );
  nnd2s1 _49759_inst ( .DIN1(_49113), .DIN2(_49114), .Q(_49112) );
  nor2s1 _49760_inst ( .DIN1(_49115), .DIN2(_49116), .Q(_49113) );
  nor2s1 _49761_inst ( .DIN1(_49117), .DIN2(_49118), .Q(_49116) );
  nor2s1 _49762_inst ( .DIN1(_49119), .DIN2(_49120), .Q(_49115) );
  nnd2s1 _49763_inst ( .DIN1(_49121), .DIN2(_49122), .Q(_49111) );
  nor2s1 _49764_inst ( .DIN1(_49123), .DIN2(_49124), .Q(_49122) );
  nor2s1 _49765_inst ( .DIN1(_49125), .DIN2(_49126), .Q(_49121) );
  nor2s1 _49766_inst ( .DIN1(_49127), .DIN2(_49128), .Q(_49125) );
  nor2s1 _49767_inst ( .DIN1(_49129), .DIN2(_49130), .Q(_49109) );
  nnd2s1 _49768_inst ( .DIN1(_49131), .DIN2(_49132), .Q(_49130) );
  hi1s1 _49769_inst ( .DIN(_49133), .Q(_49132) );
  nor2s1 _49770_inst ( .DIN1(_49134), .DIN2(_49135), .Q(_49131) );
  nnd2s1 _49771_inst ( .DIN1(_49136), .DIN2(_49137), .Q(_49129) );
  hi1s1 _49772_inst ( .DIN(_49138), .Q(_49137) );
  nor2s1 _49773_inst ( .DIN1(_49139), .DIN2(_49140), .Q(_49136) );
  nnd2s1 _49774_inst ( .DIN1(_49141), .DIN2(_49142), .Q(____0___________[8])
         );
  nor2s1 _49775_inst ( .DIN1(_49143), .DIN2(_49144), .Q(_49142) );
  nnd2s1 _49776_inst ( .DIN1(_49145), .DIN2(_49146), .Q(_49144) );
  nor2s1 _49777_inst ( .DIN1(_49147), .DIN2(_49148), .Q(_49146) );
  nor2s1 _49778_inst ( .DIN1(_49149), .DIN2(_49150), .Q(_49148) );
  nor2s1 _49779_inst ( .DIN1(_49151), .DIN2(_49152), .Q(_49147) );
  nor2s1 _49780_inst ( .DIN1(_49153), .DIN2(_49154), .Q(_49145) );
  nor2s1 _49781_inst ( .DIN1(_49155), .DIN2(_49156), .Q(_49153) );
  nnd2s1 _49782_inst ( .DIN1(_49157), .DIN2(_49158), .Q(_49143) );
  nor2s1 _49783_inst ( .DIN1(_49159), .DIN2(_49160), .Q(_49158) );
  nor2s1 _49784_inst ( .DIN1(_49161), .DIN2(_49162), .Q(_49160) );
  nor2s1 _49785_inst ( .DIN1(_49163), .DIN2(_49164), .Q(_49157) );
  nor2s1 _49786_inst ( .DIN1(_49165), .DIN2(_49166), .Q(_49164) );
  nor2s1 _49787_inst ( .DIN1(_49167), .DIN2(_49168), .Q(_49141) );
  nnd2s1 _49788_inst ( .DIN1(_49169), .DIN2(_49170), .Q(_49168) );
  nor2s1 _49789_inst ( .DIN1(_49171), .DIN2(_49172), .Q(_49169) );
  nnd2s1 _49790_inst ( .DIN1(_49173), .DIN2(_49174), .Q(_49167) );
  nor2s1 _49791_inst ( .DIN1(_49175), .DIN2(_49176), .Q(_49174) );
  nor2s1 _49792_inst ( .DIN1(_49177), .DIN2(_49178), .Q(_49173) );
  nnd2s1 _49793_inst ( .DIN1(_49179), .DIN2(_49180), .Q(____0___________[7])
         );
  nor2s1 _49794_inst ( .DIN1(_49181), .DIN2(_49182), .Q(_49180) );
  nnd2s1 _49795_inst ( .DIN1(_49183), .DIN2(_49184), .Q(_49182) );
  nor2s1 _49796_inst ( .DIN1(_49185), .DIN2(_49186), .Q(_49183) );
  nor2s1 _49797_inst ( .DIN1(_49187), .DIN2(_49188), .Q(_49186) );
  nnd2s1 _49798_inst ( .DIN1(_49189), .DIN2(_49190), .Q(_49181) );
  nor2s1 _49799_inst ( .DIN1(_49191), .DIN2(_49192), .Q(_49190) );
  nor2s1 _49800_inst ( .DIN1(_49193), .DIN2(_49194), .Q(_49189) );
  nor2s1 _49801_inst ( .DIN1(_49195), .DIN2(_49161), .Q(_49194) );
  nor2s1 _49802_inst ( .DIN1(_49196), .DIN2(_49197), .Q(_49193) );
  nor2s1 _49803_inst ( .DIN1(_49198), .DIN2(_49199), .Q(_49179) );
  nnd2s1 _49804_inst ( .DIN1(_49200), .DIN2(_49201), .Q(_49199) );
  nor2s1 _49805_inst ( .DIN1(_49202), .DIN2(_49203), .Q(_49200) );
  nnd2s1 _49806_inst ( .DIN1(_49204), .DIN2(_49205), .Q(_49198) );
  nor2s1 _49807_inst ( .DIN1(_49206), .DIN2(_49207), .Q(_49205) );
  nor2s1 _49808_inst ( .DIN1(_49208), .DIN2(_49209), .Q(_49204) );
  nnd2s1 _49809_inst ( .DIN1(_49210), .DIN2(_49211), .Q(____0___________[6])
         );
  nor2s1 _49810_inst ( .DIN1(_49212), .DIN2(_49213), .Q(_49211) );
  nnd2s1 _49811_inst ( .DIN1(_49214), .DIN2(_49215), .Q(_49213) );
  nor2s1 _49812_inst ( .DIN1(_49216), .DIN2(_49217), .Q(_49214) );
  nor2s1 _49813_inst ( .DIN1(_49218), .DIN2(_49219), .Q(_49217) );
  nnd2s1 _49814_inst ( .DIN1(_49220), .DIN2(_49221), .Q(_49212) );
  and2s1 _49815_inst ( .DIN1(_49222), .DIN2(_49223), .Q(_49221) );
  nor2s1 _49816_inst ( .DIN1(_49224), .DIN2(_49225), .Q(_49220) );
  nor2s1 _49817_inst ( .DIN1(_49226), .DIN2(_49227), .Q(_49225) );
  nor2s1 _49818_inst ( .DIN1(_49161), .DIN2(_49228), .Q(_49224) );
  nor2s1 _49819_inst ( .DIN1(_49229), .DIN2(_49230), .Q(_49210) );
  nnd2s1 _49820_inst ( .DIN1(_49231), .DIN2(_49232), .Q(_49230) );
  hi1s1 _49821_inst ( .DIN(_49233), .Q(_49232) );
  nor2s1 _49822_inst ( .DIN1(_49234), .DIN2(_49235), .Q(_49231) );
  nnd2s1 _49823_inst ( .DIN1(_49236), .DIN2(_49237), .Q(_49229) );
  hi1s1 _49824_inst ( .DIN(_49238), .Q(_49237) );
  nor2s1 _49825_inst ( .DIN1(_49177), .DIN2(_49239), .Q(_49236) );
  nnd2s1 _49826_inst ( .DIN1(_49240), .DIN2(_49241), .Q(_49177) );
  nor2s1 _49827_inst ( .DIN1(_49242), .DIN2(_49243), .Q(_49241) );
  nnd2s1 _49828_inst ( .DIN1(_49244), .DIN2(_49245), .Q(_49243) );
  nor2s1 _49829_inst ( .DIN1(_49246), .DIN2(_49247), .Q(_49244) );
  nor2s1 _49830_inst ( .DIN1(_49161), .DIN2(_49248), .Q(_49247) );
  nor2s1 _49831_inst ( .DIN1(_49249), .DIN2(_49165), .Q(_49246) );
  nnd2s1 _49832_inst ( .DIN1(_49250), .DIN2(_49251), .Q(_49242) );
  nor2s1 _49833_inst ( .DIN1(_49252), .DIN2(_49253), .Q(_49250) );
  nor2s1 _49834_inst ( .DIN1(_49254), .DIN2(_49255), .Q(_49253) );
  nor2s1 _49835_inst ( .DIN1(_49256), .DIN2(_49257), .Q(_49254) );
  hi1s1 _49836_inst ( .DIN(_49258), .Q(_49252) );
  nor2s1 _49837_inst ( .DIN1(_49259), .DIN2(_49260), .Q(_49240) );
  or2s1 _49838_inst ( .DIN1(_49261), .DIN2(_49262), .Q(_49260) );
  nnd2s1 _49839_inst ( .DIN1(_49263), .DIN2(_49264), .Q(_49259) );
  nor2s1 _49840_inst ( .DIN1(_49265), .DIN2(_49266), .Q(_49263) );
  nnd2s1 _49841_inst ( .DIN1(_49267), .DIN2(_49268), .Q(____0___________[5])
         );
  nor2s1 _49842_inst ( .DIN1(_49269), .DIN2(_49270), .Q(_49268) );
  nnd2s1 _49843_inst ( .DIN1(_49271), .DIN2(_49272), .Q(_49270) );
  nor2s1 _49844_inst ( .DIN1(_49273), .DIN2(_49274), .Q(_49272) );
  nor2s1 _49845_inst ( .DIN1(_49275), .DIN2(_49117), .Q(_49274) );
  nor2s1 _49846_inst ( .DIN1(_49276), .DIN2(_49277), .Q(_49271) );
  nor2s1 _49847_inst ( .DIN1(_49149), .DIN2(_49278), .Q(_49277) );
  nor2s1 _49848_inst ( .DIN1(_49255), .DIN2(_49279), .Q(_49276) );
  nnd2s1 _49849_inst ( .DIN1(_49280), .DIN2(_49281), .Q(_49269) );
  nor2s1 _49850_inst ( .DIN1(_49282), .DIN2(_49283), .Q(_49281) );
  and2s1 _49851_inst ( .DIN1(_49284), .DIN2(_49285), .Q(_49280) );
  nor2s1 _49852_inst ( .DIN1(_49286), .DIN2(_49287), .Q(_49267) );
  nnd2s1 _49853_inst ( .DIN1(_49288), .DIN2(_49289), .Q(_49287) );
  hi1s1 _49854_inst ( .DIN(_49290), .Q(_49289) );
  nor2s1 _49855_inst ( .DIN1(_49291), .DIN2(_49292), .Q(_49288) );
  nnd2s1 _49856_inst ( .DIN1(_49293), .DIN2(_49294), .Q(_49286) );
  nor2s1 _49857_inst ( .DIN1(_49295), .DIN2(_49296), .Q(_49294) );
  nor2s1 _49858_inst ( .DIN1(_49206), .DIN2(_49297), .Q(_49293) );
  nnd2s1 _49859_inst ( .DIN1(_49298), .DIN2(_49299), .Q(_49206) );
  nnd2s1 _49860_inst ( .DIN1(_49300), .DIN2(_49301), .Q(_49299) );
  nnd2s1 _49861_inst ( .DIN1(_49302), .DIN2(_49303), .Q(____0___________[4])
         );
  nor2s1 _49862_inst ( .DIN1(_49304), .DIN2(_49305), .Q(_49303) );
  nnd2s1 _49863_inst ( .DIN1(_49306), .DIN2(_49307), .Q(_49305) );
  nor2s1 _49864_inst ( .DIN1(_49308), .DIN2(_49309), .Q(_49307) );
  nor2s1 _49865_inst ( .DIN1(_49149), .DIN2(_49310), .Q(_49309) );
  nor2s1 _49866_inst ( .DIN1(_49311), .DIN2(_49312), .Q(_49308) );
  nor2s1 _49867_inst ( .DIN1(_49313), .DIN2(_49314), .Q(_49306) );
  nor2s1 _49868_inst ( .DIN1(_49187), .DIN2(_49315), .Q(_49313) );
  nnd2s1 _49869_inst ( .DIN1(_49316), .DIN2(_49317), .Q(_49304) );
  nor2s1 _49870_inst ( .DIN1(_49318), .DIN2(_49319), .Q(_49317) );
  nor2s1 _49871_inst ( .DIN1(_49320), .DIN2(_49321), .Q(_49316) );
  nor2s1 _49872_inst ( .DIN1(_49322), .DIN2(_49323), .Q(_49302) );
  nnd2s1 _49873_inst ( .DIN1(_49324), .DIN2(_49325), .Q(_49323) );
  hi1s1 _49874_inst ( .DIN(_49326), .Q(_49325) );
  nor2s1 _49875_inst ( .DIN1(_49327), .DIN2(_49328), .Q(_49324) );
  nnd2s1 _49876_inst ( .DIN1(_49329), .DIN2(_49330), .Q(_49322) );
  nor2s1 _49877_inst ( .DIN1(_49331), .DIN2(_49178), .Q(_49330) );
  nnd2s1 _49878_inst ( .DIN1(_49332), .DIN2(_49333), .Q(_49178) );
  nor2s1 _49879_inst ( .DIN1(_49334), .DIN2(_49335), .Q(_49333) );
  nnd2s1 _49880_inst ( .DIN1(_49336), .DIN2(_49337), .Q(_49335) );
  nor2s1 _49881_inst ( .DIN1(_49338), .DIN2(_49339), .Q(_49332) );
  nnd2s1 _49882_inst ( .DIN1(_49340), .DIN2(_49341), .Q(_49339) );
  nnd2s1 _49883_inst ( .DIN1(_49342), .DIN2(_49343), .Q(_49341) );
  nor2s1 _49884_inst ( .DIN1(_49344), .DIN2(_49345), .Q(_49338) );
  nor2s1 _49885_inst ( .DIN1(_49346), .DIN2(_49347), .Q(_49329) );
  nnd2s1 _49886_inst ( .DIN1(_49348), .DIN2(_49349), .Q(____0___________[3])
         );
  nor2s1 _49887_inst ( .DIN1(_49350), .DIN2(_49351), .Q(_49349) );
  nnd2s1 _49888_inst ( .DIN1(_49352), .DIN2(_49353), .Q(_49351) );
  nor2s1 _49889_inst ( .DIN1(_49354), .DIN2(_49355), .Q(_49352) );
  nor2s1 _49890_inst ( .DIN1(_49310), .DIN2(_49165), .Q(_49355) );
  nnd2s1 _49891_inst ( .DIN1(_49356), .DIN2(_49357), .Q(_49350) );
  nor2s1 _49892_inst ( .DIN1(_49159), .DIN2(_49320), .Q(_49357) );
  nor2s1 _49893_inst ( .DIN1(_49358), .DIN2(_49359), .Q(_49356) );
  nor2s1 _49894_inst ( .DIN1(_49360), .DIN2(_49361), .Q(_49348) );
  nnd2s1 _49895_inst ( .DIN1(_49362), .DIN2(_49363), .Q(_49361) );
  nor2s1 _49896_inst ( .DIN1(_49364), .DIN2(_49365), .Q(_49362) );
  nnd2s1 _49897_inst ( .DIN1(_49366), .DIN2(_49367), .Q(_49360) );
  nor2s1 _49898_inst ( .DIN1(_49135), .DIN2(_49235), .Q(_49367) );
  nnd2s1 _49899_inst ( .DIN1(_49368), .DIN2(_49369), .Q(_49235) );
  nor2s1 _49900_inst ( .DIN1(_49370), .DIN2(_49371), .Q(_49369) );
  nnd2s1 _49901_inst ( .DIN1(_49372), .DIN2(_49373), .Q(_49371) );
  hi1s1 _49902_inst ( .DIN(_49374), .Q(_49373) );
  nnd2s1 _49903_inst ( .DIN1(_49375), .DIN2(_49376), .Q(_49372) );
  nnd2s1 _49904_inst ( .DIN1(_49377), .DIN2(_49378), .Q(_49370) );
  nor2s1 _49905_inst ( .DIN1(_49379), .DIN2(_49380), .Q(_49368) );
  nnd2s1 _49906_inst ( .DIN1(_49381), .DIN2(_49382), .Q(_49380) );
  nnd2s1 _49907_inst ( .DIN1(_49383), .DIN2(_49343), .Q(_49382) );
  hi1s1 _49908_inst ( .DIN(_49297), .Q(_49381) );
  nnd2s1 _49909_inst ( .DIN1(_49384), .DIN2(_49385), .Q(_49297) );
  nor2s1 _49910_inst ( .DIN1(_49386), .DIN2(_49387), .Q(_49385) );
  nnd2s1 _49911_inst ( .DIN1(_49388), .DIN2(_49389), .Q(_49387) );
  hi1s1 _49912_inst ( .DIN(_49390), .Q(_49389) );
  nnd2s1 _49913_inst ( .DIN1(_49391), .DIN2(_49392), .Q(_49388) );
  nor2s1 _49914_inst ( .DIN1(_49393), .DIN2(_49127), .Q(_49386) );
  nor2s1 _49915_inst ( .DIN1(_49394), .DIN2(_49395), .Q(_49384) );
  nnd2s1 _49916_inst ( .DIN1(_49396), .DIN2(_49397), .Q(_49395) );
  nnd2s1 _49917_inst ( .DIN1(_49398), .DIN2(_49399), .Q(_49396) );
  nor2s1 _49918_inst ( .DIN1(_49400), .DIN2(_49120), .Q(_49394) );
  nnd2s1 _49919_inst ( .DIN1(_49401), .DIN2(_49402), .Q(_49135) );
  nor2s1 _49920_inst ( .DIN1(_49403), .DIN2(_49404), .Q(_49402) );
  nor2s1 _49921_inst ( .DIN1(_49155), .DIN2(_49405), .Q(_49404) );
  nor2s1 _49922_inst ( .DIN1(_49406), .DIN2(_49311), .Q(_49403) );
  nor2s1 _49923_inst ( .DIN1(_49407), .DIN2(_49408), .Q(_49406) );
  nor2s1 _49924_inst ( .DIN1(_49409), .DIN2(_49410), .Q(_49401) );
  nor2s1 _49925_inst ( .DIN1(_49411), .DIN2(_49412), .Q(_49410) );
  nor2s1 _49926_inst ( .DIN1(_49149), .DIN2(_49413), .Q(_49409) );
  nor2s1 _49927_inst ( .DIN1(_49414), .DIN2(_49415), .Q(_49366) );
  nnd2s1 _49928_inst ( .DIN1(_49416), .DIN2(_49417), .Q(____0___________[2])
         );
  nor2s1 _49929_inst ( .DIN1(_49418), .DIN2(_49419), .Q(_49417) );
  nnd2s1 _49930_inst ( .DIN1(_49264), .DIN2(_49114), .Q(_49419) );
  and2s1 _49931_inst ( .DIN1(_49420), .DIN2(_49421), .Q(_49114) );
  nor2s1 _49932_inst ( .DIN1(_49422), .DIN2(_49423), .Q(_49421) );
  nnd2s1 _49933_inst ( .DIN1(_49424), .DIN2(_49425), .Q(_49423) );
  hi1s1 _49934_inst ( .DIN(_49426), .Q(_49424) );
  nnd2s1 _49935_inst ( .DIN1(_49427), .DIN2(_49428), .Q(_49422) );
  nor2s1 _49936_inst ( .DIN1(_49429), .DIN2(_49430), .Q(_49420) );
  nnd2s1 _49937_inst ( .DIN1(_49184), .DIN2(_49215), .Q(_49430) );
  and2s1 _49938_inst ( .DIN1(_49431), .DIN2(_49432), .Q(_49215) );
  nor2s1 _49939_inst ( .DIN1(_49433), .DIN2(_49434), .Q(_49432) );
  nnd2s1 _49940_inst ( .DIN1(_49435), .DIN2(_49436), .Q(_49434) );
  or2s1 _49941_inst ( .DIN1(_49197), .DIN2(_49196), .Q(_49435) );
  nnd2s1 _49942_inst ( .DIN1(_49437), .DIN2(_49438), .Q(_49433) );
  nor2s1 _49943_inst ( .DIN1(_49439), .DIN2(_49440), .Q(_49437) );
  nor2s1 _49944_inst ( .DIN1(_49441), .DIN2(_49442), .Q(_49431) );
  or2s1 _49945_inst ( .DIN1(_49443), .DIN2(_49444), .Q(_49442) );
  or2s1 _49946_inst ( .DIN1(_49445), .DIN2(_49446), .Q(_49441) );
  and2s1 _49947_inst ( .DIN1(_49447), .DIN2(_49448), .Q(_49184) );
  nor2s1 _49948_inst ( .DIN1(_49449), .DIN2(_49450), .Q(_49448) );
  nor2s1 _49949_inst ( .DIN1(_49451), .DIN2(_49452), .Q(_49450) );
  nor2s1 _49950_inst ( .DIN1(_49295), .DIN2(_49453), .Q(_49447) );
  nnd2s1 _49951_inst ( .DIN1(_49454), .DIN2(_49455), .Q(_49295) );
  nnd2s1 _49952_inst ( .DIN1(_49456), .DIN2(_49457), .Q(_49455) );
  or2s1 _49953_inst ( .DIN1(_49458), .DIN2(_49459), .Q(_49456) );
  hi1s1 _49954_inst ( .DIN(_49154), .Q(_49454) );
  nnd2s1 _49955_inst ( .DIN1(_49460), .DIN2(_49461), .Q(_49154) );
  nnd2s1 _49956_inst ( .DIN1(_49462), .DIN2(_49463), .Q(_49461) );
  or2s1 _49957_inst ( .DIN1(_49464), .DIN2(_49465), .Q(_49460) );
  nnd2s1 _49958_inst ( .DIN1(_49466), .DIN2(_49467), .Q(_49429) );
  nor2s1 _49959_inst ( .DIN1(_49468), .DIN2(_49469), .Q(_49264) );
  or2s1 _49960_inst ( .DIN1(_49124), .DIN2(_49470), .Q(_49468) );
  nor2s1 _49961_inst ( .DIN1(_49465), .DIN2(_49471), .Q(_49470) );
  and2s1 _49962_inst ( .DIN1(_49472), .DIN2(_49473), .Q(_49471) );
  hi1s1 _49963_inst ( .DIN(_49285), .Q(_49124) );
  nnd2s1 _49964_inst ( .DIN1(_49474), .DIN2(_49475), .Q(_49418) );
  nor2s1 _49965_inst ( .DIN1(_49476), .DIN2(_49358), .Q(_49474) );
  hi1s1 _49966_inst ( .DIN(_49477), .Q(_49358) );
  nor2s1 _49967_inst ( .DIN1(_49478), .DIN2(_49479), .Q(_49416) );
  or2s1 _49968_inst ( .DIN1(_49480), .DIN2(_49481), .Q(_49479) );
  nnd2s1 _49969_inst ( .DIN1(_49482), .DIN2(_49483), .Q(_49478) );
  nor2s1 _49970_inst ( .DIN1(_49176), .DIN2(_49209), .Q(_49482) );
  nnd2s1 _49971_inst ( .DIN1(_49484), .DIN2(_49485), .Q(_49209) );
  nor2s1 _49972_inst ( .DIN1(_49486), .DIN2(_49487), .Q(_49484) );
  nnd2s1 _49973_inst ( .DIN1(_49488), .DIN2(_49489), .Q(_49176) );
  nnd2s1 _49974_inst ( .DIN1(_49490), .DIN2(_49491), .Q(____0___________[1])
         );
  nor2s1 _49975_inst ( .DIN1(_49492), .DIN2(_49493), .Q(_49491) );
  nnd2s1 _49976_inst ( .DIN1(_49494), .DIN2(_49495), .Q(_49493) );
  nor2s1 _49977_inst ( .DIN1(_49496), .DIN2(_49497), .Q(_49495) );
  nor2s1 _49978_inst ( .DIN1(_49187), .DIN2(_49498), .Q(_49497) );
  and2s1 _49979_inst ( .DIN1(_49376), .DIN2(_49499), .Q(_49496) );
  nor2s1 _49980_inst ( .DIN1(_49185), .DIN2(_49500), .Q(_49494) );
  nor2s1 _49981_inst ( .DIN1(_49501), .DIN2(_49156), .Q(_49500) );
  nor2s1 _49982_inst ( .DIN1(_49149), .DIN2(_49166), .Q(_49185) );
  nnd2s1 _49983_inst ( .DIN1(_49502), .DIN2(_49503), .Q(_49492) );
  nor2s1 _49984_inst ( .DIN1(_49504), .DIN2(_49505), .Q(_49503) );
  or2s1 _49985_inst ( .DIN1(_49506), .DIN2(_49123), .Q(_49505) );
  nor2s1 _49986_inst ( .DIN1(_49507), .DIN2(_49508), .Q(_49502) );
  nor2s1 _49987_inst ( .DIN1(_49117), .DIN2(_49509), .Q(_49508) );
  nor2s1 _49988_inst ( .DIN1(_49196), .DIN2(_49510), .Q(_49507) );
  nor2s1 _49989_inst ( .DIN1(_49511), .DIN2(_49512), .Q(_49490) );
  nnd2s1 _49990_inst ( .DIN1(_49513), .DIN2(_49514), .Q(_49512) );
  nor2s1 _49991_inst ( .DIN1(_49515), .DIN2(_49414), .Q(_49514) );
  nnd2s1 _49992_inst ( .DIN1(_49516), .DIN2(_49251), .Q(_49414) );
  nnd2s1 _49993_inst ( .DIN1(_49517), .DIN2(_49518), .Q(_49251) );
  nor2s1 _49994_inst ( .DIN1(_49519), .DIN2(_49520), .Q(_49513) );
  nnd2s1 _49995_inst ( .DIN1(_49521), .DIN2(_49522), .Q(_49511) );
  nor2s1 _49996_inst ( .DIN1(_49469), .DIN2(_49523), .Q(_49522) );
  nnd2s1 _49997_inst ( .DIN1(_49524), .DIN2(_49525), .Q(_49469) );
  nnd2s1 _49998_inst ( .DIN1(_49408), .DIN2(_49463), .Q(_49525) );
  nor2s1 _49999_inst ( .DIN1(_49292), .DIN2(_49526), .Q(_49521) );
  nnd2s1 _50000_inst ( .DIN1(_49527), .DIN2(_49528), .Q(_49292) );
  nor2s1 _50001_inst ( .DIN1(_49529), .DIN2(_49530), .Q(_49528) );
  nnd2s1 _50002_inst ( .DIN1(_49340), .DIN2(_49531), .Q(_49530) );
  nnd2s1 _50003_inst ( .DIN1(_49532), .DIN2(_49301), .Q(_49531) );
  nnd2s1 _50004_inst ( .DIN1(_49533), .DIN2(_49383), .Q(_49340) );
  nnd2s1 _50005_inst ( .DIN1(_49534), .DIN2(_49535), .Q(_49529) );
  nor2s1 _50006_inst ( .DIN1(_49159), .DIN2(_49536), .Q(_49534) );
  and2s1 _50007_inst ( .DIN1(_49537), .DIN2(_49538), .Q(_49159) );
  nor2s1 _50008_inst ( .DIN1(_49149), .DIN2(_49539), .Q(_49538) );
  or2s1 _50009_inst ( .DIN1(_49540), .DIN2(_2273), .Q(_49539) );
  nor2s1 _50010_inst ( .DIN1(_49541), .DIN2(_49542), .Q(_49527) );
  nnd2s1 _50011_inst ( .DIN1(_49543), .DIN2(_49544), .Q(_49542) );
  hi1s1 _50012_inst ( .DIN(_49207), .Q(_49543) );
  nnd2s1 _50013_inst ( .DIN1(_49545), .DIN2(_49546), .Q(_49207) );
  nnd2s1 _50014_inst ( .DIN1(_49407), .DIN2(_49392), .Q(_49546) );
  nnd2s1 _50015_inst ( .DIN1(_49547), .DIN2(_49301), .Q(_49545) );
  nnd2s1 _50016_inst ( .DIN1(_49548), .DIN2(_49549), .Q(_49541) );
  nnd2s1 _50017_inst ( .DIN1(_49550), .DIN2(_49551), .Q(_49549) );
  nnd2s1 _50018_inst ( .DIN1(_49552), .DIN2(_49553), .Q(_49548) );
  nnd2s1 _50019_inst ( .DIN1(_49554), .DIN2(_49555), .Q(____0___________[15])
         );
  nor2s1 _50020_inst ( .DIN1(_49556), .DIN2(_49557), .Q(_49555) );
  nnd2s1 _50021_inst ( .DIN1(_49558), .DIN2(_49559), .Q(_49557) );
  nor2s1 _50022_inst ( .DIN1(_49560), .DIN2(_49561), .Q(_49559) );
  nor2s1 _50023_inst ( .DIN1(_49311), .DIN2(_49562), .Q(_49561) );
  nor2s1 _50024_inst ( .DIN1(_49563), .DIN2(_49564), .Q(_49558) );
  nor2s1 _50025_inst ( .DIN1(_49565), .DIN2(_49165), .Q(_49564) );
  nor2s1 _50026_inst ( .DIN1(_49411), .DIN2(_49566), .Q(_49563) );
  nnd2s1 _50027_inst ( .DIN1(_49567), .DIN2(_49568), .Q(_49556) );
  nor2s1 _50028_inst ( .DIN1(_49439), .DIN2(_49318), .Q(_49568) );
  and2s1 _50029_inst ( .DIN1(_49517), .DIN2(_49569), .Q(_49318) );
  and2s1 _50030_inst ( .DIN1(_49436), .DIN2(_49337), .Q(_49567) );
  nor2s1 _50031_inst ( .DIN1(_49570), .DIN2(_49571), .Q(_49554) );
  nnd2s1 _50032_inst ( .DIN1(_49572), .DIN2(_49573), .Q(_49571) );
  nor2s1 _50033_inst ( .DIN1(_49480), .DIN2(_49574), .Q(_49572) );
  nnd2s1 _50034_inst ( .DIN1(_49575), .DIN2(_49576), .Q(_49480) );
  nor2s1 _50035_inst ( .DIN1(_49577), .DIN2(_49578), .Q(_49576) );
  nnd2s1 _50036_inst ( .DIN1(_49579), .DIN2(_49580), .Q(_49578) );
  nor2s1 _50037_inst ( .DIN1(_49581), .DIN2(_49249), .Q(_49577) );
  nor2s1 _50038_inst ( .DIN1(_49202), .DIN2(_49582), .Q(_49575) );
  nnd2s1 _50039_inst ( .DIN1(_49583), .DIN2(_49584), .Q(_49582) );
  nnd2s1 _50040_inst ( .DIN1(_49585), .DIN2(_49586), .Q(_49202) );
  nor2s1 _50041_inst ( .DIN1(_49587), .DIN2(_49588), .Q(_49586) );
  nnd2s1 _50042_inst ( .DIN1(_49535), .DIN2(_49589), .Q(_49588) );
  nnd2s1 _50043_inst ( .DIN1(_49590), .DIN2(_49591), .Q(_49587) );
  nor2s1 _50044_inst ( .DIN1(_49592), .DIN2(_49321), .Q(_49590) );
  nor2s1 _50045_inst ( .DIN1(_49593), .DIN2(_49594), .Q(_49585) );
  or2s1 _50046_inst ( .DIN1(_49595), .DIN2(_49596), .Q(_49594) );
  nnd2s1 _50047_inst ( .DIN1(_49597), .DIN2(_49598), .Q(_49593) );
  hi1s1 _50048_inst ( .DIN(_49171), .Q(_49598) );
  nnd2s1 _50049_inst ( .DIN1(_49599), .DIN2(_49600), .Q(_49171) );
  nor2s1 _50050_inst ( .DIN1(_49601), .DIN2(_49602), .Q(_49600) );
  nor2s1 _50051_inst ( .DIN1(_49603), .DIN2(_49604), .Q(_49599) );
  nor2s1 _50052_inst ( .DIN1(_49465), .DIN2(_49227), .Q(_49604) );
  hi1s1 _50053_inst ( .DIN(_49605), .Q(_49603) );
  nor2s1 _50054_inst ( .DIN1(_49138), .DIN2(_49261), .Q(_49597) );
  nnd2s1 _50055_inst ( .DIN1(_49606), .DIN2(_49607), .Q(_49138) );
  nnd2s1 _50056_inst ( .DIN1(_49608), .DIN2(_49609), .Q(_49607) );
  nor2s1 _50057_inst ( .DIN1(_49319), .DIN2(_49610), .Q(_49606) );
  nor2s1 _50058_inst ( .DIN1(_49465), .DIN2(_49611), .Q(_49610) );
  nor2s1 _50059_inst ( .DIN1(_49612), .DIN2(_47930), .Q(_49319) );
  nnd2s1 _50060_inst ( .DIN1(_49613), .DIN2(_49614), .Q(_49570) );
  nor2s1 _50061_inst ( .DIN1(_49140), .DIN2(_49615), .Q(_49614) );
  nnd2s1 _50062_inst ( .DIN1(_49616), .DIN2(_49617), .Q(_49140) );
  nor2s1 _50063_inst ( .DIN1(_49476), .DIN2(_49618), .Q(_49617) );
  nor2s1 _50064_inst ( .DIN1(_49619), .DIN2(_49620), .Q(_49616) );
  nor2s1 _50065_inst ( .DIN1(_49187), .DIN2(_49621), .Q(_49619) );
  nor2s1 _50066_inst ( .DIN1(_49208), .DIN2(_49364), .Q(_49613) );
  nnd2s1 _50067_inst ( .DIN1(_49622), .DIN2(_49623), .Q(_49364) );
  nor2s1 _50068_inst ( .DIN1(_49624), .DIN2(_49625), .Q(_49623) );
  nnd2s1 _50069_inst ( .DIN1(_49626), .DIN2(_49627), .Q(_49625) );
  hi1s1 _50070_inst ( .DIN(_49628), .Q(_49627) );
  or2s1 _50071_inst ( .DIN1(_49345), .DIN2(_49344), .Q(_49626) );
  nor2s1 _50072_inst ( .DIN1(_49278), .DIN2(_49165), .Q(_49624) );
  nor2s1 _50073_inst ( .DIN1(_49515), .DIN2(_49629), .Q(_49622) );
  nnd2s1 _50074_inst ( .DIN1(_49467), .DIN2(_49245), .Q(_49629) );
  and2s1 _50075_inst ( .DIN1(_49630), .DIN2(_49631), .Q(_49467) );
  nnd2s1 _50076_inst ( .DIN1(_49632), .DIN2(_49633), .Q(_49631) );
  nor2s1 _50077_inst ( .DIN1(_49282), .DIN2(_49634), .Q(_49630) );
  nnd2s1 _50078_inst ( .DIN1(_49635), .DIN2(_49636), .Q(_49515) );
  nnd2s1 _50079_inst ( .DIN1(_49637), .DIN2(_49457), .Q(_49636) );
  nnd2s1 _50080_inst ( .DIN1(_49638), .DIN2(_49639), .Q(_49208) );
  nor2s1 _50081_inst ( .DIN1(_49640), .DIN2(_49641), .Q(_49639) );
  nor2s1 _50082_inst ( .DIN1(_49642), .DIN2(_49643), .Q(_49638) );
  nor2s1 _50083_inst ( .DIN1(_49473), .DIN2(_49165), .Q(_49642) );
  nnd2s1 _50084_inst ( .DIN1(_49644), .DIN2(_49645), .Q(____0___________[14])
         );
  nor2s1 _50085_inst ( .DIN1(_49646), .DIN2(_49647), .Q(_49645) );
  nnd2s1 _50086_inst ( .DIN1(_49648), .DIN2(_49649), .Q(_49647) );
  nor2s1 _50087_inst ( .DIN1(_49650), .DIN2(_49651), .Q(_49649) );
  nor2s1 _50088_inst ( .DIN1(_49465), .DIN2(_49128), .Q(_49651) );
  nor2s1 _50089_inst ( .DIN1(_49196), .DIN2(_49498), .Q(_49650) );
  nor2s1 _50090_inst ( .DIN1(_49652), .DIN2(_49175), .Q(_49648) );
  nnd2s1 _50091_inst ( .DIN1(_49584), .DIN2(_49653), .Q(_49175) );
  nnd2s1 _50092_inst ( .DIN1(_49458), .DIN2(_49392), .Q(_49653) );
  nnd2s1 _50093_inst ( .DIN1(_49654), .DIN2(_49655), .Q(_49584) );
  nor2s1 _50094_inst ( .DIN1(_49501), .DIN2(_49656), .Q(_49652) );
  nnd2s1 _50095_inst ( .DIN1(_49657), .DIN2(_49658), .Q(_49646) );
  nor2s1 _50096_inst ( .DIN1(_49659), .DIN2(_49390), .Q(_49658) );
  nor2s1 _50097_inst ( .DIN1(_49660), .DIN2(_49661), .Q(_49657) );
  nor2s1 _50098_inst ( .DIN1(_49344), .DIN2(_49464), .Q(_49661) );
  nor2s1 _50099_inst ( .DIN1(_49127), .DIN2(_49510), .Q(_49660) );
  nor2s1 _50100_inst ( .DIN1(_49662), .DIN2(_49663), .Q(_49644) );
  nnd2s1 _50101_inst ( .DIN1(_49664), .DIN2(_49665), .Q(_49663) );
  nor2s1 _50102_inst ( .DIN1(_49666), .DIN2(_49667), .Q(_49664) );
  nnd2s1 _50103_inst ( .DIN1(_49668), .DIN2(_49669), .Q(_49662) );
  nor2s1 _50104_inst ( .DIN1(_49238), .DIN2(_49347), .Q(_49669) );
  nnd2s1 _50105_inst ( .DIN1(_49670), .DIN2(_49671), .Q(_49347) );
  nnd2s1 _50106_inst ( .DIN1(_49256), .DIN2(_49672), .Q(_49671) );
  nor2s1 _50107_inst ( .DIN1(_49673), .DIN2(_49674), .Q(_49670) );
  nor2s1 _50108_inst ( .DIN1(_49675), .DIN2(_49161), .Q(_49674) );
  nor2s1 _50109_inst ( .DIN1(_49632), .DIN2(_49676), .Q(_49675) );
  nnd2s1 _50110_inst ( .DIN1(_49677), .DIN2(_49579), .Q(_49238) );
  nnd2s1 _50111_inst ( .DIN1(_49407), .DIN2(_49463), .Q(_49579) );
  nnd2s1 _50112_inst ( .DIN1(_49678), .DIN2(_49679), .Q(_49677) );
  nor2s1 _50113_inst ( .DIN1(_49519), .DIN2(_49680), .Q(_49668) );
  nnd2s1 _50114_inst ( .DIN1(_49681), .DIN2(_49682), .Q(_49519) );
  nor2s1 _50115_inst ( .DIN1(_49683), .DIN2(_49684), .Q(_49682) );
  nnd2s1 _50116_inst ( .DIN1(_49685), .DIN2(_49489), .Q(_49684) );
  nnd2s1 _50117_inst ( .DIN1(_49686), .DIN2(_49687), .Q(_49489) );
  nor2s1 _50118_inst ( .DIN1(_49688), .DIN2(_49689), .Q(_49685) );
  nor2s1 _50119_inst ( .DIN1(_49165), .DIN2(_49472), .Q(_49689) );
  and2s1 _50120_inst ( .DIN1(_49609), .DIN2(_49608), .Q(_49688) );
  nnd2s1 _50121_inst ( .DIN1(_49690), .DIN2(_49691), .Q(_49683) );
  nor2s1 _50122_inst ( .DIN1(_49449), .DIN2(_49602), .Q(_49691) );
  and2s1 _50123_inst ( .DIN1(_49569), .DIN2(_49609), .Q(_49449) );
  nor2s1 _50124_inst ( .DIN1(_49628), .DIN2(_49692), .Q(_49690) );
  nor2s1 _50125_inst ( .DIN1(_49693), .DIN2(_49694), .Q(_49681) );
  nnd2s1 _50126_inst ( .DIN1(_49695), .DIN2(_49696), .Q(_49694) );
  nor2s1 _50127_inst ( .DIN1(_49697), .DIN2(_49379), .Q(_49695) );
  nnd2s1 _50128_inst ( .DIN1(_49698), .DIN2(_49699), .Q(_49693) );
  hi1s1 _50129_inst ( .DIN(_49445), .Q(_49699) );
  nor2s1 _50130_inst ( .DIN1(_49700), .DIN2(_49701), .Q(_49698) );
  nor2s1 _50131_inst ( .DIN1(_49218), .DIN2(_49228), .Q(_49700) );
  nnd2s1 _50132_inst ( .DIN1(_49702), .DIN2(_49703), .Q(____0___________[13])
         );
  nor2s1 _50133_inst ( .DIN1(_49704), .DIN2(_49705), .Q(_49703) );
  nnd2s1 _50134_inst ( .DIN1(_49706), .DIN2(_49707), .Q(_49705) );
  hi1s1 _50135_inst ( .DIN(_49453), .Q(_49707) );
  nor2s1 _50136_inst ( .DIN1(_49708), .DIN2(_49709), .Q(_49706) );
  nor2s1 _50137_inst ( .DIN1(_49187), .DIN2(_49710), .Q(_49709) );
  nor2s1 _50138_inst ( .DIN1(_49196), .DIN2(_49315), .Q(_49708) );
  nnd2s1 _50139_inst ( .DIN1(_49711), .DIN2(_49712), .Q(_49704) );
  nor2s1 _50140_inst ( .DIN1(_49191), .DIN2(_49506), .Q(_49712) );
  nor2s1 _50141_inst ( .DIN1(_49713), .DIN2(_49618), .Q(_49711) );
  nor2s1 _50142_inst ( .DIN1(_49117), .DIN2(_49714), .Q(_49618) );
  nor2s1 _50143_inst ( .DIN1(_49715), .DIN2(_49716), .Q(_49702) );
  nnd2s1 _50144_inst ( .DIN1(_49717), .DIN2(_49718), .Q(_49716) );
  nor2s1 _50145_inst ( .DIN1(_49415), .DIN2(_49719), .Q(_49717) );
  nnd2s1 _50146_inst ( .DIN1(_49720), .DIN2(_49721), .Q(_49415) );
  nnd2s1 _50147_inst ( .DIN1(_49722), .DIN2(_49723), .Q(_49721) );
  nor2s1 _50148_inst ( .DIN1(_49602), .DIN2(_49724), .Q(_49720) );
  nor2s1 _50149_inst ( .DIN1(_49451), .DIN2(_49279), .Q(_49724) );
  nor2s1 _50150_inst ( .DIN1(_49725), .DIN2(_49726), .Q(_49602) );
  nnd2s1 _50151_inst ( .DIN1(_49727), .DIN2(_49728), .Q(_49715) );
  hi1s1 _50152_inst ( .DIN(_49327), .Q(_49728) );
  nnd2s1 _50153_inst ( .DIN1(_49729), .DIN2(_49730), .Q(_49327) );
  nor2s1 _50154_inst ( .DIN1(_49731), .DIN2(_49732), .Q(_49730) );
  nnd2s1 _50155_inst ( .DIN1(_49733), .DIN2(_49516), .Q(_49732) );
  nnd2s1 _50156_inst ( .DIN1(_49734), .DIN2(_49687), .Q(_49516) );
  nor2s1 _50157_inst ( .DIN1(_49735), .DIN2(_49736), .Q(_49733) );
  nor2s1 _50158_inst ( .DIN1(_49393), .DIN2(_49187), .Q(_49736) );
  hi1s1 _50159_inst ( .DIN(_49737), .Q(_49393) );
  nor2s1 _50160_inst ( .DIN1(_49344), .DIN2(_49738), .Q(_49735) );
  nnd2s1 _50161_inst ( .DIN1(_49739), .DIN2(_49740), .Q(_49731) );
  nor2s1 _50162_inst ( .DIN1(_49560), .DIN2(_49390), .Q(_49739) );
  nor2s1 _50163_inst ( .DIN1(_49741), .DIN2(_49161), .Q(_49390) );
  nor2s1 _50164_inst ( .DIN1(_49742), .DIN2(_49743), .Q(_49729) );
  nnd2s1 _50165_inst ( .DIN1(_49744), .DIN2(_49745), .Q(_49743) );
  hi1s1 _50166_inst ( .DIN(_49291), .Q(_49745) );
  nnd2s1 _50167_inst ( .DIN1(_49746), .DIN2(_49747), .Q(_49291) );
  or2s1 _50168_inst ( .DIN1(_49166), .DIN2(_49165), .Q(_49747) );
  nnd2s1 _50169_inst ( .DIN1(_49748), .DIN2(_49679), .Q(_49746) );
  nnd2s1 _50170_inst ( .DIN1(_49749), .DIN2(_49544), .Q(_49742) );
  nor2s1 _50171_inst ( .DIN1(_49750), .DIN2(_49446), .Q(_49749) );
  nnd2s1 _50172_inst ( .DIN1(_49751), .DIN2(_49752), .Q(_49446) );
  nnd2s1 _50173_inst ( .DIN1(_49753), .DIN2(_49754), .Q(_49752) );
  nor2s1 _50174_inst ( .DIN1(_49536), .DIN2(_49273), .Q(_49751) );
  nor2s1 _50175_inst ( .DIN1(_49726), .DIN2(_49755), .Q(_49273) );
  nor2s1 _50176_inst ( .DIN1(_49726), .DIN2(_49756), .Q(_49536) );
  nor2s1 _50177_inst ( .DIN1(_49255), .DIN2(_49757), .Q(_49750) );
  nor2s1 _50178_inst ( .DIN1(_49443), .DIN2(_49758), .Q(_49727) );
  nnd2s1 _50179_inst ( .DIN1(_49759), .DIN2(_49760), .Q(____0___________[12])
         );
  nor2s1 _50180_inst ( .DIN1(_49761), .DIN2(_49762), .Q(_49760) );
  nnd2s1 _50181_inst ( .DIN1(_49763), .DIN2(_49764), .Q(_49762) );
  nor2s1 _50182_inst ( .DIN1(_49765), .DIN2(_49766), .Q(_49764) );
  nor2s1 _50183_inst ( .DIN1(_49451), .DIN2(_49757), .Q(_49766) );
  nor2s1 _50184_inst ( .DIN1(_49149), .DIN2(_49472), .Q(_49765) );
  nor2s1 _50185_inst ( .DIN1(_49767), .DIN2(_49133), .Q(_49763) );
  nnd2s1 _50186_inst ( .DIN1(_49768), .DIN2(_49769), .Q(_49133) );
  nor2s1 _50187_inst ( .DIN1(_49770), .DIN2(_49771), .Q(_49769) );
  nnd2s1 _50188_inst ( .DIN1(_49772), .DIN2(_49284), .Q(_49771) );
  nor2s1 _50189_inst ( .DIN1(_49149), .DIN2(_49249), .Q(_49770) );
  nor2s1 _50190_inst ( .DIN1(_49314), .DIN2(_49773), .Q(_49768) );
  nnd2s1 _50191_inst ( .DIN1(_49353), .DIN2(_49245), .Q(_49773) );
  and2s1 _50192_inst ( .DIN1(_49774), .DIN2(_49775), .Q(_49245) );
  or2s1 _50193_inst ( .DIN1(_49741), .DIN2(_49776), .Q(_49775) );
  or2s1 _50194_inst ( .DIN1(_49117), .DIN2(_49156), .Q(_49774) );
  hi1s1 _50195_inst ( .DIN(_49701), .Q(_49353) );
  nnd2s1 _50196_inst ( .DIN1(_49777), .DIN2(_49778), .Q(_49701) );
  nnd2s1 _50197_inst ( .DIN1(_49633), .DIN2(_49779), .Q(_49778) );
  nnd2s1 _50198_inst ( .DIN1(_49780), .DIN2(_49781), .Q(_49777) );
  nnd2s1 _50199_inst ( .DIN1(_49222), .DIN2(_49782), .Q(_49314) );
  nnd2s1 _50200_inst ( .DIN1(_49679), .DIN2(_49654), .Q(_49782) );
  hi1s1 _50201_inst ( .DIN(_49195), .Q(_49654) );
  nor2s1 _50202_inst ( .DIN1(_49783), .DIN2(_49784), .Q(_49767) );
  nnd2s1 _50203_inst ( .DIN1(_49785), .DIN2(_49786), .Q(_49761) );
  nor2s1 _50204_inst ( .DIN1(_49282), .DIN2(_49787), .Q(_49786) );
  or2s1 _50205_inst ( .DIN1(_49440), .DIN2(_49640), .Q(_49787) );
  nor2s1 _50206_inst ( .DIN1(_49788), .DIN2(_49789), .Q(_49785) );
  nor2s1 _50207_inst ( .DIN1(_49790), .DIN2(_49791), .Q(_49759) );
  nnd2s1 _50208_inst ( .DIN1(_49792), .DIN2(_49793), .Q(_49791) );
  nor2s1 _50209_inst ( .DIN1(_49379), .DIN2(_49523), .Q(_49793) );
  nnd2s1 _50210_inst ( .DIN1(_49794), .DIN2(_49795), .Q(_49379) );
  nnd2s1 _50211_inst ( .DIN1(_49462), .DIN2(_49392), .Q(_49795) );
  nor2s1 _50212_inst ( .DIN1(_49192), .DIN2(_49796), .Q(_49794) );
  and2s1 _50213_inst ( .DIN1(_49797), .DIN2(_49798), .Q(_49192) );
  nor2s1 _50214_inst ( .DIN1(_49365), .DIN2(_49680), .Q(_49792) );
  nnd2s1 _50215_inst ( .DIN1(_49799), .DIN2(_49800), .Q(_49680) );
  nor2s1 _50216_inst ( .DIN1(_49374), .DIN2(_49801), .Q(_49800) );
  or2s1 _50217_inst ( .DIN1(_49320), .DIN2(_49486), .Q(_49801) );
  nor2s1 _50218_inst ( .DIN1(_49405), .DIN2(_49117), .Q(_49486) );
  nor2s1 _50219_inst ( .DIN1(_49710), .DIN2(_49196), .Q(_49320) );
  nor2s1 _50220_inst ( .DIN1(_49574), .DIN2(_49802), .Q(_49799) );
  nnd2s1 _50221_inst ( .DIN1(_49803), .DIN2(_49285), .Q(_49802) );
  nnd2s1 _50222_inst ( .DIN1(_49804), .DIN2(_49805), .Q(_49285) );
  nnd2s1 _50223_inst ( .DIN1(_49806), .DIN2(_49399), .Q(_49803) );
  nnd2s1 _50224_inst ( .DIN1(_49397), .DIN2(_49807), .Q(_49574) );
  nnd2s1 _50225_inst ( .DIN1(_49459), .DIN2(_49805), .Q(_49807) );
  nnd2s1 _50226_inst ( .DIN1(_49808), .DIN2(_49798), .Q(_49397) );
  hi1s1 _50227_inst ( .DIN(_49312), .Q(_49808) );
  nnd2s1 _50228_inst ( .DIN1(_49809), .DIN2(_49810), .Q(_49365) );
  nnd2s1 _50229_inst ( .DIN1(_49748), .DIN2(_49655), .Q(_49810) );
  hi1s1 _50230_inst ( .DIN(_49228), .Q(_49748) );
  nor2s1 _50231_inst ( .DIN1(_49283), .DIN2(_49811), .Q(_49809) );
  and2s1 _50232_inst ( .DIN1(_49812), .DIN2(_49813), .Q(_49283) );
  nor2s1 _50233_inst ( .DIN1(_49726), .DIN2(_49814), .Q(_49812) );
  nnd2s1 _50234_inst ( .DIN1(_49815), .DIN2(_49816), .Q(_49790) );
  nor2s1 _50235_inst ( .DIN1(_49262), .DIN2(_49172), .Q(_49816) );
  nnd2s1 _50236_inst ( .DIN1(_49817), .DIN2(_49818), .Q(_49172) );
  nor2s1 _50237_inst ( .DIN1(_49819), .DIN2(_49820), .Q(_49818) );
  nnd2s1 _50238_inst ( .DIN1(_49821), .DIN2(_49822), .Q(_49820) );
  nnd2s1 _50239_inst ( .DIN1(_49823), .DIN2(_49612), .Q(_49819) );
  nor2s1 _50240_inst ( .DIN1(_49476), .DIN2(_49824), .Q(_49823) );
  nor2s1 _50241_inst ( .DIN1(_49825), .DIN2(_49826), .Q(_49817) );
  or2s1 _50242_inst ( .DIN1(_49296), .DIN2(_49615), .Q(_49826) );
  nnd2s1 _50243_inst ( .DIN1(_49827), .DIN2(_49828), .Q(_49615) );
  nnd2s1 _50244_inst ( .DIN1(_49391), .DIN2(_49798), .Q(_49828) );
  hi1s1 _50245_inst ( .DIN(_49738), .Q(_49391) );
  or2s1 _50246_inst ( .DIN1(_49498), .DIN2(_49187), .Q(_49827) );
  nnd2s1 _50247_inst ( .DIN1(_49829), .DIN2(_49830), .Q(_49296) );
  or2s1 _50248_inst ( .DIN1(_49315), .DIN2(_49196), .Q(_49830) );
  nor2s1 _50249_inst ( .DIN1(_49321), .DIN2(_49628), .Q(_49829) );
  nor2s1 _50250_inst ( .DIN1(_49197), .DIN2(_49187), .Q(_49628) );
  and2s1 _50251_inst ( .DIN1(_49831), .DIN2(_49399), .Q(_49321) );
  nnd2s1 _50252_inst ( .DIN1(_49832), .DIN2(_49833), .Q(_49825) );
  hi1s1 _50253_inst ( .DIN(_49697), .Q(_49833) );
  nnd2s1 _50254_inst ( .DIN1(_49834), .DIN2(_49835), .Q(_49697) );
  nnd2s1 _50255_inst ( .DIN1(_49398), .DIN2(_49457), .Q(_49835) );
  nor2s1 _50256_inst ( .DIN1(_49487), .DIN2(_49836), .Q(_49832) );
  nor2s1 _50257_inst ( .DIN1(_49255), .DIN2(_48130), .Q(_49836) );
  nor2s1 _50258_inst ( .DIN1(_49155), .DIN2(_49118), .Q(_49487) );
  or2s1 _50259_inst ( .DIN1(_49837), .DIN2(_49331), .Q(_49262) );
  nnd2s1 _50260_inst ( .DIN1(_49838), .DIN2(_49839), .Q(_49331) );
  or2s1 _50261_inst ( .DIN1(_49840), .DIN2(_49218), .Q(_49839) );
  nnd2s1 _50262_inst ( .DIN1(_49841), .DIN2(_49780), .Q(_49838) );
  or2s1 _50263_inst ( .DIN1(_49842), .DIN2(_49641), .Q(_49837) );
  nor2s1 _50264_inst ( .DIN1(_49501), .DIN2(_49275), .Q(_49641) );
  nor2s1 _50265_inst ( .DIN1(_49465), .DIN2(_49843), .Q(_49842) );
  nor2s1 _50266_inst ( .DIN1(_49844), .DIN2(_49845), .Q(_49815) );
  nnd2s1 _50267_inst ( .DIN1(_49846), .DIN2(_49847), .Q(____0___________[11])
         );
  nor2s1 _50268_inst ( .DIN1(_49848), .DIN2(_49849), .Q(_49847) );
  nnd2s1 _50269_inst ( .DIN1(_49850), .DIN2(_49851), .Q(_49849) );
  hi1s1 _50270_inst ( .DIN(_49203), .Q(_49851) );
  nnd2s1 _50271_inst ( .DIN1(_49852), .DIN2(_49853), .Q(_49203) );
  nor2s1 _50272_inst ( .DIN1(_49854), .DIN2(_49855), .Q(_49853) );
  nnd2s1 _50273_inst ( .DIN1(_49856), .DIN2(_49857), .Q(_49855) );
  or2s1 _50274_inst ( .DIN1(_49560), .DIN2(_49824), .Q(_49854) );
  hi1s1 _50275_inst ( .DIN(_49772), .Q(_49560) );
  nnd2s1 _50276_inst ( .DIN1(_49553), .DIN2(_49686), .Q(_49772) );
  nor2s1 _50277_inst ( .DIN1(_49844), .DIN2(_49858), .Q(_49852) );
  nnd2s1 _50278_inst ( .DIN1(_49466), .DIN2(_49859), .Q(_49858) );
  hi1s1 _50279_inst ( .DIN(_49443), .Q(_49859) );
  nnd2s1 _50280_inst ( .DIN1(_49860), .DIN2(_49861), .Q(_49443) );
  nnd2s1 _50281_inst ( .DIN1(_49537), .DIN2(_49862), .Q(_49861) );
  nor2s1 _50282_inst ( .DIN1(_49540), .DIN2(_49863), .Q(_49862) );
  nnd2s1 _50283_inst ( .DIN1(_49754), .DIN2(_49864), .Q(_49863) );
  nor2s1 _50284_inst ( .DIN1(_49865), .DIN2(_49866), .Q(_49537) );
  nnd2s1 _50285_inst ( .DIN1(_49867), .DIN2(_49813), .Q(_49860) );
  hi1s1 _50286_inst ( .DIN(_49868), .Q(_49813) );
  nor2s1 _50287_inst ( .DIN1(_49465), .DIN2(_49814), .Q(_49867) );
  hi1s1 _50288_inst ( .DIN(_49869), .Q(_49814) );
  and2s1 _50289_inst ( .DIN1(_49870), .DIN2(_49871), .Q(_49466) );
  nnd2s1 _50290_inst ( .DIN1(_49737), .DIN2(_49687), .Q(_49871) );
  nnd2s1 _50291_inst ( .DIN1(_49498), .DIN2(_49510), .Q(_49737) );
  nnd2s1 _50292_inst ( .DIN1(_49872), .DIN2(_26210), .Q(_49510) );
  nnd2s1 _50293_inst ( .DIN1(_49873), .DIN2(_49874), .Q(_49872) );
  nnd2s1 _50294_inst ( .DIN1(_49875), .DIN2(_49876), .Q(_49874) );
  nor2s1 _50295_inst ( .DIN1(_2175), .DIN2(_49877), .Q(_49876) );
  nnd2s1 _50296_inst ( .DIN1(_26223), .DIN2(_49864), .Q(_49877) );
  nor2s1 _50297_inst ( .DIN1(_49878), .DIN2(_49879), .Q(_49875) );
  nnd2s1 _50298_inst ( .DIN1(_49880), .DIN2(_49881), .Q(_49873) );
  nor2s1 _50299_inst ( .DIN1(_49882), .DIN2(_49883), .Q(_49880) );
  nor2s1 _50300_inst ( .DIN1(_49506), .DIN2(_49692), .Q(_49870) );
  nor2s1 _50301_inst ( .DIN1(_49884), .DIN2(_49738), .Q(_49692) );
  nnd2s1 _50302_inst ( .DIN1(_49885), .DIN2(_49886), .Q(_49738) );
  nor2s1 _50303_inst ( .DIN1(_26210), .DIN2(_49887), .Q(_49885) );
  nor2s1 _50304_inst ( .DIN1(_49312), .DIN2(_49884), .Q(_49506) );
  nnd2s1 _50305_inst ( .DIN1(_49888), .DIN2(_49889), .Q(_49312) );
  nor2s1 _50306_inst ( .DIN1(_2175), .DIN2(_49890), .Q(_49889) );
  nnd2s1 _50307_inst ( .DIN1(_26223), .DIN2(_26210), .Q(_49890) );
  nor2s1 _50308_inst ( .DIN1(_49887), .DIN2(_49891), .Q(_49888) );
  nnd2s1 _50309_inst ( .DIN1(_2273), .DIN2(_49892), .Q(_49891) );
  nor2s1 _50310_inst ( .DIN1(_49620), .DIN2(_49596), .Q(_49850) );
  hi1s1 _50311_inst ( .DIN(_49893), .Q(_49596) );
  nnd2s1 _50312_inst ( .DIN1(_49894), .DIN2(_49895), .Q(_49620) );
  or2s1 _50313_inst ( .DIN1(_49344), .DIN2(_49896), .Q(_49895) );
  nnd2s1 _50314_inst ( .DIN1(_49672), .DIN2(_49841), .Q(_49894) );
  nnd2s1 _50315_inst ( .DIN1(_49897), .DIN2(_49898), .Q(_49848) );
  nor2s1 _50316_inst ( .DIN1(_49440), .DIN2(_49123), .Q(_49898) );
  nor2s1 _50317_inst ( .DIN1(_49634), .DIN2(_49899), .Q(_49897) );
  nor2s1 _50318_inst ( .DIN1(_49451), .DIN2(_49900), .Q(_49899) );
  nor2s1 _50319_inst ( .DIN1(_49901), .DIN2(_49902), .Q(_49846) );
  nnd2s1 _50320_inst ( .DIN1(_49903), .DIN2(_49718), .Q(_49902) );
  and2s1 _50321_inst ( .DIN1(_49904), .DIN2(_49905), .Q(_49718) );
  nor2s1 _50322_inst ( .DIN1(_49906), .DIN2(_49907), .Q(_49905) );
  nnd2s1 _50323_inst ( .DIN1(_49908), .DIN2(_49909), .Q(_49907) );
  nnd2s1 _50324_inst ( .DIN1(_49910), .DIN2(_49911), .Q(_49909) );
  nnd2s1 _50325_inst ( .DIN1(_49128), .DIN2(_49197), .Q(_49911) );
  nnd2s1 _50326_inst ( .DIN1(_49912), .DIN2(_49913), .Q(_49197) );
  nor2s1 _50327_inst ( .DIN1(_49914), .DIN2(_49915), .Q(_49913) );
  nor2s1 _50328_inst ( .DIN1(_49866), .DIN2(_49868), .Q(_49912) );
  nnd2s1 _50329_inst ( .DIN1(_2273), .DIN2(_49916), .Q(_49868) );
  nnd2s1 _50330_inst ( .DIN1(_49462), .DIN2(_49798), .Q(_49908) );
  hi1s1 _50331_inst ( .DIN(_49562), .Q(_49462) );
  nnd2s1 _50332_inst ( .DIN1(_49917), .DIN2(_49918), .Q(_49562) );
  nor2s1 _50333_inst ( .DIN1(_49311), .DIN2(_49464), .Q(_49906) );
  nnd2s1 _50334_inst ( .DIN1(_49886), .DIN2(_49919), .Q(_49464) );
  and2s1 _50335_inst ( .DIN1(_49920), .DIN2(_49921), .Q(_49886) );
  nor2s1 _50336_inst ( .DIN1(_26419), .DIN2(_26223), .Q(_49921) );
  nor2s1 _50337_inst ( .DIN1(_49878), .DIN2(_49864), .Q(_49920) );
  nor2s1 _50338_inst ( .DIN1(_49922), .DIN2(_49923), .Q(_49904) );
  nnd2s1 _50339_inst ( .DIN1(_49524), .DIN2(_49924), .Q(_49923) );
  nnd2s1 _50340_inst ( .DIN1(_49925), .DIN2(_49301), .Q(_49924) );
  nnd2s1 _50341_inst ( .DIN1(_49300), .DIN2(_49754), .Q(_49524) );
  nor2s1 _50342_inst ( .DIN1(_49328), .DIN2(_49666), .Q(_49903) );
  nnd2s1 _50343_inst ( .DIN1(_49926), .DIN2(_49927), .Q(_49666) );
  hi1s1 _50344_inst ( .DIN(_49928), .Q(_49927) );
  nor2s1 _50345_inst ( .DIN1(_49929), .DIN2(_49930), .Q(_49926) );
  nor2s1 _50346_inst ( .DIN1(_49931), .DIN2(_49165), .Q(_49930) );
  nor2s1 _50347_inst ( .DIN1(_49532), .DIN2(_49753), .Q(_49931) );
  hi1s1 _50348_inst ( .DIN(_49278), .Q(_49753) );
  nnd2s1 _50349_inst ( .DIN1(_49932), .DIN2(_49933), .Q(_49328) );
  nor2s1 _50350_inst ( .DIN1(_49354), .DIN2(_49934), .Q(_49933) );
  nnd2s1 _50351_inst ( .DIN1(_49258), .DIN2(_49935), .Q(_49934) );
  nor2s1 _50352_inst ( .DIN1(_49255), .DIN2(_49755), .Q(_49354) );
  nor2s1 _50353_inst ( .DIN1(_49126), .DIN2(_49216), .Q(_49932) );
  nor2s1 _50354_inst ( .DIN1(_49581), .DIN2(_49150), .Q(_49216) );
  nor2s1 _50355_inst ( .DIN1(_49149), .DIN2(_49473), .Q(_49126) );
  nnd2s1 _50356_inst ( .DIN1(_49936), .DIN2(_49744), .Q(_49901) );
  and2s1 _50357_inst ( .DIN1(_49822), .DIN2(_49937), .Q(_49744) );
  nnd2s1 _50358_inst ( .DIN1(_49398), .DIN2(_49551), .Q(_49937) );
  hi1s1 _50359_inst ( .DIN(_49611), .Q(_49398) );
  nnd2s1 _50360_inst ( .DIN1(_49938), .DIN2(_49881), .Q(_49611) );
  nor2s1 _50361_inst ( .DIN1(_26210), .DIN2(_49865), .Q(_49938) );
  nnd2s1 _50362_inst ( .DIN1(_49722), .DIN2(_49608), .Q(_49822) );
  hi1s1 _50363_inst ( .DIN(_49400), .Q(_49608) );
  nnd2s1 _50364_inst ( .DIN1(_49939), .DIN2(_49940), .Q(_49400) );
  nor2s1 _50365_inst ( .DIN1(_49864), .DIN2(_49941), .Q(_49940) );
  nnd2s1 _50366_inst ( .DIN1(_49942), .DIN2(_26294), .Q(_49941) );
  nor2s1 _50367_inst ( .DIN1(_49943), .DIN2(_49944), .Q(_49939) );
  nnd2s1 _50368_inst ( .DIN1(_49945), .DIN2(_2216), .Q(_49944) );
  nor2s1 _50369_inst ( .DIN1(_49233), .DIN2(_49290), .Q(_49936) );
  nnd2s1 _50370_inst ( .DIN1(_49946), .DIN2(_49947), .Q(_49290) );
  nor2s1 _50371_inst ( .DIN1(_49948), .DIN2(_49949), .Q(_49947) );
  nnd2s1 _50372_inst ( .DIN1(_49950), .DIN2(_49201), .Q(_49949) );
  nor2s1 _50373_inst ( .DIN1(_49951), .DIN2(_49758), .Q(_49201) );
  nnd2s1 _50374_inst ( .DIN1(_49952), .DIN2(_49953), .Q(_49758) );
  nnd2s1 _50375_inst ( .DIN1(_49408), .DIN2(_49392), .Q(_49953) );
  hi1s1 _50376_inst ( .DIN(_49311), .Q(_49392) );
  nnd2s1 _50377_inst ( .DIN1(_49954), .DIN2(_49955), .Q(_49952) );
  nnd2s1 _50378_inst ( .DIN1(_49336), .DIN2(_49488), .Q(_49951) );
  and2s1 _50379_inst ( .DIN1(_49956), .DIN2(_49957), .Q(_49488) );
  nnd2s1 _50380_inst ( .DIN1(_49722), .DIN2(_49958), .Q(_49957) );
  nor2s1 _50381_inst ( .DIN1(_49453), .DIN2(_49445), .Q(_49950) );
  nnd2s1 _50382_inst ( .DIN1(_49959), .DIN2(_49960), .Q(_49445) );
  nnd2s1 _50383_inst ( .DIN1(_49961), .DIN2(_49533), .Q(_49960) );
  nnd2s1 _50384_inst ( .DIN1(_49257), .DIN2(_49672), .Q(_49959) );
  nnd2s1 _50385_inst ( .DIN1(_49962), .DIN2(_49963), .Q(_49453) );
  nnd2s1 _50386_inst ( .DIN1(_49964), .DIN2(_49457), .Q(_49963) );
  nnd2s1 _50387_inst ( .DIN1(_49518), .DIN2(_49609), .Q(_49962) );
  hi1s1 _50388_inst ( .DIN(_49965), .Q(_49518) );
  nnd2s1 _50389_inst ( .DIN1(_49966), .DIN2(_49967), .Q(_49948) );
  nnd2s1 _50390_inst ( .DIN1(_49968), .DIN2(_49533), .Q(_49967) );
  and2s1 _50391_inst ( .DIN1(_49969), .DIN2(_49377), .Q(_49966) );
  nnd2s1 _50392_inst ( .DIN1(_49722), .DIN2(_49569), .Q(_49377) );
  and2s1 _50393_inst ( .DIN1(_49970), .DIN2(_49881), .Q(_49569) );
  and2s1 _50394_inst ( .DIN1(_49971), .DIN2(_49972), .Q(_49881) );
  nor2s1 _50395_inst ( .DIN1(_49973), .DIN2(_49864), .Q(_49972) );
  nor2s1 _50396_inst ( .DIN1(_49540), .DIN2(_49974), .Q(_49971) );
  nor2s1 _50397_inst ( .DIN1(_2216), .DIN2(_49943), .Q(_49970) );
  nor2s1 _50398_inst ( .DIN1(_49975), .DIN2(_49976), .Q(_49946) );
  or2s1 _50399_inst ( .DIN1(_49977), .DIN2(_49523), .Q(_49976) );
  nnd2s1 _50400_inst ( .DIN1(_49580), .DIN2(_49978), .Q(_49523) );
  nnd2s1 _50401_inst ( .DIN1(_49678), .DIN2(_49633), .Q(_49978) );
  nnd2s1 _50402_inst ( .DIN1(_49979), .DIN2(_49635), .Q(_49975) );
  and2s1 _50403_inst ( .DIN1(_49980), .DIN2(_49981), .Q(_49635) );
  nnd2s1 _50404_inst ( .DIN1(_49256), .DIN2(_49780), .Q(_49981) );
  hi1s1 _50405_inst ( .DIN(_49452), .Q(_49256) );
  nnd2s1 _50406_inst ( .DIN1(_49982), .DIN2(_49919), .Q(_49452) );
  nor2s1 _50407_inst ( .DIN1(_2273), .DIN2(_49943), .Q(_49982) );
  nnd2s1 _50408_inst ( .DIN1(_49676), .DIN2(_49655), .Q(_49980) );
  nor2s1 _50409_inst ( .DIN1(_49983), .DIN2(_49346), .Q(_49979) );
  nnd2s1 _50410_inst ( .DIN1(_49984), .DIN2(_49985), .Q(_49346) );
  or2s1 _50411_inst ( .DIN1(_49725), .DIN2(_49451), .Q(_49985) );
  nnd2s1 _50412_inst ( .DIN1(_49954), .DIN2(_49637), .Q(_49984) );
  nnd2s1 _50413_inst ( .DIN1(_49986), .DIN2(_49987), .Q(_49233) );
  or2s1 _50414_inst ( .DIN1(_49988), .DIN2(_49152), .Q(_49987) );
  nnd2s1 _50415_inst ( .DIN1(_49550), .DIN2(_49399), .Q(_49986) );
  nnd2s1 _50416_inst ( .DIN1(_49989), .DIN2(_49990), .Q(____0___________[10])
         );
  nor2s1 _50417_inst ( .DIN1(_49991), .DIN2(_49992), .Q(_49990) );
  nnd2s1 _50418_inst ( .DIN1(_49993), .DIN2(_49994), .Q(_49992) );
  nor2s1 _50419_inst ( .DIN1(_49995), .DIN2(_49163), .Q(_49994) );
  nor2s1 _50420_inst ( .DIN1(_49344), .DIN2(_49996), .Q(_49163) );
  hi1s1 _50421_inst ( .DIN(_49407), .Q(_49996) );
  nor2s1 _50422_inst ( .DIN1(_49943), .DIN2(_49997), .Q(_49407) );
  nor2s1 _50423_inst ( .DIN1(_49465), .DIN2(_49998), .Q(_49995) );
  nor2s1 _50424_inst ( .DIN1(_49925), .DIN2(_49806), .Q(_49998) );
  hi1s1 _50425_inst ( .DIN(_49714), .Q(_49806) );
  hi1s1 _50426_inst ( .DIN(_49472), .Q(_49925) );
  nnd2s1 _50427_inst ( .DIN1(_49918), .DIN2(_49999), .Q(_49472) );
  nor2s1 _50428_inst ( .DIN1(_50000), .DIN2(_50001), .Q(_49993) );
  nor2s1 _50429_inst ( .DIN1(_49127), .DIN2(_49498), .Q(_50001) );
  nnd2s1 _50430_inst ( .DIN1(_50002), .DIN2(_49869), .Q(_49498) );
  nor2s1 _50431_inst ( .DIN1(_50003), .DIN2(_49879), .Q(_49869) );
  nnd2s1 _50432_inst ( .DIN1(_50004), .DIN2(_2216), .Q(_50003) );
  nor2s1 _50433_inst ( .DIN1(_2273), .DIN2(_50005), .Q(_50002) );
  nor2s1 _50434_inst ( .DIN1(_49965), .DIN2(_49152), .Q(_50000) );
  nnd2s1 _50435_inst ( .DIN1(_50006), .DIN2(_49917), .Q(_49965) );
  hi1s1 _50436_inst ( .DIN(_50007), .Q(_49917) );
  nor2s1 _50437_inst ( .DIN1(_49882), .DIN2(_49914), .Q(_50006) );
  nnd2s1 _50438_inst ( .DIN1(_50008), .DIN2(_50009), .Q(_49991) );
  nor2s1 _50439_inst ( .DIN1(_49788), .DIN2(_50010), .Q(_50009) );
  nnd2s1 _50440_inst ( .DIN1(_49834), .DIN2(_49956), .Q(_50010) );
  hi1s1 _50441_inst ( .DIN(_49592), .Q(_49834) );
  and2s1 _50442_inst ( .DIN1(_49553), .DIN2(_50011), .Q(_49788) );
  nnd2s1 _50443_inst ( .DIN1(_49128), .DIN2(_49188), .Q(_50011) );
  nor2s1 _50444_inst ( .DIN1(_50012), .DIN2(_50013), .Q(_50008) );
  nor2s1 _50445_inst ( .DIN1(_50014), .DIN2(_49776), .Q(_50013) );
  nor2s1 _50446_inst ( .DIN1(_49964), .DIN2(_49632), .Q(_50014) );
  hi1s1 _50447_inst ( .DIN(_49162), .Q(_49964) );
  nnd2s1 _50448_inst ( .DIN1(_50015), .DIN2(_50016), .Q(_49162) );
  nor2s1 _50449_inst ( .DIN1(_49864), .DIN2(_49540), .Q(_50016) );
  nor2s1 _50450_inst ( .DIN1(_49943), .DIN2(_49866), .Q(_50015) );
  nnd2s1 _50451_inst ( .DIN1(_50017), .DIN2(_50018), .Q(_49866) );
  nor2s1 _50452_inst ( .DIN1(_49973), .DIN2(_50019), .Q(_50018) );
  nnd2s1 _50453_inst ( .DIN1(_26433), .DIN2(_26217), .Q(_50019) );
  nor2s1 _50454_inst ( .DIN1(_26646), .DIN2(_50020), .Q(_50017) );
  nnd2s1 _50455_inst ( .DIN1(_2216), .DIN2(_50021), .Q(_50020) );
  nor2s1 _50456_inst ( .DIN1(_50022), .DIN2(_49783), .Q(_50012) );
  nor2s1 _50457_inst ( .DIN1(_49342), .DIN2(_49968), .Q(_50022) );
  hi1s1 _50458_inst ( .DIN(_49227), .Q(_49968) );
  nor2s1 _50459_inst ( .DIN1(_50023), .DIN2(_50024), .Q(_49989) );
  nnd2s1 _50460_inst ( .DIN1(_50025), .DIN2(_50026), .Q(_50024) );
  nor2s1 _50461_inst ( .DIN1(_50027), .DIN2(_50028), .Q(_50026) );
  hi1s1 _50462_inst ( .DIN(_49573), .Q(_50028) );
  nor2s1 _50463_inst ( .DIN1(_50029), .DIN2(_50030), .Q(_49573) );
  or2s1 _50464_inst ( .DIN1(_50031), .DIN2(_49444), .Q(_50029) );
  nor2s1 _50465_inst ( .DIN1(_49117), .DIN2(_49656), .Q(_50031) );
  nor2s1 _50466_inst ( .DIN1(_49667), .DIN2(_49922), .Q(_50025) );
  nnd2s1 _50467_inst ( .DIN1(_50032), .DIN2(_50033), .Q(_49922) );
  nnd2s1 _50468_inst ( .DIN1(_49459), .DIN2(_49533), .Q(_50033) );
  nor2s1 _50469_inst ( .DIN1(_49865), .DIN2(_49997), .Q(_49459) );
  nnd2s1 _50470_inst ( .DIN1(_49458), .DIN2(_49798), .Q(_50032) );
  and2s1 _50471_inst ( .DIN1(_50034), .DIN2(_50035), .Q(_49458) );
  nor2s1 _50472_inst ( .DIN1(_2179), .DIN2(_2175), .Q(_50035) );
  nor2s1 _50473_inst ( .DIN1(_49878), .DIN2(_50007), .Q(_50034) );
  nnd2s1 _50474_inst ( .DIN1(_50036), .DIN2(_50037), .Q(_50007) );
  hi1s1 _50475_inst ( .DIN(_49892), .Q(_49878) );
  nnd2s1 _50476_inst ( .DIN1(_50038), .DIN2(_50039), .Q(_49667) );
  nor2s1 _50477_inst ( .DIN1(_50040), .DIN2(_50041), .Q(_50039) );
  nnd2s1 _50478_inst ( .DIN1(_49336), .DIN2(_49475), .Q(_50041) );
  hi1s1 _50479_inst ( .DIN(_49811), .Q(_49475) );
  nor2s1 _50480_inst ( .DIN1(_50042), .DIN2(_49161), .Q(_49811) );
  or2s1 _50481_inst ( .DIN1(_49621), .DIN2(_49196), .Q(_49336) );
  nnd2s1 _50482_inst ( .DIN1(_50043), .DIN2(_49222), .Q(_50040) );
  nnd2s1 _50483_inst ( .DIN1(_49301), .DIN2(_49955), .Q(_49222) );
  nor2s1 _50484_inst ( .DIN1(_49440), .DIN2(_49191), .Q(_50043) );
  and2s1 _50485_inst ( .DIN1(_50044), .DIN2(_50045), .Q(_49191) );
  nor2s1 _50486_inst ( .DIN1(_29741), .DIN2(_49161), .Q(_50044) );
  nor2s1 _50487_inst ( .DIN1(_50046), .DIN2(_50047), .Q(_50038) );
  nnd2s1 _50488_inst ( .DIN1(_50048), .DIN2(_50049), .Q(_50047) );
  nnd2s1 _50489_inst ( .DIN1(_49547), .DIN2(_49754), .Q(_50049) );
  hi1s1 _50490_inst ( .DIN(_49249), .Q(_49547) );
  nnd2s1 _50491_inst ( .DIN1(_50050), .DIN2(_49919), .Q(_49249) );
  hi1s1 _50492_inst ( .DIN(_50051), .Q(_49919) );
  and2s1 _50493_inst ( .DIN1(_2273), .DIN2(_49918), .Q(_50050) );
  nor2s1 _50494_inst ( .DIN1(_49883), .DIN2(_50005), .Q(_49918) );
  hi1s1 _50495_inst ( .DIN(_49265), .Q(_50048) );
  nnd2s1 _50496_inst ( .DIN1(_50052), .DIN2(_50053), .Q(_49265) );
  nnd2s1 _50497_inst ( .DIN1(_49552), .DIN2(_49910), .Q(_50053) );
  hi1s1 _50498_inst ( .DIN(_50054), .Q(_49552) );
  nor2s1 _50499_inst ( .DIN1(_50055), .DIN2(_50056), .Q(_50052) );
  nnd2s1 _50500_inst ( .DIN1(_50057), .DIN2(_49605), .Q(_50046) );
  nnd2s1 _50501_inst ( .DIN1(_49408), .DIN2(_49798), .Q(_50057) );
  and2s1 _50502_inst ( .DIN1(_50058), .DIN2(_50059), .Q(_49408) );
  nor2s1 _50503_inst ( .DIN1(_2273), .DIN2(_49882), .Q(_50059) );
  nor2s1 _50504_inst ( .DIN1(_49883), .DIN2(_50051), .Q(_50058) );
  nnd2s1 _50505_inst ( .DIN1(_50060), .DIN2(_50061), .Q(_50051) );
  nor2s1 _50506_inst ( .DIN1(_50062), .DIN2(_50063), .Q(_50061) );
  nnd2s1 _50507_inst ( .DIN1(_26248), .DIN2(_26210), .Q(_50063) );
  nnd2s1 _50508_inst ( .DIN1(_26294), .DIN2(_26217), .Q(_50062) );
  nor2s1 _50509_inst ( .DIN1(_50064), .DIN2(_50065), .Q(_50060) );
  nnd2s1 _50510_inst ( .DIN1(_2274), .DIN2(_2217), .Q(_50065) );
  nnd2s1 _50511_inst ( .DIN1(_2214), .DIN2(_49942), .Q(_50064) );
  nnd2s1 _50512_inst ( .DIN1(_50066), .DIN2(_50067), .Q(_50023) );
  nor2s1 _50513_inst ( .DIN1(_49261), .DIN2(_50068), .Q(_50067) );
  nnd2s1 _50514_inst ( .DIN1(_50069), .DIN2(_50070), .Q(_50068) );
  nnd2s1 _50515_inst ( .DIN1(_49954), .DIN2(_49300), .Q(_50070) );
  hi1s1 _50516_inst ( .DIN(_49413), .Q(_49300) );
  nnd2s1 _50517_inst ( .DIN1(_50071), .DIN2(_50072), .Q(_49413) );
  nor2s1 _50518_inst ( .DIN1(_2216), .DIN2(_49864), .Q(_50072) );
  nor2s1 _50519_inst ( .DIN1(_49879), .DIN2(_49865), .Q(_50071) );
  nnd2s1 _50520_inst ( .DIN1(_50004), .DIN2(_50073), .Q(_49865) );
  hi1s1 _50521_inst ( .DIN(_49165), .Q(_49954) );
  hi1s1 _50522_inst ( .DIN(_49134), .Q(_50069) );
  nnd2s1 _50523_inst ( .DIN1(_50074), .DIN2(_50075), .Q(_49134) );
  nor2s1 _50524_inst ( .DIN1(_49824), .DIN2(_49713), .Q(_50074) );
  nor2s1 _50525_inst ( .DIN1(_49161), .DIN2(_49840), .Q(_49713) );
  nor2s1 _50526_inst ( .DIN1(_49756), .DIN2(_49255), .Q(_49824) );
  nnd2s1 _50527_inst ( .DIN1(_49544), .DIN2(_50076), .Q(_49261) );
  and2s1 _50528_inst ( .DIN1(_50077), .DIN2(_50078), .Q(_49544) );
  nnd2s1 _50529_inst ( .DIN1(_49779), .DIN2(_49679), .Q(_50078) );
  hi1s1 _50530_inst ( .DIN(_49161), .Q(_49679) );
  nnd2s1 _50531_inst ( .DIN1(_49672), .DIN2(_49781), .Q(_50077) );
  nor2s1 _50532_inst ( .DIN1(_49234), .DIN2(_49326), .Q(_50066) );
  nnd2s1 _50533_inst ( .DIN1(_50079), .DIN2(_50080), .Q(_49326) );
  nor2s1 _50534_inst ( .DIN1(_50081), .DIN2(_50082), .Q(_50080) );
  or2s1 _50535_inst ( .DIN1(_49796), .DIN2(_49123), .Q(_50082) );
  nor2s1 _50536_inst ( .DIN1(_49155), .DIN2(_49275), .Q(_49123) );
  hi1s1 _50537_inst ( .DIN(_49428), .Q(_49796) );
  nnd2s1 _50538_inst ( .DIN1(_50083), .DIN2(_49798), .Q(_49428) );
  or2s1 _50539_inst ( .DIN1(_49282), .DIN2(_49601), .Q(_50081) );
  nor2s1 _50540_inst ( .DIN1(_50084), .DIN2(_49161), .Q(_49282) );
  nor2s1 _50541_inst ( .DIN1(_50085), .DIN2(_50086), .Q(_50079) );
  or2s1 _50542_inst ( .DIN1(_49239), .DIN2(_49266), .Q(_50086) );
  nnd2s1 _50543_inst ( .DIN1(_49969), .DIN2(_50087), .Q(_49266) );
  nnd2s1 _50544_inst ( .DIN1(_50088), .DIN2(_49722), .Q(_50087) );
  hi1s1 _50545_inst ( .DIN(_49152), .Q(_49722) );
  nnd2s1 _50546_inst ( .DIN1(_49284), .DIN2(_49856), .Q(_49239) );
  nnd2s1 _50547_inst ( .DIN1(_49533), .DIN2(_49804), .Q(_49856) );
  hi1s1 _50548_inst ( .DIN(_49783), .Q(_49533) );
  nnd2s1 _50549_inst ( .DIN1(_49723), .DIN2(_49609), .Q(_49284) );
  nnd2s1 _50550_inst ( .DIN1(_49298), .DIN2(_49535), .Q(_50085) );
  nnd2s1 _50551_inst ( .DIN1(_49375), .DIN2(_49780), .Q(_49298) );
  nnd2s1 _50552_inst ( .DIN1(_50089), .DIN2(_50090), .Q(_49234) );
  nnd2s1 _50553_inst ( .DIN1(_49910), .DIN2(_49686), .Q(_50090) );
  and2s1 _50554_inst ( .DIN1(_50091), .DIN2(_49999), .Q(_49686) );
  hi1s1 _50555_inst ( .DIN(_49997), .Q(_49999) );
  nnd2s1 _50556_inst ( .DIN1(_50092), .DIN2(_50037), .Q(_49997) );
  hi1s1 _50557_inst ( .DIN(_49887), .Q(_50037) );
  nnd2s1 _50558_inst ( .DIN1(_50093), .DIN2(_49945), .Q(_49887) );
  nor2s1 _50559_inst ( .DIN1(_49915), .DIN2(_49973), .Q(_50093) );
  nor2s1 _50560_inst ( .DIN1(_2273), .DIN2(_2216), .Q(_50092) );
  nor2s1 _50561_inst ( .DIN1(_50005), .DIN2(_50094), .Q(_50091) );
  nor2s1 _50562_inst ( .DIN1(_49504), .DIN2(_50095), .Q(_50089) );
  nor2s1 _50563_inst ( .DIN1(_49195), .DIN2(_49776), .Q(_50095) );
  nnd2s1 _50564_inst ( .DIN1(_50096), .DIN2(_50036), .Q(_49195) );
  nor2s1 _50565_inst ( .DIN1(_2273), .DIN2(_26210), .Q(_50036) );
  nor2s1 _50566_inst ( .DIN1(_49943), .DIN2(_49879), .Q(_50096) );
  nnd2s1 _50567_inst ( .DIN1(_50097), .DIN2(_49945), .Q(_49879) );
  hi1s1 _50568_inst ( .DIN(_49974), .Q(_49945) );
  nnd2s1 _50569_inst ( .DIN1(_50098), .DIN2(_50099), .Q(_49974) );
  nor2s1 _50570_inst ( .DIN1(_2214), .DIN2(_50100), .Q(_50099) );
  nnd2s1 _50571_inst ( .DIN1(_26370), .DIN2(_26217), .Q(_50100) );
  nor2s1 _50572_inst ( .DIN1(_26248), .DIN2(_26646), .Q(_50098) );
  nor2s1 _50573_inst ( .DIN1(_50101), .DIN2(_49540), .Q(_50097) );
  nnd2s1 _50574_inst ( .DIN1(_50102), .DIN2(_49916), .Q(_49943) );
  hi1s1 _50575_inst ( .DIN(_49857), .Q(_49504) );
  nnd2s1 _50576_inst ( .DIN1(_50103), .DIN2(_49551), .Q(_49857) );
  hi1s1 _50577_inst ( .DIN(_49117), .Q(_49551) );
  nnd2s1 _50578_inst ( .DIN1(_50104), .DIN2(_50105), .Q(____0___________[0])
         );
  nor2s1 _50579_inst ( .DIN1(_50106), .DIN2(_50107), .Q(_50105) );
  nnd2s1 _50580_inst ( .DIN1(_50108), .DIN2(_50109), .Q(_50107) );
  nor2s1 _50581_inst ( .DIN1(_50110), .DIN2(_50111), .Q(_50109) );
  nnd2s1 _50582_inst ( .DIN1(_50112), .DIN2(_50113), .Q(_50111) );
  nnd2s1 _50583_inst ( .DIN1(_49805), .DIN2(_50114), .Q(_50113) );
  nnd2s1 _50584_inst ( .DIN1(_50115), .DIN2(_50116), .Q(_50114) );
  nnd2s1 _50585_inst ( .DIN1(_49633), .DIN2(_50117), .Q(_50112) );
  nnd2s1 _50586_inst ( .DIN1(_50118), .DIN2(_50119), .Q(_50117) );
  nor2s1 _50587_inst ( .DIN1(_49884), .DIN2(_50120), .Q(_50110) );
  nor2s1 _50588_inst ( .DIN1(_49797), .DIN2(_50083), .Q(_50120) );
  and2s1 _50589_inst ( .DIN1(_50121), .DIN2(_50122), .Q(_50083) );
  nor2s1 _50590_inst ( .DIN1(_34413), .DIN2(_44324), .Q(_50121) );
  and2s1 _50591_inst ( .DIN1(_50123), .DIN2(_50124), .Q(_49797) );
  nor2s1 _50592_inst ( .DIN1(_32091), .DIN2(_32820), .Q(_50123) );
  hi1s1 _50593_inst ( .DIN(_49463), .Q(_49884) );
  nnd2s1 _50594_inst ( .DIN1(_49311), .DIN2(_49344), .Q(_49463) );
  nor2s1 _50595_inst ( .DIN1(_50125), .DIN2(_50126), .Q(_50108) );
  nor2s1 _50596_inst ( .DIN1(_49218), .DIN2(_50127), .Q(_50126) );
  nor2s1 _50597_inst ( .DIN1(_49779), .DIN2(_50128), .Q(_50127) );
  nnd2s1 _50598_inst ( .DIN1(_50084), .DIN2(_50042), .Q(_50128) );
  nnd2s1 _50599_inst ( .DIN1(_50129), .DIN2(_50130), .Q(_50042) );
  nor2s1 _50600_inst ( .DIN1(_32824), .DIN2(_37299), .Q(_50129) );
  nnd2s1 _50601_inst ( .DIN1(_50131), .DIN2(_27308), .Q(_50084) );
  and2s1 _50602_inst ( .DIN1(_30771), .DIN2(_50132), .Q(_50131) );
  hi1s1 _50603_inst ( .DIN(_34855), .Q(_30771) );
  and2s1 _50604_inst ( .DIN1(_50133), .DIN2(_50134), .Q(_49779) );
  nor2s1 _50605_inst ( .DIN1(_38682), .DIN2(_45434), .Q(_50133) );
  hi1s1 _50606_inst ( .DIN(_49655), .Q(_49218) );
  nor2s1 _50607_inst ( .DIN1(_49451), .DIN2(_50135), .Q(_50125) );
  nor2s1 _50608_inst ( .DIN1(_49781), .DIN2(_50136), .Q(_50135) );
  nnd2s1 _50609_inst ( .DIN1(_49756), .DIN2(_49725), .Q(_50136) );
  nnd2s1 _50610_inst ( .DIN1(_50137), .DIN2(_50138), .Q(_49725) );
  nor2s1 _50611_inst ( .DIN1(_30939), .DIN2(_50139), .Q(_50137) );
  nnd2s1 _50612_inst ( .DIN1(_31400), .DIN2(_50140), .Q(_49756) );
  hi1s1 _50613_inst ( .DIN(_32821), .Q(_31400) );
  and2s1 _50614_inst ( .DIN1(_50141), .DIN2(_50142), .Q(_49781) );
  nor2s1 _50615_inst ( .DIN1(_30434), .DIN2(_35720), .Q(_50142) );
  nor2s1 _50616_inst ( .DIN1(_37983), .DIN2(_27446), .Q(_50141) );
  hi1s1 _50617_inst ( .DIN(_49376), .Q(_49451) );
  nnd2s1 _50618_inst ( .DIN1(_49726), .DIN2(_49255), .Q(_49376) );
  nnd2s1 _50619_inst ( .DIN1(_50143), .DIN2(_50144), .Q(_50106) );
  nor2s1 _50620_inst ( .DIN1(_49374), .DIN2(_50145), .Q(_50144) );
  nnd2s1 _50621_inst ( .DIN1(_49591), .DIN2(_49969), .Q(_50145) );
  or2s1 _50622_inst ( .DIN1(_49405), .DIN2(_49501), .Q(_49969) );
  nnd2s1 _50623_inst ( .DIN1(_50140), .DIN2(_27430), .Q(_49405) );
  hi1s1 _50624_inst ( .DIN(_50146), .Q(_27430) );
  hi1s1 _50625_inst ( .DIN(_49359), .Q(_49591) );
  nor2s1 _50626_inst ( .DIN1(_49840), .DIN2(_49776), .Q(_49359) );
  nnd2s1 _50627_inst ( .DIN1(_50147), .DIN2(_50148), .Q(_49840) );
  nor2s1 _50628_inst ( .DIN1(_29741), .DIN2(_33293), .Q(_50148) );
  nor2s1 _50629_inst ( .DIN1(_35721), .DIN2(_30940), .Q(_50147) );
  nor2s1 _50630_inst ( .DIN1(_49166), .DIN2(_49581), .Q(_49374) );
  nnd2s1 _50631_inst ( .DIN1(_50149), .DIN2(_50150), .Q(_49166) );
  nor2s1 _50632_inst ( .DIN1(_35723), .DIN2(_39111), .Q(_50150) );
  nor2s1 _50633_inst ( .DIN1(_50146), .DIN2(_27828), .Q(_50149) );
  nnd2s1 _50634_inst ( .DIN1(_50151), .DIN2(_50073), .Q(_50146) );
  nor2s1 _50635_inst ( .DIN1(_50152), .DIN2(_50153), .Q(_50143) );
  nor2s1 _50636_inst ( .DIN1(_49411), .DIN2(_50154), .Q(_50153) );
  nor2s1 _50637_inst ( .DIN1(_49804), .DIN2(_49961), .Q(_50154) );
  hi1s1 _50638_inst ( .DIN(_49784), .Q(_49961) );
  nnd2s1 _50639_inst ( .DIN1(_50155), .DIN2(_50156), .Q(_49784) );
  nor2s1 _50640_inst ( .DIN1(_39117), .DIN2(_27441), .Q(_50155) );
  and2s1 _50641_inst ( .DIN1(_50157), .DIN2(_50158), .Q(_49804) );
  nor2s1 _50642_inst ( .DIN1(_34870), .DIN2(_50139), .Q(_50157) );
  hi1s1 _50643_inst ( .DIN(_49343), .Q(_49411) );
  nnd2s1 _50644_inst ( .DIN1(_49226), .DIN2(_49783), .Q(_49343) );
  nor2s1 _50645_inst ( .DIN1(_50159), .DIN2(_50160), .Q(_50152) );
  nnd2s1 _50646_inst ( .DIN1(_29288), .DIN2(_50161), .Q(_50160) );
  nnd2s1 _50647_inst ( .DIN1(_49517), .DIN2(_31195), .Q(_50159) );
  nor2s1 _50648_inst ( .DIN1(_50162), .DIN2(_50163), .Q(_50104) );
  nnd2s1 _50649_inst ( .DIN1(_50164), .DIN2(_50165), .Q(_50163) );
  nor2s1 _50650_inst ( .DIN1(_49481), .DIN2(_49520), .Q(_50165) );
  nnd2s1 _50651_inst ( .DIN1(_50166), .DIN2(_50167), .Q(_49520) );
  nor2s1 _50652_inst ( .DIN1(_49634), .DIN2(_50168), .Q(_50167) );
  nnd2s1 _50653_inst ( .DIN1(_49477), .DIN2(_49956), .Q(_50168) );
  or2s1 _50654_inst ( .DIN1(_49710), .DIN2(_49127), .Q(_49956) );
  nnd2s1 _50655_inst ( .DIN1(_50169), .DIN2(_27821), .Q(_49710) );
  nor2s1 _50656_inst ( .DIN1(_29741), .DIN2(_50170), .Q(_50169) );
  nnd2s1 _50657_inst ( .DIN1(_49955), .DIN2(_49754), .Q(_49477) );
  hi1s1 _50658_inst ( .DIN(_49565), .Q(_49955) );
  nnd2s1 _50659_inst ( .DIN1(_50171), .DIN2(_50172), .Q(_49565) );
  nor2s1 _50660_inst ( .DIN1(_37982), .DIN2(_27445), .Q(_50171) );
  nor2s1 _50661_inst ( .DIN1(_49315), .DIN2(_49127), .Q(_49634) );
  nnd2s1 _50662_inst ( .DIN1(_50173), .DIN2(_50174), .Q(_49315) );
  nor2s1 _50663_inst ( .DIN1(_35723), .DIN2(_34870), .Q(_50174) );
  nor2s1 _50664_inst ( .DIN1(_37984), .DIN2(_32809), .Q(_50173) );
  nor2s1 _50665_inst ( .DIN1(_50175), .DIN2(_50176), .Q(_50166) );
  nor2s1 _50666_inst ( .DIN1(_49581), .DIN2(_49278), .Q(_50176) );
  nnd2s1 _50667_inst ( .DIN1(_50177), .DIN2(_50178), .Q(_49278) );
  nor2s1 _50668_inst ( .DIN1(_36248), .DIN2(_39117), .Q(_50178) );
  nor2s1 _50669_inst ( .DIN1(_43422), .DIN2(_37299), .Q(_50177) );
  hi1s1 _50670_inst ( .DIN(_49754), .Q(_49581) );
  nnd2s1 _50671_inst ( .DIN1(_49149), .DIN2(_49165), .Q(_49754) );
  nnd2s1 _50672_inst ( .DIN1(_50179), .DIN2(_50180), .Q(_49165) );
  nor2s1 _50673_inst ( .DIN1(_49776), .DIN2(_49741), .Q(_50175) );
  nnd2s1 _50674_inst ( .DIN1(_50181), .DIN2(_50182), .Q(_49741) );
  nor2s1 _50675_inst ( .DIN1(_35300), .DIN2(_30939), .Q(_50182) );
  nor2s1 _50676_inst ( .DIN1(_37984), .DIN2(_32825), .Q(_50181) );
  nnd2s1 _50677_inst ( .DIN1(_49378), .DIN2(_49223), .Q(_49481) );
  hi1s1 _50678_inst ( .DIN(_49789), .Q(_49223) );
  nor2s1 _50679_inst ( .DIN1(_49127), .DIN2(_49621), .Q(_49789) );
  nnd2s1 _50680_inst ( .DIN1(_50183), .DIN2(_50184), .Q(_49621) );
  nor2s1 _50681_inst ( .DIN1(_36832), .DIN2(_35300), .Q(_50184) );
  nor2s1 _50682_inst ( .DIN1(_34870), .DIN2(_29742), .Q(_50183) );
  nnd2s1 _50683_inst ( .DIN1(_50185), .DIN2(_49457), .Q(_49378) );
  nnd2s1 _50684_inst ( .DIN1(_49714), .DIN2(_49128), .Q(_50185) );
  nnd2s1 _50685_inst ( .DIN1(_50186), .DIN2(_45421), .Q(_49128) );
  hi1s1 _50686_inst ( .DIN(_44326), .Q(_45421) );
  nnd2s1 _50687_inst ( .DIN1(_50186), .DIN2(_27310), .Q(_49714) );
  hi1s1 _50688_inst ( .DIN(_43422), .Q(_27310) );
  nor2s1 _50689_inst ( .DIN1(_34855), .DIN2(_50187), .Q(_50186) );
  nor2s1 _50690_inst ( .DIN1(_49928), .DIN2(_49719), .Q(_50164) );
  nnd2s1 _50691_inst ( .DIN1(_50188), .DIN2(_50189), .Q(_49719) );
  nor2s1 _50692_inst ( .DIN1(_50190), .DIN2(_50191), .Q(_50189) );
  nnd2s1 _50693_inst ( .DIN1(_50192), .DIN2(_50076), .Q(_50191) );
  nnd2s1 _50694_inst ( .DIN1(_49532), .DIN2(_49457), .Q(_50076) );
  hi1s1 _50695_inst ( .DIN(_49310), .Q(_49532) );
  nnd2s1 _50696_inst ( .DIN1(_50193), .DIN2(_50194), .Q(_49310) );
  nor2s1 _50697_inst ( .DIN1(_39117), .DIN2(_50195), .Q(_50193) );
  nnd2s1 _50698_inst ( .DIN1(_49632), .DIN2(_49655), .Q(_50192) );
  hi1s1 _50699_inst ( .DIN(_49219), .Q(_49632) );
  nnd2s1 _50700_inst ( .DIN1(_50196), .DIN2(_37987), .Q(_49219) );
  nnd2s1 _50701_inst ( .DIN1(_50197), .DIN2(_49580), .Q(_50190) );
  nnd2s1 _50702_inst ( .DIN1(_49342), .DIN2(_49805), .Q(_49580) );
  hi1s1 _50703_inst ( .DIN(_49412), .Q(_49342) );
  nnd2s1 _50704_inst ( .DIN1(_50198), .DIN2(_50199), .Q(_49412) );
  nor2s1 _50705_inst ( .DIN1(_35300), .DIN2(_34870), .Q(_50199) );
  nnd2s1 _50706_inst ( .DIN1(_49659), .DIN2(_47930), .Q(_50197) );
  nnd2s1 _50707_inst ( .DIN1(_50200), .DIN2(_46247), .Q(_47930) );
  and2s1 _50708_inst ( .DIN1(_50201), .DIN2(_50202), .Q(_46247) );
  nor2s1 _50709_inst ( .DIN1(_46705), .DIN2(_50203), .Q(_50202) );
  nnd2s1 _50710_inst ( .DIN1(_46271), .DIN2(_46360), .Q(_50203) );
  nnd2s1 _50711_inst ( .DIN1(_50204), .DIN2(_46312), .Q(_46360) );
  nor2s1 _50712_inst ( .DIN1(_46859), .DIN2(_46813), .Q(_50204) );
  nor2s1 _50713_inst ( .DIN1(_46828), .DIN2(_45547), .Q(_46705) );
  hi1s1 _50714_inst ( .DIN(_46615), .Q(_45547) );
  nnd2s1 _50715_inst ( .DIN1(_46879), .DIN2(_26468), .Q(_46828) );
  nor2s1 _50716_inst ( .DIN1(_50205), .DIN2(_46892), .Q(_46879) );
  nnd2s1 _50717_inst ( .DIN1(_26225), .DIN2(_26363), .Q(_50205) );
  nor2s1 _50718_inst ( .DIN1(_46629), .DIN2(_46790), .Q(_50201) );
  nnd2s1 _50719_inst ( .DIN1(_46499), .DIN2(_50206), .Q(_46790) );
  nnd2s1 _50720_inst ( .DIN1(_45212), .DIN2(_46757), .Q(_50206) );
  hi1s1 _50721_inst ( .DIN(_46368), .Q(_46757) );
  hi1s1 _50722_inst ( .DIN(_45553), .Q(_45212) );
  nnd2s1 _50723_inst ( .DIN1(_46853), .DIN2(_46884), .Q(_45553) );
  hi1s1 _50724_inst ( .DIN(_46795), .Q(_46884) );
  nnd2s1 _50725_inst ( .DIN1(_46655), .DIN2(_39514), .Q(_46499) );
  hi1s1 _50726_inst ( .DIN(_46728), .Q(_39514) );
  nnd2s1 _50727_inst ( .DIN1(_45207), .DIN2(_46866), .Q(_46728) );
  nor2s1 _50728_inst ( .DIN1(_50207), .DIN2(_2711), .Q(_46866) );
  and2s1 _50729_inst ( .DIN1(_50208), .DIN2(_46905), .Q(_46655) );
  hi1s1 _50730_inst ( .DIN(_46796), .Q(_46905) );
  nnd2s1 _50731_inst ( .DIN1(_50209), .DIN2(_2684), .Q(_46796) );
  nor2s1 _50732_inst ( .DIN1(_26225), .DIN2(_26363), .Q(_50209) );
  nor2s1 _50733_inst ( .DIN1(_28976), .DIN2(_26328), .Q(_50208) );
  nnd2s1 _50734_inst ( .DIN1(_50210), .DIN2(_46469), .Q(_46629) );
  nnd2s1 _50735_inst ( .DIN1(_46797), .DIN2(_39521), .Q(_46469) );
  hi1s1 _50736_inst ( .DIN(_46647), .Q(_39521) );
  nnd2s1 _50737_inst ( .DIN1(_46920), .DIN2(_46853), .Q(_46647) );
  hi1s1 _50738_inst ( .DIN(_46812), .Q(_46853) );
  nnd2s1 _50739_inst ( .DIN1(_2722), .DIN2(_2724), .Q(_46812) );
  and2s1 _50740_inst ( .DIN1(_50211), .DIN2(_28218), .Q(_46797) );
  nor2s1 _50741_inst ( .DIN1(_26225), .DIN2(_46923), .Q(_50211) );
  nnd2s1 _50742_inst ( .DIN1(_50212), .DIN2(_2697), .Q(_46923) );
  nor2s1 _50743_inst ( .DIN1(_2684), .DIN2(_26328), .Q(_50212) );
  nor2s1 _50744_inst ( .DIN1(_46389), .DIN2(_46473), .Q(_50210) );
  and2s1 _50745_inst ( .DIN1(_46717), .DIN2(_46529), .Q(_46473) );
  and2s1 _50746_inst ( .DIN1(_50213), .DIN2(_2698), .Q(_46529) );
  nor2s1 _50747_inst ( .DIN1(_28976), .DIN2(_46893), .Q(_50213) );
  nnd2s1 _50748_inst ( .DIN1(_2731), .DIN2(_2730), .Q(_28976) );
  hi1s1 _50749_inst ( .DIN(_45533), .Q(_46717) );
  nnd2s1 _50750_inst ( .DIN1(_46920), .DIN2(_46844), .Q(_45533) );
  hi1s1 _50751_inst ( .DIN(_46821), .Q(_46844) );
  and2s1 _50752_inst ( .DIN1(_46615), .DIN2(_46701), .Q(_46389) );
  and2s1 _50753_inst ( .DIN1(_50214), .DIN2(_50215), .Q(_46701) );
  nor2s1 _50754_inst ( .DIN1(_2684), .DIN2(_26225), .Q(_50215) );
  nor2s1 _50755_inst ( .DIN1(_46892), .DIN2(_26363), .Q(_50214) );
  nnd2s1 _50756_inst ( .DIN1(_28717), .DIN2(_26328), .Q(_46892) );
  hi1s1 _50757_inst ( .DIN(_37006), .Q(_28717) );
  nnd2s1 _50758_inst ( .DIN1(_2730), .DIN2(_26724), .Q(_37006) );
  nor2s1 _50759_inst ( .DIN1(_46813), .DIN2(_46821), .Q(_46615) );
  nnd2s1 _50760_inst ( .DIN1(_50216), .DIN2(_53521), .Q(_46813) );
  nor2s1 _50761_inst ( .DIN1(_2718), .DIN2(_2711), .Q(_50216) );
  nor2s1 _50762_inst ( .DIN1(_50217), .DIN2(_50218), .Q(_50200) );
  nor2s1 _50763_inst ( .DIN1(_46346), .DIN2(_46123), .Q(_50218) );
  nnd2s1 _50764_inst ( .DIN1(_50219), .DIN2(_46271), .Q(_46123) );
  nnd2s1 _50765_inst ( .DIN1(_46312), .DIN2(_46341), .Q(_46271) );
  nor2s1 _50766_inst ( .DIN1(_46859), .DIN2(_46795), .Q(_46341) );
  hi1s1 _50767_inst ( .DIN(_46664), .Q(_50219) );
  nnd2s1 _50768_inst ( .DIN1(_50220), .DIN2(_50221), .Q(_46664) );
  nnd2s1 _50769_inst ( .DIN1(_46312), .DIN2(_46770), .Q(_50221) );
  hi1s1 _50770_inst ( .DIN(_46313), .Q(_46770) );
  nnd2s1 _50771_inst ( .DIN1(_45207), .DIN2(_46920), .Q(_46313) );
  and2s1 _50772_inst ( .DIN1(_46906), .DIN2(_26692), .Q(_46920) );
  nor2s1 _50773_inst ( .DIN1(_53521), .DIN2(_2711), .Q(_46906) );
  hi1s1 _50774_inst ( .DIN(_46859), .Q(_45207) );
  and2s1 _50775_inst ( .DIN1(_50222), .DIN2(_50223), .Q(_46312) );
  nor2s1 _50776_inst ( .DIN1(_2731), .DIN2(_2730), .Q(_50223) );
  nor2s1 _50777_inst ( .DIN1(_2684), .DIN2(_46847), .Q(_50222) );
  nnd2s1 _50778_inst ( .DIN1(_50224), .DIN2(_2697), .Q(_46847) );
  nor2s1 _50779_inst ( .DIN1(_2699), .DIN2(_2698), .Q(_50224) );
  nor2s1 _50780_inst ( .DIN1(_46368), .DIN2(_45203), .Q(_46346) );
  hi1s1 _50781_inst ( .DIN(_39523), .Q(_45203) );
  nor2s1 _50782_inst ( .DIN1(_46821), .DIN2(_46795), .Q(_39523) );
  nnd2s1 _50783_inst ( .DIN1(_2711), .DIN2(_50225), .Q(_46795) );
  hi1s1 _50784_inst ( .DIN(_50207), .Q(_50225) );
  nnd2s1 _50785_inst ( .DIN1(_53521), .DIN2(_2718), .Q(_50207) );
  nnd2s1 _50786_inst ( .DIN1(_2724), .DIN2(_26575), .Q(_46821) );
  nnd2s1 _50787_inst ( .DIN1(_50226), .DIN2(_28218), .Q(_46368) );
  hi1s1 _50788_inst ( .DIN(_29221), .Q(_28218) );
  nnd2s1 _50789_inst ( .DIN1(_2731), .DIN2(_26315), .Q(_29221) );
  nor2s1 _50790_inst ( .DIN1(_46893), .DIN2(_26328), .Q(_50226) );
  nnd2s1 _50791_inst ( .DIN1(_50227), .DIN2(_2699), .Q(_46893) );
  nor2s1 _50792_inst ( .DIN1(_2697), .DIN2(_2684), .Q(_50227) );
  hi1s1 _50793_inst ( .DIN(_50220), .Q(_50217) );
  nnd2s1 _50794_inst ( .DIN1(_46776), .DIN2(_46771), .Q(_50220) );
  hi1s1 _50795_inst ( .DIN(_46854), .Q(_46771) );
  nnd2s1 _50796_inst ( .DIN1(_50228), .DIN2(_50229), .Q(_46854) );
  nor2s1 _50797_inst ( .DIN1(_2698), .DIN2(_46909), .Q(_50229) );
  nnd2s1 _50798_inst ( .DIN1(_26315), .DIN2(_26724), .Q(_46909) );
  nor2s1 _50799_inst ( .DIN1(_26468), .DIN2(_50230), .Q(_50228) );
  nnd2s1 _50800_inst ( .DIN1(_2699), .DIN2(_26363), .Q(_50230) );
  nor2s1 _50801_inst ( .DIN1(_46820), .DIN2(_46859), .Q(_46776) );
  nnd2s1 _50802_inst ( .DIN1(_2722), .DIN2(_26249), .Q(_46859) );
  nnd2s1 _50803_inst ( .DIN1(_50231), .DIN2(_2711), .Q(_46820) );
  nor2s1 _50804_inst ( .DIN1(_53521), .DIN2(_2718), .Q(_50231) );
  hi1s1 _50805_inst ( .DIN(_49612), .Q(_49659) );
  nnd2s1 _50806_inst ( .DIN1(_50232), .DIN2(_50196), .Q(_49612) );
  nor2s1 _50807_inst ( .DIN1(_49465), .DIN2(_37984), .Q(_50232) );
  nor2s1 _50808_inst ( .DIN1(_50233), .DIN2(_50234), .Q(_50188) );
  nnd2s1 _50809_inst ( .DIN1(_49665), .DIN2(_49483), .Q(_50234) );
  and2s1 _50810_inst ( .DIN1(_50075), .DIN2(_50235), .Q(_49483) );
  or2s1 _50811_inst ( .DIN1(_49117), .DIN2(_49275), .Q(_50235) );
  nnd2s1 _50812_inst ( .DIN1(_50236), .DIN2(_50237), .Q(_49275) );
  nor2s1 _50813_inst ( .DIN1(_29741), .DIN2(_35300), .Q(_50237) );
  nor2s1 _50814_inst ( .DIN1(_30939), .DIN2(_33293), .Q(_50236) );
  nnd2s1 _50815_inst ( .DIN1(_49383), .DIN2(_49805), .Q(_50075) );
  hi1s1 _50816_inst ( .DIN(_49226), .Q(_49805) );
  nnd2s1 _50817_inst ( .DIN1(_49457), .DIN2(_50238), .Q(_49226) );
  nnd2s1 _50818_inst ( .DIN1(_50239), .DIN2(______[6]), .Q(_50238) );
  hi1s1 _50819_inst ( .DIN(_49566), .Q(_49383) );
  nnd2s1 _50820_inst ( .DIN1(_50240), .DIN2(_27316), .Q(_49566) );
  nor2s1 _50821_inst ( .DIN1(_36832), .DIN2(_50170), .Q(_50240) );
  and2s1 _50822_inst ( .DIN1(_49427), .DIN2(_50241), .Q(_49665) );
  nnd2s1 _50823_inst ( .DIN1(_26806), .DIN2(_49780), .Q(_50241) );
  nnd2s1 _50824_inst ( .DIN1(_49375), .DIN2(_49672), .Q(_49427) );
  hi1s1 _50825_inst ( .DIN(_49900), .Q(_49375) );
  nnd2s1 _50826_inst ( .DIN1(_50242), .DIN2(_50243), .Q(_49900) );
  nor2s1 _50827_inst ( .DIN1(_36832), .DIN2(_32809), .Q(_50242) );
  nnd2s1 _50828_inst ( .DIN1(_49363), .DIN2(_49485), .Q(_50233) );
  nnd2s1 _50829_inst ( .DIN1(_49676), .DIN2(_49633), .Q(_49485) );
  hi1s1 _50830_inst ( .DIN(_49776), .Q(_49633) );
  hi1s1 _50831_inst ( .DIN(_49248), .Q(_49676) );
  nnd2s1 _50832_inst ( .DIN1(_50244), .DIN2(_50245), .Q(_49248) );
  nor2s1 _50833_inst ( .DIN1(_35721), .DIN2(_32825), .Q(_50245) );
  nor2s1 _50834_inst ( .DIN1(_27828), .DIN2(_30940), .Q(_50244) );
  and2s1 _50835_inst ( .DIN1(_50246), .DIN2(_50247), .Q(_49363) );
  nor2s1 _50836_inst ( .DIN1(_50248), .DIN2(_50249), .Q(_50247) );
  nnd2s1 _50837_inst ( .DIN1(_49821), .DIN2(_49605), .Q(_50249) );
  nnd2s1 _50838_inst ( .DIN1(_49457), .DIN2(_50250), .Q(_49605) );
  nnd2s1 _50839_inst ( .DIN1(_49988), .DIN2(_50251), .Q(_50250) );
  nnd2s1 _50840_inst ( .DIN1(_50252), .DIN2(_50161), .Q(_50251) );
  nnd2s1 _50841_inst ( .DIN1(_50253), .DIN2(_50132), .Q(_49988) );
  nor2s1 _50842_inst ( .DIN1(_39117), .DIN2(_44324), .Q(_50253) );
  nor2s1 _50843_inst ( .DIN1(_50254), .DIN2(_49673), .Q(_49821) );
  and2s1 _50844_inst ( .DIN1(_50103), .DIN2(_50255), .Q(_49673) );
  and2s1 _50845_inst ( .DIN1(_50256), .DIN2(_50257), .Q(_50103) );
  nor2s1 _50846_inst ( .DIN1(_39110), .DIN2(_35721), .Q(_50257) );
  nor2s1 _50847_inst ( .DIN1(_32825), .DIN2(_27828), .Q(_50256) );
  hi1s1 _50848_inst ( .DIN(_49535), .Q(_50254) );
  nnd2s1 _50849_inst ( .DIN1(_50258), .DIN2(_50259), .Q(_49535) );
  nor2s1 _50850_inst ( .DIN1(_34855), .DIN2(_49344), .Q(_50259) );
  nor2s1 _50851_inst ( .DIN1(_44324), .DIN2(_50260), .Q(_50258) );
  nnd2s1 _50852_inst ( .DIN1(_50261), .DIN2(_49438), .Q(_50248) );
  hi1s1 _50853_inst ( .DIN(_49929), .Q(_49438) );
  nor2s1 _50854_inst ( .DIN1(_50118), .DIN2(_49161), .Q(_49929) );
  nnd2s1 _50855_inst ( .DIN1(_50262), .DIN2(_50172), .Q(_50118) );
  nor2s1 _50856_inst ( .DIN1(_30434), .DIN2(_36248), .Q(_50172) );
  nor2s1 _50857_inst ( .DIN1(_38682), .DIN2(_45435), .Q(_50262) );
  nnd2s1 _50858_inst ( .DIN1(_50073), .DIN2(_50263), .Q(_45435) );
  nor2s1 _50859_inst ( .DIN1(_49592), .DIN2(_49440), .Q(_50261) );
  nor2s1 _50860_inst ( .DIN1(_49345), .DIN2(_49311), .Q(_49440) );
  nnd2s1 _50861_inst ( .DIN1(_50264), .DIN2(_50243), .Q(_49345) );
  nor2s1 _50862_inst ( .DIN1(_33293), .DIN2(_50139), .Q(_50264) );
  nor2s1 _50863_inst ( .DIN1(_49155), .DIN2(_50265), .Q(_49592) );
  nor2s1 _50864_inst ( .DIN1(_50266), .DIN2(_50267), .Q(_50246) );
  nnd2s1 _50865_inst ( .DIN1(_50268), .DIN2(_49696), .Q(_50267) );
  and2s1 _50866_inst ( .DIN1(_50269), .DIN2(_50270), .Q(_49696) );
  nor2s1 _50867_inst ( .DIN1(_50271), .DIN2(_50272), .Q(_50270) );
  nnd2s1 _50868_inst ( .DIN1(_49170), .DIN2(_49425), .Q(_50272) );
  and2s1 _50869_inst ( .DIN1(_49258), .DIN2(_50273), .Q(_49425) );
  or2s1 _50870_inst ( .DIN1(_49150), .DIN2(_49149), .Q(_50273) );
  nnd2s1 _50871_inst ( .DIN1(_50274), .DIN2(_50158), .Q(_49150) );
  nor2s1 _50872_inst ( .DIN1(_35300), .DIN2(_50275), .Q(_50158) );
  nor2s1 _50873_inst ( .DIN1(_39111), .DIN2(_32821), .Q(_50274) );
  nnd2s1 _50874_inst ( .DIN1(_50263), .DIN2(_50276), .Q(_32821) );
  nnd2s1 _50875_inst ( .DIN1(_50277), .DIN2(_50278), .Q(_49258) );
  nor2s1 _50876_inst ( .DIN1(_32824), .DIN2(_49344), .Q(_50278) );
  hi1s1 _50877_inst ( .DIN(_49643), .Q(_49170) );
  nnd2s1 _50878_inst ( .DIN1(_50279), .DIN2(_50280), .Q(_49643) );
  or2s1 _50879_inst ( .DIN1(_49509), .DIN2(_49155), .Q(_50280) );
  nor2s1 _50880_inst ( .DIN1(_50281), .DIN2(_50282), .Q(_50279) );
  nor2s1 _50881_inst ( .DIN1(_49187), .DIN2(_50283), .Q(_50282) );
  nor2s1 _50882_inst ( .DIN1(_50284), .DIN2(_50285), .Q(_50281) );
  nnd2s1 _50883_inst ( .DIN1(_29433), .DIN2(_49780), .Q(_50285) );
  nnd2s1 _50884_inst ( .DIN1(_50286), .DIN2(_49935), .Q(_50271) );
  hi1s1 _50885_inst ( .DIN(_49439), .Q(_49935) );
  nor2s1 _50886_inst ( .DIN1(_49783), .DIN2(_50116), .Q(_49439) );
  nnd2s1 _50887_inst ( .DIN1(_50287), .DIN2(_50288), .Q(_50116) );
  hi1s1 _50888_inst ( .DIN(_50187), .Q(_50288) );
  nor2s1 _50889_inst ( .DIN1(_30434), .DIN2(_27446), .Q(_50287) );
  nnd2s1 _50890_inst ( .DIN1(_50289), .DIN2(_49457), .Q(_50286) );
  nnd2s1 _50891_inst ( .DIN1(_49473), .DIN2(_49227), .Q(_50289) );
  nnd2s1 _50892_inst ( .DIN1(_50290), .DIN2(_30026), .Q(_49227) );
  nor2s1 _50893_inst ( .DIN1(_45434), .DIN2(_50187), .Q(_50290) );
  nnd2s1 _50894_inst ( .DIN1(_50291), .DIN2(_49916), .Q(_45434) );
  nnd2s1 _50895_inst ( .DIN1(_50292), .DIN2(_34414), .Q(_49473) );
  nor2s1 _50896_inst ( .DIN1(_50293), .DIN2(_32820), .Q(_50292) );
  nor2s1 _50897_inst ( .DIN1(_50030), .DIN2(_50294), .Q(_50269) );
  or2s1 _50898_inst ( .DIN1(_49983), .DIN2(_49844), .Q(_50294) );
  nnd2s1 _50899_inst ( .DIN1(_50295), .DIN2(_50296), .Q(_49844) );
  nnd2s1 _50900_inst ( .DIN1(_50088), .DIN2(_49609), .Q(_50296) );
  and2s1 _50901_inst ( .DIN1(_50297), .DIN2(_50298), .Q(_50088) );
  nor2s1 _50902_inst ( .DIN1(_35720), .DIN2(_34413), .Q(_50298) );
  nor2s1 _50903_inst ( .DIN1(_37299), .DIN2(_32826), .Q(_50297) );
  nnd2s1 _50904_inst ( .DIN1(_49399), .DIN2(_50299), .Q(_50295) );
  or2s1 _50905_inst ( .DIN1(_49601), .DIN2(_49334), .Q(_49983) );
  hi1s1 _50906_inst ( .DIN(_49589), .Q(_49334) );
  nnd2s1 _50907_inst ( .DIN1(_50300), .DIN2(_49553), .Q(_49589) );
  hi1s1 _50908_inst ( .DIN(_49187), .Q(_49553) );
  nor2s1 _50909_inst ( .DIN1(_50119), .DIN2(_49161), .Q(_49601) );
  nnd2s1 _50910_inst ( .DIN1(_50301), .DIN2(_30026), .Q(_50119) );
  hi1s1 _50911_inst ( .DIN(_30433), .Q(_30026) );
  nor2s1 _50912_inst ( .DIN1(_43422), .DIN2(_50260), .Q(_50301) );
  nnd2s1 _50913_inst ( .DIN1(_50302), .DIN2(_50303), .Q(_50030) );
  nnd2s1 _50914_inst ( .DIN1(_49958), .DIN2(_49609), .Q(_50303) );
  nnd2s1 _50915_inst ( .DIN1(_49120), .DIN2(_49152), .Q(_49609) );
  hi1s1 _50916_inst ( .DIN(_49119), .Q(_49958) );
  nnd2s1 _50917_inst ( .DIN1(_50304), .DIN2(_27308), .Q(_49119) );
  hi1s1 _50918_inst ( .DIN(_32820), .Q(_27308) );
  or2s1 _50919_inst ( .DIN1(_49118), .DIN2(_49501), .Q(_50302) );
  hi1s1 _50920_inst ( .DIN(_50255), .Q(_49501) );
  nnd2s1 _50921_inst ( .DIN1(_50305), .DIN2(_50194), .Q(_49118) );
  nor2s1 _50922_inst ( .DIN1(_36248), .DIN2(_27446), .Q(_50194) );
  nor2s1 _50923_inst ( .DIN1(_32091), .DIN2(_50306), .Q(_50305) );
  hi1s1 _50924_inst ( .DIN(_49526), .Q(_50268) );
  nnd2s1 _50925_inst ( .DIN1(_50307), .DIN2(_50308), .Q(_49526) );
  nor2s1 _50926_inst ( .DIN1(_49640), .DIN2(_50309), .Q(_50308) );
  nor2s1 _50927_inst ( .DIN1(_49896), .DIN2(_49344), .Q(_50309) );
  nor2s1 _50928_inst ( .DIN1(_50115), .DIN2(_49783), .Q(_49640) );
  nnd2s1 _50929_inst ( .DIN1(_50310), .DIN2(_50239), .Q(_49783) );
  nnd2s1 _50930_inst ( .DIN1(_50311), .DIN2(_50124), .Q(_50115) );
  nor2s1 _50931_inst ( .DIN1(_30434), .DIN2(_32826), .Q(_50311) );
  nor2s1 _50932_inst ( .DIN1(_49977), .DIN2(_50027), .Q(_50307) );
  nnd2s1 _50933_inst ( .DIN1(_50312), .DIN2(_50313), .Q(_50027) );
  nnd2s1 _50934_inst ( .DIN1(_49831), .DIN2(_50255), .Q(_50313) );
  and2s1 _50935_inst ( .DIN1(_50314), .DIN2(_50315), .Q(_49831) );
  nor2s1 _50936_inst ( .DIN1(_36248), .DIN2(_38682), .Q(_50315) );
  nor2s1 _50937_inst ( .DIN1(_32091), .DIN2(_50316), .Q(_50314) );
  nnd2s1 _50938_inst ( .DIN1(_49798), .DIN2(_50317), .Q(_50312) );
  hi1s1 _50939_inst ( .DIN(_49344), .Q(_49798) );
  nnd2s1 _50940_inst ( .DIN1(_50318), .DIN2(_50319), .Q(_49344) );
  or2s1 _50941_inst ( .DIN1(_49595), .DIN2(_49476), .Q(_49977) );
  nor2s1 _50942_inst ( .DIN1(_50320), .DIN2(_49187), .Q(_49476) );
  nnd2s1 _50943_inst ( .DIN1(_50321), .DIN2(_50322), .Q(_49595) );
  nnd2s1 _50944_inst ( .DIN1(_50323), .DIN2(_50324), .Q(_50322) );
  nor2s1 _50945_inst ( .DIN1(_50306), .DIN2(_49152), .Q(_50324) );
  nnd2s1 _50946_inst ( .DIN1(_50310), .DIN2(_50180), .Q(_49152) );
  nor2s1 _50947_inst ( .DIN1(_49465), .DIN2(_26846), .Q(_50310) );
  and2s1 _50948_inst ( .DIN1(_50161), .DIN2(_29288), .Q(_50323) );
  hi1s1 _50949_inst ( .DIN(_29408), .Q(_29288) );
  nnd2s1 _50950_inst ( .DIN1(_50073), .DIN2(_50325), .Q(_29408) );
  nnd2s1 _50951_inst ( .DIN1(_50326), .DIN2(_49780), .Q(_50321) );
  hi1s1 _50952_inst ( .DIN(_49255), .Q(_49780) );
  nnd2s1 _50953_inst ( .DIN1(_50179), .DIN2(_50239), .Q(_49255) );
  nor2s1 _50954_inst ( .DIN1(______[6]), .DIN2(_49465), .Q(_50179) );
  nnd2s1 _50955_inst ( .DIN1(_50327), .DIN2(_49893), .Q(_50266) );
  nor2s1 _50956_inst ( .DIN1(_50328), .DIN2(_49845), .Q(_49893) );
  nnd2s1 _50957_inst ( .DIN1(_50329), .DIN2(_50330), .Q(_49845) );
  nnd2s1 _50958_inst ( .DIN1(_50331), .DIN2(_50332), .Q(_50330) );
  nor2s1 _50959_inst ( .DIN1(_27442), .DIN2(_49127), .Q(_50331) );
  nnd2s1 _50960_inst ( .DIN1(_50333), .DIN2(_50045), .Q(_50329) );
  and2s1 _50961_inst ( .DIN1(_50334), .DIN2(_27821), .Q(_50045) );
  hi1s1 _50962_inst ( .DIN(_27828), .Q(_27821) );
  nor2s1 _50963_inst ( .DIN1(_30939), .DIN2(_35721), .Q(_50334) );
  nnd2s1 _50964_inst ( .DIN1(_50335), .DIN2(_2216), .Q(_30939) );
  nor2s1 _50965_inst ( .DIN1(_50336), .DIN2(_26433), .Q(_50335) );
  nor2s1 _50966_inst ( .DIN1(_29741), .DIN2(_49776), .Q(_50333) );
  or2s1 _50967_inst ( .DIN1(_50055), .DIN2(_50337), .Q(_50328) );
  nor2s1 _50968_inst ( .DIN1(_49196), .DIN2(_50054), .Q(_50337) );
  nnd2s1 _50969_inst ( .DIN1(_50338), .DIN2(_29433), .Q(_50054) );
  hi1s1 _50970_inst ( .DIN(_27441), .Q(_29433) );
  nor2s1 _50971_inst ( .DIN1(_39117), .DIN2(_50293), .Q(_50338) );
  hi1s1 _50972_inst ( .DIN(_49687), .Q(_49196) );
  nnd2s1 _50973_inst ( .DIN1(_49127), .DIN2(_49187), .Q(_49687) );
  and2s1 _50974_inst ( .DIN1(_50339), .DIN2(_49399), .Q(_50055) );
  nor2s1 _50975_inst ( .DIN1(_49444), .DIN2(_49426), .Q(_50327) );
  nnd2s1 _50976_inst ( .DIN1(_49337), .DIN2(_50340), .Q(_49426) );
  nnd2s1 _50977_inst ( .DIN1(_49550), .DIN2(_50255), .Q(_50340) );
  nnd2s1 _50978_inst ( .DIN1(_49117), .DIN2(_49155), .Q(_50255) );
  hi1s1 _50979_inst ( .DIN(_49656), .Q(_49550) );
  nnd2s1 _50980_inst ( .DIN1(_50341), .DIN2(_50342), .Q(_49656) );
  nor2s1 _50981_inst ( .DIN1(_35720), .DIN2(_27446), .Q(_50342) );
  nor2s1 _50982_inst ( .DIN1(_37942), .DIN2(_39114), .Q(_50341) );
  nnd2s1 _50983_inst ( .DIN1(_49678), .DIN2(_49655), .Q(_49337) );
  nnd2s1 _50984_inst ( .DIN1(_49776), .DIN2(_49161), .Q(_49655) );
  nnd2s1 _50985_inst ( .DIN1(_50343), .DIN2(_50319), .Q(_49161) );
  and2s1 _50986_inst ( .DIN1(_50344), .DIN2(_50130), .Q(_49678) );
  nor2s1 _50987_inst ( .DIN1(_27445), .DIN2(_50195), .Q(_50344) );
  nnd2s1 _50988_inst ( .DIN1(_50345), .DIN2(_50346), .Q(_49444) );
  nnd2s1 _50989_inst ( .DIN1(_50347), .DIN2(_49399), .Q(_50346) );
  hi1s1 _50990_inst ( .DIN(_49155), .Q(_49399) );
  nnd2s1 _50991_inst ( .DIN1(_50343), .DIN2(_50348), .Q(_49155) );
  nor2s1 _50992_inst ( .DIN1(_49465), .DIN2(_27066), .Q(_50343) );
  nnd2s1 _50993_inst ( .DIN1(_48332), .DIN2(_49672), .Q(_50345) );
  nnd2s1 _50994_inst ( .DIN1(_50349), .DIN2(_50138), .Q(_48130) );
  nor2s1 _50995_inst ( .DIN1(_36832), .DIN2(_35723), .Q(_50138) );
  nnd2s1 _50996_inst ( .DIN1(_49436), .DIN2(_49583), .Q(_49928) );
  nnd2s1 _50997_inst ( .DIN1(_49517), .DIN2(_49723), .Q(_49583) );
  hi1s1 _50998_inst ( .DIN(_49151), .Q(_49723) );
  nnd2s1 _50999_inst ( .DIN1(_50350), .DIN2(_50351), .Q(_49151) );
  nor2s1 _51000_inst ( .DIN1(_39111), .DIN2(_35721), .Q(_50351) );
  nnd2s1 _51001_inst ( .DIN1(_50352), .DIN2(_50021), .Q(_39111) );
  hi1s1 _51002_inst ( .DIN(_50336), .Q(_50021) );
  nor2s1 _51003_inst ( .DIN1(_2216), .DIN2(_2214), .Q(_50352) );
  nor2s1 _51004_inst ( .DIN1(_37984), .DIN2(_45436), .Q(_50350) );
  nnd2s1 _51005_inst ( .DIN1(_50151), .DIN2(_45431), .Q(_45436) );
  hi1s1 _51006_inst ( .DIN(_49120), .Q(_49517) );
  nnd2s1 _51007_inst ( .DIN1(_49457), .DIN2(_50353), .Q(_49120) );
  nnd2s1 _51008_inst ( .DIN1(_50180), .DIN2(______[6]), .Q(_50353) );
  nnd2s1 _51009_inst ( .DIN1(_49910), .DIN2(_49734), .Q(_49436) );
  hi1s1 _51010_inst ( .DIN(_49188), .Q(_49734) );
  nnd2s1 _51011_inst ( .DIN1(_50196), .DIN2(_36829), .Q(_49188) );
  hi1s1 _51012_inst ( .DIN(_36832), .Q(_36829) );
  nnd2s1 _51013_inst ( .DIN1(_50354), .DIN2(_50355), .Q(_36832) );
  and2s1 _51014_inst ( .DIN1(_50356), .DIN2(_27316), .Q(_50196) );
  hi1s1 _51015_inst ( .DIN(_27442), .Q(_27316) );
  nor2s1 _51016_inst ( .DIN1(_34870), .DIN2(_35721), .Q(_50356) );
  nnd2s1 _51017_inst ( .DIN1(_50357), .DIN2(_50358), .Q(_50162) );
  nor2s1 _51018_inst ( .DIN1(_50359), .DIN2(_50360), .Q(_50358) );
  nnd2s1 _51019_inst ( .DIN1(_50361), .DIN2(_50362), .Q(_50360) );
  nnd2s1 _51020_inst ( .DIN1(_49910), .DIN2(_50363), .Q(_50362) );
  nnd2s1 _51021_inst ( .DIN1(_50364), .DIN2(_50320), .Q(_50363) );
  nnd2s1 _51022_inst ( .DIN1(_50122), .DIN2(_50365), .Q(_50320) );
  nor2s1 _51023_inst ( .DIN1(_27445), .DIN2(_39117), .Q(_50365) );
  nnd2s1 _51024_inst ( .DIN1(_50366), .DIN2(_50367), .Q(_39117) );
  nor2s1 _51025_inst ( .DIN1(_2216), .DIN2(_26248), .Q(_50366) );
  nnd2s1 _51026_inst ( .DIN1(_50073), .DIN2(_45430), .Q(_27445) );
  nor2s1 _51027_inst ( .DIN1(_50300), .DIN2(_50368), .Q(_50364) );
  hi1s1 _51028_inst ( .DIN(_50283), .Q(_50368) );
  nnd2s1 _51029_inst ( .DIN1(_50369), .DIN2(_50370), .Q(_50283) );
  nor2s1 _51030_inst ( .DIN1(_39282), .DIN2(_32091), .Q(_50370) );
  nor2s1 _51031_inst ( .DIN1(_50195), .DIN2(_32826), .Q(_50369) );
  and2s1 _51032_inst ( .DIN1(_50371), .DIN2(_50372), .Q(_50300) );
  nor2s1 _51033_inst ( .DIN1(_43422), .DIN2(_30433), .Q(_50371) );
  nnd2s1 _51034_inst ( .DIN1(_50373), .DIN2(_50374), .Q(_30433) );
  nor2s1 _51035_inst ( .DIN1(_2203), .DIN2(_26433), .Q(_50374) );
  nor2s1 _51036_inst ( .DIN1(_26370), .DIN2(_26210), .Q(_50373) );
  hi1s1 _51037_inst ( .DIN(_49127), .Q(_49910) );
  nnd2s1 _51038_inst ( .DIN1(_49457), .DIN2(_50375), .Q(_49127) );
  nnd2s1 _51039_inst ( .DIN1(_50348), .DIN2(_26854), .Q(_50375) );
  nnd2s1 _51040_inst ( .DIN1(_49672), .DIN2(_50376), .Q(_50361) );
  nnd2s1 _51041_inst ( .DIN1(_50377), .DIN2(_50378), .Q(_50376) );
  nor2s1 _51042_inst ( .DIN1(_50326), .DIN2(_49257), .Q(_50378) );
  hi1s1 _51043_inst ( .DIN(_49757), .Q(_49257) );
  nnd2s1 _51044_inst ( .DIN1(_45424), .DIN2(_50140), .Q(_49757) );
  hi1s1 _51045_inst ( .DIN(_29742), .Q(_45424) );
  nnd2s1 _51046_inst ( .DIN1(_45430), .DIN2(_50276), .Q(_29742) );
  and2s1 _51047_inst ( .DIN1(_50252), .DIN2(_50130), .Q(_50326) );
  nor2s1 _51048_inst ( .DIN1(_39114), .DIN2(_36248), .Q(_50130) );
  hi1s1 _51049_inst ( .DIN(_34414), .Q(_39114) );
  nor2s1 _51050_inst ( .DIN1(_37983), .DIN2(_32820), .Q(_50252) );
  nnd2s1 _51051_inst ( .DIN1(_50276), .DIN2(_50379), .Q(_32820) );
  nor2s1 _51052_inst ( .DIN1(_50380), .DIN2(_49499), .Q(_50377) );
  nnd2s1 _51053_inst ( .DIN1(_49279), .DIN2(_49755), .Q(_49499) );
  nnd2s1 _51054_inst ( .DIN1(_50198), .DIN2(_50243), .Q(_49755) );
  nor2s1 _51055_inst ( .DIN1(_30940), .DIN2(_35300), .Q(_50243) );
  nnd2s1 _51056_inst ( .DIN1(_50381), .DIN2(_50367), .Q(_30940) );
  hi1s1 _51057_inst ( .DIN(_50382), .Q(_50367) );
  nor2s1 _51058_inst ( .DIN1(_2216), .DIN2(_2203), .Q(_50381) );
  nor2s1 _51059_inst ( .DIN1(_50139), .DIN2(_27828), .Q(_50198) );
  nnd2s1 _51060_inst ( .DIN1(_50355), .DIN2(_50383), .Q(_27828) );
  hi1s1 _51061_inst ( .DIN(_50101), .Q(_50355) );
  hi1s1 _51062_inst ( .DIN(_49841), .Q(_49279) );
  nor2s1 _51063_inst ( .DIN1(_50384), .DIN2(_50170), .Q(_49841) );
  or2s1 _51064_inst ( .DIN1(_33293), .DIN2(_32825), .Q(_50384) );
  nnd2s1 _51065_inst ( .DIN1(_49916), .DIN2(_50325), .Q(_32825) );
  nor2s1 _51066_inst ( .DIN1(_27441), .DIN2(_50284), .Q(_50380) );
  nnd2s1 _51067_inst ( .DIN1(_50372), .DIN2(_30925), .Q(_50284) );
  nor2s1 _51068_inst ( .DIN1(_36248), .DIN2(_50306), .Q(_50372) );
  nnd2s1 _51069_inst ( .DIN1(_50385), .DIN2(_49892), .Q(_27441) );
  nor2s1 _51070_inst ( .DIN1(_2175), .DIN2(_26223), .Q(_50385) );
  hi1s1 _51071_inst ( .DIN(_49726), .Q(_49672) );
  nnd2s1 _51072_inst ( .DIN1(_49457), .DIN2(_50386), .Q(_49726) );
  nnd2s1 _51073_inst ( .DIN1(_50239), .DIN2(_28646), .Q(_50386) );
  nor2s1 _51074_inst ( .DIN1(_28100), .DIN2(_27066), .Q(_50239) );
  nor2s1 _51075_inst ( .DIN1(_50387), .DIN2(_49311), .Q(_50359) );
  nnd2s1 _51076_inst ( .DIN1(_49457), .DIN2(_50388), .Q(_49311) );
  nnd2s1 _51077_inst ( .DIN1(_50319), .DIN2(_26854), .Q(_50388) );
  nor2s1 _51078_inst ( .DIN1(_50389), .DIN2(_50390), .Q(_50387) );
  nnd2s1 _51079_inst ( .DIN1(_50391), .DIN2(_50392), .Q(_50390) );
  nnd2s1 _51080_inst ( .DIN1(_50393), .DIN2(_50124), .Q(_50392) );
  hi1s1 _51081_inst ( .DIN(_50260), .Q(_50124) );
  nor2s1 _51082_inst ( .DIN1(_34855), .DIN2(_44324), .Q(_50393) );
  nnd2s1 _51083_inst ( .DIN1(_49916), .DIN2(_50379), .Q(_44324) );
  and2s1 _51084_inst ( .DIN1(_50394), .DIN2(_26223), .Q(_50379) );
  hi1s1 _51085_inst ( .DIN(_50317), .Q(_50391) );
  nnd2s1 _51086_inst ( .DIN1(_50395), .DIN2(_50396), .Q(_50317) );
  nnd2s1 _51087_inst ( .DIN1(_50304), .DIN2(_32813), .Q(_50396) );
  hi1s1 _51088_inst ( .DIN(_50316), .Q(_32813) );
  nnd2s1 _51089_inst ( .DIN1(_50277), .DIN2(_42131), .Q(_50395) );
  hi1s1 _51090_inst ( .DIN(_32826), .Q(_42131) );
  nnd2s1 _51091_inst ( .DIN1(_50397), .DIN2(_49892), .Q(_32826) );
  nor2s1 _51092_inst ( .DIN1(_50398), .DIN2(_2180), .Q(_49892) );
  or2s1 _51093_inst ( .DIN1(_2182), .DIN2(_2181), .Q(_50398) );
  nor2s1 _51094_inst ( .DIN1(_2179), .DIN2(_26419), .Q(_50397) );
  nor2s1 _51095_inst ( .DIN1(_50187), .DIN2(_34413), .Q(_50277) );
  nnd2s1 _51096_inst ( .DIN1(_50399), .DIN2(_49896), .Q(_50389) );
  nnd2s1 _51097_inst ( .DIN1(_50304), .DIN2(_31397), .Q(_49896) );
  hi1s1 _51098_inst ( .DIN(_32824), .Q(_31397) );
  nor2s1 _51099_inst ( .DIN1(_50293), .DIN2(_32091), .Q(_50304) );
  or2s1 _51100_inst ( .DIN1(_35720), .DIN2(_37982), .Q(_50293) );
  nnd2s1 _51101_inst ( .DIN1(_50354), .DIN2(_50400), .Q(_37982) );
  nnd2s1 _51102_inst ( .DIN1(_50401), .DIN2(_30925), .Q(_50399) );
  hi1s1 _51103_inst ( .DIN(_34413), .Q(_30925) );
  nor2s1 _51104_inst ( .DIN1(_32824), .DIN2(_50187), .Q(_50401) );
  nnd2s1 _51105_inst ( .DIN1(_50073), .DIN2(_50291), .Q(_32824) );
  nor2s1 _51106_inst ( .DIN1(_2175), .DIN2(_2181), .Q(_50073) );
  nor2s1 _51107_inst ( .DIN1(_50402), .DIN2(_49139), .Q(_50357) );
  nnd2s1 _51108_inst ( .DIN1(_50403), .DIN2(_50404), .Q(_49139) );
  nnd2s1 _51109_inst ( .DIN1(_49637), .DIN2(_49301), .Q(_50404) );
  hi1s1 _51110_inst ( .DIN(_49149), .Q(_49301) );
  nnd2s1 _51111_inst ( .DIN1(_49457), .DIN2(_50405), .Q(_49149) );
  nnd2s1 _51112_inst ( .DIN1(_50180), .DIN2(_28646), .Q(_50405) );
  nor2s1 _51113_inst ( .DIN1(_28100), .DIN2(______[8]), .Q(_50180) );
  hi1s1 _51114_inst ( .DIN(_49843), .Q(_49637) );
  nnd2s1 _51115_inst ( .DIN1(_50406), .DIN2(_50349), .Q(_49843) );
  nor2s1 _51116_inst ( .DIN1(_39110), .DIN2(_29741), .Q(_50349) );
  nnd2s1 _51117_inst ( .DIN1(_50151), .DIN2(_49916), .Q(_29741) );
  hi1s1 _51118_inst ( .DIN(_50094), .Q(_50151) );
  nnd2s1 _51119_inst ( .DIN1(_50407), .DIN2(_2180), .Q(_50094) );
  nor2s1 _51120_inst ( .DIN1(_2182), .DIN2(_26223), .Q(_50407) );
  nor2s1 _51121_inst ( .DIN1(_50275), .DIN2(_35721), .Q(_50406) );
  nnd2s1 _51122_inst ( .DIN1(_50408), .DIN2(_53522), .Q(_35721) );
  nor2s1 _51123_inst ( .DIN1(_2274), .DIN2(_49864), .Q(_50408) );
  hi1s1 _51124_inst ( .DIN(_36828), .Q(_50275) );
  nor2s1 _51125_inst ( .DIN1(_49540), .DIN2(_50409), .Q(_36828) );
  nnd2s1 _51126_inst ( .DIN1(_2238), .DIN2(_2253), .Q(_49540) );
  nor2s1 _51127_inst ( .DIN1(_50056), .DIN2(_50410), .Q(_50403) );
  nor2s1 _51128_inst ( .DIN1(_49776), .DIN2(_49228), .Q(_50410) );
  nnd2s1 _51129_inst ( .DIN1(_50140), .DIN2(_27309), .Q(_49228) );
  hi1s1 _51130_inst ( .DIN(_50139), .Q(_27309) );
  nnd2s1 _51131_inst ( .DIN1(_50291), .DIN2(_45431), .Q(_50139) );
  and2s1 _51132_inst ( .DIN1(_50411), .DIN2(_29940), .Q(_50140) );
  hi1s1 _51133_inst ( .DIN(_34870), .Q(_29940) );
  nnd2s1 _51134_inst ( .DIN1(_50412), .DIN2(_2217), .Q(_34870) );
  nor2s1 _51135_inst ( .DIN1(_2216), .DIN2(_50413), .Q(_50412) );
  nor2s1 _51136_inst ( .DIN1(_35723), .DIN2(_33293), .Q(_50411) );
  nnd2s1 _51137_inst ( .DIN1(_49457), .DIN2(_50414), .Q(_49776) );
  nnd2s1 _51138_inst ( .DIN1(_50319), .DIN2(______[8]), .Q(_50414) );
  nor2s1 _51139_inst ( .DIN1(_28646), .DIN2(______[30]), .Q(_50319) );
  hi1s1 _51140_inst ( .DIN(_49740), .Q(_50056) );
  nnd2s1 _51141_inst ( .DIN1(_50415), .DIN2(_50332), .Q(_49740) );
  nor2s1 _51142_inst ( .DIN1(_33293), .DIN2(_50416), .Q(_50332) );
  nnd2s1 _51143_inst ( .DIN1(_30772), .DIN2(_50417), .Q(_50416) );
  hi1s1 _51144_inst ( .DIN(_35723), .Q(_50417) );
  nnd2s1 _51145_inst ( .DIN1(_50418), .DIN2(_2274), .Q(_35723) );
  nor2s1 _51146_inst ( .DIN1(_2273), .DIN2(_26217), .Q(_50418) );
  hi1s1 _51147_inst ( .DIN(_37987), .Q(_33293) );
  nor2s1 _51148_inst ( .DIN1(_50409), .DIN2(_49915), .Q(_37987) );
  hi1s1 _51149_inst ( .DIN(_50400), .Q(_50409) );
  nor2s1 _51150_inst ( .DIN1(_49187), .DIN2(_27442), .Q(_50415) );
  nnd2s1 _51151_inst ( .DIN1(_50325), .DIN2(_45431), .Q(_27442) );
  nnd2s1 _51152_inst ( .DIN1(_50318), .DIN2(_50348), .Q(_49187) );
  nor2s1 _51153_inst ( .DIN1(______[8]), .DIN2(_49465), .Q(_50318) );
  nor2s1 _51154_inst ( .DIN1(_50419), .DIN2(_49117), .Q(_50402) );
  nnd2s1 _51155_inst ( .DIN1(_49457), .DIN2(_50420), .Q(_49117) );
  nnd2s1 _51156_inst ( .DIN1(_50348), .DIN2(______[8]), .Q(_50420) );
  nor2s1 _51157_inst ( .DIN1(______[30]), .DIN2(______[6]), .Q(_50348) );
  nor2s1 _51158_inst ( .DIN1(_50421), .DIN2(_50422), .Q(_50419) );
  nnd2s1 _51159_inst ( .DIN1(_50423), .DIN2(_50265), .Q(_50422) );
  and2s1 _51160_inst ( .DIN1(_50424), .DIN2(_50425), .Q(_50265) );
  nnd2s1 _51161_inst ( .DIN1(_50426), .DIN2(_50156), .Q(_50425) );
  nor2s1 _51162_inst ( .DIN1(_35720), .DIN2(_37983), .Q(_50156) );
  nnd2s1 _51163_inst ( .DIN1(_50354), .DIN2(_50427), .Q(_37983) );
  nor2s1 _51164_inst ( .DIN1(_34413), .DIN2(_44326), .Q(_50426) );
  nnd2s1 _51165_inst ( .DIN1(_50102), .DIN2(_50276), .Q(_44326) );
  and2s1 _51166_inst ( .DIN1(_50394), .DIN2(_2179), .Q(_50102) );
  nor2s1 _51167_inst ( .DIN1(_2182), .DIN2(_2180), .Q(_50394) );
  nnd2s1 _51168_inst ( .DIN1(_50428), .DIN2(_34414), .Q(_50424) );
  nor2s1 _51169_inst ( .DIN1(_50429), .DIN2(_50413), .Q(_34414) );
  nnd2s1 _51170_inst ( .DIN1(_26370), .DIN2(_26210), .Q(_50429) );
  nor2s1 _51171_inst ( .DIN1(_27446), .DIN2(_50187), .Q(_50428) );
  nnd2s1 _51172_inst ( .DIN1(_31195), .DIN2(_39319), .Q(_50187) );
  hi1s1 _51173_inst ( .DIN(_39282), .Q(_39319) );
  hi1s1 _51174_inst ( .DIN(_50306), .Q(_31195) );
  nnd2s1 _51175_inst ( .DIN1(_50430), .DIN2(_50354), .Q(_50306) );
  nor2s1 _51176_inst ( .DIN1(_26294), .DIN2(_2253), .Q(_50354) );
  nnd2s1 _51177_inst ( .DIN1(_50325), .DIN2(_50276), .Q(_27446) );
  and2s1 _51178_inst ( .DIN1(_50431), .DIN2(_2182), .Q(_50325) );
  nor2s1 _51179_inst ( .DIN1(_2180), .DIN2(_2179), .Q(_50431) );
  nor2s1 _51180_inst ( .DIN1(_50432), .DIN2(_50299), .Q(_50423) );
  nnd2s1 _51181_inst ( .DIN1(_50433), .DIN2(_50434), .Q(_50299) );
  nnd2s1 _51182_inst ( .DIN1(_50435), .DIN2(_50122), .Q(_50434) );
  nor2s1 _51183_inst ( .DIN1(_39282), .DIN2(_37942), .Q(_50122) );
  nnd2s1 _51184_inst ( .DIN1(_50436), .DIN2(_53522), .Q(_39282) );
  nor2s1 _51185_inst ( .DIN1(_2274), .DIN2(_2273), .Q(_50436) );
  nor2s1 _51186_inst ( .DIN1(_43422), .DIN2(_34413), .Q(_50435) );
  nnd2s1 _51187_inst ( .DIN1(_50437), .DIN2(_2216), .Q(_34413) );
  nor2s1 _51188_inst ( .DIN1(_2217), .DIN2(_50413), .Q(_50437) );
  nnd2s1 _51189_inst ( .DIN1(_50438), .DIN2(_50161), .Q(_50433) );
  nor2s1 _51190_inst ( .DIN1(_32091), .DIN2(_35720), .Q(_50161) );
  nnd2s1 _51191_inst ( .DIN1(_50439), .DIN2(_2214), .Q(_32091) );
  nor2s1 _51192_inst ( .DIN1(_2216), .DIN2(_50336), .Q(_50439) );
  nnd2s1 _51193_inst ( .DIN1(_26370), .DIN2(_26248), .Q(_50336) );
  nor2s1 _51194_inst ( .DIN1(_38682), .DIN2(_43497), .Q(_50438) );
  nnd2s1 _51195_inst ( .DIN1(_50400), .DIN2(_50383), .Q(_38682) );
  nor2s1 _51196_inst ( .DIN1(_2252), .DIN2(_2251), .Q(_50400) );
  nor2s1 _51197_inst ( .DIN1(_53266), .DIN2(_49509), .Q(_50432) );
  nnd2s1 _51198_inst ( .DIN1(_50440), .DIN2(_42750), .Q(_49509) );
  hi1s1 _51199_inst ( .DIN(_43497), .Q(_42750) );
  nnd2s1 _51200_inst ( .DIN1(_50291), .DIN2(_50276), .Q(_43497) );
  hi1s1 _51201_inst ( .DIN(_50005), .Q(_50276) );
  nnd2s1 _51202_inst ( .DIN1(_2181), .DIN2(_26419), .Q(_50005) );
  and2s1 _51203_inst ( .DIN1(_50441), .DIN2(_2179), .Q(_50291) );
  nor2s1 _51204_inst ( .DIN1(_2180), .DIN2(_26509), .Q(_50441) );
  nor2s1 _51205_inst ( .DIN1(_30434), .DIN2(_50260), .Q(_50440) );
  nnd2s1 _51206_inst ( .DIN1(_27822), .DIN2(_35301), .Q(_50260) );
  hi1s1 _51207_inst ( .DIN(_36248), .Q(_35301) );
  nnd2s1 _51208_inst ( .DIN1(_50442), .DIN2(_2273), .Q(_36248) );
  hi1s1 _51209_inst ( .DIN(_37942), .Q(_27822) );
  nnd2s1 _51210_inst ( .DIN1(_50443), .DIN2(_2252), .Q(_37942) );
  nor2s1 _51211_inst ( .DIN1(_49915), .DIN2(_26311), .Q(_50443) );
  nnd2s1 _51212_inst ( .DIN1(_50444), .DIN2(_49156), .Q(_50421) );
  nnd2s1 _51213_inst ( .DIN1(_50445), .DIN2(_29767), .Q(_49156) );
  hi1s1 _51214_inst ( .DIN(_32809), .Q(_29767) );
  nnd2s1 _51215_inst ( .DIN1(_49916), .DIN2(_45430), .Q(_32809) );
  and2s1 _51216_inst ( .DIN1(_50446), .DIN2(_2180), .Q(_45430) );
  nor2s1 _51217_inst ( .DIN1(_26509), .DIN2(_26223), .Q(_50446) );
  hi1s1 _51218_inst ( .DIN(_49882), .Q(_49916) );
  nnd2s1 _51219_inst ( .DIN1(_2175), .DIN2(_2181), .Q(_49882) );
  nor2s1 _51220_inst ( .DIN1(_37984), .DIN2(_50170), .Q(_50445) );
  nnd2s1 _51221_inst ( .DIN1(_35724), .DIN2(_30772), .Q(_50170) );
  hi1s1 _51222_inst ( .DIN(_39110), .Q(_30772) );
  nnd2s1 _51223_inst ( .DIN1(_50447), .DIN2(_2216), .Q(_39110) );
  nor2s1 _51224_inst ( .DIN1(_50413), .DIN2(_26370), .Q(_50447) );
  nnd2s1 _51225_inst ( .DIN1(_2203), .DIN2(_2214), .Q(_50413) );
  hi1s1 _51226_inst ( .DIN(_35300), .Q(_35724) );
  nnd2s1 _51227_inst ( .DIN1(_50448), .DIN2(_2274), .Q(_35300) );
  nor2s1 _51228_inst ( .DIN1(_49864), .DIN2(_26217), .Q(_50448) );
  nnd2s1 _51229_inst ( .DIN1(_2238), .DIN2(_49942), .Q(_37984) );
  and2s1 _51230_inst ( .DIN1(_50430), .DIN2(_2253), .Q(_49942) );
  nor2s1 _51231_inst ( .DIN1(_26311), .DIN2(_26706), .Q(_50430) );
  nor2s1 _51232_inst ( .DIN1(_50339), .DIN2(_50347), .Q(_50444) );
  and2s1 _51233_inst ( .DIN1(_50449), .DIN2(_50132), .Q(_50347) );
  nor2s1 _51234_inst ( .DIN1(_50195), .DIN2(_35720), .Q(_50132) );
  hi1s1 _51235_inst ( .DIN(_37931), .Q(_50195) );
  nor2s1 _51236_inst ( .DIN1(_50101), .DIN2(_49915), .Q(_37931) );
  nnd2s1 _51237_inst ( .DIN1(_26709), .DIN2(_26294), .Q(_49915) );
  nnd2s1 _51238_inst ( .DIN1(_2251), .DIN2(_26706), .Q(_50101) );
  nor2s1 _51239_inst ( .DIN1(_30434), .DIN2(_43422), .Q(_50449) );
  nnd2s1 _51240_inst ( .DIN1(_50004), .DIN2(_45431), .Q(_43422) );
  hi1s1 _51241_inst ( .DIN(_49883), .Q(_50004) );
  nnd2s1 _51242_inst ( .DIN1(_50450), .DIN2(_2180), .Q(_49883) );
  nor2s1 _51243_inst ( .DIN1(_2179), .DIN2(_26509), .Q(_50450) );
  nnd2s1 _51244_inst ( .DIN1(_50451), .DIN2(_2216), .Q(_30434) );
  nor2s1 _51245_inst ( .DIN1(_2203), .DIN2(_50382), .Q(_50451) );
  and2s1 _51246_inst ( .DIN1(_50452), .DIN2(_50134), .Q(_50339) );
  nor2s1 _51247_inst ( .DIN1(_35720), .DIN2(_34855), .Q(_50134) );
  nnd2s1 _51248_inst ( .DIN1(_50453), .DIN2(_2216), .Q(_34855) );
  nor2s1 _51249_inst ( .DIN1(_26248), .DIN2(_50382), .Q(_50453) );
  nnd2s1 _51250_inst ( .DIN1(_2217), .DIN2(_26433), .Q(_50382) );
  nnd2s1 _51251_inst ( .DIN1(_50442), .DIN2(_49864), .Q(_35720) );
  hi1s1 _51252_inst ( .DIN(_2273), .Q(_49864) );
  nor2s1 _51253_inst ( .DIN1(_53522), .DIN2(_2274), .Q(_50442) );
  nor2s1 _51254_inst ( .DIN1(_37299), .DIN2(_50316), .Q(_50452) );
  nnd2s1 _51255_inst ( .DIN1(_50263), .DIN2(_45431), .Q(_50316) );
  nor2s1 _51256_inst ( .DIN1(_26419), .DIN2(_2181), .Q(_45431) );
  hi1s1 _51257_inst ( .DIN(_49914), .Q(_50263) );
  nnd2s1 _51258_inst ( .DIN1(_50454), .DIN2(_2180), .Q(_49914) );
  nor2s1 _51259_inst ( .DIN1(_2182), .DIN2(_2179), .Q(_50454) );
  nnd2s1 _51260_inst ( .DIN1(_50427), .DIN2(_50383), .Q(_37299) );
  nor2s1 _51261_inst ( .DIN1(_26709), .DIN2(_2238), .Q(_50383) );
  hi1s1 _51262_inst ( .DIN(_49973), .Q(_50427) );
  nnd2s1 _51263_inst ( .DIN1(_2252), .DIN2(_26311), .Q(_49973) );
  nnd2s1 _51264_inst ( .DIN1(_50455), .DIN2(_50456), .Q(____1___________0[9])
         );
  nor2s1 _51265_inst ( .DIN1(_50457), .DIN2(_50458), .Q(_50456) );
  nnd2s1 _51266_inst ( .DIN1(_50459), .DIN2(_50460), .Q(_50458) );
  nor2s1 _51267_inst ( .DIN1(_50461), .DIN2(_50462), .Q(_50459) );
  nnd2s1 _51268_inst ( .DIN1(_50463), .DIN2(_50464), .Q(_50457) );
  nor2s1 _51269_inst ( .DIN1(_50465), .DIN2(_50466), .Q(_50464) );
  nor2s1 _51270_inst ( .DIN1(_50467), .DIN2(_50468), .Q(_50463) );
  nor2s1 _51271_inst ( .DIN1(_50469), .DIN2(_50470), .Q(_50468) );
  nor2s1 _51272_inst ( .DIN1(_50471), .DIN2(_50472), .Q(_50467) );
  nor2s1 _51273_inst ( .DIN1(_49465), .DIN2(_50473), .Q(_50472) );
  nor2s1 _51274_inst ( .DIN1(_50474), .DIN2(_50475), .Q(_50455) );
  nnd2s1 _51275_inst ( .DIN1(_50476), .DIN2(_50477), .Q(_50475) );
  nor2s1 _51276_inst ( .DIN1(_50478), .DIN2(_50479), .Q(_50476) );
  nnd2s1 _51277_inst ( .DIN1(_50480), .DIN2(_50481), .Q(_50474) );
  nor2s1 _51278_inst ( .DIN1(_50482), .DIN2(_50483), .Q(_50481) );
  nor2s1 _51279_inst ( .DIN1(_50484), .DIN2(_50485), .Q(_50480) );
  nnd2s1 _51280_inst ( .DIN1(_50486), .DIN2(_50487), .Q(____1___________0[8])
         );
  nor2s1 _51281_inst ( .DIN1(_50488), .DIN2(_50489), .Q(_50487) );
  nnd2s1 _51282_inst ( .DIN1(_50490), .DIN2(_50491), .Q(_50489) );
  nor2s1 _51283_inst ( .DIN1(_50492), .DIN2(_50493), .Q(_50491) );
  nor2s1 _51284_inst ( .DIN1(_50494), .DIN2(_50495), .Q(_50493) );
  nor2s1 _51285_inst ( .DIN1(_50496), .DIN2(_50497), .Q(_50490) );
  nor2s1 _51286_inst ( .DIN1(_50498), .DIN2(_50499), .Q(_50497) );
  nor2s1 _51287_inst ( .DIN1(_50500), .DIN2(_50501), .Q(_50496) );
  nnd2s1 _51288_inst ( .DIN1(_50502), .DIN2(_50503), .Q(_50488) );
  nor2s1 _51289_inst ( .DIN1(_50504), .DIN2(_50505), .Q(_50503) );
  or2s1 _51290_inst ( .DIN1(_50506), .DIN2(_50507), .Q(_50505) );
  nor2s1 _51291_inst ( .DIN1(_50508), .DIN2(_50509), .Q(_50502) );
  nor2s1 _51292_inst ( .DIN1(_50510), .DIN2(_50511), .Q(_50509) );
  and2s1 _51293_inst ( .DIN1(_50512), .DIN2(_50513), .Q(_50510) );
  nor2s1 _51294_inst ( .DIN1(_50514), .DIN2(_50515), .Q(_50486) );
  nnd2s1 _51295_inst ( .DIN1(_50516), .DIN2(_50517), .Q(_50515) );
  nor2s1 _51296_inst ( .DIN1(_50518), .DIN2(_50519), .Q(_50517) );
  nor2s1 _51297_inst ( .DIN1(_50520), .DIN2(_50521), .Q(_50516) );
  nnd2s1 _51298_inst ( .DIN1(_50522), .DIN2(_50523), .Q(_50514) );
  nor2s1 _51299_inst ( .DIN1(_50524), .DIN2(_50525), .Q(_50523) );
  nor2s1 _51300_inst ( .DIN1(_50526), .DIN2(_50527), .Q(_50522) );
  nnd2s1 _51301_inst ( .DIN1(_50528), .DIN2(_50529), .Q(____1___________0[7])
         );
  nor2s1 _51302_inst ( .DIN1(_50530), .DIN2(_50531), .Q(_50529) );
  nnd2s1 _51303_inst ( .DIN1(_50532), .DIN2(_50533), .Q(_50531) );
  hi1s1 _51304_inst ( .DIN(_50534), .Q(_50532) );
  nnd2s1 _51305_inst ( .DIN1(_50535), .DIN2(_50536), .Q(_50530) );
  nnd2s1 _51306_inst ( .DIN1(_50537), .DIN2(_50538), .Q(_50536) );
  nor2s1 _51307_inst ( .DIN1(_50539), .DIN2(_50540), .Q(_50535) );
  nor2s1 _51308_inst ( .DIN1(_50541), .DIN2(_50542), .Q(_50528) );
  or2s1 _51309_inst ( .DIN1(_50543), .DIN2(_50544), .Q(_50542) );
  nnd2s1 _51310_inst ( .DIN1(_50545), .DIN2(_50546), .Q(_50541) );
  hi1s1 _51311_inst ( .DIN(_50547), .Q(_50546) );
  nor2s1 _51312_inst ( .DIN1(_50548), .DIN2(_50549), .Q(_50545) );
  nnd2s1 _51313_inst ( .DIN1(_50550), .DIN2(_50551), .Q(____1___________0[6])
         );
  nor2s1 _51314_inst ( .DIN1(_50552), .DIN2(_50553), .Q(_50551) );
  nnd2s1 _51315_inst ( .DIN1(_50554), .DIN2(_50555), .Q(_50553) );
  nor2s1 _51316_inst ( .DIN1(_50556), .DIN2(_50557), .Q(_50555) );
  nor2s1 _51317_inst ( .DIN1(_50558), .DIN2(_50559), .Q(_50554) );
  nor2s1 _51318_inst ( .DIN1(_50560), .DIN2(_50561), .Q(_50559) );
  nor2s1 _51319_inst ( .DIN1(_50562), .DIN2(_50563), .Q(_50558) );
  nnd2s1 _51320_inst ( .DIN1(_50564), .DIN2(_50565), .Q(_50552) );
  nor2s1 _51321_inst ( .DIN1(_50504), .DIN2(_50566), .Q(_50565) );
  nor2s1 _51322_inst ( .DIN1(_50567), .DIN2(_50568), .Q(_50564) );
  nor2s1 _51323_inst ( .DIN1(_50569), .DIN2(_50570), .Q(_50550) );
  nnd2s1 _51324_inst ( .DIN1(_50571), .DIN2(_50572), .Q(_50570) );
  nor2s1 _51325_inst ( .DIN1(_50573), .DIN2(_50574), .Q(_50571) );
  nnd2s1 _51326_inst ( .DIN1(_50575), .DIN2(_50576), .Q(_50569) );
  nor2s1 _51327_inst ( .DIN1(_50577), .DIN2(_50578), .Q(_50576) );
  nor2s1 _51328_inst ( .DIN1(_50547), .DIN2(_50579), .Q(_50575) );
  nnd2s1 _51329_inst ( .DIN1(_50580), .DIN2(_50581), .Q(_50547) );
  nor2s1 _51330_inst ( .DIN1(_50582), .DIN2(_50583), .Q(_50581) );
  nnd2s1 _51331_inst ( .DIN1(_50584), .DIN2(_50585), .Q(_50583) );
  nnd2s1 _51332_inst ( .DIN1(_50586), .DIN2(_50587), .Q(_50585) );
  nnd2s1 _51333_inst ( .DIN1(_50588), .DIN2(_50589), .Q(_50584) );
  nor2s1 _51334_inst ( .DIN1(_50590), .DIN2(_50591), .Q(_50582) );
  nor2s1 _51335_inst ( .DIN1(_50592), .DIN2(_50593), .Q(_50580) );
  nnd2s1 _51336_inst ( .DIN1(_50594), .DIN2(_50595), .Q(____1___________0[5])
         );
  nor2s1 _51337_inst ( .DIN1(_50596), .DIN2(_50597), .Q(_50595) );
  nnd2s1 _51338_inst ( .DIN1(_50598), .DIN2(_50599), .Q(_50597) );
  hi1s1 _51339_inst ( .DIN(_50482), .Q(_50599) );
  nnd2s1 _51340_inst ( .DIN1(_50600), .DIN2(_50601), .Q(_50482) );
  nnd2s1 _51341_inst ( .DIN1(_50602), .DIN2(_50537), .Q(_50601) );
  nor2s1 _51342_inst ( .DIN1(_50603), .DIN2(_50604), .Q(_50600) );
  nor2s1 _51343_inst ( .DIN1(_50605), .DIN2(_50606), .Q(_50604) );
  nor2s1 _51344_inst ( .DIN1(_50607), .DIN2(_50608), .Q(_50598) );
  nnd2s1 _51345_inst ( .DIN1(_50609), .DIN2(_50610), .Q(_50596) );
  nor2s1 _51346_inst ( .DIN1(_50568), .DIN2(_50611), .Q(_50609) );
  nor2s1 _51347_inst ( .DIN1(_50469), .DIN2(_50612), .Q(_50611) );
  nor2s1 _51348_inst ( .DIN1(_50613), .DIN2(_50614), .Q(_50594) );
  or2s1 _51349_inst ( .DIN1(_50615), .DIN2(_50616), .Q(_50614) );
  nnd2s1 _51350_inst ( .DIN1(_50617), .DIN2(_50618), .Q(_50613) );
  nor2s1 _51351_inst ( .DIN1(_50619), .DIN2(_50620), .Q(_50617) );
  nnd2s1 _51352_inst ( .DIN1(_50621), .DIN2(_50622), .Q(____1___________0[4])
         );
  nor2s1 _51353_inst ( .DIN1(_50623), .DIN2(_50624), .Q(_50622) );
  nnd2s1 _51354_inst ( .DIN1(_50625), .DIN2(_50626), .Q(_50624) );
  nor2s1 _51355_inst ( .DIN1(_50627), .DIN2(_50628), .Q(_50626) );
  nor2s1 _51356_inst ( .DIN1(_50629), .DIN2(_50630), .Q(_50627) );
  nor2s1 _51357_inst ( .DIN1(_50631), .DIN2(_50478), .Q(_50625) );
  nnd2s1 _51358_inst ( .DIN1(_50632), .DIN2(_50633), .Q(_50623) );
  nor2s1 _51359_inst ( .DIN1(_50508), .DIN2(_50634), .Q(_50633) );
  nor2s1 _51360_inst ( .DIN1(_50635), .DIN2(_50636), .Q(_50632) );
  nor2s1 _51361_inst ( .DIN1(_50637), .DIN2(_50638), .Q(_50636) );
  nor2s1 _51362_inst ( .DIN1(_50639), .DIN2(_50640), .Q(_50621) );
  nnd2s1 _51363_inst ( .DIN1(_50641), .DIN2(_50642), .Q(_50640) );
  hi1s1 _51364_inst ( .DIN(_50643), .Q(_50642) );
  nor2s1 _51365_inst ( .DIN1(_50644), .DIN2(_50645), .Q(_50641) );
  nnd2s1 _51366_inst ( .DIN1(_50646), .DIN2(_50647), .Q(_50639) );
  nor2s1 _51367_inst ( .DIN1(_50648), .DIN2(_50574), .Q(_50647) );
  nor2s1 _51368_inst ( .DIN1(_50620), .DIN2(_50649), .Q(_50646) );
  nnd2s1 _51369_inst ( .DIN1(_50650), .DIN2(_50651), .Q(_50620) );
  nor2s1 _51370_inst ( .DIN1(_50539), .DIN2(_50567), .Q(_50650) );
  nnd2s1 _51371_inst ( .DIN1(_50652), .DIN2(_50653), .Q(____1___________0[3])
         );
  nor2s1 _51372_inst ( .DIN1(_50654), .DIN2(_50655), .Q(_50653) );
  nnd2s1 _51373_inst ( .DIN1(_50656), .DIN2(_50657), .Q(_50655) );
  nor2s1 _51374_inst ( .DIN1(_50492), .DIN2(_50658), .Q(_50657) );
  nor2s1 _51375_inst ( .DIN1(_50637), .DIN2(_50659), .Q(_50658) );
  nor2s1 _51376_inst ( .DIN1(_50660), .DIN2(_50661), .Q(_50492) );
  nor2s1 _51377_inst ( .DIN1(_50662), .DIN2(_50663), .Q(_50656) );
  nor2s1 _51378_inst ( .DIN1(_50591), .DIN2(_50664), .Q(_50663) );
  nor2s1 _51379_inst ( .DIN1(_50665), .DIN2(_50666), .Q(_50662) );
  nnd2s1 _51380_inst ( .DIN1(_50667), .DIN2(_50668), .Q(_50654) );
  nor2s1 _51381_inst ( .DIN1(_50669), .DIN2(_50635), .Q(_50668) );
  nor2s1 _51382_inst ( .DIN1(_50670), .DIN2(_50671), .Q(_50635) );
  nor2s1 _51383_inst ( .DIN1(_50672), .DIN2(_50673), .Q(_50667) );
  nor2s1 _51384_inst ( .DIN1(_50562), .DIN2(_50612), .Q(_50673) );
  nor2s1 _51385_inst ( .DIN1(_50674), .DIN2(_50675), .Q(_50652) );
  nnd2s1 _51386_inst ( .DIN1(_50676), .DIN2(_50677), .Q(_50675) );
  nor2s1 _51387_inst ( .DIN1(_50678), .DIN2(_50679), .Q(_50676) );
  nnd2s1 _51388_inst ( .DIN1(_50680), .DIN2(_50681), .Q(_50674) );
  nor2s1 _51389_inst ( .DIN1(_50682), .DIN2(_50593), .Q(_50681) );
  nnd2s1 _51390_inst ( .DIN1(_50683), .DIN2(_50684), .Q(_50593) );
  nor2s1 _51391_inst ( .DIN1(_50685), .DIN2(_50686), .Q(_50684) );
  nor2s1 _51392_inst ( .DIN1(_50687), .DIN2(_50513), .Q(_50686) );
  nor2s1 _51393_inst ( .DIN1(_50560), .DIN2(_50688), .Q(_50685) );
  nor2s1 _51394_inst ( .DIN1(_50689), .DIN2(_50690), .Q(_50683) );
  nor2s1 _51395_inst ( .DIN1(_50471), .DIN2(_50691), .Q(_50690) );
  nor2s1 _51396_inst ( .DIN1(_50692), .DIN2(_50511), .Q(_50689) );
  nor2s1 _51397_inst ( .DIN1(_50693), .DIN2(_50694), .Q(_50680) );
  nnd2s1 _51398_inst ( .DIN1(_50695), .DIN2(_50696), .Q(____1___________0[2])
         );
  nor2s1 _51399_inst ( .DIN1(_50697), .DIN2(_50698), .Q(_50696) );
  nnd2s1 _51400_inst ( .DIN1(_50699), .DIN2(_50700), .Q(_50698) );
  nor2s1 _51401_inst ( .DIN1(_50701), .DIN2(_50461), .Q(_50700) );
  nor2s1 _51402_inst ( .DIN1(_50494), .DIN2(_50702), .Q(_50461) );
  nor2s1 _51403_inst ( .DIN1(_50703), .DIN2(_50704), .Q(_50701) );
  nor2s1 _51404_inst ( .DIN1(_50705), .DIN2(_50706), .Q(_50699) );
  nor2s1 _51405_inst ( .DIN1(_50707), .DIN2(_50708), .Q(_50705) );
  nnd2s1 _51406_inst ( .DIN1(_50709), .DIN2(_50710), .Q(_50697) );
  nor2s1 _51407_inst ( .DIN1(_50603), .DIN2(_50711), .Q(_50710) );
  or2s1 _51408_inst ( .DIN1(_50669), .DIN2(_50567), .Q(_50711) );
  nor2s1 _51409_inst ( .DIN1(_50470), .DIN2(_50670), .Q(_50567) );
  nor2s1 _51410_inst ( .DIN1(_50712), .DIN2(_50713), .Q(_50709) );
  nor2s1 _51411_inst ( .DIN1(_50714), .DIN2(_50715), .Q(_50695) );
  nnd2s1 _51412_inst ( .DIN1(_50716), .DIN2(_50717), .Q(_50715) );
  nor2s1 _51413_inst ( .DIN1(_50527), .DIN2(_50549), .Q(_50717) );
  nnd2s1 _51414_inst ( .DIN1(_50718), .DIN2(_50719), .Q(_50549) );
  nor2s1 _51415_inst ( .DIN1(_50720), .DIN2(_50721), .Q(_50719) );
  nnd2s1 _51416_inst ( .DIN1(_50722), .DIN2(_50723), .Q(_50721) );
  nor2s1 _51417_inst ( .DIN1(_50724), .DIN2(_50725), .Q(_50723) );
  and2s1 _51418_inst ( .DIN1(_50726), .DIN2(_50727), .Q(_50724) );
  nor2s1 _51419_inst ( .DIN1(_50728), .DIN2(_50729), .Q(_50722) );
  nor2s1 _51420_inst ( .DIN1(_50605), .DIN2(_50660), .Q(_50729) );
  nor2s1 _51421_inst ( .DIN1(_50562), .DIN2(_50730), .Q(_50728) );
  nnd2s1 _51422_inst ( .DIN1(_50731), .DIN2(_50732), .Q(_50720) );
  nor2s1 _51423_inst ( .DIN1(_50733), .DIN2(_50734), .Q(_50732) );
  nor2s1 _51424_inst ( .DIN1(_50735), .DIN2(_50736), .Q(_50731) );
  nor2s1 _51425_inst ( .DIN1(_50737), .DIN2(_50738), .Q(_50736) );
  or2s1 _51426_inst ( .DIN1(_50739), .DIN2(_50740), .Q(_50738) );
  nnd2s1 _51427_inst ( .DIN1(_50741), .DIN2(_44570), .Q(_50737) );
  hi1s1 _51428_inst ( .DIN(_50742), .Q(_44570) );
  nor2s1 _51429_inst ( .DIN1(_50469), .DIN2(_50743), .Q(_50741) );
  nor2s1 _51430_inst ( .DIN1(_50744), .DIN2(_50745), .Q(_50718) );
  nnd2s1 _51431_inst ( .DIN1(_50746), .DIN2(_50747), .Q(_50745) );
  nor2s1 _51432_inst ( .DIN1(_50648), .DIN2(_50748), .Q(_50746) );
  nnd2s1 _51433_inst ( .DIN1(_50749), .DIN2(_50750), .Q(_50648) );
  nnd2s1 _51434_inst ( .DIN1(_50751), .DIN2(_50752), .Q(_50750) );
  nnd2s1 _51435_inst ( .DIN1(_50753), .DIN2(_50754), .Q(_50749) );
  nnd2s1 _51436_inst ( .DIN1(_50755), .DIN2(_50756), .Q(_50744) );
  nor2s1 _51437_inst ( .DIN1(_50607), .DIN2(_50526), .Q(_50756) );
  nnd2s1 _51438_inst ( .DIN1(_50757), .DIN2(_50758), .Q(_50526) );
  nor2s1 _51439_inst ( .DIN1(_50759), .DIN2(_50760), .Q(_50758) );
  nnd2s1 _51440_inst ( .DIN1(_50761), .DIN2(_50762), .Q(_50760) );
  nnd2s1 _51441_inst ( .DIN1(_50763), .DIN2(_50764), .Q(_50761) );
  nnd2s1 _51442_inst ( .DIN1(_50765), .DIN2(_50766), .Q(_50759) );
  nor2s1 _51443_inst ( .DIN1(_50767), .DIN2(_50768), .Q(_50757) );
  nnd2s1 _51444_inst ( .DIN1(_50769), .DIN2(_50770), .Q(_50768) );
  nnd2s1 _51445_inst ( .DIN1(_50771), .DIN2(_50772), .Q(_50770) );
  hi1s1 _51446_inst ( .DIN(_50773), .Q(_50769) );
  nnd2s1 _51447_inst ( .DIN1(_50774), .DIN2(_50775), .Q(_50767) );
  nnd2s1 _51448_inst ( .DIN1(_50776), .DIN2(_50777), .Q(_50775) );
  nor2s1 _51449_inst ( .DIN1(_50778), .DIN2(_50779), .Q(_50755) );
  nnd2s1 _51450_inst ( .DIN1(_50780), .DIN2(_50781), .Q(_50527) );
  nor2s1 _51451_inst ( .DIN1(_50782), .DIN2(_50783), .Q(_50781) );
  nor2s1 _51452_inst ( .DIN1(_50784), .DIN2(_50785), .Q(_50780) );
  nor2s1 _51453_inst ( .DIN1(_50786), .DIN2(_50787), .Q(_50785) );
  nor2s1 _51454_inst ( .DIN1(_50788), .DIN2(_50789), .Q(_50716) );
  nnd2s1 _51455_inst ( .DIN1(_50790), .DIN2(_50791), .Q(_50714) );
  nor2s1 _51456_inst ( .DIN1(_50792), .DIN2(_50793), .Q(_50791) );
  nnd2s1 _51457_inst ( .DIN1(_50794), .DIN2(_50795), .Q(_50793) );
  nnd2s1 _51458_inst ( .DIN1(_50796), .DIN2(_50797), .Q(_50795) );
  nor2s1 _51459_inst ( .DIN1(_50665), .DIN2(_50798), .Q(_50792) );
  nor2s1 _51460_inst ( .DIN1(_50799), .DIN2(_50800), .Q(_50790) );
  nnd2s1 _51461_inst ( .DIN1(_50801), .DIN2(_50802), .Q(____1___________0[1])
         );
  nor2s1 _51462_inst ( .DIN1(_50803), .DIN2(_50804), .Q(_50802) );
  nnd2s1 _51463_inst ( .DIN1(_50805), .DIN2(_50806), .Q(_50804) );
  or2s1 _51464_inst ( .DIN1(_50495), .DIN2(_50494), .Q(_50806) );
  nnd2s1 _51465_inst ( .DIN1(_50807), .DIN2(_50808), .Q(_50803) );
  nor2s1 _51466_inst ( .DIN1(_50809), .DIN2(_50810), .Q(_50807) );
  nor2s1 _51467_inst ( .DIN1(_50562), .DIN2(_50811), .Q(_50810) );
  hi1s1 _51468_inst ( .DIN(_50812), .Q(_50809) );
  nor2s1 _51469_inst ( .DIN1(_50813), .DIN2(_50814), .Q(_50801) );
  nnd2s1 _51470_inst ( .DIN1(_50815), .DIN2(_50618), .Q(_50814) );
  and2s1 _51471_inst ( .DIN1(_50816), .DIN2(_50817), .Q(_50618) );
  nor2s1 _51472_inst ( .DIN1(_50818), .DIN2(_50819), .Q(_50817) );
  nnd2s1 _51473_inst ( .DIN1(_50820), .DIN2(_50821), .Q(_50819) );
  nnd2s1 _51474_inst ( .DIN1(_50822), .DIN2(_50823), .Q(_50821) );
  nnd2s1 _51475_inst ( .DIN1(_50824), .DIN2(_50825), .Q(_50820) );
  nnd2s1 _51476_inst ( .DIN1(_50826), .DIN2(_50827), .Q(_50818) );
  nnd2s1 _51477_inst ( .DIN1(_50537), .DIN2(_50828), .Q(_50827) );
  nnd2s1 _51478_inst ( .DIN1(_50829), .DIN2(_50830), .Q(_50828) );
  nor2s1 _51479_inst ( .DIN1(_50831), .DIN2(_50832), .Q(_50816) );
  nnd2s1 _51480_inst ( .DIN1(_50833), .DIN2(_50834), .Q(_50832) );
  nnd2s1 _51481_inst ( .DIN1(_50835), .DIN2(_50836), .Q(_50834) );
  nor2s1 _51482_inst ( .DIN1(_50605), .DIN2(_50837), .Q(_50831) );
  hi1s1 _51483_inst ( .DIN(_50645), .Q(_50815) );
  nnd2s1 _51484_inst ( .DIN1(_50838), .DIN2(_50839), .Q(_50645) );
  nor2s1 _51485_inst ( .DIN1(_50840), .DIN2(_50841), .Q(_50839) );
  nor2s1 _51486_inst ( .DIN1(_50498), .DIN2(_50842), .Q(_50841) );
  and2s1 _51487_inst ( .DIN1(_50727), .DIN2(_50843), .Q(_50840) );
  nor2s1 _51488_inst ( .DIN1(_50844), .DIN2(_50845), .Q(_50838) );
  nor2s1 _51489_inst ( .DIN1(_50511), .DIN2(_50512), .Q(_50845) );
  or2s1 _51490_inst ( .DIN1(_50579), .DIN2(_50483), .Q(_50813) );
  nnd2s1 _51491_inst ( .DIN1(_50846), .DIN2(_50847), .Q(_50483) );
  nor2s1 _51492_inst ( .DIN1(_50848), .DIN2(_50849), .Q(_50847) );
  nnd2s1 _51493_inst ( .DIN1(_50850), .DIN2(_50851), .Q(_50849) );
  nor2s1 _51494_inst ( .DIN1(_50852), .DIN2(_50853), .Q(_50850) );
  nor2s1 _51495_inst ( .DIN1(_50665), .DIN2(_50854), .Q(_50853) );
  nnd2s1 _51496_inst ( .DIN1(_50855), .DIN2(_50856), .Q(_50848) );
  nor2s1 _51497_inst ( .DIN1(_50540), .DIN2(_50735), .Q(_50855) );
  hi1s1 _51498_inst ( .DIN(_50857), .Q(_50540) );
  nor2s1 _51499_inst ( .DIN1(_50858), .DIN2(_50859), .Q(_50846) );
  or2s1 _51500_inst ( .DIN1(_50860), .DIN2(_50861), .Q(_50859) );
  nnd2s1 _51501_inst ( .DIN1(_50862), .DIN2(_50863), .Q(_50858) );
  nor2s1 _51502_inst ( .DIN1(_50608), .DIN2(_50631), .Q(_50862) );
  nnd2s1 _51503_inst ( .DIN1(_50864), .DIN2(_50865), .Q(_50631) );
  hi1s1 _51504_inst ( .DIN(_50866), .Q(_50865) );
  nor2s1 _51505_inst ( .DIN1(_50867), .DIN2(_50868), .Q(_50864) );
  nor2s1 _51506_inst ( .DIN1(_50869), .DIN2(_50664), .Q(_50867) );
  nnd2s1 _51507_inst ( .DIN1(_50870), .DIN2(_50871), .Q(_50608) );
  nor2s1 _51508_inst ( .DIN1(_50872), .DIN2(_50873), .Q(_50870) );
  nor2s1 _51509_inst ( .DIN1(_50874), .DIN2(_50666), .Q(_50872) );
  nnd2s1 _51510_inst ( .DIN1(_50875), .DIN2(_50876), .Q(_50579) );
  nor2s1 _51511_inst ( .DIN1(_50783), .DIN2(_50524), .Q(_50875) );
  nor2s1 _51512_inst ( .DIN1(_50877), .DIN2(_50664), .Q(_50524) );
  hi1s1 _51513_inst ( .DIN(_50878), .Q(_50783) );
  nnd2s1 _51514_inst ( .DIN1(_50879), .DIN2(_50880), .Q(____1___________0[15])
         );
  nor2s1 _51515_inst ( .DIN1(_50881), .DIN2(_50882), .Q(_50880) );
  nnd2s1 _51516_inst ( .DIN1(_50883), .DIN2(_50884), .Q(_50882) );
  nor2s1 _51517_inst ( .DIN1(_50885), .DIN2(_50886), .Q(_50884) );
  nor2s1 _51518_inst ( .DIN1(_50687), .DIN2(_50887), .Q(_50886) );
  nor2s1 _51519_inst ( .DIN1(_50888), .DIN2(_50889), .Q(_50883) );
  nor2s1 _51520_inst ( .DIN1(_50471), .DIN2(_50499), .Q(_50889) );
  hi1s1 _51521_inst ( .DIN(_50824), .Q(_50499) );
  nnd2s1 _51522_inst ( .DIN1(_50890), .DIN2(_50891), .Q(_50881) );
  nor2s1 _51523_inst ( .DIN1(_50466), .DIN2(_50782), .Q(_50891) );
  nor2s1 _51524_inst ( .DIN1(_50556), .DIN2(_50892), .Q(_50890) );
  nor2s1 _51525_inst ( .DIN1(_50562), .DIN2(_50893), .Q(_50892) );
  nor2s1 _51526_inst ( .DIN1(_50894), .DIN2(_50895), .Q(_50879) );
  nnd2s1 _51527_inst ( .DIN1(_50896), .DIN2(_50897), .Q(_50895) );
  nor2s1 _51528_inst ( .DIN1(_50574), .DIN2(_50788), .Q(_50897) );
  nnd2s1 _51529_inst ( .DIN1(_50898), .DIN2(_50856), .Q(_50788) );
  nnd2s1 _51530_inst ( .DIN1(_50899), .DIN2(_50900), .Q(_50574) );
  or2s1 _51531_inst ( .DIN1(_50811), .DIN2(_50562), .Q(_50900) );
  nor2s1 _51532_inst ( .DIN1(_50901), .DIN2(_50902), .Q(_50899) );
  nor2s1 _51533_inst ( .DIN1(_50874), .DIN2(_50903), .Q(_50902) );
  hi1s1 _51534_inst ( .DIN(_50766), .Q(_50901) );
  nor2s1 _51535_inst ( .DIN1(_50904), .DIN2(_50905), .Q(_50896) );
  nnd2s1 _51536_inst ( .DIN1(_50906), .DIN2(_50907), .Q(_50894) );
  nor2s1 _51537_inst ( .DIN1(_50908), .DIN2(_50909), .Q(_50907) );
  nor2s1 _51538_inst ( .DIN1(_50664), .DIN2(_50910), .Q(_50908) );
  nor2s1 _51539_inst ( .DIN1(_50779), .DIN2(_50548), .Q(_50906) );
  nnd2s1 _51540_inst ( .DIN1(_50911), .DIN2(_50912), .Q(_50548) );
  nnd2s1 _51541_inst ( .DIN1(_50913), .DIN2(_50764), .Q(_50912) );
  hi1s1 _51542_inst ( .DIN(_50914), .Q(_50764) );
  nnd2s1 _51543_inst ( .DIN1(_50915), .DIN2(_50916), .Q(_50911) );
  nnd2s1 _51544_inst ( .DIN1(_50917), .DIN2(_50918), .Q(_50779) );
  nnd2s1 _51545_inst ( .DIN1(_50919), .DIN2(_50920), .Q(_50918) );
  nor2s1 _51546_inst ( .DIN1(_50921), .DIN2(_50922), .Q(_50917) );
  hi1s1 _51547_inst ( .DIN(_50923), .Q(_50922) );
  nnd2s1 _51548_inst ( .DIN1(_50924), .DIN2(_50925), .Q(____1___________0[14])
         );
  nor2s1 _51549_inst ( .DIN1(_50926), .DIN2(_50927), .Q(_50925) );
  nnd2s1 _51550_inst ( .DIN1(_50928), .DIN2(_50929), .Q(_50927) );
  nor2s1 _51551_inst ( .DIN1(_50930), .DIN2(_50931), .Q(_50929) );
  nor2s1 _51552_inst ( .DIN1(_50471), .DIN2(_50932), .Q(_50931) );
  nor2s1 _51553_inst ( .DIN1(_50501), .DIN2(_50933), .Q(_50930) );
  nor2s1 _51554_inst ( .DIN1(_50934), .DIN2(_50935), .Q(_50928) );
  nor2s1 _51555_inst ( .DIN1(_50605), .DIN2(_50798), .Q(_50935) );
  nor2s1 _51556_inst ( .DIN1(_50874), .DIN2(_50936), .Q(_50934) );
  nnd2s1 _51557_inst ( .DIN1(_50937), .DIN2(_50938), .Q(_50926) );
  nor2s1 _51558_inst ( .DIN1(_50939), .DIN2(_50508), .Q(_50938) );
  and2s1 _51559_inst ( .DIN1(_50940), .DIN2(_50941), .Q(_50508) );
  hi1s1 _51560_inst ( .DIN(_50942), .Q(_50939) );
  nor2s1 _51561_inst ( .DIN1(_50943), .DIN2(_50944), .Q(_50937) );
  nor2s1 _51562_inst ( .DIN1(_50945), .DIN2(_50562), .Q(_50944) );
  nor2s1 _51563_inst ( .DIN1(_50946), .DIN2(_50947), .Q(_50945) );
  nnd2s1 _51564_inst ( .DIN1(_50671), .DIN2(_50563), .Q(_50947) );
  nor2s1 _51565_inst ( .DIN1(_50948), .DIN2(_50949), .Q(_50924) );
  nnd2s1 _51566_inst ( .DIN1(_50950), .DIN2(_50951), .Q(_50949) );
  hi1s1 _51567_inst ( .DIN(_50952), .Q(_50951) );
  nor2s1 _51568_inst ( .DIN1(_50694), .DIN2(_50904), .Q(_50950) );
  nnd2s1 _51569_inst ( .DIN1(_50953), .DIN2(_50954), .Q(_50904) );
  nor2s1 _51570_inst ( .DIN1(_50955), .DIN2(_50956), .Q(_50954) );
  nnd2s1 _51571_inst ( .DIN1(_50957), .DIN2(_50958), .Q(_50956) );
  nnd2s1 _51572_inst ( .DIN1(_50959), .DIN2(_50960), .Q(_50958) );
  nor2s1 _51573_inst ( .DIN1(_50961), .DIN2(_50844), .Q(_50957) );
  nor2s1 _51574_inst ( .DIN1(_50962), .DIN2(_50963), .Q(_50844) );
  nor2s1 _51575_inst ( .DIN1(_50605), .DIN2(_50842), .Q(_50961) );
  nnd2s1 _51576_inst ( .DIN1(_50964), .DIN2(_50965), .Q(_50955) );
  nor2s1 _51577_inst ( .DIN1(_50465), .DIN2(_50966), .Q(_50965) );
  nor2s1 _51578_inst ( .DIN1(_50967), .DIN2(_50852), .Q(_50964) );
  hi1s1 _51579_inst ( .DIN(_50765), .Q(_50852) );
  nor2s1 _51580_inst ( .DIN1(_50968), .DIN2(_50969), .Q(_50953) );
  nnd2s1 _51581_inst ( .DIN1(_50970), .DIN2(_50971), .Q(_50969) );
  nor2s1 _51582_inst ( .DIN1(_50789), .DIN2(_50972), .Q(_50970) );
  hi1s1 _51583_inst ( .DIN(_50973), .Q(_50972) );
  nnd2s1 _51584_inst ( .DIN1(_50863), .DIN2(_50974), .Q(_50789) );
  or2s1 _51585_inst ( .DIN1(_50854), .DIN2(_50703), .Q(_50974) );
  and2s1 _51586_inst ( .DIN1(_50975), .DIN2(_50976), .Q(_50863) );
  or2s1 _51587_inst ( .DIN1(_50977), .DIN2(_50665), .Q(_50976) );
  nor2s1 _51588_inst ( .DIN1(_50978), .DIN2(_50979), .Q(_50975) );
  nor2s1 _51589_inst ( .DIN1(_50980), .DIN2(_50981), .Q(_50979) );
  or2s1 _51590_inst ( .DIN1(_50982), .DIN2(_50562), .Q(_50981) );
  nor2s1 _51591_inst ( .DIN1(_50983), .DIN2(_50984), .Q(_50978) );
  nnd2s1 _51592_inst ( .DIN1(_50960), .DIN2(_50985), .Q(_50984) );
  nnd2s1 _51593_inst ( .DIN1(_50986), .DIN2(_50987), .Q(_50983) );
  nor2s1 _51594_inst ( .DIN1(_50743), .DIN2(_50988), .Q(_50986) );
  nnd2s1 _51595_inst ( .DIN1(_50989), .DIN2(_50572), .Q(_50968) );
  and2s1 _51596_inst ( .DIN1(_50990), .DIN2(_50991), .Q(_50572) );
  nor2s1 _51597_inst ( .DIN1(_50992), .DIN2(_50672), .Q(_50990) );
  nor2s1 _51598_inst ( .DIN1(_50993), .DIN2(_50787), .Q(_50672) );
  hi1s1 _51599_inst ( .DIN(_50994), .Q(_50787) );
  nor2s1 _51600_inst ( .DIN1(_50995), .DIN2(_50702), .Q(_50992) );
  nor2s1 _51601_inst ( .DIN1(_50996), .DIN2(_50534), .Q(_50989) );
  nnd2s1 _51602_inst ( .DIN1(_50997), .DIN2(_50998), .Q(_50534) );
  nnd2s1 _51603_inst ( .DIN1(_50999), .DIN2(_50797), .Q(_50998) );
  nor2s1 _51604_inst ( .DIN1(_50590), .DIN2(_51000), .Q(_50996) );
  nnd2s1 _51605_inst ( .DIN1(_51001), .DIN2(_51002), .Q(_50694) );
  nor2s1 _51606_inst ( .DIN1(_50504), .DIN2(_50706), .Q(_51001) );
  nor2s1 _51607_inst ( .DIN1(_50687), .DIN2(_50512), .Q(_50706) );
  and2s1 _51608_inst ( .DIN1(_51003), .DIN2(_51004), .Q(_50504) );
  nnd2s1 _51609_inst ( .DIN1(_51005), .DIN2(_51006), .Q(_50948) );
  nor2s1 _51610_inst ( .DIN1(_51007), .DIN2(_50748), .Q(_51006) );
  nnd2s1 _51611_inst ( .DIN1(_51008), .DIN2(_51009), .Q(_50748) );
  nor2s1 _51612_inst ( .DIN1(_51010), .DIN2(_51011), .Q(_51009) );
  nor2s1 _51613_inst ( .DIN1(_50670), .DIN2(_50893), .Q(_51011) );
  hi1s1 _51614_inst ( .DIN(_51012), .Q(_50893) );
  hi1s1 _51615_inst ( .DIN(_51013), .Q(_51010) );
  nor2s1 _51616_inst ( .DIN1(_51014), .DIN2(_51015), .Q(_51008) );
  nor2s1 _51617_inst ( .DIN1(_50471), .DIN2(_51016), .Q(_51015) );
  nor2s1 _51618_inst ( .DIN1(_50544), .DIN2(_51017), .Q(_51005) );
  nnd2s1 _51619_inst ( .DIN1(_51018), .DIN2(_51019), .Q(_50544) );
  nor2s1 _51620_inst ( .DIN1(_51020), .DIN2(_51021), .Q(_51019) );
  nor2s1 _51621_inst ( .DIN1(_51022), .DIN2(_51023), .Q(_51018) );
  nnd2s1 _51622_inst ( .DIN1(_51024), .DIN2(_51025), .Q(____1___________0[13])
         );
  nor2s1 _51623_inst ( .DIN1(_51026), .DIN2(_51027), .Q(_51025) );
  nnd2s1 _51624_inst ( .DIN1(_51028), .DIN2(_51029), .Q(_51027) );
  nor2s1 _51625_inst ( .DIN1(_50868), .DIN2(_51030), .Q(_51028) );
  nnd2s1 _51626_inst ( .DIN1(_51013), .DIN2(_51031), .Q(_50868) );
  or2s1 _51627_inst ( .DIN1(_51016), .DIN2(_50498), .Q(_51031) );
  nnd2s1 _51628_inst ( .DIN1(_51032), .DIN2(_51033), .Q(_51013) );
  nor2s1 _51629_inst ( .DIN1(_51034), .DIN2(_50494), .Q(_51033) );
  nor2s1 _51630_inst ( .DIN1(_51035), .DIN2(_51036), .Q(_51032) );
  nnd2s1 _51631_inst ( .DIN1(_51037), .DIN2(_51038), .Q(_51026) );
  nor2s1 _51632_inst ( .DIN1(_50507), .DIN2(_50943), .Q(_51038) );
  and2s1 _51633_inst ( .DIN1(_51039), .DIN2(_50923), .Q(_51037) );
  nor2s1 _51634_inst ( .DIN1(_51040), .DIN2(_51041), .Q(_51024) );
  nnd2s1 _51635_inst ( .DIN1(_51042), .DIN2(_51043), .Q(_51041) );
  hi1s1 _51636_inst ( .DIN(_51044), .Q(_51043) );
  nor2s1 _51637_inst ( .DIN1(_51045), .DIN2(_51046), .Q(_51042) );
  nnd2s1 _51638_inst ( .DIN1(_51047), .DIN2(_50973), .Q(_51040) );
  nor2s1 _51639_inst ( .DIN1(_50778), .DIN2(_51048), .Q(_50973) );
  nnd2s1 _51640_inst ( .DIN1(_51049), .DIN2(_51050), .Q(_50778) );
  hi1s1 _51641_inst ( .DIN(_51051), .Q(_51050) );
  nor2s1 _51642_inst ( .DIN1(_51052), .DIN2(_51053), .Q(_51049) );
  nor2s1 _51643_inst ( .DIN1(_51054), .DIN2(_51055), .Q(_51053) );
  or2s1 _51644_inst ( .DIN1(_50560), .DIN2(_44572), .Q(_51055) );
  or2s1 _51645_inst ( .DIN1(_51056), .DIN2(_51057), .Q(_51054) );
  nor2s1 _51646_inst ( .DIN1(_50615), .DIN2(_50678), .Q(_51047) );
  nnd2s1 _51647_inst ( .DIN1(_51058), .DIN2(_51059), .Q(_50678) );
  nor2s1 _51648_inst ( .DIN1(_51060), .DIN2(_51061), .Q(_51059) );
  nnd2s1 _51649_inst ( .DIN1(_51062), .DIN2(_51063), .Q(_51061) );
  nor2s1 _51650_inst ( .DIN1(_51064), .DIN2(_50888), .Q(_51062) );
  nor2s1 _51651_inst ( .DIN1(_50670), .DIN2(_51065), .Q(_50888) );
  hi1s1 _51652_inst ( .DIN(_51066), .Q(_51064) );
  nnd2s1 _51653_inst ( .DIN1(_51067), .DIN2(_51068), .Q(_51060) );
  nor2s1 _51654_inst ( .DIN1(_51069), .DIN2(_50713), .Q(_51067) );
  hi1s1 _51655_inst ( .DIN(_51070), .Q(_51069) );
  nor2s1 _51656_inst ( .DIN1(_51071), .DIN2(_51072), .Q(_51058) );
  nnd2s1 _51657_inst ( .DIN1(_51073), .DIN2(_51074), .Q(_51072) );
  nor2s1 _51658_inst ( .DIN1(_50616), .DIN2(_50649), .Q(_51073) );
  nnd2s1 _51659_inst ( .DIN1(_50898), .DIN2(_51075), .Q(_50649) );
  nnd2s1 _51660_inst ( .DIN1(_51076), .DIN2(_50771), .Q(_51075) );
  and2s1 _51661_inst ( .DIN1(_51077), .DIN2(_51078), .Q(_50898) );
  nnd2s1 _51662_inst ( .DIN1(_50602), .DIN2(_50916), .Q(_51078) );
  nnd2s1 _51663_inst ( .DIN1(_51079), .DIN2(_51080), .Q(_50616) );
  nor2s1 _51664_inst ( .DIN1(_51020), .DIN2(_50556), .Q(_51080) );
  hi1s1 _51665_inst ( .DIN(_50762), .Q(_50556) );
  nnd2s1 _51666_inst ( .DIN1(_51081), .DIN2(_51082), .Q(_50762) );
  nor2s1 _51667_inst ( .DIN1(_51083), .DIN2(_51084), .Q(_51082) );
  hi1s1 _51668_inst ( .DIN(_51085), .Q(_51020) );
  nor2s1 _51669_inst ( .DIN1(_51086), .DIN2(_51087), .Q(_51079) );
  nnd2s1 _51670_inst ( .DIN1(_51088), .DIN2(_51089), .Q(_51071) );
  nor2s1 _51671_inst ( .DIN1(_50866), .DIN2(_50861), .Q(_51088) );
  nnd2s1 _51672_inst ( .DIN1(_51090), .DIN2(_51091), .Q(_50615) );
  nor2s1 _51673_inst ( .DIN1(_50885), .DIN2(_51092), .Q(_51091) );
  nnd2s1 _51674_inst ( .DIN1(_50997), .DIN2(_50766), .Q(_51092) );
  nnd2s1 _51675_inst ( .DIN1(_50946), .DIN2(_51093), .Q(_50766) );
  nnd2s1 _51676_inst ( .DIN1(_50588), .DIN2(_50843), .Q(_50997) );
  nor2s1 _51677_inst ( .DIN1(_50786), .DIN2(_51094), .Q(_50885) );
  nor2s1 _51678_inst ( .DIN1(_51095), .DIN2(_50484), .Q(_51090) );
  nnd2s1 _51679_inst ( .DIN1(_51096), .DIN2(_51097), .Q(_50484) );
  nor2s1 _51680_inst ( .DIN1(_51098), .DIN2(_51099), .Q(_51097) );
  nnd2s1 _51681_inst ( .DIN1(_51100), .DIN2(_50774), .Q(_51099) );
  nnd2s1 _51682_inst ( .DIN1(_51101), .DIN2(_51102), .Q(_50774) );
  nor2s1 _51683_inst ( .DIN1(_50967), .DIN2(_51103), .Q(_51100) );
  nor2s1 _51684_inst ( .DIN1(_50914), .DIN2(_50665), .Q(_51103) );
  nnd2s1 _51685_inst ( .DIN1(_51104), .DIN2(_51105), .Q(_51098) );
  hi1s1 _51686_inst ( .DIN(_51106), .Q(_51105) );
  nor2s1 _51687_inst ( .DIN1(_50506), .DIN2(_50712), .Q(_51104) );
  nor2s1 _51688_inst ( .DIN1(_51107), .DIN2(_51108), .Q(_51096) );
  nnd2s1 _51689_inst ( .DIN1(_51109), .DIN2(_51110), .Q(_51108) );
  nnd2s1 _51690_inst ( .DIN1(_51111), .DIN2(_50805), .Q(_51107) );
  and2s1 _51691_inst ( .DIN1(_51112), .DIN2(_51113), .Q(_50805) );
  nor2s1 _51692_inst ( .DIN1(_51114), .DIN2(_51115), .Q(_51113) );
  nnd2s1 _51693_inst ( .DIN1(_51116), .DIN2(_51117), .Q(_51115) );
  nnd2s1 _51694_inst ( .DIN1(_51118), .DIN2(_51102), .Q(_51117) );
  or2s1 _51695_inst ( .DIN1(_50936), .DIN2(_50874), .Q(_51116) );
  nor2s1 _51696_inst ( .DIN1(_50471), .DIN2(_51119), .Q(_51114) );
  nor2s1 _51697_inst ( .DIN1(_51120), .DIN2(_51121), .Q(_51112) );
  nor2s1 _51698_inst ( .DIN1(_50661), .DIN2(_50691), .Q(_51120) );
  nor2s1 _51699_inst ( .DIN1(_51122), .DIN2(_50682), .Q(_51111) );
  or2s1 _51700_inst ( .DIN1(_51123), .DIN2(_51124), .Q(_50682) );
  nnd2s1 _51701_inst ( .DIN1(_51125), .DIN2(_51126), .Q(____1___________0[12])
         );
  nor2s1 _51702_inst ( .DIN1(_51127), .DIN2(_51128), .Q(_51126) );
  nnd2s1 _51703_inst ( .DIN1(_51129), .DIN2(_51130), .Q(_51128) );
  nor2s1 _51704_inst ( .DIN1(_50557), .DIN2(_51131), .Q(_51130) );
  nor2s1 _51705_inst ( .DIN1(_50562), .DIN2(_50671), .Q(_51131) );
  nor2s1 _51706_inst ( .DIN1(_50661), .DIN2(_50842), .Q(_50557) );
  nor2s1 _51707_inst ( .DIN1(_51132), .DIN2(_51133), .Q(_51129) );
  nor2s1 _51708_inst ( .DIN1(_50659), .DIN2(_50995), .Q(_51133) );
  nnd2s1 _51709_inst ( .DIN1(_51134), .DIN2(_51135), .Q(_51127) );
  nor2s1 _51710_inst ( .DIN1(_50465), .DIN2(_51136), .Q(_51135) );
  nnd2s1 _51711_inst ( .DIN1(_51085), .DIN2(_51070), .Q(_51136) );
  nnd2s1 _51712_inst ( .DIN1(_51137), .DIN2(_51138), .Q(_51085) );
  nor2s1 _51713_inst ( .DIN1(_44998), .DIN2(_50874), .Q(_51137) );
  nor2s1 _51714_inst ( .DIN1(_50962), .DIN2(_50708), .Q(_50465) );
  nor2s1 _51715_inst ( .DIN1(_50784), .DIN2(_51014), .Q(_51134) );
  nor2s1 _51716_inst ( .DIN1(_51094), .DIN2(_50560), .Q(_51014) );
  nor2s1 _51717_inst ( .DIN1(_50469), .DIN2(_50811), .Q(_50784) );
  hi1s1 _51718_inst ( .DIN(_51139), .Q(_50469) );
  nor2s1 _51719_inst ( .DIN1(_51140), .DIN2(_51141), .Q(_51125) );
  nnd2s1 _51720_inst ( .DIN1(_51142), .DIN2(_51143), .Q(_51141) );
  nor2s1 _51721_inst ( .DIN1(_50679), .DIN2(_51046), .Q(_51143) );
  nnd2s1 _51722_inst ( .DIN1(_51144), .DIN2(_51145), .Q(_51046) );
  nor2s1 _51723_inst ( .DIN1(_51022), .DIN2(_51146), .Q(_51145) );
  nnd2s1 _51724_inst ( .DIN1(_50856), .DIN2(_51147), .Q(_51146) );
  hi1s1 _51725_inst ( .DIN(_50566), .Q(_51147) );
  nnd2s1 _51726_inst ( .DIN1(_51148), .DIN2(_51093), .Q(_50856) );
  nor2s1 _51727_inst ( .DIN1(_50874), .DIN2(_50977), .Q(_51022) );
  nnd2s1 _51728_inst ( .DIN1(_51149), .DIN2(_51150), .Q(_50977) );
  nor2s1 _51729_inst ( .DIN1(_51151), .DIN2(_50742), .Q(_51150) );
  nor2s1 _51730_inst ( .DIN1(_51152), .DIN2(_51153), .Q(_51149) );
  nor2s1 _51731_inst ( .DIN1(_51154), .DIN2(_51155), .Q(_51144) );
  nnd2s1 _51732_inst ( .DIN1(_51156), .DIN2(_51157), .Q(_51155) );
  or2s1 _51733_inst ( .DIN1(_50702), .DIN2(_50995), .Q(_51157) );
  nnd2s1 _51734_inst ( .DIN1(_51158), .DIN2(_50537), .Q(_51156) );
  nor2s1 _51735_inst ( .DIN1(_50605), .DIN2(_50563), .Q(_51154) );
  nnd2s1 _51736_inst ( .DIN1(_51159), .DIN2(_51160), .Q(_50679) );
  nor2s1 _51737_inst ( .DIN1(_51161), .DIN2(_51162), .Q(_51160) );
  nnd2s1 _51738_inst ( .DIN1(_51163), .DIN2(_50878), .Q(_51162) );
  nnd2s1 _51739_inst ( .DIN1(_51164), .DIN2(_51165), .Q(_50878) );
  nor2s1 _51740_inst ( .DIN1(_50562), .DIN2(_50988), .Q(_51165) );
  nor2s1 _51741_inst ( .DIN1(_51166), .DIN2(_45000), .Q(_51164) );
  nnd2s1 _51742_inst ( .DIN1(_51012), .DIN2(_51093), .Q(_51163) );
  or2s1 _51743_inst ( .DIN1(_51167), .DIN2(_50603), .Q(_51161) );
  nor2s1 _51744_inst ( .DIN1(_51168), .DIN2(_50995), .Q(_50603) );
  nor2s1 _51745_inst ( .DIN1(_50525), .DIN2(_51169), .Q(_51159) );
  nnd2s1 _51746_inst ( .DIN1(_51170), .DIN2(_51171), .Q(_51169) );
  nnd2s1 _51747_inst ( .DIN1(_50772), .DIN2(_50836), .Q(_51170) );
  hi1s1 _51748_inst ( .DIN(_50869), .Q(_50772) );
  nnd2s1 _51749_inst ( .DIN1(_51172), .DIN2(_51173), .Q(_50525) );
  nnd2s1 _51750_inst ( .DIN1(_50999), .DIN2(_51139), .Q(_51173) );
  hi1s1 _51751_inst ( .DIN(_50470), .Q(_50999) );
  nnd2s1 _51752_inst ( .DIN1(_51174), .DIN2(_51175), .Q(_50470) );
  nor2s1 _51753_inst ( .DIN1(_51176), .DIN2(_51177), .Q(_51175) );
  nnd2s1 _51754_inst ( .DIN1(_2022), .DIN2(_26326), .Q(_51177) );
  nor2s1 _51755_inst ( .DIN1(_51178), .DIN2(_44572), .Q(_51174) );
  nnd2s1 _51756_inst ( .DIN1(_51179), .DIN2(_50537), .Q(_51172) );
  nor2s1 _51757_inst ( .DIN1(_51180), .DIN2(_51181), .Q(_51142) );
  nnd2s1 _51758_inst ( .DIN1(_51182), .DIN2(_51183), .Q(_51140) );
  nor2s1 _51759_inst ( .DIN1(_51184), .DIN2(_51185), .Q(_51183) );
  nor2s1 _51760_inst ( .DIN1(_50829), .DIN2(_50501), .Q(_51185) );
  nor2s1 _51761_inst ( .DIN1(_50629), .DIN2(_51186), .Q(_51184) );
  nor2s1 _51762_inst ( .DIN1(_51187), .DIN2(_50643), .Q(_51182) );
  nnd2s1 _51763_inst ( .DIN1(_51188), .DIN2(_51189), .Q(_50643) );
  nor2s1 _51764_inst ( .DIN1(_51190), .DIN2(_51191), .Q(_51189) );
  nnd2s1 _51765_inst ( .DIN1(_51192), .DIN2(_51193), .Q(_51191) );
  nnd2s1 _51766_inst ( .DIN1(_51194), .DIN2(_50913), .Q(_51192) );
  nor2s1 _51767_inst ( .DIN1(_50498), .DIN2(_51195), .Q(_51190) );
  nor2s1 _51768_inst ( .DIN1(_51196), .DIN2(_51197), .Q(_51188) );
  or2s1 _51769_inst ( .DIN1(_51017), .DIN2(_50518), .Q(_51197) );
  nnd2s1 _51770_inst ( .DIN1(_51198), .DIN2(_51199), .Q(_50518) );
  nor2s1 _51771_inst ( .DIN1(_51200), .DIN2(_51201), .Q(_51199) );
  nnd2s1 _51772_inst ( .DIN1(_50876), .DIN2(_50851), .Q(_51201) );
  nor2s1 _51773_inst ( .DIN1(_51202), .DIN2(_51203), .Q(_50851) );
  nor2s1 _51774_inst ( .DIN1(_50561), .DIN2(_50993), .Q(_51203) );
  nor2s1 _51775_inst ( .DIN1(_50909), .DIN2(_51204), .Q(_50876) );
  and2s1 _51776_inst ( .DIN1(_50919), .DIN2(_50754), .Q(_51204) );
  nnd2s1 _51777_inst ( .DIN1(_51205), .DIN2(_51206), .Q(_50909) );
  nor2s1 _51778_inst ( .DIN1(_51207), .DIN2(_50733), .Q(_51206) );
  and2s1 _51779_inst ( .DIN1(_51208), .DIN2(_51209), .Q(_50733) );
  nor2s1 _51780_inst ( .DIN1(_51210), .DIN2(_51211), .Q(_51209) );
  nor2s1 _51781_inst ( .DIN1(_50560), .DIN2(_44577), .Q(_51208) );
  hi1s1 _51782_inst ( .DIN(_51212), .Q(_51207) );
  nor2s1 _51783_inst ( .DIN1(_51213), .DIN2(_50800), .Q(_51205) );
  nnd2s1 _51784_inst ( .DIN1(_51214), .DIN2(_51215), .Q(_50800) );
  nnd2s1 _51785_inst ( .DIN1(_51216), .DIN2(_51138), .Q(_51215) );
  nor2s1 _51786_inst ( .DIN1(_44998), .DIN2(_50665), .Q(_51216) );
  nor2s1 _51787_inst ( .DIN1(_51217), .DIN2(_51218), .Q(_51214) );
  nor2s1 _51788_inst ( .DIN1(_51219), .DIN2(_51220), .Q(_51218) );
  or2s1 _51789_inst ( .DIN1(_51221), .DIN2(_50687), .Q(_51220) );
  nnd2s1 _51790_inst ( .DIN1(_51222), .DIN2(_51223), .Q(_51219) );
  nor2s1 _51791_inst ( .DIN1(_51224), .DIN2(_51225), .Q(_51217) );
  nnd2s1 _51792_inst ( .DIN1(_50537), .DIN2(_51226), .Q(_51225) );
  nnd2s1 _51793_inst ( .DIN1(_51227), .DIN2(_50985), .Q(_51224) );
  nor2s1 _51794_inst ( .DIN1(_51035), .DIN2(_51228), .Q(_51227) );
  nor2s1 _51795_inst ( .DIN1(_50605), .DIN2(_50730), .Q(_51213) );
  nnd2s1 _51796_inst ( .DIN1(_50610), .DIN2(_51066), .Q(_51200) );
  nnd2s1 _51797_inst ( .DIN1(_51229), .DIN2(_50754), .Q(_50610) );
  nor2s1 _51798_inst ( .DIN1(_51051), .DIN2(_51230), .Q(_51198) );
  or2s1 _51799_inst ( .DIN1(_51030), .DIN2(_51231), .Q(_51230) );
  nor2s1 _51800_inst ( .DIN1(_50707), .DIN2(_51232), .Q(_51187) );
  nnd2s1 _51801_inst ( .DIN1(_51233), .DIN2(_51234), .Q(____1___________0[11])
         );
  nor2s1 _51802_inst ( .DIN1(_51235), .DIN2(_51236), .Q(_51234) );
  nnd2s1 _51803_inst ( .DIN1(_51237), .DIN2(_50826), .Q(_51236) );
  nnd2s1 _51804_inst ( .DIN1(_51238), .DIN2(_51093), .Q(_50826) );
  hi1s1 _51805_inst ( .DIN(_50563), .Q(_51238) );
  nor2s1 _51806_inst ( .DIN1(_50966), .DIN2(_51239), .Q(_51237) );
  nor2s1 _51807_inst ( .DIN1(_51240), .DIN2(_50962), .Q(_51239) );
  nor2s1 _51808_inst ( .DIN1(_50915), .DIN2(_51241), .Q(_51240) );
  hi1s1 _51809_inst ( .DIN(_51242), .Q(_50966) );
  nnd2s1 _51810_inst ( .DIN1(_51243), .DIN2(_51244), .Q(_51235) );
  nor2s1 _51811_inst ( .DIN1(_50539), .DIN2(_50712), .Q(_51244) );
  nor2s1 _51812_inst ( .DIN1(_50995), .DIN2(_50638), .Q(_50712) );
  nor2s1 _51813_inst ( .DIN1(_50702), .DIN2(_50637), .Q(_50539) );
  nnd2s1 _51814_inst ( .DIN1(_51245), .DIN2(_51246), .Q(_50702) );
  nor2s1 _51815_inst ( .DIN1(_50743), .DIN2(_51247), .Q(_51246) );
  nor2s1 _51816_inst ( .DIN1(_50739), .DIN2(_45000), .Q(_51245) );
  nor2s1 _51817_inst ( .DIN1(_50782), .DIN2(_51123), .Q(_51243) );
  nor2s1 _51818_inst ( .DIN1(_51248), .DIN2(_51249), .Q(_51233) );
  nnd2s1 _51819_inst ( .DIN1(_51250), .DIN2(_51251), .Q(_51249) );
  hi1s1 _51820_inst ( .DIN(_51180), .Q(_51251) );
  nnd2s1 _51821_inst ( .DIN1(_51252), .DIN2(_51253), .Q(_51180) );
  nor2s1 _51822_inst ( .DIN1(_51254), .DIN2(_51255), .Q(_51253) );
  nnd2s1 _51823_inst ( .DIN1(_50651), .DIN2(_51077), .Q(_51255) );
  hi1s1 _51824_inst ( .DIN(_51256), .Q(_51077) );
  nnd2s1 _51825_inst ( .DIN1(_50588), .DIN2(_51003), .Q(_50651) );
  hi1s1 _51826_inst ( .DIN(_50995), .Q(_50588) );
  nnd2s1 _51827_inst ( .DIN1(_51257), .DIN2(_50812), .Q(_51254) );
  nor2s1 _51828_inst ( .DIN1(_50466), .DIN2(_50921), .Q(_51257) );
  nor2s1 _51829_inst ( .DIN1(_50590), .DIN2(_50877), .Q(_50466) );
  nor2s1 _51830_inst ( .DIN1(_51258), .DIN2(_51259), .Q(_51252) );
  nnd2s1 _51831_inst ( .DIN1(_50677), .DIN2(_51260), .Q(_51259) );
  hi1s1 _51832_inst ( .DIN(_50861), .Q(_51260) );
  nnd2s1 _51833_inst ( .DIN1(_51261), .DIN2(_51262), .Q(_50861) );
  nnd2s1 _51834_inst ( .DIN1(_51263), .DIN2(_51093), .Q(_51262) );
  nor2s1 _51835_inst ( .DIN1(_51021), .DIN2(_51264), .Q(_51261) );
  nor2s1 _51836_inst ( .DIN1(_51265), .DIN2(_51266), .Q(_51264) );
  or2s1 _51837_inst ( .DIN1(_44577), .DIN2(_50993), .Q(_51266) );
  and2s1 _51838_inst ( .DIN1(_51267), .DIN2(_51268), .Q(_51021) );
  nor2s1 _51839_inst ( .DIN1(_51269), .DIN2(_51270), .Q(_51268) );
  nnd2s1 _51840_inst ( .DIN1(_51271), .DIN2(_51272), .Q(_51270) );
  nor2s1 _51841_inst ( .DIN1(_42876), .DIN2(_50560), .Q(_51267) );
  and2s1 _51842_inst ( .DIN1(_51273), .DIN2(_51274), .Q(_50677) );
  nnd2s1 _51843_inst ( .DIN1(_50771), .DIN2(_51275), .Q(_51274) );
  nnd2s1 _51844_inst ( .DIN1(_50910), .DIN2(_51000), .Q(_51275) );
  nor2s1 _51845_inst ( .DIN1(_51276), .DIN2(_50506), .Q(_51273) );
  nor2s1 _51846_inst ( .DIN1(_50903), .DIN2(_50665), .Q(_50506) );
  nnd2s1 _51847_inst ( .DIN1(_51277), .DIN2(_51278), .Q(_51258) );
  hi1s1 _51848_inst ( .DIN(_51122), .Q(_51278) );
  nnd2s1 _51849_inst ( .DIN1(_50942), .DIN2(_51279), .Q(_51122) );
  nnd2s1 _51850_inst ( .DIN1(_50994), .DIN2(_50941), .Q(_51279) );
  nnd2s1 _51851_inst ( .DIN1(_51280), .DIN2(_51281), .Q(_50942) );
  nnd2s1 _51852_inst ( .DIN1(_51282), .DIN2(_51283), .Q(_51280) );
  nor2s1 _51853_inst ( .DIN1(_51086), .DIN2(_51284), .Q(_51277) );
  nor2s1 _51854_inst ( .DIN1(_50605), .DIN2(_51065), .Q(_51284) );
  nor2s1 _51855_inst ( .DIN1(_50963), .DIN2(_50501), .Q(_51086) );
  nor2s1 _51856_inst ( .DIN1(_50952), .DIN2(_51045), .Q(_51250) );
  nnd2s1 _51857_inst ( .DIN1(_51285), .DIN2(_51286), .Q(_51045) );
  nnd2s1 _51858_inst ( .DIN1(_51179), .DIN2(_50916), .Q(_51286) );
  nnd2s1 _51859_inst ( .DIN1(_51194), .DIN2(_50763), .Q(_51285) );
  hi1s1 _51860_inst ( .DIN(_50798), .Q(_51194) );
  nnd2s1 _51861_inst ( .DIN1(_51287), .DIN2(_51288), .Q(_50952) );
  nor2s1 _51862_inst ( .DIN1(_51289), .DIN2(_51290), .Q(_51288) );
  nnd2s1 _51863_inst ( .DIN1(_51291), .DIN2(_51292), .Q(_51290) );
  nnd2s1 _51864_inst ( .DIN1(_50919), .DIN2(_50960), .Q(_51292) );
  and2s1 _51865_inst ( .DIN1(_51293), .DIN2(_51294), .Q(_50919) );
  nor2s1 _51866_inst ( .DIN1(_51035), .DIN2(_45587), .Q(_51294) );
  nnd2s1 _51867_inst ( .DIN1(_51295), .DIN2(_51296), .Q(_45587) );
  nnd2s1 _51868_inst ( .DIN1(_51148), .DIN2(_51139), .Q(_51291) );
  nor2s1 _51869_inst ( .DIN1(_50513), .DIN2(_50511), .Q(_51289) );
  nor2s1 _51870_inst ( .DIN1(_50485), .DIN2(_51297), .Q(_51287) );
  nnd2s1 _51871_inst ( .DIN1(_50833), .DIN2(_51298), .Q(_51297) );
  nnd2s1 _51872_inst ( .DIN1(_51299), .DIN2(_50916), .Q(_51298) );
  nnd2s1 _51873_inst ( .DIN1(_50473), .DIN2(_50777), .Q(_50833) );
  nnd2s1 _51874_inst ( .DIN1(_51300), .DIN2(_51301), .Q(_50485) );
  hi1s1 _51875_inst ( .DIN(_50628), .Q(_51301) );
  nnd2s1 _51876_inst ( .DIN1(_51039), .DIN2(_50794), .Q(_50628) );
  nnd2s1 _51877_inst ( .DIN1(_50586), .DIN2(_50916), .Q(_50794) );
  hi1s1 _51878_inst ( .DIN(_50830), .Q(_50586) );
  nor2s1 _51879_inst ( .DIN1(_51302), .DIN2(_51303), .Q(_51300) );
  nor2s1 _51880_inst ( .DIN1(_50665), .DIN2(_50837), .Q(_51303) );
  nor2s1 _51881_inst ( .DIN1(_50914), .DIN2(_50874), .Q(_51302) );
  nnd2s1 _51882_inst ( .DIN1(_51304), .DIN2(_51305), .Q(_50914) );
  nor2s1 _51883_inst ( .DIN1(_26326), .DIN2(_51178), .Q(_51304) );
  nnd2s1 _51884_inst ( .DIN1(_51306), .DIN2(_51307), .Q(_51248) );
  hi1s1 _51885_inst ( .DIN(_50573), .Q(_51307) );
  nnd2s1 _51886_inst ( .DIN1(_51308), .DIN2(_51309), .Q(_50573) );
  nor2s1 _51887_inst ( .DIN1(_51310), .DIN2(_51311), .Q(_51309) );
  nnd2s1 _51888_inst ( .DIN1(_51312), .DIN2(_51313), .Q(_51311) );
  hi1s1 _51889_inst ( .DIN(_51314), .Q(_51313) );
  nor2s1 _51890_inst ( .DIN1(_51315), .DIN2(_51023), .Q(_51312) );
  nor2s1 _51891_inst ( .DIN1(_50664), .DIN2(_50630), .Q(_51023) );
  nor2s1 _51892_inst ( .DIN1(_50471), .DIN2(_49457), .Q(_51315) );
  hi1s1 _51893_inst ( .DIN(_51316), .Q(_50471) );
  nnd2s1 _51894_inst ( .DIN1(_51317), .DIN2(_51002), .Q(_51310) );
  nnd2s1 _51895_inst ( .DIN1(_51229), .DIN2(_50920), .Q(_51002) );
  nor2s1 _51896_inst ( .DIN1(_51318), .DIN2(_51319), .Q(_51317) );
  nor2s1 _51897_inst ( .DIN1(_50590), .DIN2(_50869), .Q(_51319) );
  nor2s1 _51898_inst ( .DIN1(_51320), .DIN2(_51321), .Q(_51308) );
  nnd2s1 _51899_inst ( .DIN1(_51322), .DIN2(_51323), .Q(_51321) );
  hi1s1 _51900_inst ( .DIN(_50619), .Q(_51322) );
  nnd2s1 _51901_inst ( .DIN1(_51324), .DIN2(_51325), .Q(_50619) );
  nor2s1 _51902_inst ( .DIN1(_51326), .DIN2(_51327), .Q(_51325) );
  nnd2s1 _51903_inst ( .DIN1(_51171), .DIN2(_51328), .Q(_51327) );
  nnd2s1 _51904_inst ( .DIN1(_51158), .DIN2(_50916), .Q(_51328) );
  hi1s1 _51905_inst ( .DIN(_50962), .Q(_50916) );
  hi1s1 _51906_inst ( .DIN(_50933), .Q(_51158) );
  nnd2s1 _51907_inst ( .DIN1(_51329), .DIN2(_51330), .Q(_50933) );
  nnd2s1 _51908_inst ( .DIN1(_50940), .DIN2(_50823), .Q(_51171) );
  nnd2s1 _51909_inst ( .DIN1(_51331), .DIN2(_51066), .Q(_51326) );
  nnd2s1 _51910_inst ( .DIN1(_51332), .DIN2(_51333), .Q(_51066) );
  nor2s1 _51911_inst ( .DIN1(_50740), .DIN2(_51334), .Q(_51333) );
  or2s1 _51912_inst ( .DIN1(_50742), .DIN2(_50743), .Q(_51334) );
  nor2s1 _51913_inst ( .DIN1(_50670), .DIN2(_50739), .Q(_51332) );
  nnd2s1 _51914_inst ( .DIN1(_51335), .DIN2(_50771), .Q(_51331) );
  hi1s1 _51915_inst ( .DIN(_50664), .Q(_50771) );
  nor2s1 _51916_inst ( .DIN1(_51336), .DIN2(_51337), .Q(_51324) );
  nnd2s1 _51917_inst ( .DIN1(_51029), .DIN2(_51338), .Q(_51337) );
  hi1s1 _51918_inst ( .DIN(_51196), .Q(_51338) );
  nnd2s1 _51919_inst ( .DIN1(_50857), .DIN2(_51339), .Q(_51196) );
  nnd2s1 _51920_inst ( .DIN1(_50776), .DIN2(_50825), .Q(_51339) );
  hi1s1 _51921_inst ( .DIN(_50498), .Q(_50825) );
  hi1s1 _51922_inst ( .DIN(_50932), .Q(_50776) );
  nnd2s1 _51923_inst ( .DIN1(_51340), .DIN2(_51341), .Q(_50932) );
  nnd2s1 _51924_inst ( .DIN1(_50754), .DIN2(_50959), .Q(_50857) );
  hi1s1 _51925_inst ( .DIN(_50511), .Q(_50754) );
  and2s1 _51926_inst ( .DIN1(_51342), .DIN2(_51343), .Q(_51029) );
  nnd2s1 _51927_inst ( .DIN1(_51012), .DIN2(_51139), .Q(_51343) );
  nnd2s1 _51928_inst ( .DIN1(_50670), .DIN2(_50562), .Q(_51139) );
  or2s1 _51929_inst ( .DIN1(_50660), .DIN2(_50605), .Q(_51342) );
  or2s1 _51930_inst ( .DIN1(_51017), .DIN2(_51051), .Q(_51336) );
  nnd2s1 _51931_inst ( .DIN1(_51344), .DIN2(_51345), .Q(_51051) );
  nnd2s1 _51932_inst ( .DIN1(_51346), .DIN2(_51347), .Q(_51345) );
  nor2s1 _51933_inst ( .DIN1(_51247), .DIN2(_50687), .Q(_51347) );
  nor2s1 _51934_inst ( .DIN1(_40395), .DIN2(_51348), .Q(_51346) );
  nnd2s1 _51935_inst ( .DIN1(_51349), .DIN2(_51350), .Q(_51344) );
  nor2s1 _51936_inst ( .DIN1(_51351), .DIN2(_50494), .Q(_51350) );
  nor2s1 _51937_inst ( .DIN1(_51352), .DIN2(_51353), .Q(_51349) );
  nnd2s1 _51938_inst ( .DIN1(_51354), .DIN2(_51355), .Q(_51017) );
  nnd2s1 _51939_inst ( .DIN1(_51356), .DIN2(_51357), .Q(_51355) );
  nor2s1 _51940_inst ( .DIN1(_50494), .DIN2(_51358), .Q(_51357) );
  nnd2s1 _51941_inst ( .DIN1(_51359), .DIN2(_1986), .Q(_51358) );
  nor2s1 _51942_inst ( .DIN1(_51178), .DIN2(_45000), .Q(_51356) );
  nnd2s1 _51943_inst ( .DIN1(_51360), .DIN2(_51361), .Q(_45000) );
  nnd2s1 _51944_inst ( .DIN1(_51362), .DIN2(_51138), .Q(_51354) );
  and2s1 _51945_inst ( .DIN1(_51363), .DIN2(_51364), .Q(_51138) );
  nor2s1 _51946_inst ( .DIN1(_50742), .DIN2(_50670), .Q(_51362) );
  nnd2s1 _51947_inst ( .DIN1(_51365), .DIN2(_51366), .Q(_51320) );
  hi1s1 _51948_inst ( .DIN(_50519), .Q(_51366) );
  nnd2s1 _51949_inst ( .DIN1(_51367), .DIN2(_51368), .Q(_50519) );
  nor2s1 _51950_inst ( .DIN1(_51124), .DIN2(_51369), .Q(_51368) );
  or2s1 _51951_inst ( .DIN1(_51106), .DIN2(_50634), .Q(_51369) );
  hi1s1 _51952_inst ( .DIN(_51370), .Q(_51124) );
  nor2s1 _51953_inst ( .DIN1(_51007), .DIN2(_51371), .Q(_51367) );
  or2s1 _51954_inst ( .DIN1(_51087), .DIN2(_50866), .Q(_51371) );
  nnd2s1 _51955_inst ( .DIN1(_51372), .DIN2(_51373), .Q(_50866) );
  nnd2s1 _51956_inst ( .DIN1(_51374), .DIN2(_51271), .Q(_51373) );
  nor2s1 _51957_inst ( .DIN1(_51375), .DIN2(_51210), .Q(_51374) );
  nor2s1 _51958_inst ( .DIN1(_51376), .DIN2(_51377), .Q(_51375) );
  nor2s1 _51959_inst ( .DIN1(_45001), .DIN2(_51378), .Q(_51377) );
  nnd2s1 _51960_inst ( .DIN1(_50537), .DIN2(_51330), .Q(_51378) );
  nor2s1 _51961_inst ( .DIN1(_51379), .DIN2(_51380), .Q(_51376) );
  nnd2s1 _51962_inst ( .DIN1(_50960), .DIN2(_50987), .Q(_51380) );
  or2s1 _51963_inst ( .DIN1(_51381), .DIN2(_50874), .Q(_51372) );
  nnd2s1 _51964_inst ( .DIN1(_51382), .DIN2(_51383), .Q(_51087) );
  nnd2s1 _51965_inst ( .DIN1(_50538), .DIN2(_50587), .Q(_51383) );
  hi1s1 _51966_inst ( .DIN(_50708), .Q(_50538) );
  nnd2s1 _51967_inst ( .DIN1(_51384), .DIN2(_51385), .Q(_50708) );
  nor2s1 _51968_inst ( .DIN1(_51386), .DIN2(_51387), .Q(_51385) );
  nor2s1 _51969_inst ( .DIN1(_51152), .DIN2(_44620), .Q(_51384) );
  nnd2s1 _51970_inst ( .DIN1(_50727), .DIN2(_50726), .Q(_51382) );
  nnd2s1 _51971_inst ( .DIN1(_51388), .DIN2(_51389), .Q(_50726) );
  nnd2s1 _51972_inst ( .DIN1(_51390), .DIN2(_51391), .Q(_51389) );
  nor2s1 _51973_inst ( .DIN1(_51392), .DIN2(_51393), .Q(_51391) );
  nor2s1 _51974_inst ( .DIN1(_51394), .DIN2(_44626), .Q(_51390) );
  nnd2s1 _51975_inst ( .DIN1(_45588), .DIN2(_51296), .Q(_44626) );
  nnd2s1 _51976_inst ( .DIN1(_51081), .DIN2(_51395), .Q(_51388) );
  nor2s1 _51977_inst ( .DIN1(_50743), .DIN2(_51152), .Q(_51395) );
  nor2s1 _51978_inst ( .DIN1(_51396), .DIN2(_44999), .Q(_51081) );
  nnd2s1 _51979_inst ( .DIN1(_51109), .DIN2(_51397), .Q(_51007) );
  nnd2s1 _51980_inst ( .DIN1(_51398), .DIN2(_50777), .Q(_51397) );
  nor2s1 _51981_inst ( .DIN1(_51399), .DIN2(_50860), .Q(_51365) );
  nnd2s1 _51982_inst ( .DIN1(_51400), .DIN2(_51401), .Q(_50860) );
  hi1s1 _51983_inst ( .DIN(_51048), .Q(_51401) );
  nor2s1 _51984_inst ( .DIN1(_50704), .DIN2(_50665), .Q(_51048) );
  nor2s1 _51985_inst ( .DIN1(_51052), .DIN2(_51402), .Q(_51400) );
  nor2s1 _51986_inst ( .DIN1(_50873), .DIN2(_50478), .Q(_51306) );
  nnd2s1 _51987_inst ( .DIN1(_51403), .DIN2(_51404), .Q(_50478) );
  hi1s1 _51988_inst ( .DIN(_50607), .Q(_51403) );
  nnd2s1 _51989_inst ( .DIN1(_51405), .DIN2(_51406), .Q(_50607) );
  nnd2s1 _51990_inst ( .DIN1(_51407), .DIN2(_51408), .Q(_51406) );
  nor2s1 _51991_inst ( .DIN1(_50670), .DIN2(_50982), .Q(_51407) );
  nnd2s1 _51992_inst ( .DIN1(_51409), .DIN2(_51410), .Q(_50982) );
  nor2s1 _51993_inst ( .DIN1(_26415), .DIN2(_51411), .Q(_51410) );
  nnd2s1 _51994_inst ( .DIN1(_2025), .DIN2(_2064), .Q(_51411) );
  nor2s1 _51995_inst ( .DIN1(_51412), .DIN2(_42877), .Q(_51409) );
  nnd2s1 _51996_inst ( .DIN1(_51263), .DIN2(_50797), .Q(_51405) );
  and2s1 _51997_inst ( .DIN1(_51413), .DIN2(_51414), .Q(_51263) );
  nor2s1 _51998_inst ( .DIN1(_51152), .DIN2(_26326), .Q(_51414) );
  nor2s1 _51999_inst ( .DIN1(_51178), .DIN2(_44994), .Q(_51413) );
  nor2s1 _52000_inst ( .DIN1(_50590), .DIN2(_51186), .Q(_50873) );
  nnd2s1 _52001_inst ( .DIN1(_51415), .DIN2(_51416), .Q(____1___________0[10])
         );
  nor2s1 _52002_inst ( .DIN1(_51417), .DIN2(_51418), .Q(_51416) );
  nnd2s1 _52003_inst ( .DIN1(_51419), .DIN2(_51420), .Q(_51418) );
  nor2s1 _52004_inst ( .DIN1(_51421), .DIN2(_50725), .Q(_51420) );
  nor2s1 _52005_inst ( .DIN1(_50703), .DIN2(_50903), .Q(_50725) );
  nnd2s1 _52006_inst ( .DIN1(_51422), .DIN2(_51423), .Q(_50903) );
  nor2s1 _52007_inst ( .DIN1(_51424), .DIN2(_50664), .Q(_51421) );
  nor2s1 _52008_inst ( .DIN1(_51101), .DIN2(_50835), .Q(_51424) );
  hi1s1 _52009_inst ( .DIN(_51000), .Q(_51101) );
  nnd2s1 _52010_inst ( .DIN1(_51425), .DIN2(_51422), .Q(_51000) );
  hi1s1 _52011_inst ( .DIN(_44997), .Q(_51422) );
  nor2s1 _52012_inst ( .DIN1(_51426), .DIN2(_50479), .Q(_51419) );
  nnd2s1 _52013_inst ( .DIN1(_51427), .DIN2(_51428), .Q(_50479) );
  nor2s1 _52014_inst ( .DIN1(_51429), .DIN2(_51430), .Q(_51428) );
  nnd2s1 _52015_inst ( .DIN1(_51242), .DIN2(_50923), .Q(_51430) );
  nnd2s1 _52016_inst ( .DIN1(_50727), .DIN2(_51003), .Q(_50923) );
  and2s1 _52017_inst ( .DIN1(_51431), .DIN2(_51432), .Q(_51003) );
  nor2s1 _52018_inst ( .DIN1(_44995), .DIN2(_50740), .Q(_51431) );
  nnd2s1 _52019_inst ( .DIN1(_51433), .DIN2(_51364), .Q(_51242) );
  nor2s1 _52020_inst ( .DIN1(_50742), .DIN2(_51434), .Q(_51433) );
  nor2s1 _52021_inst ( .DIN1(_51435), .DIN2(_50562), .Q(_51429) );
  nor2s1 _52022_inst ( .DIN1(_51012), .DIN2(_50796), .Q(_51435) );
  nor2s1 _52023_inst ( .DIN1(_51436), .DIN2(_51437), .Q(_51012) );
  or2s1 _52024_inst ( .DIN1(_42877), .DIN2(_51269), .Q(_51436) );
  nor2s1 _52025_inst ( .DIN1(_50773), .DIN2(_51314), .Q(_51427) );
  nnd2s1 _52026_inst ( .DIN1(_51438), .DIN2(_51439), .Q(_51314) );
  nnd2s1 _52027_inst ( .DIN1(_50843), .DIN2(_51004), .Q(_51439) );
  nor2s1 _52028_inst ( .DIN1(_51265), .DIN2(_42877), .Q(_50843) );
  nnd2s1 _52029_inst ( .DIN1(_51272), .DIN2(_51440), .Q(_51265) );
  or2s1 _52030_inst ( .DIN1(_50993), .DIN2(_51094), .Q(_51438) );
  nnd2s1 _52031_inst ( .DIN1(_51441), .DIN2(_51432), .Q(_51094) );
  nor2s1 _52032_inst ( .DIN1(_51412), .DIN2(_51442), .Q(_51432) );
  nnd2s1 _52033_inst ( .DIN1(_51222), .DIN2(_26415), .Q(_51442) );
  nor2s1 _52034_inst ( .DIN1(_44995), .DIN2(_51443), .Q(_51441) );
  nnd2s1 _52035_inst ( .DIN1(_51444), .DIN2(_51445), .Q(_50773) );
  nnd2s1 _52036_inst ( .DIN1(_51446), .DIN2(_51281), .Q(_51445) );
  nnd2s1 _52037_inst ( .DIN1(_50563), .DIN2(_50842), .Q(_51446) );
  nnd2s1 _52038_inst ( .DIN1(_51425), .DIN2(_44628), .Q(_50842) );
  nor2s1 _52039_inst ( .DIN1(_51447), .DIN2(_51211), .Q(_51425) );
  hi1s1 _52040_inst ( .DIN(_51440), .Q(_51211) );
  nor2s1 _52041_inst ( .DIN1(_51057), .DIN2(_51448), .Q(_51440) );
  nnd2s1 _52042_inst ( .DIN1(_51449), .DIN2(_51450), .Q(_50563) );
  nor2s1 _52043_inst ( .DIN1(_51443), .DIN2(_44998), .Q(_51449) );
  or2s1 _52044_inst ( .DIN1(_50963), .DIN2(_50707), .Q(_51444) );
  nnd2s1 _52045_inst ( .DIN1(_51451), .DIN2(_51452), .Q(_50963) );
  nor2s1 _52046_inst ( .DIN1(_51210), .DIN2(_42877), .Q(_51452) );
  nor2s1 _52047_inst ( .DIN1(_51035), .DIN2(_50988), .Q(_51451) );
  nor2s1 _52048_inst ( .DIN1(_50993), .DIN2(_50688), .Q(_51426) );
  nnd2s1 _52049_inst ( .DIN1(_51453), .DIN2(_51454), .Q(_51417) );
  nor2s1 _52050_inst ( .DIN1(_51052), .DIN2(_50713), .Q(_51454) );
  and2s1 _52051_inst ( .DIN1(_50959), .DIN2(_50920), .Q(_50713) );
  and2s1 _52052_inst ( .DIN1(_51293), .DIN2(_51455), .Q(_50959) );
  nor2s1 _52053_inst ( .DIN1(_51035), .DIN2(_42875), .Q(_51455) );
  and2s1 _52054_inst ( .DIN1(_51456), .DIN2(_51457), .Q(_51052) );
  nor2s1 _52055_inst ( .DIN1(_50605), .DIN2(_44994), .Q(_51457) );
  nor2s1 _52056_inst ( .DIN1(_50739), .DIN2(_51166), .Q(_51456) );
  nor2s1 _52057_inst ( .DIN1(_51106), .DIN2(_51458), .Q(_51453) );
  nor2s1 _52058_inst ( .DIN1(_51459), .DIN2(_50874), .Q(_51458) );
  nor2s1 _52059_inst ( .DIN1(_51460), .DIN2(_51461), .Q(_51459) );
  nor2s1 _52060_inst ( .DIN1(_50671), .DIN2(_50605), .Q(_51106) );
  nnd2s1 _52061_inst ( .DIN1(_51462), .DIN2(_51463), .Q(_50671) );
  nor2s1 _52062_inst ( .DIN1(_51210), .DIN2(_42876), .Q(_51463) );
  nor2s1 _52063_inst ( .DIN1(_51396), .DIN2(_51247), .Q(_51462) );
  nor2s1 _52064_inst ( .DIN1(_51464), .DIN2(_51465), .Q(_51415) );
  nnd2s1 _52065_inst ( .DIN1(_51466), .DIN2(_51467), .Q(_51465) );
  nor2s1 _52066_inst ( .DIN1(_51468), .DIN2(_50905), .Q(_51467) );
  nnd2s1 _52067_inst ( .DIN1(_51469), .DIN2(_51470), .Q(_50905) );
  nor2s1 _52068_inst ( .DIN1(_50735), .DIN2(_51471), .Q(_51470) );
  or2s1 _52069_inst ( .DIN1(_50669), .DIN2(_50566), .Q(_51471) );
  nor2s1 _52070_inst ( .DIN1(_50512), .DIN2(_50605), .Q(_50566) );
  nnd2s1 _52071_inst ( .DIN1(_51293), .DIN2(_51472), .Q(_50512) );
  nor2s1 _52072_inst ( .DIN1(_50988), .DIN2(_51473), .Q(_51293) );
  nor2s1 _52073_inst ( .DIN1(_50936), .DIN2(_50665), .Q(_50669) );
  and2s1 _52074_inst ( .DIN1(_50752), .DIN2(_50940), .Q(_50735) );
  and2s1 _52075_inst ( .DIN1(_51474), .DIN2(_51475), .Q(_50940) );
  nor2s1 _52076_inst ( .DIN1(_51448), .DIN2(_51443), .Q(_51475) );
  hi1s1 _52077_inst ( .DIN(_51330), .Q(_51443) );
  nor2s1 _52078_inst ( .DIN1(_51476), .DIN2(_2025), .Q(_51330) );
  nor2s1 _52079_inst ( .DIN1(_51228), .DIN2(_40395), .Q(_51474) );
  nnd2s1 _52080_inst ( .DIN1(_51477), .DIN2(_45588), .Q(_40395) );
  nor2s1 _52081_inst ( .DIN1(_51318), .DIN2(_51095), .Q(_51469) );
  nor2s1 _52082_inst ( .DIN1(_50498), .DIN2(_49457), .Q(_51095) );
  nor2s1 _52083_inst ( .DIN1(_50661), .DIN2(_51016), .Q(_51318) );
  nnd2s1 _52084_inst ( .DIN1(_51478), .DIN2(_51450), .Q(_51016) );
  nor2s1 _52085_inst ( .DIN1(_50742), .DIN2(_51479), .Q(_51478) );
  hi1s1 _52086_inst ( .DIN(_50971), .Q(_51468) );
  nor2s1 _52087_inst ( .DIN1(_51276), .DIN2(_51480), .Q(_50971) );
  nor2s1 _52088_inst ( .DIN1(_50869), .DIN2(_50629), .Q(_51480) );
  nnd2s1 _52089_inst ( .DIN1(_51481), .DIN2(_51329), .Q(_50869) );
  and2s1 _52090_inst ( .DIN1(_51482), .DIN2(_51483), .Q(_51329) );
  nor2s1 _52091_inst ( .DIN1(_51153), .DIN2(_44998), .Q(_51482) );
  nor2s1 _52092_inst ( .DIN1(_26413), .DIN2(_51484), .Q(_51481) );
  nor2s1 _52093_inst ( .DIN1(_51485), .DIN2(_51486), .Q(_51276) );
  nnd2s1 _52094_inst ( .DIN1(_44628), .DIN2(_50763), .Q(_51485) );
  nor2s1 _52095_inst ( .DIN1(_51044), .DIN2(_51181), .Q(_51466) );
  nnd2s1 _52096_inst ( .DIN1(_51487), .DIN2(_51109), .Q(_51181) );
  and2s1 _52097_inst ( .DIN1(_51488), .DIN2(_51489), .Q(_51109) );
  nnd2s1 _52098_inst ( .DIN1(_51490), .DIN2(_51491), .Q(_51489) );
  nor2s1 _52099_inst ( .DIN1(_51057), .DIN2(_50993), .Q(_51491) );
  nor2s1 _52100_inst ( .DIN1(_51056), .DIN2(_44572), .Q(_51490) );
  nnd2s1 _52101_inst ( .DIN1(_44030), .DIN2(_51295), .Q(_44572) );
  hi1s1 _52102_inst ( .DIN(_51450), .Q(_51056) );
  nor2s1 _52103_inst ( .DIN1(_51492), .DIN2(_51493), .Q(_51488) );
  nor2s1 _52104_inst ( .DIN1(_51494), .DIN2(_51495), .Q(_51493) );
  or2s1 _52105_inst ( .DIN1(_50739), .DIN2(_51083), .Q(_51495) );
  nnd2s1 _52106_inst ( .DIN1(_51496), .DIN2(_51364), .Q(_51494) );
  nor2s1 _52107_inst ( .DIN1(_44620), .DIN2(_50494), .Q(_51496) );
  nor2s1 _52108_inst ( .DIN1(_51497), .DIN2(_51498), .Q(_51492) );
  nnd2s1 _52109_inst ( .DIN1(_51499), .DIN2(_50985), .Q(_51498) );
  hi1s1 _52110_inst ( .DIN(_45002), .Q(_50985) );
  nnd2s1 _52111_inst ( .DIN1(_45585), .DIN2(_51296), .Q(_45002) );
  nor2s1 _52112_inst ( .DIN1(_51412), .DIN2(_50562), .Q(_51499) );
  nnd2s1 _52113_inst ( .DIN1(_51500), .DIN2(_51222), .Q(_51497) );
  nor2s1 _52114_inst ( .DIN1(_51501), .DIN2(_26415), .Q(_51500) );
  nor2s1 _52115_inst ( .DIN1(_50734), .DIN2(_51502), .Q(_51487) );
  nor2s1 _52116_inst ( .DIN1(_50590), .DIN2(_50630), .Q(_51502) );
  hi1s1 _52117_inst ( .DIN(_51068), .Q(_50734) );
  nnd2s1 _52118_inst ( .DIN1(_50777), .DIN2(_50824), .Q(_51068) );
  nnd2s1 _52119_inst ( .DIN1(_51212), .DIN2(_51503), .Q(_51044) );
  or2s1 _52120_inst ( .DIN1(_50730), .DIN2(_50670), .Q(_51503) );
  nnd2s1 _52121_inst ( .DIN1(_51504), .DIN2(_51505), .Q(_50730) );
  nor2s1 _52122_inst ( .DIN1(_51501), .DIN2(_42877), .Q(_51504) );
  nnd2s1 _52123_inst ( .DIN1(_51506), .DIN2(_51507), .Q(_51212) );
  and2s1 _52124_inst ( .DIN1(_51508), .DIN2(_50727), .Q(_51507) );
  nor2s1 _52125_inst ( .DIN1(_40394), .DIN2(_51394), .Q(_51506) );
  nnd2s1 _52126_inst ( .DIN1(_51509), .DIN2(_51226), .Q(_51394) );
  nor2s1 _52127_inst ( .DIN1(_51510), .DIN2(_51210), .Q(_51509) );
  nnd2s1 _52128_inst ( .DIN1(_51511), .DIN2(_51512), .Q(_51464) );
  nor2s1 _52129_inst ( .DIN1(_51231), .DIN2(_50520), .Q(_51512) );
  nnd2s1 _52130_inst ( .DIN1(_51513), .DIN2(_51514), .Q(_50520) );
  hi1s1 _52131_inst ( .DIN(_50577), .Q(_51514) );
  nnd2s1 _52132_inst ( .DIN1(_51515), .DIN2(_51516), .Q(_50577) );
  nnd2s1 _52133_inst ( .DIN1(_50751), .DIN2(_50823), .Q(_51516) );
  hi1s1 _52134_inst ( .DIN(_50993), .Q(_50823) );
  hi1s1 _52135_inst ( .DIN(_51283), .Q(_50751) );
  nnd2s1 _52136_inst ( .DIN1(_51517), .DIN2(_51518), .Q(_51283) );
  nor2s1 _52137_inst ( .DIN1(_51151), .DIN2(_51476), .Q(_51518) );
  nor2s1 _52138_inst ( .DIN1(_51353), .DIN2(_44573), .Q(_51517) );
  nnd2s1 _52139_inst ( .DIN1(_50753), .DIN2(_50960), .Q(_51515) );
  hi1s1 _52140_inst ( .DIN(_51282), .Q(_50753) );
  nnd2s1 _52141_inst ( .DIN1(_51519), .DIN2(_51520), .Q(_51282) );
  nor2s1 _52142_inst ( .DIN1(_51448), .DIN2(_51476), .Q(_51520) );
  nor2s1 _52143_inst ( .DIN1(_42876), .DIN2(_51353), .Q(_51519) );
  nor2s1 _52144_inst ( .DIN1(_50943), .DIN2(_51521), .Q(_51513) );
  nor2s1 _52145_inst ( .DIN1(_50830), .DIN2(_50501), .Q(_51521) );
  nor2s1 _52146_inst ( .DIN1(_50659), .DIN2(_50494), .Q(_50943) );
  or2s1 _52147_inst ( .DIN1(_50568), .DIN2(_51522), .Q(_51231) );
  nor2s1 _52148_inst ( .DIN1(_50692), .DIN2(_50687), .Q(_51522) );
  nor2s1 _52149_inst ( .DIN1(_50704), .DIN2(_50874), .Q(_50568) );
  nnd2s1 _52150_inst ( .DIN1(_51523), .DIN2(_44578), .Q(_50704) );
  hi1s1 _52151_inst ( .DIN(_40394), .Q(_44578) );
  nnd2s1 _52152_inst ( .DIN1(_51361), .DIN2(_51524), .Q(_40394) );
  nor2s1 _52153_inst ( .DIN1(_51437), .DIN2(_51247), .Q(_51523) );
  nor2s1 _52154_inst ( .DIN1(_50543), .DIN2(_50644), .Q(_51511) );
  nnd2s1 _52155_inst ( .DIN1(_51525), .DIN2(_51526), .Q(_50644) );
  nor2s1 _52156_inst ( .DIN1(_51527), .DIN2(_51528), .Q(_51526) );
  nnd2s1 _52157_inst ( .DIN1(_50765), .DIN2(_51370), .Q(_51528) );
  nnd2s1 _52158_inst ( .DIN1(_50796), .DIN2(_51093), .Q(_51370) );
  hi1s1 _52159_inst ( .DIN(_50670), .Q(_51093) );
  and2s1 _52160_inst ( .DIN1(_51423), .DIN2(_44628), .Q(_50796) );
  and2s1 _52161_inst ( .DIN1(_51529), .DIN2(_51364), .Q(_51423) );
  hi1s1 _52162_inst ( .DIN(_51153), .Q(_51364) );
  nor2s1 _52163_inst ( .DIN1(_51448), .DIN2(_51035), .Q(_51529) );
  nnd2s1 _52164_inst ( .DIN1(_51530), .DIN2(_51531), .Q(_50765) );
  nor2s1 _52165_inst ( .DIN1(_51057), .DIN2(_51084), .Q(_51531) );
  nnd2s1 _52166_inst ( .DIN1(_50727), .DIN2(_51272), .Q(_51084) );
  nor2s1 _52167_inst ( .DIN1(_50739), .DIN2(_44577), .Q(_51530) );
  nnd2s1 _52168_inst ( .DIN1(_45584), .DIN2(_45588), .Q(_44577) );
  nnd2s1 _52169_inst ( .DIN1(_51532), .DIN2(_51533), .Q(_51527) );
  nor2s1 _52170_inst ( .DIN1(_51402), .DIN2(_50782), .Q(_51532) );
  nor2s1 _52171_inst ( .DIN1(_50691), .DIN2(_50498), .Q(_50782) );
  hi1s1 _52172_inst ( .DIN(_51534), .Q(_50691) );
  and2s1 _52173_inst ( .DIN1(_51535), .DIN2(_51536), .Q(_51402) );
  nor2s1 _52174_inst ( .DIN1(_51151), .DIN2(_42877), .Q(_51536) );
  nor2s1 _52175_inst ( .DIN1(_50687), .DIN2(_51166), .Q(_51535) );
  nnd2s1 _52176_inst ( .DIN1(_51537), .DIN2(_51538), .Q(_51166) );
  hi1s1 _52177_inst ( .DIN(_51353), .Q(_51538) );
  nnd2s1 _52178_inst ( .DIN1(_51539), .DIN2(_2025), .Q(_51353) );
  nor2s1 _52179_inst ( .DIN1(_51540), .DIN2(_51541), .Q(_51525) );
  nnd2s1 _52180_inst ( .DIN1(_50747), .DIN2(_50477), .Q(_51541) );
  and2s1 _52181_inst ( .DIN1(_51542), .DIN2(_51543), .Q(_50477) );
  nnd2s1 _52182_inst ( .DIN1(_51299), .DIN2(_51281), .Q(_51543) );
  hi1s1 _52183_inst ( .DIN(_50829), .Q(_51299) );
  nor2s1 _52184_inst ( .DIN1(_50921), .DIN2(_51544), .Q(_51542) );
  nor2s1 _52185_inst ( .DIN1(_50660), .DIN2(_50498), .Q(_51544) );
  nnd2s1 _52186_inst ( .DIN1(_51545), .DIN2(_51546), .Q(_50660) );
  nor2s1 _52187_inst ( .DIN1(_51152), .DIN2(_45001), .Q(_51546) );
  nnd2s1 _52188_inst ( .DIN1(_51360), .DIN2(_45588), .Q(_45001) );
  nor2s1 _52189_inst ( .DIN1(_51547), .DIN2(_51548), .Q(_51545) );
  and2s1 _52190_inst ( .DIN1(_51110), .DIN2(_51549), .Q(_50747) );
  hi1s1 _52191_inst ( .DIN(_51399), .Q(_51110) );
  nnd2s1 _52192_inst ( .DIN1(_51550), .DIN2(_51551), .Q(_51399) );
  nnd2s1 _52193_inst ( .DIN1(_51552), .DIN2(_44627), .Q(_51551) );
  hi1s1 _52194_inst ( .DIN(_44999), .Q(_44627) );
  nnd2s1 _52195_inst ( .DIN1(_45585), .DIN2(_51477), .Q(_44999) );
  nor2s1 _52196_inst ( .DIN1(_51210), .DIN2(_51434), .Q(_51552) );
  nor2s1 _52197_inst ( .DIN1(_51553), .DIN2(_51554), .Q(_51550) );
  nor2s1 _52198_inst ( .DIN1(_51555), .DIN2(_51556), .Q(_51554) );
  nnd2s1 _52199_inst ( .DIN1(_50960), .DIN2(_51341), .Q(_51556) );
  nnd2s1 _52200_inst ( .DIN1(_51557), .DIN2(_51271), .Q(_51555) );
  hi1s1 _52201_inst ( .DIN(_50988), .Q(_51271) );
  nnd2s1 _52202_inst ( .DIN1(_51558), .DIN2(_51559), .Q(_50988) );
  nor2s1 _52203_inst ( .DIN1(_51152), .DIN2(_42877), .Q(_51557) );
  nnd2s1 _52204_inst ( .DIN1(_51360), .DIN2(_51295), .Q(_42877) );
  hi1s1 _52205_inst ( .DIN(_51560), .Q(_51360) );
  nor2s1 _52206_inst ( .DIN1(_51561), .DIN2(_51562), .Q(_51553) );
  nnd2s1 _52207_inst ( .DIN1(_50777), .DIN2(_44625), .Q(_51562) );
  hi1s1 _52208_inst ( .DIN(_44994), .Q(_44625) );
  nnd2s1 _52209_inst ( .DIN1(_51563), .DIN2(_51359), .Q(_51561) );
  nnd2s1 _52210_inst ( .DIN1(_51564), .DIN2(_51063), .Q(_51540) );
  nnd2s1 _52211_inst ( .DIN1(_51241), .DIN2(_50537), .Q(_51063) );
  hi1s1 _52212_inst ( .DIN(_50501), .Q(_50537) );
  nor2s1 _52213_inst ( .DIN1(_51132), .DIN2(_50799), .Q(_51564) );
  nor2s1 _52214_inst ( .DIN1(_50590), .DIN2(_50910), .Q(_50799) );
  nor2s1 _52215_inst ( .DIN1(_50498), .DIN2(_51119), .Q(_51132) );
  nnd2s1 _52216_inst ( .DIN1(_51565), .DIN2(_51566), .Q(_50543) );
  nor2s1 _52217_inst ( .DIN1(_51567), .DIN2(_51568), .Q(_51566) );
  nnd2s1 _52218_inst ( .DIN1(_51569), .DIN2(_50808), .Q(_51568) );
  nnd2s1 _52219_inst ( .DIN1(_50752), .DIN2(_50994), .Q(_50808) );
  nor2s1 _52220_inst ( .DIN1(_51221), .DIN2(_51386), .Q(_50994) );
  nnd2s1 _52221_inst ( .DIN1(_51570), .DIN2(_51571), .Q(_51221) );
  nor2s1 _52222_inst ( .DIN1(_44994), .DIN2(_51247), .Q(_51570) );
  nnd2s1 _52223_inst ( .DIN1(_45585), .DIN2(_51572), .Q(_44994) );
  hi1s1 _52224_inst ( .DIN(_50560), .Q(_50752) );
  or2s1 _52225_inst ( .DIN1(_50561), .DIN2(_50786), .Q(_51569) );
  hi1s1 _52226_inst ( .DIN(_50941), .Q(_50786) );
  nnd2s1 _52227_inst ( .DIN1(_50993), .DIN2(_50560), .Q(_50941) );
  nnd2s1 _52228_inst ( .DIN1(_51281), .DIN2(_51573), .Q(_50993) );
  nnd2s1 _52229_inst ( .DIN1(_51574), .DIN2(______[16]), .Q(_51573) );
  nnd2s1 _52230_inst ( .DIN1(_51575), .DIN2(_51576), .Q(_50561) );
  nor2s1 _52231_inst ( .DIN1(_51057), .DIN2(_51577), .Q(_51576) );
  nnd2s1 _52232_inst ( .DIN1(_51578), .DIN2(_51222), .Q(_51577) );
  and2s1 _52233_inst ( .DIN1(_44628), .DIN2(_51579), .Q(_51575) );
  nnd2s1 _52234_inst ( .DIN1(_51580), .DIN2(_51581), .Q(_51567) );
  nnd2s1 _52235_inst ( .DIN1(_51229), .DIN2(_50960), .Q(_51581) );
  hi1s1 _52236_inst ( .DIN(_50687), .Q(_50960) );
  hi1s1 _52237_inst ( .DIN(_50887), .Q(_51229) );
  nnd2s1 _52238_inst ( .DIN1(_51582), .DIN2(_51583), .Q(_50887) );
  nor2s1 _52239_inst ( .DIN1(_51386), .DIN2(_51035), .Q(_51583) );
  nnd2s1 _52240_inst ( .DIN1(_51558), .DIN2(_51223), .Q(_51386) );
  nor2s1 _52241_inst ( .DIN1(_2030), .DIN2(_26321), .Q(_51558) );
  nor2s1 _52242_inst ( .DIN1(_51473), .DIN2(_44576), .Q(_51582) );
  nnd2s1 _52243_inst ( .DIN1(_51572), .DIN2(_51295), .Q(_44576) );
  nor2s1 _52244_inst ( .DIN1(_50507), .DIN2(_51123), .Q(_51580) );
  nor2s1 _52245_inst ( .DIN1(_50811), .DIN2(_50670), .Q(_51123) );
  nnd2s1 _52246_inst ( .DIN1(_51281), .DIN2(_51584), .Q(_50670) );
  nnd2s1 _52247_inst ( .DIN1(_51574), .DIN2(_26772), .Q(_51584) );
  nnd2s1 _52248_inst ( .DIN1(_51585), .DIN2(_51586), .Q(_50811) );
  nor2s1 _52249_inst ( .DIN1(_51393), .DIN2(_26415), .Q(_51586) );
  nor2s1 _52250_inst ( .DIN1(_51412), .DIN2(_51352), .Q(_51585) );
  nnd2s1 _52251_inst ( .DIN1(_51587), .DIN2(_51588), .Q(_51352) );
  hi1s1 _52252_inst ( .DIN(_42876), .Q(_51588) );
  nor2s1 _52253_inst ( .DIN1(_26321), .DIN2(_50980), .Q(_51587) );
  nor2s1 _52254_inst ( .DIN1(_50854), .DIN2(_50874), .Q(_50507) );
  nnd2s1 _52255_inst ( .DIN1(_51340), .DIN2(_51571), .Q(_50854) );
  and2s1 _52256_inst ( .DIN1(_51589), .DIN2(_51590), .Q(_51340) );
  nor2s1 _52257_inst ( .DIN1(_50742), .DIN2(_51510), .Q(_51590) );
  nor2s1 _52258_inst ( .DIN1(_51176), .DIN2(_51448), .Q(_51589) );
  nnd2s1 _52259_inst ( .DIN1(_1986), .DIN2(_51591), .Q(_51448) );
  nor2s1 _52260_inst ( .DIN1(_51592), .DIN2(_51593), .Q(_51565) );
  nnd2s1 _52261_inst ( .DIN1(_51594), .DIN2(_50991), .Q(_51593) );
  and2s1 _52262_inst ( .DIN1(_51070), .DIN2(_51595), .Q(_50991) );
  nnd2s1 _52263_inst ( .DIN1(_51179), .DIN2(_51281), .Q(_51595) );
  hi1s1 _52264_inst ( .DIN(_50606), .Q(_51179) );
  nnd2s1 _52265_inst ( .DIN1(_51596), .DIN2(_51597), .Q(_50606) );
  nor2s1 _52266_inst ( .DIN1(_50743), .DIN2(_51598), .Q(_51597) );
  or2s1 _52267_inst ( .DIN1(_51151), .DIN2(_2022), .Q(_51598) );
  nor2s1 _52268_inst ( .DIN1(_51176), .DIN2(_44998), .Q(_51596) );
  nnd2s1 _52269_inst ( .DIN1(_45584), .DIN2(_51361), .Q(_44998) );
  nnd2s1 _52270_inst ( .DIN1(_51335), .DIN2(_50836), .Q(_51070) );
  hi1s1 _52271_inst ( .DIN(_50590), .Q(_50836) );
  and2s1 _52272_inst ( .DIN1(_51472), .DIN2(_51450), .Q(_51335) );
  nor2s1 _52273_inst ( .DIN1(_51412), .DIN2(_51599), .Q(_51450) );
  nnd2s1 _52274_inst ( .DIN1(_51578), .DIN2(_26326), .Q(_51412) );
  nor2s1 _52275_inst ( .DIN1(_50742), .DIN2(_51152), .Q(_51472) );
  hi1s1 _52276_inst ( .DIN(_50578), .Q(_51594) );
  nnd2s1 _52277_inst ( .DIN1(_51600), .DIN2(_51601), .Q(_50578) );
  or2s1 _52278_inst ( .DIN1(_50638), .DIN2(_50637), .Q(_51601) );
  hi1s1 _52279_inst ( .DIN(_51004), .Q(_50637) );
  nnd2s1 _52280_inst ( .DIN1(_51602), .DIN2(_51563), .Q(_50638) );
  nor2s1 _52281_inst ( .DIN1(_51501), .DIN2(_44997), .Q(_51602) );
  nnd2s1 _52282_inst ( .DIN1(_51603), .DIN2(_51361), .Q(_44997) );
  nnd2s1 _52283_inst ( .DIN1(_51148), .DIN2(_50797), .Q(_51600) );
  hi1s1 _52284_inst ( .DIN(_50612), .Q(_51148) );
  nnd2s1 _52285_inst ( .DIN1(_51604), .DIN2(_51605), .Q(_50612) );
  nor2s1 _52286_inst ( .DIN1(_51510), .DIN2(_51606), .Q(_51605) );
  nnd2s1 _52287_inst ( .DIN1(_51508), .DIN2(_26326), .Q(_51606) );
  nor2s1 _52288_inst ( .DIN1(_44995), .DIN2(_51178), .Q(_51604) );
  nnd2s1 _52289_inst ( .DIN1(_51607), .DIN2(_51591), .Q(_51178) );
  nnd2s1 _52290_inst ( .DIN1(_51361), .DIN2(_51477), .Q(_44995) );
  nnd2s1 _52291_inst ( .DIN1(_51608), .DIN2(_51323), .Q(_51592) );
  nor2s1 _52292_inst ( .DIN1(_50967), .DIN2(_51609), .Q(_51323) );
  and2s1 _52293_inst ( .DIN1(_50946), .DIN2(_50797), .Q(_51609) );
  and2s1 _52294_inst ( .DIN1(_51610), .DIN2(_51505), .Q(_50946) );
  hi1s1 _52295_inst ( .DIN(_51348), .Q(_51505) );
  nnd2s1 _52296_inst ( .DIN1(_51571), .DIN2(_51226), .Q(_51348) );
  hi1s1 _52297_inst ( .DIN(_50739), .Q(_51226) );
  hi1s1 _52298_inst ( .DIN(_51473), .Q(_51571) );
  nnd2s1 _52299_inst ( .DIN1(_51611), .DIN2(_2026), .Q(_51473) );
  nor2s1 _52300_inst ( .DIN1(_26277), .DIN2(_26641), .Q(_51611) );
  nor2s1 _52301_inst ( .DIN1(_51152), .DIN2(_42875), .Q(_51610) );
  nnd2s1 _52302_inst ( .DIN1(_2022), .DIN2(_51612), .Q(_51152) );
  nor2s1 _52303_inst ( .DIN1(_51613), .DIN2(_51434), .Q(_50967) );
  nnd2s1 _52304_inst ( .DIN1(_51363), .DIN2(_50797), .Q(_51434) );
  hi1s1 _52305_inst ( .DIN(_50562), .Q(_50797) );
  nnd2s1 _52306_inst ( .DIN1(_51614), .DIN2(_51574), .Q(_50562) );
  nor2s1 _52307_inst ( .DIN1(_51151), .DIN2(_51035), .Q(_51363) );
  nnd2s1 _52308_inst ( .DIN1(_51615), .DIN2(_51393), .Q(_51035) );
  or2s1 _52309_inst ( .DIN1(_44620), .DIN2(_51210), .Q(_51613) );
  nor2s1 _52310_inst ( .DIN1(_50462), .DIN2(_51202), .Q(_51608) );
  nnd2s1 _52311_inst ( .DIN1(_51616), .DIN2(_51617), .Q(_51202) );
  nnd2s1 _52312_inst ( .DIN1(_50727), .DIN2(_51618), .Q(_51617) );
  nnd2s1 _52313_inst ( .DIN1(_51168), .DIN2(_51619), .Q(_51618) );
  nnd2s1 _52314_inst ( .DIN1(_51620), .DIN2(_51621), .Q(_51619) );
  nor2s1 _52315_inst ( .DIN1(_51393), .DIN2(_51476), .Q(_51621) );
  nor2s1 _52316_inst ( .DIN1(_51437), .DIN2(_44573), .Q(_51620) );
  nnd2s1 _52317_inst ( .DIN1(_51295), .DIN2(_51524), .Q(_44573) );
  nnd2s1 _52318_inst ( .DIN1(_51622), .DIN2(_51579), .Q(_51437) );
  nor2s1 _52319_inst ( .DIN1(_51548), .DIN2(_51153), .Q(_51622) );
  nnd2s1 _52320_inst ( .DIN1(_51623), .DIN2(_51624), .Q(_51168) );
  nor2s1 _52321_inst ( .DIN1(_51210), .DIN2(_51379), .Q(_51624) );
  nnd2s1 _52322_inst ( .DIN1(_45585), .DIN2(_44030), .Q(_51379) );
  nor2s1 _52323_inst ( .DIN1(_51057), .DIN2(_51396), .Q(_51623) );
  hi1s1 _52324_inst ( .DIN(_50494), .Q(_50727) );
  nor2s1 _52325_inst ( .DIN1(_51625), .DIN2(_51626), .Q(_51616) );
  nor2s1 _52326_inst ( .DIN1(_51486), .DIN2(_51627), .Q(_51626) );
  nnd2s1 _52327_inst ( .DIN1(_50913), .DIN2(_44628), .Q(_51627) );
  hi1s1 _52328_inst ( .DIN(_42875), .Q(_44628) );
  nnd2s1 _52329_inst ( .DIN1(_45584), .DIN2(_51295), .Q(_42875) );
  and2s1 _52330_inst ( .DIN1(_51628), .DIN2(_2057), .Q(_45584) );
  nor2s1 _52331_inst ( .DIN1(_26280), .DIN2(_26647), .Q(_51628) );
  nnd2s1 _52332_inst ( .DIN1(_51629), .DIN2(_51483), .Q(_51486) );
  hi1s1 _52333_inst ( .DIN(_51396), .Q(_51483) );
  nnd2s1 _52334_inst ( .DIN1(_51630), .DIN2(_51222), .Q(_51396) );
  nor2s1 _52335_inst ( .DIN1(_2006), .DIN2(_1986), .Q(_51630) );
  nor2s1 _52336_inst ( .DIN1(_50740), .DIN2(_51228), .Q(_51629) );
  nnd2s1 _52337_inst ( .DIN1(_51631), .DIN2(_2027), .Q(_50740) );
  nor2s1 _52338_inst ( .DIN1(_51632), .DIN2(_51633), .Q(_51625) );
  or2s1 _52339_inst ( .DIN1(_51036), .DIN2(_50560), .Q(_51633) );
  nnd2s1 _52340_inst ( .DIN1(_51574), .DIN2(_51634), .Q(_50560) );
  nor2s1 _52341_inst ( .DIN1(______[20]), .DIN2(______[25]), .Q(_51574) );
  nnd2s1 _52342_inst ( .DIN1(_51635), .DIN2(_51222), .Q(_51036) );
  nor2s1 _52343_inst ( .DIN1(_44620), .DIN2(_51210), .Q(_51635) );
  nnd2s1 _52344_inst ( .DIN1(_51603), .DIN2(_51295), .Q(_44620) );
  hi1s1 _52345_inst ( .DIN(_51636), .Q(_51603) );
  nnd2s1 _52346_inst ( .DIN1(_51579), .DIN2(_51637), .Q(_51632) );
  nor2s1 _52347_inst ( .DIN1(_50995), .DIN2(_50495), .Q(_50462) );
  nnd2s1 _52348_inst ( .DIN1(_51638), .DIN2(_51639), .Q(____1___________0[0])
         );
  nor2s1 _52349_inst ( .DIN1(_51640), .DIN2(_51641), .Q(_51639) );
  nnd2s1 _52350_inst ( .DIN1(_51642), .DIN2(_51404), .Q(_51641) );
  and2s1 _52351_inst ( .DIN1(_51643), .DIN2(_51644), .Q(_51404) );
  nnd2s1 _52352_inst ( .DIN1(_50824), .DIN2(_51316), .Q(_51644) );
  nor2s1 _52353_inst ( .DIN1(_51645), .DIN2(_51646), .Q(_50824) );
  nnd2s1 _52354_inst ( .DIN1(_50589), .DIN2(_51004), .Q(_51643) );
  nnd2s1 _52355_inst ( .DIN1(_50995), .DIN2(_50494), .Q(_51004) );
  nnd2s1 _52356_inst ( .DIN1(_51647), .DIN2(_51634), .Q(_50494) );
  nnd2s1 _52357_inst ( .DIN1(_51281), .DIN2(_51648), .Q(_50995) );
  nnd2s1 _52358_inst ( .DIN1(_51647), .DIN2(______[16]), .Q(_51648) );
  hi1s1 _52359_inst ( .DIN(_50659), .Q(_50589) );
  nnd2s1 _52360_inst ( .DIN1(_51649), .DIN2(_51650), .Q(_50659) );
  nor2s1 _52361_inst ( .DIN1(_26327), .DIN2(_51479), .Q(_51650) );
  nor2s1 _52362_inst ( .DIN1(_51651), .DIN2(_51652), .Q(_51649) );
  hi1s1 _52363_inst ( .DIN(_51121), .Q(_51642) );
  nnd2s1 _52364_inst ( .DIN1(_51653), .DIN2(_51654), .Q(_51121) );
  nnd2s1 _52365_inst ( .DIN1(_51655), .DIN2(_50920), .Q(_51654) );
  nnd2s1 _52366_inst ( .DIN1(_50511), .DIN2(_50687), .Q(_50920) );
  nnd2s1 _52367_inst ( .DIN1(_51614), .DIN2(_51647), .Q(_50687) );
  nnd2s1 _52368_inst ( .DIN1(_51281), .DIN2(_51656), .Q(_50511) );
  nnd2s1 _52369_inst ( .DIN1(_51647), .DIN2(_26772), .Q(_51656) );
  nor2s1 _52370_inst ( .DIN1(_51657), .DIN2(______[20]), .Q(_51647) );
  hi1s1 _52371_inst ( .DIN(_50692), .Q(_51655) );
  nnd2s1 _52372_inst ( .DIN1(_51658), .DIN2(_50987), .Q(_50692) );
  nor2s1 _52373_inst ( .DIN1(_51659), .DIN2(_51660), .Q(_51658) );
  nor2s1 _52374_inst ( .DIN1(_51167), .DIN2(_51661), .Q(_51653) );
  nor2s1 _52375_inst ( .DIN1(_50605), .DIN2(_50513), .Q(_51661) );
  nnd2s1 _52376_inst ( .DIN1(_51662), .DIN2(_51663), .Q(_50513) );
  nor2s1 _52377_inst ( .DIN1(_51636), .DIN2(_51664), .Q(_51663) );
  nnd2s1 _52378_inst ( .DIN1(_51510), .DIN2(_26254), .Q(_51664) );
  nor2s1 _52379_inst ( .DIN1(_51665), .DIN2(_51547), .Q(_51662) );
  hi1s1 _52380_inst ( .DIN(_51533), .Q(_51167) );
  nnd2s1 _52381_inst ( .DIN1(_50915), .DIN2(_51281), .Q(_51533) );
  hi1s1 _52382_inst ( .DIN(_50500), .Q(_50915) );
  nnd2s1 _52383_inst ( .DIN1(_51666), .DIN2(_51667), .Q(_50500) );
  nor2s1 _52384_inst ( .DIN1(_51659), .DIN2(_51510), .Q(_51667) );
  nor2s1 _52385_inst ( .DIN1(_51034), .DIN2(_51668), .Q(_51666) );
  nnd2s1 _52386_inst ( .DIN1(_51669), .DIN2(_51670), .Q(_51640) );
  nnd2s1 _52387_inst ( .DIN1(_51534), .DIN2(_51316), .Q(_51670) );
  nor2s1 _52388_inst ( .DIN1(_51671), .DIN2(_51672), .Q(_51534) );
  or2s1 _52389_inst ( .DIN1(_2063), .DIN2(_51673), .Q(_51671) );
  nor2s1 _52390_inst ( .DIN1(_51256), .DIN2(_51674), .Q(_51669) );
  nor2s1 _52391_inst ( .DIN1(_51381), .DIN2(_51675), .Q(_51674) );
  nnd2s1 _52392_inst ( .DIN1(_50913), .DIN2(_53523), .Q(_51675) );
  nnd2s1 _52393_inst ( .DIN1(_51676), .DIN2(_51677), .Q(_51381) );
  nor2s1 _52394_inst ( .DIN1(_50743), .DIN2(_51057), .Q(_51677) );
  nnd2s1 _52395_inst ( .DIN1(_51612), .DIN2(_51510), .Q(_51057) );
  and2s1 _52396_inst ( .DIN1(_51678), .DIN2(_2031), .Q(_51612) );
  nor2s1 _52397_inst ( .DIN1(_51393), .DIN2(_26413), .Q(_51678) );
  nor2s1 _52398_inst ( .DIN1(_42876), .DIN2(_50739), .Q(_51676) );
  nnd2s1 _52399_inst ( .DIN1(_51222), .DIN2(_51559), .Q(_50739) );
  hi1s1 _52400_inst ( .DIN(_51548), .Q(_51222) );
  nnd2s1 _52401_inst ( .DIN1(_2030), .DIN2(_2064), .Q(_51548) );
  nnd2s1 _52402_inst ( .DIN1(_44030), .DIN2(_51361), .Q(_42876) );
  hi1s1 _52403_inst ( .DIN(_40397), .Q(_44030) );
  nnd2s1 _52404_inst ( .DIN1(_51679), .DIN2(_2057), .Q(_40397) );
  nor2s1 _52405_inst ( .DIN1(_2062), .DIN2(_2056), .Q(_51679) );
  nor2s1 _52406_inst ( .DIN1(_50495), .DIN2(_50605), .Q(_51256) );
  nnd2s1 _52407_inst ( .DIN1(_51680), .DIN2(_51681), .Q(_50495) );
  nor2s1 _52408_inst ( .DIN1(_2022), .DIN2(_51560), .Q(_51681) );
  nor2s1 _52409_inst ( .DIN1(_50743), .DIN2(_51682), .Q(_51680) );
  nor2s1 _52410_inst ( .DIN1(_51683), .DIN2(_51684), .Q(_51638) );
  nnd2s1 _52411_inst ( .DIN1(_51074), .DIN2(_50533), .Q(_51684) );
  nor2s1 _52412_inst ( .DIN1(_50693), .DIN2(_50634), .Q(_50533) );
  nor2s1 _52413_inst ( .DIN1(_50936), .DIN2(_50703), .Q(_50634) );
  nnd2s1 _52414_inst ( .DIN1(_51685), .DIN2(_51686), .Q(_50936) );
  nor2s1 _52415_inst ( .DIN1(_51393), .DIN2(_51687), .Q(_51686) );
  nnd2s1 _52416_inst ( .DIN1(_45585), .DIN2(_51524), .Q(_51687) );
  hi1s1 _52417_inst ( .DIN(_51688), .Q(_45585) );
  nor2s1 _52418_inst ( .DIN1(_50980), .DIN2(_51652), .Q(_51685) );
  nnd2s1 _52419_inst ( .DIN1(_51689), .DIN2(_51193), .Q(_50693) );
  nnd2s1 _52420_inst ( .DIN1(_49465), .DIN2(_50777), .Q(_51193) );
  hi1s1 _52421_inst ( .DIN(_50661), .Q(_50777) );
  hi1s1 _52422_inst ( .DIN(_49457), .Q(_49465) );
  nnd2s1 _52423_inst ( .DIN1(_51305), .DIN2(_51563), .Q(_49457) );
  nor2s1 _52424_inst ( .DIN1(_51151), .DIN2(_50743), .Q(_51563) );
  nnd2s1 _52425_inst ( .DIN1(_51690), .DIN2(_2023), .Q(_50743) );
  nor2s1 _52426_inst ( .DIN1(_2026), .DIN2(_26277), .Q(_51690) );
  nnd2s1 _52427_inst ( .DIN1(_51591), .DIN2(_26326), .Q(_51151) );
  hi1s1 _52428_inst ( .DIN(_51599), .Q(_51591) );
  nnd2s1 _52429_inst ( .DIN1(_51691), .DIN2(_2064), .Q(_51599) );
  nor2s1 _52430_inst ( .DIN1(_2030), .DIN2(_2006), .Q(_51691) );
  nor2s1 _52431_inst ( .DIN1(_51501), .DIN2(_50742), .Q(_51305) );
  nnd2s1 _52432_inst ( .DIN1(_51477), .DIN2(_51295), .Q(_50742) );
  nor2s1 _52433_inst ( .DIN1(_26444), .DIN2(_26254), .Q(_51295) );
  and2s1 _52434_inst ( .DIN1(_51692), .DIN2(_2057), .Q(_51477) );
  nor2s1 _52435_inst ( .DIN1(_2062), .DIN2(_26280), .Q(_51692) );
  nnd2s1 _52436_inst ( .DIN1(_51398), .DIN2(_51316), .Q(_51689) );
  hi1s1 _52437_inst ( .DIN(_51119), .Q(_51398) );
  nnd2s1 _52438_inst ( .DIN1(_51693), .DIN2(_51694), .Q(_51119) );
  nor2s1 _52439_inst ( .DIN1(_2063), .DIN2(_51695), .Q(_51694) );
  nor2s1 _52440_inst ( .DIN1(_51696), .DIN2(_51673), .Q(_51693) );
  and2s1 _52441_inst ( .DIN1(_51697), .DIN2(_51549), .Q(_51074) );
  nnd2s1 _52442_inst ( .DIN1(_51698), .DIN2(_51102), .Q(_51549) );
  hi1s1 _52443_inst ( .DIN(_50877), .Q(_51698) );
  nnd2s1 _52444_inst ( .DIN1(_51699), .DIN2(_51359), .Q(_50877) );
  hi1s1 _52445_inst ( .DIN(_51479), .Q(_51359) );
  nnd2s1 _52446_inst ( .DIN1(_51631), .DIN2(_26413), .Q(_51479) );
  and2s1 _52447_inst ( .DIN1(_51700), .DIN2(_2022), .Q(_51631) );
  and2s1 _52448_inst ( .DIN1(_51393), .DIN2(_2031), .Q(_51700) );
  nor2s1 _52449_inst ( .DIN1(_51560), .DIN2(_51660), .Q(_51699) );
  nnd2s1 _52450_inst ( .DIN1(_51701), .DIN2(_2030), .Q(_51660) );
  nor2s1 _52451_inst ( .DIN1(_51688), .DIN2(_51646), .Q(_51701) );
  nnd2s1 _52452_inst ( .DIN1(_51702), .DIN2(_26280), .Q(_51560) );
  nor2s1 _52453_inst ( .DIN1(_50921), .DIN2(_51703), .Q(_51697) );
  nor2s1 _52454_inst ( .DIN1(_50707), .DIN2(_50830), .Q(_51703) );
  nnd2s1 _52455_inst ( .DIN1(_51704), .DIN2(_51705), .Q(_50830) );
  nor2s1 _52456_inst ( .DIN1(_51636), .DIN2(_51706), .Q(_51705) );
  nnd2s1 _52457_inst ( .DIN1(_45588), .DIN2(_26327), .Q(_51706) );
  nor2s1 _52458_inst ( .DIN1(_51646), .DIN2(_51083), .Q(_51704) );
  hi1s1 _52459_inst ( .DIN(_50587), .Q(_50707) );
  and2s1 _52460_inst ( .DIN1(_51707), .DIN2(_51708), .Q(_50921) );
  nor2s1 _52461_inst ( .DIN1(_51034), .DIN2(_51709), .Q(_51708) );
  nnd2s1 _52462_inst ( .DIN1(_51281), .DIN2(_51510), .Q(_51709) );
  nor2s1 _52463_inst ( .DIN1(_51665), .DIN2(_51710), .Q(_51707) );
  nnd2s1 _52464_inst ( .DIN1(_51711), .DIN2(_51539), .Q(_51710) );
  and2s1 _52465_inst ( .DIN1(_51712), .DIN2(_2026), .Q(_51539) );
  nor2s1 _52466_inst ( .DIN1(_2023), .DIN2(_2015), .Q(_51712) );
  hi1s1 _52467_inst ( .DIN(_51695), .Q(_51711) );
  or2s1 _52468_inst ( .DIN1(_50521), .DIN2(_51030), .Q(_51683) );
  nnd2s1 _52469_inst ( .DIN1(_50460), .DIN2(_51713), .Q(_51030) );
  or2s1 _52470_inst ( .DIN1(_50666), .DIN2(_50703), .Q(_51713) );
  nor2s1 _52471_inst ( .DIN1(_50913), .DIN2(_50763), .Q(_50703) );
  hi1s1 _52472_inst ( .DIN(_50874), .Q(_50763) );
  nnd2s1 _52473_inst ( .DIN1(_51614), .DIN2(_51714), .Q(_50874) );
  hi1s1 _52474_inst ( .DIN(_50665), .Q(_50913) );
  nnd2s1 _52475_inst ( .DIN1(_51281), .DIN2(_51715), .Q(_50665) );
  nnd2s1 _52476_inst ( .DIN1(_51714), .DIN2(_26772), .Q(_51715) );
  hi1s1 _52477_inst ( .DIN(_51460), .Q(_50666) );
  nor2s1 _52478_inst ( .DIN1(_51716), .DIN2(_51645), .Q(_51460) );
  nnd2s1 _52479_inst ( .DIN1(_51717), .DIN2(_51718), .Q(_51645) );
  nor2s1 _52480_inst ( .DIN1(_40396), .DIN2(_51659), .Q(_51717) );
  or2s1 _52481_inst ( .DIN1(_2064), .DIN2(_51547), .Q(_51716) );
  nnd2s1 _52482_inst ( .DIN1(_50822), .DIN2(_51281), .Q(_50460) );
  hi1s1 _52483_inst ( .DIN(_50688), .Q(_50822) );
  nnd2s1 _52484_inst ( .DIN1(_51719), .DIN2(_51720), .Q(_50688) );
  nor2s1 _52485_inst ( .DIN1(_51393), .DIN2(_51652), .Q(_51719) );
  nnd2s1 _52486_inst ( .DIN1(_51721), .DIN2(_51722), .Q(_50521) );
  nor2s1 _52487_inst ( .DIN1(_51723), .DIN2(_51724), .Q(_51722) );
  nnd2s1 _52488_inst ( .DIN1(_51039), .DIN2(_50812), .Q(_51724) );
  nnd2s1 _52489_inst ( .DIN1(_50602), .DIN2(_50587), .Q(_50812) );
  and2s1 _52490_inst ( .DIN1(_51725), .DIN2(_51726), .Q(_50602) );
  nor2s1 _52491_inst ( .DIN1(_51688), .DIN2(_51727), .Q(_51726) );
  nnd2s1 _52492_inst ( .DIN1(_51524), .DIN2(_26327), .Q(_51727) );
  nnd2s1 _52493_inst ( .DIN1(_2061), .DIN2(_26444), .Q(_51688) );
  nor2s1 _52494_inst ( .DIN1(_51153), .DIN2(_51728), .Q(_51725) );
  nnd2s1 _52495_inst ( .DIN1(_51729), .DIN2(_51637), .Q(_51728) );
  hi1s1 _52496_inst ( .DIN(_51501), .Q(_51637) );
  nnd2s1 _52497_inst ( .DIN1(_51508), .DIN2(_51510), .Q(_51501) );
  nor2s1 _52498_inst ( .DIN1(_51392), .DIN2(_2025), .Q(_51508) );
  nnd2s1 _52499_inst ( .DIN1(_50835), .DIN2(_51102), .Q(_51039) );
  hi1s1 _52500_inst ( .DIN(_50591), .Q(_50835) );
  nnd2s1 _52501_inst ( .DIN1(_51730), .DIN2(_51731), .Q(_50591) );
  nor2s1 _52502_inst ( .DIN1(_51176), .DIN2(_51732), .Q(_51731) );
  nnd2s1 _52503_inst ( .DIN1(_2030), .DIN2(_51510), .Q(_51732) );
  nor2s1 _52504_inst ( .DIN1(_51651), .DIN2(_51673), .Q(_51730) );
  nor2s1 _52505_inst ( .DIN1(_50629), .DIN2(_51733), .Q(_51723) );
  nor2s1 _52506_inst ( .DIN1(_51076), .DIN2(_51118), .Q(_51733) );
  nnd2s1 _52507_inst ( .DIN1(_50910), .DIN2(_50630), .Q(_51118) );
  nnd2s1 _52508_inst ( .DIN1(_51734), .DIN2(_51720), .Q(_50630) );
  and2s1 _52509_inst ( .DIN1(_51735), .DIN2(_51408), .Q(_51720) );
  nor2s1 _52510_inst ( .DIN1(_40396), .DIN2(_51636), .Q(_51735) );
  nor2s1 _52511_inst ( .DIN1(_2025), .DIN2(_51673), .Q(_51734) );
  nnd2s1 _52512_inst ( .DIN1(_51578), .DIN2(_51729), .Q(_51673) );
  hi1s1 _52513_inst ( .DIN(_51447), .Q(_51578) );
  nnd2s1 _52514_inst ( .DIN1(_51736), .DIN2(_2026), .Q(_51447) );
  nor2s1 _52515_inst ( .DIN1(_2015), .DIN2(_26641), .Q(_51736) );
  nnd2s1 _52516_inst ( .DIN1(_51737), .DIN2(_51738), .Q(_50910) );
  nor2s1 _52517_inst ( .DIN1(_2030), .DIN2(_51646), .Q(_51738) );
  nor2s1 _52518_inst ( .DIN1(_51651), .DIN2(_51247), .Q(_51737) );
  nnd2s1 _52519_inst ( .DIN1(_51537), .DIN2(_2025), .Q(_51247) );
  nor2s1 _52520_inst ( .DIN1(_2022), .DIN2(_51392), .Q(_51537) );
  hi1s1 _52521_inst ( .DIN(_51186), .Q(_51076) );
  nnd2s1 _52522_inst ( .DIN1(_51739), .DIN2(_51740), .Q(_51186) );
  nor2s1 _52523_inst ( .DIN1(_51034), .DIN2(_51741), .Q(_51740) );
  nor2s1 _52524_inst ( .DIN1(_51153), .DIN2(_51672), .Q(_51739) );
  nnd2s1 _52525_inst ( .DIN1(_51742), .DIN2(_51408), .Q(_51672) );
  hi1s1 _52526_inst ( .DIN(_50980), .Q(_51408) );
  nnd2s1 _52527_inst ( .DIN1(_51743), .DIN2(_2022), .Q(_50980) );
  nor2s1 _52528_inst ( .DIN1(_2030), .DIN2(_51392), .Q(_51743) );
  or2s1 _52529_inst ( .DIN1(_2027), .DIN2(_2031), .Q(_51392) );
  nor2s1 _52530_inst ( .DIN1(_2025), .DIN2(_51695), .Q(_51742) );
  nnd2s1 _52531_inst ( .DIN1(_51744), .DIN2(_2026), .Q(_51153) );
  nor2s1 _52532_inst ( .DIN1(_2023), .DIN2(_26277), .Q(_51744) );
  hi1s1 _52533_inst ( .DIN(_51102), .Q(_50629) );
  nnd2s1 _52534_inst ( .DIN1(_50664), .DIN2(_50590), .Q(_51102) );
  nnd2s1 _52535_inst ( .DIN1(_51634), .DIN2(_51745), .Q(_50590) );
  nnd2s1 _52536_inst ( .DIN1(_51281), .DIN2(_51746), .Q(_50664) );
  nnd2s1 _52537_inst ( .DIN1(_51745), .DIN2(______[16]), .Q(_51746) );
  and2s1 _52538_inst ( .DIN1(_50871), .DIN2(_51089), .Q(_51721) );
  nor2s1 _52539_inst ( .DIN1(_50592), .DIN2(_51747), .Q(_51089) );
  nor2s1 _52540_inst ( .DIN1(_50829), .DIN2(_50605), .Q(_51747) );
  nnd2s1 _52541_inst ( .DIN1(_51748), .DIN2(_51749), .Q(_50829) );
  nor2s1 _52542_inst ( .DIN1(_51695), .DIN2(_51741), .Q(_51749) );
  nnd2s1 _52543_inst ( .DIN1(_2063), .DIN2(_26321), .Q(_51741) );
  nor2s1 _52544_inst ( .DIN1(_51547), .DIN2(_51696), .Q(_51748) );
  hi1s1 _52545_inst ( .DIN(_51718), .Q(_51696) );
  nor2s1 _52546_inst ( .DIN1(_51750), .DIN2(_51484), .Q(_51718) );
  nnd2s1 _52547_inst ( .DIN1(_26327), .DIN2(_2027), .Q(_51750) );
  nnd2s1 _52548_inst ( .DIN1(_51272), .DIN2(_51223), .Q(_51547) );
  hi1s1 _52549_inst ( .DIN(_51034), .Q(_51223) );
  nnd2s1 _52550_inst ( .DIN1(_2006), .DIN2(_26326), .Q(_51034) );
  hi1s1 _52551_inst ( .DIN(_51210), .Q(_51272) );
  nnd2s1 _52552_inst ( .DIN1(_51751), .DIN2(_51752), .Q(_50592) );
  nnd2s1 _52553_inst ( .DIN1(_50473), .DIN2(_51316), .Q(_51752) );
  nnd2s1 _52554_inst ( .DIN1(_50498), .DIN2(_50661), .Q(_51316) );
  nnd2s1 _52555_inst ( .DIN1(_51714), .DIN2(_51634), .Q(_50661) );
  nor2s1 _52556_inst ( .DIN1(_26771), .DIN2(_50605), .Q(_51634) );
  nnd2s1 _52557_inst ( .DIN1(_51281), .DIN2(_51753), .Q(_50498) );
  nnd2s1 _52558_inst ( .DIN1(_51714), .DIN2(______[16]), .Q(_51753) );
  nor2s1 _52559_inst ( .DIN1(_51657), .DIN2(_27448), .Q(_51714) );
  hi1s1 _52560_inst ( .DIN(______[25]), .Q(_51657) );
  hi1s1 _52561_inst ( .DIN(_51195), .Q(_50473) );
  nnd2s1 _52562_inst ( .DIN1(_51754), .DIN2(_51755), .Q(_51195) );
  nor2s1 _52563_inst ( .DIN1(_51646), .DIN2(_51756), .Q(_51755) );
  nnd2s1 _52564_inst ( .DIN1(_51524), .DIN2(_45588), .Q(_51756) );
  hi1s1 _52565_inst ( .DIN(_40396), .Q(_45588) );
  nnd2s1 _52566_inst ( .DIN1(_26254), .DIN2(_26444), .Q(_40396) );
  hi1s1 _52567_inst ( .DIN(_51659), .Q(_51524) );
  nnd2s1 _52568_inst ( .DIN1(_51757), .DIN2(_2062), .Q(_51659) );
  nor2s1 _52569_inst ( .DIN1(_2057), .DIN2(_2056), .Q(_51757) );
  nnd2s1 _52570_inst ( .DIN1(_51729), .DIN2(_51607), .Q(_51646) );
  hi1s1 _52571_inst ( .DIN(_51387), .Q(_51607) );
  nnd2s1 _52572_inst ( .DIN1(_51758), .DIN2(_2023), .Q(_51387) );
  nor2s1 _52573_inst ( .DIN1(_2026), .DIN2(_2015), .Q(_51758) );
  hi1s1 _52574_inst ( .DIN(_51759), .Q(_51729) );
  nor2s1 _52575_inst ( .DIN1(_26327), .DIN2(_51269), .Q(_51754) );
  hi1s1 _52576_inst ( .DIN(_50987), .Q(_51269) );
  nor2s1 _52577_inst ( .DIN1(_51484), .DIN2(_2027), .Q(_50987) );
  nnd2s1 _52578_inst ( .DIN1(_51760), .DIN2(_2031), .Q(_51484) );
  nor2s1 _52579_inst ( .DIN1(_2025), .DIN2(_2022), .Q(_51760) );
  nnd2s1 _52580_inst ( .DIN1(_51461), .DIN2(_51281), .Q(_51751) );
  hi1s1 _52581_inst ( .DIN(_50837), .Q(_51461) );
  nnd2s1 _52582_inst ( .DIN1(_51761), .DIN2(_51762), .Q(_50837) );
  nor2s1 _52583_inst ( .DIN1(_2022), .DIN2(_51636), .Q(_51762) );
  nor2s1 _52584_inst ( .DIN1(_51351), .DIN2(_51668), .Q(_51761) );
  nnd2s1 _52585_inst ( .DIN1(_51763), .DIN2(_51341), .Q(_51668) );
  hi1s1 _52586_inst ( .DIN(_51228), .Q(_51341) );
  and2s1 _52587_inst ( .DIN1(_51764), .DIN2(_51765), .Q(_50871) );
  nnd2s1 _52588_inst ( .DIN1(_51766), .DIN2(_51281), .Q(_51765) );
  nnd2s1 _52589_inst ( .DIN1(_50798), .DIN2(_51065), .Q(_51766) );
  nnd2s1 _52590_inst ( .DIN1(_51767), .DIN2(_51768), .Q(_51065) );
  nor2s1 _52591_inst ( .DIN1(_51636), .DIN2(_51510), .Q(_51768) );
  hi1s1 _52592_inst ( .DIN(_2022), .Q(_51510) );
  nnd2s1 _52593_inst ( .DIN1(_51769), .DIN2(_2057), .Q(_51636) );
  nor2s1 _52594_inst ( .DIN1(_2056), .DIN2(_26647), .Q(_51769) );
  nor2s1 _52595_inst ( .DIN1(_51210), .DIN2(_51682), .Q(_51767) );
  nnd2s1 _52596_inst ( .DIN1(_51763), .DIN2(_51579), .Q(_51682) );
  nor2s1 _52597_inst ( .DIN1(_26254), .DIN2(_51665), .Q(_51763) );
  nnd2s1 _52598_inst ( .DIN1(_51770), .DIN2(_51771), .Q(_51665) );
  nor2s1 _52599_inst ( .DIN1(_2064), .DIN2(_2063), .Q(_51771) );
  nor2s1 _52600_inst ( .DIN1(_26327), .DIN2(_51176), .Q(_51770) );
  nnd2s1 _52601_inst ( .DIN1(_51772), .DIN2(_2031), .Q(_51176) );
  nor2s1 _52602_inst ( .DIN1(_2027), .DIN2(_51393), .Q(_51772) );
  hi1s1 _52603_inst ( .DIN(_2025), .Q(_51393) );
  nnd2s1 _52604_inst ( .DIN1(_51773), .DIN2(_51774), .Q(_50798) );
  nor2s1 _52605_inst ( .DIN1(_51759), .DIN2(_51775), .Q(_51774) );
  nnd2s1 _52606_inst ( .DIN1(_2025), .DIN2(_26327), .Q(_51775) );
  nnd2s1 _52607_inst ( .DIN1(_51559), .DIN2(_26321), .Q(_51759) );
  hi1s1 _52608_inst ( .DIN(_51351), .Q(_51559) );
  nnd2s1 _52609_inst ( .DIN1(_1986), .DIN2(_2006), .Q(_51351) );
  nor2s1 _52610_inst ( .DIN1(_51228), .DIN2(_51776), .Q(_51773) );
  or2s1 _52611_inst ( .DIN1(_51651), .DIN2(_51476), .Q(_51776) );
  nnd2s1 _52612_inst ( .DIN1(_51777), .DIN2(_2027), .Q(_51476) );
  nor2s1 _52613_inst ( .DIN1(_2031), .DIN2(_2022), .Q(_51777) );
  nnd2s1 _52614_inst ( .DIN1(_51361), .DIN2(_51296), .Q(_51651) );
  and2s1 _52615_inst ( .DIN1(_51778), .DIN2(_2062), .Q(_51296) );
  nor2s1 _52616_inst ( .DIN1(_2057), .DIN2(_26280), .Q(_51778) );
  nor2s1 _52617_inst ( .DIN1(_26444), .DIN2(_2061), .Q(_51361) );
  nnd2s1 _52618_inst ( .DIN1(_51779), .DIN2(_2015), .Q(_51228) );
  nnd2s1 _52619_inst ( .DIN1(_51241), .DIN2(_50587), .Q(_51764) );
  nnd2s1 _52620_inst ( .DIN1(_50962), .DIN2(_50501), .Q(_50587) );
  nnd2s1 _52621_inst ( .DIN1(_51614), .DIN2(_51745), .Q(_50501) );
  nor2s1 _52622_inst ( .DIN1(_50605), .DIN2(______[16]), .Q(_51614) );
  nnd2s1 _52623_inst ( .DIN1(_51281), .DIN2(_51780), .Q(_50962) );
  nnd2s1 _52624_inst ( .DIN1(_51745), .DIN2(_26772), .Q(_51780) );
  nor2s1 _52625_inst ( .DIN1(_27448), .DIN2(______[25]), .Q(_51745) );
  hi1s1 _52626_inst ( .DIN(_51232), .Q(_51241) );
  nnd2s1 _52627_inst ( .DIN1(_51781), .DIN2(_51782), .Q(_51232) );
  nor2s1 _52628_inst ( .DIN1(_51695), .DIN2(_51783), .Q(_51782) );
  nnd2s1 _52629_inst ( .DIN1(_2063), .DIN2(_26327), .Q(_51783) );
  nnd2s1 _52630_inst ( .DIN1(_51572), .DIN2(_26254), .Q(_51695) );
  and2s1 _52631_inst ( .DIN1(_51702), .DIN2(_2056), .Q(_51572) );
  nor2s1 _52632_inst ( .DIN1(_2062), .DIN2(_2057), .Q(_51702) );
  nor2s1 _52633_inst ( .DIN1(_51652), .DIN2(_51083), .Q(_51781) );
  nnd2s1 _52634_inst ( .DIN1(_51615), .DIN2(_2025), .Q(_51083) );
  and2s1 _52635_inst ( .DIN1(_51784), .DIN2(_2022), .Q(_51615) );
  nor2s1 _52636_inst ( .DIN1(_2031), .DIN2(_26413), .Q(_51784) );
  nnd2s1 _52637_inst ( .DIN1(_51785), .DIN2(_51579), .Q(_51652) );
  nor2s1 _52638_inst ( .DIN1(_26326), .DIN2(_2006), .Q(_51579) );
  nor2s1 _52639_inst ( .DIN1(_2064), .DIN2(_51210), .Q(_51785) );
  nnd2s1 _52640_inst ( .DIN1(_51779), .DIN2(_26277), .Q(_51210) );
  nor2s1 _52641_inst ( .DIN1(_2026), .DIN2(_2023), .Q(_51779) );
  nnd2s1 _52642_inst ( .DIN1(_51786), .DIN2(_51787), .Q(____0___________0[9])
         );
  nor2s1 _52643_inst ( .DIN1(_51788), .DIN2(_51789), .Q(_51787) );
  nnd2s1 _52644_inst ( .DIN1(_51790), .DIN2(_51791), .Q(_51789) );
  nor2s1 _52645_inst ( .DIN1(_51792), .DIN2(_51793), .Q(_51791) );
  nor2s1 _52646_inst ( .DIN1(_51794), .DIN2(_51795), .Q(_51793) );
  nor2s1 _52647_inst ( .DIN1(_51796), .DIN2(_51797), .Q(_51792) );
  nor2s1 _52648_inst ( .DIN1(_51798), .DIN2(_51799), .Q(_51797) );
  nor2s1 _52649_inst ( .DIN1(_51800), .DIN2(_51801), .Q(_51790) );
  nor2s1 _52650_inst ( .DIN1(_51802), .DIN2(_51803), .Q(_51800) );
  nnd2s1 _52651_inst ( .DIN1(_51804), .DIN2(_51805), .Q(_51788) );
  nor2s1 _52652_inst ( .DIN1(_51806), .DIN2(_51807), .Q(_51805) );
  nor2s1 _52653_inst ( .DIN1(_51808), .DIN2(_51809), .Q(_51804) );
  nor2s1 _52654_inst ( .DIN1(_51810), .DIN2(_51811), .Q(_51786) );
  nnd2s1 _52655_inst ( .DIN1(_51812), .DIN2(_51813), .Q(_51811) );
  nor2s1 _52656_inst ( .DIN1(_51814), .DIN2(_51815), .Q(_51813) );
  nor2s1 _52657_inst ( .DIN1(_26807), .DIN2(_51817), .Q(_51815) );
  nor2s1 _52658_inst ( .DIN1(_51818), .DIN2(_51819), .Q(_51814) );
  nor2s1 _52659_inst ( .DIN1(_51820), .DIN2(_51821), .Q(_51812) );
  nnd2s1 _52660_inst ( .DIN1(_51822), .DIN2(_51823), .Q(_51810) );
  nor2s1 _52661_inst ( .DIN1(_51824), .DIN2(_51825), .Q(_51823) );
  nor2s1 _52662_inst ( .DIN1(_51826), .DIN2(_51827), .Q(_51822) );
  nnd2s1 _52663_inst ( .DIN1(_51828), .DIN2(_51829), .Q(____0___________0[8])
         );
  nor2s1 _52664_inst ( .DIN1(_51830), .DIN2(_51831), .Q(_51829) );
  nnd2s1 _52665_inst ( .DIN1(_51832), .DIN2(_51833), .Q(_51831) );
  nor2s1 _52666_inst ( .DIN1(_51834), .DIN2(_51835), .Q(_51833) );
  hi1s1 _52667_inst ( .DIN(_51836), .Q(_51835) );
  nor2s1 _52668_inst ( .DIN1(_51837), .DIN2(_51838), .Q(_51832) );
  nnd2s1 _52669_inst ( .DIN1(_51839), .DIN2(_51840), .Q(_51830) );
  nor2s1 _52670_inst ( .DIN1(_51841), .DIN2(_51842), .Q(_51840) );
  nnd2s1 _52671_inst ( .DIN1(_51817), .DIN2(_51843), .Q(_51842) );
  nor2s1 _52672_inst ( .DIN1(_51844), .DIN2(_51845), .Q(_51839) );
  nor2s1 _52673_inst ( .DIN1(_51818), .DIN2(_51846), .Q(_51844) );
  nor2s1 _52674_inst ( .DIN1(_51847), .DIN2(_51848), .Q(_51828) );
  nnd2s1 _52675_inst ( .DIN1(_51849), .DIN2(_51850), .Q(_51848) );
  nor2s1 _52676_inst ( .DIN1(_51851), .DIN2(_51852), .Q(_51850) );
  nor2s1 _52677_inst ( .DIN1(_51853), .DIN2(_51854), .Q(_51849) );
  nnd2s1 _52678_inst ( .DIN1(_51855), .DIN2(_51856), .Q(_51854) );
  nnd2s1 _52679_inst ( .DIN1(_51857), .DIN2(_51794), .Q(_51856) );
  nnd2s1 _52680_inst ( .DIN1(_51858), .DIN2(_51859), .Q(_51855) );
  nnd2s1 _52681_inst ( .DIN1(_51860), .DIN2(_51861), .Q(_51859) );
  nnd2s1 _52682_inst ( .DIN1(_51862), .DIN2(_51863), .Q(_51847) );
  nor2s1 _52683_inst ( .DIN1(_51864), .DIN2(_51865), .Q(_51863) );
  nor2s1 _52684_inst ( .DIN1(_51866), .DIN2(_51867), .Q(_51862) );
  nnd2s1 _52685_inst ( .DIN1(_51868), .DIN2(_51869), .Q(____0___________0[7])
         );
  nor2s1 _52686_inst ( .DIN1(_51870), .DIN2(_51871), .Q(_51869) );
  nnd2s1 _52687_inst ( .DIN1(_51872), .DIN2(_51873), .Q(_51871) );
  nnd2s1 _52688_inst ( .DIN1(_51874), .DIN2(_26807), .Q(_51872) );
  nnd2s1 _52689_inst ( .DIN1(_51875), .DIN2(_51876), .Q(_51870) );
  nor2s1 _52690_inst ( .DIN1(_51877), .DIN2(_51809), .Q(_51875) );
  nor2s1 _52691_inst ( .DIN1(_51878), .DIN2(_51879), .Q(_51868) );
  nnd2s1 _52692_inst ( .DIN1(_51880), .DIN2(_51881), .Q(_51879) );
  hi1s1 _52693_inst ( .DIN(_51882), .Q(_51881) );
  nnd2s1 _52694_inst ( .DIN1(_51883), .DIN2(_51884), .Q(_51878) );
  hi1s1 _52695_inst ( .DIN(_51885), .Q(_51884) );
  nor2s1 _52696_inst ( .DIN1(_51886), .DIN2(_51887), .Q(_51883) );
  nor2s1 _52697_inst ( .DIN1(_51888), .DIN2(_51889), .Q(_51886) );
  nnd2s1 _52698_inst ( .DIN1(_51890), .DIN2(_51891), .Q(____0___________0[6])
         );
  nor2s1 _52699_inst ( .DIN1(_51892), .DIN2(_51893), .Q(_51891) );
  nnd2s1 _52700_inst ( .DIN1(_51894), .DIN2(_51895), .Q(_51893) );
  nor2s1 _52701_inst ( .DIN1(_51896), .DIN2(_51897), .Q(_51895) );
  nor2s1 _52702_inst ( .DIN1(_26807), .DIN2(_51898), .Q(_51897) );
  nor2s1 _52703_inst ( .DIN1(_51888), .DIN2(_51899), .Q(_51896) );
  nor2s1 _52704_inst ( .DIN1(_51900), .DIN2(_51901), .Q(_51899) );
  nor2s1 _52705_inst ( .DIN1(_51902), .DIN2(_51824), .Q(_51894) );
  nnd2s1 _52706_inst ( .DIN1(_51903), .DIN2(_51904), .Q(_51824) );
  nor2s1 _52707_inst ( .DIN1(_51905), .DIN2(_51906), .Q(_51904) );
  nnd2s1 _52708_inst ( .DIN1(_51907), .DIN2(_51908), .Q(_51906) );
  nnd2s1 _52709_inst ( .DIN1(_51909), .DIN2(_51858), .Q(_51908) );
  hi1s1 _52710_inst ( .DIN(_51910), .Q(_51907) );
  nnd2s1 _52711_inst ( .DIN1(_51911), .DIN2(_51912), .Q(_51905) );
  nnd2s1 _52712_inst ( .DIN1(_50605), .DIN2(_26835), .Q(_51912) );
  nor2s1 _52713_inst ( .DIN1(_51913), .DIN2(_51914), .Q(_51911) );
  nor2s1 _52714_inst ( .DIN1(_51915), .DIN2(_51916), .Q(_51903) );
  nnd2s1 _52715_inst ( .DIN1(_51917), .DIN2(_51918), .Q(_51916) );
  hi1s1 _52716_inst ( .DIN(_51919), .Q(_51918) );
  nor2s1 _52717_inst ( .DIN1(_51920), .DIN2(_51921), .Q(_51917) );
  nor2s1 _52718_inst ( .DIN1(_26847), .DIN2(_51922), .Q(_51921) );
  nor2s1 _52719_inst ( .DIN1(_51796), .DIN2(_51923), .Q(_51920) );
  nnd2s1 _52720_inst ( .DIN1(_51924), .DIN2(_51925), .Q(_51915) );
  nor2s1 _52721_inst ( .DIN1(_51858), .DIN2(_51860), .Q(_51902) );
  nnd2s1 _52722_inst ( .DIN1(_51926), .DIN2(_51927), .Q(_51892) );
  nor2s1 _52723_inst ( .DIN1(_51928), .DIN2(_51929), .Q(_51927) );
  nor2s1 _52724_inst ( .DIN1(_51930), .DIN2(_51931), .Q(_51926) );
  nor2s1 _52725_inst ( .DIN1(_51932), .DIN2(_51933), .Q(_51890) );
  nnd2s1 _52726_inst ( .DIN1(_51934), .DIN2(_51935), .Q(_51933) );
  nor2s1 _52727_inst ( .DIN1(_51936), .DIN2(_51937), .Q(_51935) );
  nor2s1 _52728_inst ( .DIN1(_51938), .DIN2(_51939), .Q(_51934) );
  nnd2s1 _52729_inst ( .DIN1(_51940), .DIN2(_51941), .Q(_51939) );
  nnd2s1 _52730_inst ( .DIN1(_51942), .DIN2(_26847), .Q(_51941) );
  nnd2s1 _52731_inst ( .DIN1(_51943), .DIN2(_51944), .Q(_51932) );
  nor2s1 _52732_inst ( .DIN1(_51945), .DIN2(_51946), .Q(_51944) );
  nor2s1 _52733_inst ( .DIN1(_51947), .DIN2(_51948), .Q(_51943) );
  nnd2s1 _52734_inst ( .DIN1(_51949), .DIN2(_51950), .Q(____0___________0[5])
         );
  nor2s1 _52735_inst ( .DIN1(_51951), .DIN2(_51952), .Q(_51950) );
  nnd2s1 _52736_inst ( .DIN1(_51953), .DIN2(_51954), .Q(_51952) );
  nor2s1 _52737_inst ( .DIN1(_51955), .DIN2(_51956), .Q(_51954) );
  nor2s1 _52738_inst ( .DIN1(_51957), .DIN2(_51825), .Q(_51953) );
  nnd2s1 _52739_inst ( .DIN1(_51958), .DIN2(_51959), .Q(_51825) );
  nor2s1 _52740_inst ( .DIN1(_51960), .DIN2(_51961), .Q(_51959) );
  nor2s1 _52741_inst ( .DIN1(_26289), .DIN2(_51962), .Q(_51961) );
  nor2s1 _52742_inst ( .DIN1(_51796), .DIN2(_51963), .Q(_51960) );
  nor2s1 _52743_inst ( .DIN1(_51964), .DIN2(_51965), .Q(_51958) );
  nor2s1 _52744_inst ( .DIN1(_26807), .DIN2(_51966), .Q(_51965) );
  nor2s1 _52745_inst ( .DIN1(_26847), .DIN2(_51967), .Q(_51957) );
  nnd2s1 _52746_inst ( .DIN1(_51968), .DIN2(_51969), .Q(_51951) );
  nor2s1 _52747_inst ( .DIN1(_51970), .DIN2(_51971), .Q(_51969) );
  nor2s1 _52748_inst ( .DIN1(_51972), .DIN2(_51914), .Q(_51968) );
  nor2s1 _52749_inst ( .DIN1(_51973), .DIN2(_51974), .Q(_51949) );
  nnd2s1 _52750_inst ( .DIN1(_51975), .DIN2(_51976), .Q(_51974) );
  hi1s1 _52751_inst ( .DIN(_51977), .Q(_51976) );
  nor2s1 _52752_inst ( .DIN1(_51978), .DIN2(_51979), .Q(_51975) );
  nnd2s1 _52753_inst ( .DIN1(_51980), .DIN2(_51981), .Q(_51973) );
  nor2s1 _52754_inst ( .DIN1(_51982), .DIN2(_51983), .Q(_51981) );
  nor2s1 _52755_inst ( .DIN1(_51984), .DIN2(_51985), .Q(_51980) );
  nnd2s1 _52756_inst ( .DIN1(_51986), .DIN2(_51987), .Q(____0___________0[4])
         );
  nor2s1 _52757_inst ( .DIN1(_51988), .DIN2(_51989), .Q(_51987) );
  nnd2s1 _52758_inst ( .DIN1(_51990), .DIN2(_51991), .Q(_51989) );
  hi1s1 _52759_inst ( .DIN(_51992), .Q(_51991) );
  nnd2s1 _52760_inst ( .DIN1(_51993), .DIN2(_51994), .Q(_51988) );
  nnd2s1 _52761_inst ( .DIN1(_51995), .DIN2(_26848), .Q(_51994) );
  nor2s1 _52762_inst ( .DIN1(_51996), .DIN2(_51930), .Q(_51993) );
  nor2s1 _52763_inst ( .DIN1(_51997), .DIN2(_51998), .Q(_51986) );
  nnd2s1 _52764_inst ( .DIN1(_51999), .DIN2(_52000), .Q(_51998) );
  nor2s1 _52765_inst ( .DIN1(_52001), .DIN2(_52002), .Q(_51999) );
  nor2s1 _52766_inst ( .DIN1(_51818), .DIN2(_52003), .Q(_52002) );
  nor2s1 _52767_inst ( .DIN1(_52004), .DIN2(_51985), .Q(_52003) );
  nnd2s1 _52768_inst ( .DIN1(_52005), .DIN2(_52006), .Q(_51985) );
  hi1s1 _52769_inst ( .DIN(_51843), .Q(_52004) );
  nor2s1 _52770_inst ( .DIN1(_52007), .DIN2(_26807), .Q(_52001) );
  nnd2s1 _52771_inst ( .DIN1(_52008), .DIN2(_52009), .Q(_51997) );
  hi1s1 _52772_inst ( .DIN(_51979), .Q(_52009) );
  nnd2s1 _52773_inst ( .DIN1(_52010), .DIN2(_52011), .Q(_51979) );
  nor2s1 _52774_inst ( .DIN1(_52012), .DIN2(_52013), .Q(_52011) );
  nnd2s1 _52775_inst ( .DIN1(_52014), .DIN2(_52015), .Q(_52013) );
  nor2s1 _52776_inst ( .DIN1(_51802), .DIN2(_52016), .Q(_52012) );
  nor2s1 _52777_inst ( .DIN1(_52017), .DIN2(_52018), .Q(_52010) );
  nnd2s1 _52778_inst ( .DIN1(_52019), .DIN2(_52020), .Q(_52018) );
  nnd2s1 _52779_inst ( .DIN1(_52021), .DIN2(_51818), .Q(_52020) );
  nnd2s1 _52780_inst ( .DIN1(_52022), .DIN2(_26807), .Q(_52019) );
  nnd2s1 _52781_inst ( .DIN1(_52023), .DIN2(_52024), .Q(_52022) );
  nnd2s1 _52782_inst ( .DIN1(_52025), .DIN2(_52026), .Q(____0___________0[3])
         );
  nor2s1 _52783_inst ( .DIN1(_52027), .DIN2(_52028), .Q(_52026) );
  nnd2s1 _52784_inst ( .DIN1(_52029), .DIN2(_52030), .Q(_52028) );
  nor2s1 _52785_inst ( .DIN1(_52031), .DIN2(_51865), .Q(_52029) );
  nnd2s1 _52786_inst ( .DIN1(_52032), .DIN2(_52033), .Q(_51865) );
  nor2s1 _52787_inst ( .DIN1(_52034), .DIN2(_52035), .Q(_52033) );
  nnd2s1 _52788_inst ( .DIN1(_52036), .DIN2(_52037), .Q(_52035) );
  nnd2s1 _52789_inst ( .DIN1(_52038), .DIN2(_26835), .Q(_52037) );
  nnd2s1 _52790_inst ( .DIN1(_52039), .DIN2(_52040), .Q(_52038) );
  nnd2s1 _52791_inst ( .DIN1(_52041), .DIN2(_26807), .Q(_52036) );
  nnd2s1 _52792_inst ( .DIN1(_52042), .DIN2(_52043), .Q(_52034) );
  nor2s1 _52793_inst ( .DIN1(_51806), .DIN2(_52044), .Q(_52042) );
  nor2s1 _52794_inst ( .DIN1(_52045), .DIN2(_52046), .Q(_52032) );
  nnd2s1 _52795_inst ( .DIN1(_52047), .DIN2(_52048), .Q(_52046) );
  hi1s1 _52796_inst ( .DIN(_52049), .Q(_52048) );
  nor2s1 _52797_inst ( .DIN1(_52050), .DIN2(_52051), .Q(_52047) );
  nor2s1 _52798_inst ( .DIN1(_51796), .DIN2(_52052), .Q(_52051) );
  and2s1 _52799_inst ( .DIN1(_52053), .DIN2(_52054), .Q(_52052) );
  nor2s1 _52800_inst ( .DIN1(_26289), .DIN2(_52055), .Q(_52050) );
  nnd2s1 _52801_inst ( .DIN1(_52056), .DIN2(_52057), .Q(_52045) );
  hi1s1 _52802_inst ( .DIN(_52058), .Q(_52057) );
  nor2s1 _52803_inst ( .DIN1(_52059), .DIN2(_52060), .Q(_52056) );
  nor2s1 _52804_inst ( .DIN1(_52061), .DIN2(_51794), .Q(_52031) );
  nnd2s1 _52805_inst ( .DIN1(_52062), .DIN2(_52063), .Q(_52027) );
  nor2s1 _52806_inst ( .DIN1(_51964), .DIN2(_51900), .Q(_52063) );
  and2s1 _52807_inst ( .DIN1(_51846), .DIN2(_52064), .Q(_52062) );
  nor2s1 _52808_inst ( .DIN1(_52065), .DIN2(_52066), .Q(_52025) );
  nnd2s1 _52809_inst ( .DIN1(_52067), .DIN2(_52068), .Q(_52066) );
  nor2s1 _52810_inst ( .DIN1(_52069), .DIN2(_52070), .Q(_52068) );
  nor2s1 _52811_inst ( .DIN1(_51818), .DIN2(_52071), .Q(_52070) );
  nor2s1 _52812_inst ( .DIN1(_52072), .DIN2(_52073), .Q(_52071) );
  nnd2s1 _52813_inst ( .DIN1(_51836), .DIN2(_52074), .Q(_52073) );
  nor2s1 _52814_inst ( .DIN1(_52075), .DIN2(_52076), .Q(_51836) );
  hi1s1 _52815_inst ( .DIN(_52077), .Q(_52072) );
  nor2s1 _52816_inst ( .DIN1(_52078), .DIN2(_26807), .Q(_52069) );
  nor2s1 _52817_inst ( .DIN1(_51834), .DIN2(_52079), .Q(_52078) );
  nnd2s1 _52818_inst ( .DIN1(_52023), .DIN2(_51876), .Q(_52079) );
  nnd2s1 _52819_inst ( .DIN1(_52080), .DIN2(_52006), .Q(_51834) );
  nor2s1 _52820_inst ( .DIN1(_52081), .DIN2(_52082), .Q(_52067) );
  nnd2s1 _52821_inst ( .DIN1(_52083), .DIN2(_52084), .Q(_52082) );
  or2s1 _52822_inst ( .DIN1(_51923), .DIN2(_26848), .Q(_52084) );
  nnd2s1 _52823_inst ( .DIN1(_52085), .DIN2(_26848), .Q(_52083) );
  nnd2s1 _52824_inst ( .DIN1(_52086), .DIN2(_52087), .Q(_52065) );
  nor2s1 _52825_inst ( .DIN1(_51882), .DIN2(_52088), .Q(_52087) );
  nnd2s1 _52826_inst ( .DIN1(_52089), .DIN2(_52090), .Q(_51882) );
  nor2s1 _52827_inst ( .DIN1(_52091), .DIN2(_52092), .Q(_52090) );
  nor2s1 _52828_inst ( .DIN1(_52093), .DIN2(_51983), .Q(_52089) );
  nnd2s1 _52829_inst ( .DIN1(_52094), .DIN2(_52095), .Q(_51983) );
  nor2s1 _52830_inst ( .DIN1(_51888), .DIN2(_51803), .Q(_52093) );
  nor2s1 _52831_inst ( .DIN1(_51947), .DIN2(_52096), .Q(_52086) );
  nnd2s1 _52832_inst ( .DIN1(_52097), .DIN2(_52098), .Q(_51947) );
  nnd2s1 _52833_inst ( .DIN1(_51857), .DIN2(_51858), .Q(_52098) );
  hi1s1 _52834_inst ( .DIN(_52099), .Q(_51857) );
  nnd2s1 _52835_inst ( .DIN1(_52100), .DIN2(_52101), .Q(____0___________0[2])
         );
  nor2s1 _52836_inst ( .DIN1(_52102), .DIN2(_52103), .Q(_52101) );
  nnd2s1 _52837_inst ( .DIN1(_52104), .DIN2(_52105), .Q(_52103) );
  nnd2s1 _52838_inst ( .DIN1(_51818), .DIN2(_52106), .Q(_52105) );
  nnd2s1 _52839_inst ( .DIN1(_52107), .DIN2(_52108), .Q(_52106) );
  nor2s1 _52840_inst ( .DIN1(_51930), .DIN2(_52109), .Q(_52104) );
  nor2s1 _52841_inst ( .DIN1(_52110), .DIN2(_26847), .Q(_52109) );
  nor2s1 _52842_inst ( .DIN1(_52111), .DIN2(_52112), .Q(_52110) );
  nnd2s1 _52843_inst ( .DIN1(_52113), .DIN2(_51922), .Q(_52102) );
  nor2s1 _52844_inst ( .DIN1(_52114), .DIN2(_51964), .Q(_52113) );
  nor2s1 _52845_inst ( .DIN1(_52115), .DIN2(_52116), .Q(_52100) );
  nnd2s1 _52846_inst ( .DIN1(_52117), .DIN2(_52118), .Q(_52116) );
  hi1s1 _52847_inst ( .DIN(_52119), .Q(_52118) );
  nnd2s1 _52848_inst ( .DIN1(_52120), .DIN2(_52121), .Q(_52115) );
  hi1s1 _52849_inst ( .DIN(_52122), .Q(_52121) );
  nor2s1 _52850_inst ( .DIN1(_52123), .DIN2(_52124), .Q(_52120) );
  nnd2s1 _52851_inst ( .DIN1(_52125), .DIN2(_52126), .Q(____0___________0[1])
         );
  nor2s1 _52852_inst ( .DIN1(_52127), .DIN2(_52128), .Q(_52126) );
  nnd2s1 _52853_inst ( .DIN1(_52129), .DIN2(_51889), .Q(_52128) );
  nnd2s1 _52854_inst ( .DIN1(_51885), .DIN2(_26807), .Q(_52129) );
  nnd2s1 _52855_inst ( .DIN1(_52130), .DIN2(_52024), .Q(_51885) );
  nor2s1 _52856_inst ( .DIN1(_52131), .DIN2(_52041), .Q(_52130) );
  nnd2s1 _52857_inst ( .DIN1(_52132), .DIN2(_52133), .Q(_52127) );
  nor2s1 _52858_inst ( .DIN1(_52134), .DIN2(_52135), .Q(_52125) );
  nnd2s1 _52859_inst ( .DIN1(_52136), .DIN2(_51880), .Q(_52135) );
  and2s1 _52860_inst ( .DIN1(_52137), .DIN2(_52138), .Q(_51880) );
  nor2s1 _52861_inst ( .DIN1(_52139), .DIN2(_52140), .Q(_52138) );
  nnd2s1 _52862_inst ( .DIN1(_52141), .DIN2(_52142), .Q(_52140) );
  nor2s1 _52863_inst ( .DIN1(_52143), .DIN2(_52144), .Q(_52141) );
  nnd2s1 _52864_inst ( .DIN1(_52145), .DIN2(_52146), .Q(_52139) );
  nor2s1 _52865_inst ( .DIN1(_51929), .DIN2(_52147), .Q(_52146) );
  nor2s1 _52866_inst ( .DIN1(_52148), .DIN2(_52149), .Q(_52145) );
  nor2s1 _52867_inst ( .DIN1(_52150), .DIN2(_52151), .Q(_52137) );
  nnd2s1 _52868_inst ( .DIN1(_52152), .DIN2(_52030), .Q(_52151) );
  and2s1 _52869_inst ( .DIN1(_52153), .DIN2(_52154), .Q(_52030) );
  nor2s1 _52870_inst ( .DIN1(_52155), .DIN2(_52156), .Q(_52154) );
  nor2s1 _52871_inst ( .DIN1(_52157), .DIN2(_52158), .Q(_52153) );
  nor2s1 _52872_inst ( .DIN1(_51827), .DIN2(_51982), .Q(_52152) );
  nnd2s1 _52873_inst ( .DIN1(_52159), .DIN2(_52160), .Q(_51982) );
  nor2s1 _52874_inst ( .DIN1(_52044), .DIN2(_51826), .Q(_52160) );
  nnd2s1 _52875_inst ( .DIN1(_52161), .DIN2(_52162), .Q(_51826) );
  nor2s1 _52876_inst ( .DIN1(_52163), .DIN2(_52164), .Q(_52162) );
  nnd2s1 _52877_inst ( .DIN1(_52074), .DIN2(_52165), .Q(_52164) );
  nnd2s1 _52878_inst ( .DIN1(_51843), .DIN2(_52166), .Q(_52163) );
  nor2s1 _52879_inst ( .DIN1(_52167), .DIN2(_52168), .Q(_52161) );
  nnd2s1 _52880_inst ( .DIN1(_52169), .DIN2(_52170), .Q(_52168) );
  nnd2s1 _52881_inst ( .DIN1(_26848), .DIN2(_52171), .Q(_52170) );
  nnd2s1 _52882_inst ( .DIN1(_52172), .DIN2(_52173), .Q(_52171) );
  or2s1 _52883_inst ( .DIN1(_52040), .DIN2(_51888), .Q(_52169) );
  nor2s1 _52884_inst ( .DIN1(_51818), .DIN2(_51898), .Q(_52167) );
  hi1s1 _52885_inst ( .DIN(_52174), .Q(_52044) );
  nor2s1 _52886_inst ( .DIN1(_51992), .DIN2(_52175), .Q(_52159) );
  nnd2s1 _52887_inst ( .DIN1(_52176), .DIN2(_52177), .Q(_51992) );
  nor2s1 _52888_inst ( .DIN1(_52178), .DIN2(_52179), .Q(_52177) );
  nnd2s1 _52889_inst ( .DIN1(_52180), .DIN2(_52181), .Q(_52179) );
  nnd2s1 _52890_inst ( .DIN1(_52182), .DIN2(_51817), .Q(_52178) );
  nor2s1 _52891_inst ( .DIN1(_52183), .DIN2(_52184), .Q(_52176) );
  nnd2s1 _52892_inst ( .DIN1(_52185), .DIN2(_52186), .Q(_52184) );
  nnd2s1 _52893_inst ( .DIN1(_52187), .DIN2(_26289), .Q(_52186) );
  hi1s1 _52894_inst ( .DIN(_52188), .Q(_52185) );
  nnd2s1 _52895_inst ( .DIN1(_52189), .DIN2(_52190), .Q(_51827) );
  nor2s1 _52896_inst ( .DIN1(_52191), .DIN2(_52192), .Q(_52190) );
  nnd2s1 _52897_inst ( .DIN1(_52039), .DIN2(_52193), .Q(_52192) );
  hi1s1 _52898_inst ( .DIN(_52194), .Q(_52039) );
  nnd2s1 _52899_inst ( .DIN1(_52195), .DIN2(_52196), .Q(_52191) );
  nor2s1 _52900_inst ( .DIN1(_52197), .DIN2(_52198), .Q(_52189) );
  or2s1 _52901_inst ( .DIN1(_52199), .DIN2(_52059), .Q(_52198) );
  nnd2s1 _52902_inst ( .DIN1(_52200), .DIN2(_52201), .Q(_52059) );
  and2s1 _52903_inst ( .DIN1(_52202), .DIN2(_52203), .Q(_52200) );
  nnd2s1 _52904_inst ( .DIN1(_52054), .DIN2(_52204), .Q(_52197) );
  nnd2s1 _52905_inst ( .DIN1(_52205), .DIN2(_26835), .Q(_52204) );
  nnd2s1 _52906_inst ( .DIN1(_52206), .DIN2(_52043), .Q(_52205) );
  nor2s1 _52907_inst ( .DIN1(_52207), .DIN2(_52111), .Q(_52054) );
  hi1s1 _52908_inst ( .DIN(_52208), .Q(_52111) );
  nnd2s1 _52909_inst ( .DIN1(_52209), .DIN2(_52210), .Q(_52150) );
  nor2s1 _52910_inst ( .DIN1(_52211), .DIN2(_52212), .Q(_52210) );
  and2s1 _52911_inst ( .DIN1(_26835), .DIN2(_51845), .Q(_52212) );
  nnd2s1 _52912_inst ( .DIN1(_52015), .DIN2(_52213), .Q(_51845) );
  hi1s1 _52913_inst ( .DIN(_52006), .Q(_52211) );
  nor2s1 _52914_inst ( .DIN1(_52214), .DIN2(_51996), .Q(_52209) );
  nor2s1 _52915_inst ( .DIN1(_51818), .DIN2(_52215), .Q(_52214) );
  hi1s1 _52916_inst ( .DIN(_51874), .Q(_52136) );
  nnd2s1 _52917_inst ( .DIN1(_52007), .DIN2(_52107), .Q(_51874) );
  nor2s1 _52918_inst ( .DIN1(_51964), .DIN2(_51971), .Q(_52007) );
  nnd2s1 _52919_inst ( .DIN1(_52216), .DIN2(_51925), .Q(_52134) );
  and2s1 _52920_inst ( .DIN1(_52217), .DIN2(_52014), .Q(_51925) );
  nnd2s1 _52921_inst ( .DIN1(_52218), .DIN2(_26847), .Q(_52014) );
  nnd2s1 _52922_inst ( .DIN1(_52091), .DIN2(_26835), .Q(_52217) );
  hi1s1 _52923_inst ( .DIN(_52016), .Q(_52091) );
  hi1s1 _52924_inst ( .DIN(_51866), .Q(_52216) );
  nnd2s1 _52925_inst ( .DIN1(_52219), .DIN2(_52220), .Q(_51866) );
  nor2s1 _52926_inst ( .DIN1(_52221), .DIN2(_52222), .Q(_52220) );
  nnd2s1 _52927_inst ( .DIN1(_51803), .DIN2(_52223), .Q(_52222) );
  nor2s1 _52928_inst ( .DIN1(_52224), .DIN2(_52225), .Q(_52219) );
  nor2s1 _52929_inst ( .DIN1(_51796), .DIN2(_52226), .Q(_52225) );
  nor2s1 _52930_inst ( .DIN1(_51995), .DIN2(_52092), .Q(_52226) );
  nnd2s1 _52931_inst ( .DIN1(_52227), .DIN2(_52228), .Q(____0___________0[13])
         );
  nor2s1 _52932_inst ( .DIN1(_52229), .DIN2(_52230), .Q(_52228) );
  nnd2s1 _52933_inst ( .DIN1(_52231), .DIN2(_52232), .Q(_52230) );
  nor2s1 _52934_inst ( .DIN1(_52233), .DIN2(_52234), .Q(_52232) );
  nor2s1 _52935_inst ( .DIN1(_51888), .DIN2(_52235), .Q(_52234) );
  nor2s1 _52936_inst ( .DIN1(_26847), .DIN2(_52201), .Q(_52233) );
  nor2s1 _52937_inst ( .DIN1(_51820), .DIN2(_51910), .Q(_52231) );
  nnd2s1 _52938_inst ( .DIN1(_52180), .DIN2(_52236), .Q(_51910) );
  nnd2s1 _52939_inst ( .DIN1(_52131), .DIN2(_26807), .Q(_52236) );
  nnd2s1 _52940_inst ( .DIN1(_52237), .DIN2(_51818), .Q(_52180) );
  nnd2s1 _52941_inst ( .DIN1(_52238), .DIN2(_52239), .Q(_51820) );
  nor2s1 _52942_inst ( .DIN1(_52240), .DIN2(_52241), .Q(_52239) );
  nnd2s1 _52943_inst ( .DIN1(_52242), .DIN2(_52243), .Q(_52241) );
  nor2s1 _52944_inst ( .DIN1(_52244), .DIN2(_52245), .Q(_52238) );
  nnd2s1 _52945_inst ( .DIN1(_52246), .DIN2(_52247), .Q(_52245) );
  or2s1 _52946_inst ( .DIN1(_52061), .DIN2(_51858), .Q(_52246) );
  nnd2s1 _52947_inst ( .DIN1(_52248), .DIN2(_52249), .Q(_52244) );
  nnd2s1 _52948_inst ( .DIN1(_52075), .DIN2(_26807), .Q(_52249) );
  nnd2s1 _52949_inst ( .DIN1(_51818), .DIN2(_52250), .Q(_52248) );
  nnd2s1 _52950_inst ( .DIN1(_52023), .DIN2(_52174), .Q(_52250) );
  nnd2s1 _52951_inst ( .DIN1(_52251), .DIN2(_52252), .Q(_52229) );
  nor2s1 _52952_inst ( .DIN1(_51901), .DIN2(_51909), .Q(_52252) );
  hi1s1 _52953_inst ( .DIN(_52253), .Q(_51909) );
  nor2s1 _52954_inst ( .DIN1(_52218), .DIN2(_52254), .Q(_52251) );
  hi1s1 _52955_inst ( .DIN(_51873), .Q(_52218) );
  nor2s1 _52956_inst ( .DIN1(_52255), .DIN2(_52256), .Q(_52227) );
  nnd2s1 _52957_inst ( .DIN1(_52257), .DIN2(_52258), .Q(_52256) );
  nor2s1 _52958_inst ( .DIN1(_52259), .DIN2(_52260), .Q(_52258) );
  nor2s1 _52959_inst ( .DIN1(_52077), .DIN2(_26807), .Q(_52260) );
  nor2s1 _52960_inst ( .DIN1(_52261), .DIN2(_52262), .Q(_52077) );
  nor2s1 _52961_inst ( .DIN1(_51818), .DIN2(_52202), .Q(_52259) );
  nor2s1 _52962_inst ( .DIN1(_52263), .DIN2(_52264), .Q(_52257) );
  nnd2s1 _52963_inst ( .DIN1(_52265), .DIN2(_52266), .Q(_52255) );
  nor2s1 _52964_inst ( .DIN1(_52267), .DIN2(_51978), .Q(_52266) );
  nnd2s1 _52965_inst ( .DIN1(_52268), .DIN2(_52269), .Q(_51978) );
  nor2s1 _52966_inst ( .DIN1(_52270), .DIN2(_52149), .Q(_52269) );
  nor2s1 _52967_inst ( .DIN1(_52224), .DIN2(_52271), .Q(_52268) );
  nor2s1 _52968_inst ( .DIN1(_52122), .DIN2(_52272), .Q(_52265) );
  nnd2s1 _52969_inst ( .DIN1(_52273), .DIN2(_52274), .Q(_52122) );
  nnd2s1 _52970_inst ( .DIN1(_52275), .DIN2(_51858), .Q(_52274) );
  nor2s1 _52971_inst ( .DIN1(_51928), .DIN2(_51942), .Q(_52273) );
  nnd2s1 _52972_inst ( .DIN1(_52276), .DIN2(_52277), .Q(____0___________0[12])
         );
  nor2s1 _52973_inst ( .DIN1(_52278), .DIN2(_52279), .Q(_52277) );
  nnd2s1 _52974_inst ( .DIN1(_52280), .DIN2(_52281), .Q(_52279) );
  hi1s1 _52975_inst ( .DIN(_51837), .Q(_52281) );
  nnd2s1 _52976_inst ( .DIN1(_52282), .DIN2(_52283), .Q(_51837) );
  nnd2s1 _52977_inst ( .DIN1(_50605), .DIN2(_51888), .Q(_52283) );
  or2s1 _52978_inst ( .DIN1(_52064), .DIN2(_26807), .Q(_52282) );
  nor2s1 _52979_inst ( .DIN1(_51801), .DIN2(_52049), .Q(_52280) );
  nnd2s1 _52980_inst ( .DIN1(_52284), .DIN2(_52285), .Q(_52049) );
  nnd2s1 _52981_inst ( .DIN1(_52286), .DIN2(_52287), .Q(_52285) );
  nor2s1 _52982_inst ( .DIN1(_52148), .DIN2(_52288), .Q(_52284) );
  nnd2s1 _52983_inst ( .DIN1(_52289), .DIN2(_52290), .Q(_51801) );
  nor2s1 _52984_inst ( .DIN1(_52187), .DIN2(_51900), .Q(_52290) );
  hi1s1 _52985_inst ( .DIN(_51889), .Q(_51900) );
  nor2s1 _52986_inst ( .DIN1(_51841), .DIN2(_52291), .Q(_52289) );
  nor2s1 _52987_inst ( .DIN1(_26289), .DIN2(_52292), .Q(_52291) );
  nor2s1 _52988_inst ( .DIN1(_51888), .DIN2(_52293), .Q(_51841) );
  nnd2s1 _52989_inst ( .DIN1(_52294), .DIN2(_52295), .Q(_52278) );
  nor2s1 _52990_inst ( .DIN1(_52296), .DIN2(_52021), .Q(_52295) );
  hi1s1 _52991_inst ( .DIN(_52107), .Q(_52021) );
  nor2s1 _52992_inst ( .DIN1(_52297), .DIN2(_52298), .Q(_52294) );
  nor2s1 _52993_inst ( .DIN1(_51818), .DIN2(_52174), .Q(_52298) );
  nor2s1 _52994_inst ( .DIN1(_51802), .DIN2(_52040), .Q(_52297) );
  nor2s1 _52995_inst ( .DIN1(_52299), .DIN2(_52300), .Q(_52276) );
  nnd2s1 _52996_inst ( .DIN1(_52301), .DIN2(_52302), .Q(_52300) );
  hi1s1 _52997_inst ( .DIN(_52303), .Q(_52302) );
  nor2s1 _52998_inst ( .DIN1(_52096), .DIN2(_52272), .Q(_52301) );
  nnd2s1 _52999_inst ( .DIN1(_52304), .DIN2(_52305), .Q(_52272) );
  nor2s1 _53000_inst ( .DIN1(_52306), .DIN2(_52307), .Q(_52305) );
  nnd2s1 _53001_inst ( .DIN1(_52099), .DIN2(_51846), .Q(_52307) );
  nor2s1 _53002_inst ( .DIN1(_51858), .DIN2(_52308), .Q(_52306) );
  nor2s1 _53003_inst ( .DIN1(_52309), .DIN2(_52310), .Q(_52304) );
  nor2s1 _53004_inst ( .DIN1(_26807), .DIN2(_52080), .Q(_52309) );
  nnd2s1 _53005_inst ( .DIN1(_51860), .DIN2(_52311), .Q(_52096) );
  nnd2s1 _53006_inst ( .DIN1(_51818), .DIN2(_52312), .Q(_52311) );
  nnd2s1 _53007_inst ( .DIN1(_51819), .DIN2(_51843), .Q(_52312) );
  nnd2s1 _53008_inst ( .DIN1(_52313), .DIN2(_52000), .Q(_52299) );
  and2s1 _53009_inst ( .DIN1(_52314), .DIN2(_52315), .Q(_52000) );
  nor2s1 _53010_inst ( .DIN1(_52316), .DIN2(_52317), .Q(_52315) );
  nnd2s1 _53011_inst ( .DIN1(_52318), .DIN2(_52319), .Q(_52317) );
  nnd2s1 _53012_inst ( .DIN1(_26848), .DIN2(_52320), .Q(_52319) );
  nnd2s1 _53013_inst ( .DIN1(_52321), .DIN2(_52053), .Q(_52320) );
  nor2s1 _53014_inst ( .DIN1(_52322), .DIN2(_52092), .Q(_52321) );
  or2s1 _53015_inst ( .DIN1(_52074), .DIN2(_26807), .Q(_52318) );
  nnd2s1 _53016_inst ( .DIN1(_52055), .DIN2(_52166), .Q(_52316) );
  nor2s1 _53017_inst ( .DIN1(_51984), .DIN2(_52323), .Q(_52314) );
  nnd2s1 _53018_inst ( .DIN1(_52324), .DIN2(_52325), .Q(_52323) );
  nnd2s1 _53019_inst ( .DIN1(_51914), .DIN2(_26835), .Q(_52325) );
  hi1s1 _53020_inst ( .DIN(_52213), .Q(_51914) );
  hi1s1 _53021_inst ( .DIN(_51867), .Q(_52324) );
  nnd2s1 _53022_inst ( .DIN1(_52326), .DIN2(_52327), .Q(_51867) );
  nor2s1 _53023_inst ( .DIN1(_52328), .DIN2(_52329), .Q(_52327) );
  nor2s1 _53024_inst ( .DIN1(_52330), .DIN2(_52331), .Q(_52329) );
  nor2s1 _53025_inst ( .DIN1(_52332), .DIN2(_26289), .Q(_52328) );
  and2s1 _53026_inst ( .DIN1(_52173), .DIN2(_51923), .Q(_52332) );
  nor2s1 _53027_inst ( .DIN1(_52333), .DIN2(_51956), .Q(_52326) );
  nor2s1 _53028_inst ( .DIN1(_51858), .DIN2(_51795), .Q(_51956) );
  nor2s1 _53029_inst ( .DIN1(_51924), .DIN2(_26807), .Q(_52333) );
  nor2s1 _53030_inst ( .DIN1(_51955), .DIN2(_52262), .Q(_51924) );
  nnd2s1 _53031_inst ( .DIN1(_51876), .DIN2(_52334), .Q(_51984) );
  nnd2s1 _53032_inst ( .DIN1(_51901), .DIN2(_51888), .Q(_52334) );
  hi1s1 _53033_inst ( .DIN(_52206), .Q(_51901) );
  nor2s1 _53034_inst ( .DIN1(_51937), .DIN2(_51977), .Q(_52313) );
  nnd2s1 _53035_inst ( .DIN1(_52335), .DIN2(_52336), .Q(_51977) );
  nor2s1 _53036_inst ( .DIN1(_52337), .DIN2(_52338), .Q(_52336) );
  nor2s1 _53037_inst ( .DIN1(_26807), .DIN2(_52247), .Q(_52338) );
  nor2s1 _53038_inst ( .DIN1(_52339), .DIN2(_51802), .Q(_52337) );
  nor2s1 _53039_inst ( .DIN1(_51928), .DIN2(_52194), .Q(_52339) );
  nor2s1 _53040_inst ( .DIN1(_52340), .DIN2(_52341), .Q(_52335) );
  nor2s1 _53041_inst ( .DIN1(_26847), .DIN2(_52208), .Q(_52341) );
  nor2s1 _53042_inst ( .DIN1(_51858), .DIN2(_52142), .Q(_52340) );
  nnd2s1 _53043_inst ( .DIN1(_52342), .DIN2(_52343), .Q(_51937) );
  nor2s1 _53044_inst ( .DIN1(_52344), .DIN2(_52345), .Q(_52343) );
  nnd2s1 _53045_inst ( .DIN1(_52346), .DIN2(_52347), .Q(_52345) );
  hi1s1 _53046_inst ( .DIN(_51821), .Q(_52347) );
  nnd2s1 _53047_inst ( .DIN1(_52348), .DIN2(_52349), .Q(_51821) );
  nnd2s1 _53048_inst ( .DIN1(_51818), .DIN2(_52157), .Q(_52349) );
  hi1s1 _53049_inst ( .DIN(_52350), .Q(_52157) );
  nor2s1 _53050_inst ( .DIN1(_52351), .DIN2(_52352), .Q(_52348) );
  nor2s1 _53051_inst ( .DIN1(_51802), .DIN2(_52353), .Q(_52352) );
  and2s1 _53052_inst ( .DIN1(_52155), .DIN2(_26848), .Q(_52351) );
  nor2s1 _53053_inst ( .DIN1(_52261), .DIN2(_52354), .Q(_52346) );
  nor2s1 _53054_inst ( .DIN1(_51818), .DIN2(_52355), .Q(_52354) );
  nor2s1 _53055_inst ( .DIN1(_51964), .DIN2(_52356), .Q(_52355) );
  nnd2s1 _53056_inst ( .DIN1(_52357), .DIN2(_52006), .Q(_52344) );
  nnd2s1 _53057_inst ( .DIN1(_52358), .DIN2(_46019), .Q(_52006) );
  nor2s1 _53058_inst ( .DIN1(_52359), .DIN2(_52085), .Q(_52357) );
  hi1s1 _53059_inst ( .DIN(_52360), .Q(_52085) );
  nor2s1 _53060_inst ( .DIN1(_52361), .DIN2(_52362), .Q(_52342) );
  nnd2s1 _53061_inst ( .DIN1(_52363), .DIN2(_52364), .Q(_52362) );
  nor2s1 _53062_inst ( .DIN1(_52365), .DIN2(_52366), .Q(_52364) );
  nor2s1 _53063_inst ( .DIN1(_51796), .DIN2(_52094), .Q(_52366) );
  and2s1 _53064_inst ( .DIN1(_51799), .DIN2(_26848), .Q(_52365) );
  nnd2s1 _53065_inst ( .DIN1(_52367), .DIN2(_52368), .Q(_51799) );
  nor2s1 _53066_inst ( .DIN1(_52267), .DIN2(_52088), .Q(_52363) );
  nnd2s1 _53067_inst ( .DIN1(_52369), .DIN2(_52370), .Q(_52088) );
  nor2s1 _53068_inst ( .DIN1(_52371), .DIN2(_52372), .Q(_52370) );
  nnd2s1 _53069_inst ( .DIN1(_52373), .DIN2(_52195), .Q(_52372) );
  nor2s1 _53070_inst ( .DIN1(_51802), .DIN2(_52015), .Q(_52371) );
  nor2s1 _53071_inst ( .DIN1(_52199), .DIN2(_52374), .Q(_52369) );
  nnd2s1 _53072_inst ( .DIN1(_52375), .DIN2(_52376), .Q(_52374) );
  nnd2s1 _53073_inst ( .DIN1(_52143), .DIN2(_26848), .Q(_52375) );
  nnd2s1 _53074_inst ( .DIN1(_52377), .DIN2(_52378), .Q(_52199) );
  nnd2s1 _53075_inst ( .DIN1(_52379), .DIN2(_52380), .Q(_52378) );
  hi1s1 _53076_inst ( .DIN(_52381), .Q(_52380) );
  nor2s1 _53077_inst ( .DIN1(_42924), .DIN2(_51794), .Q(_52379) );
  nor2s1 _53078_inst ( .DIN1(_52114), .DIN2(_52382), .Q(_52377) );
  nor2s1 _53079_inst ( .DIN1(_46022), .DIN2(_52383), .Q(_52382) );
  nnd2s1 _53080_inst ( .DIN1(_52384), .DIN2(_26848), .Q(_52383) );
  hi1s1 _53081_inst ( .DIN(_52385), .Q(_52114) );
  nnd2s1 _53082_inst ( .DIN1(_52386), .DIN2(_52387), .Q(_52267) );
  hi1s1 _53083_inst ( .DIN(_52388), .Q(_52387) );
  nor2s1 _53084_inst ( .DIN1(_52389), .DIN2(_52390), .Q(_52386) );
  nor2s1 _53085_inst ( .DIN1(_51858), .DIN2(_52391), .Q(_52390) );
  nor2s1 _53086_inst ( .DIN1(_51802), .DIN2(_52392), .Q(_52389) );
  nnd2s1 _53087_inst ( .DIN1(_52393), .DIN2(_51990), .Q(_52361) );
  and2s1 _53088_inst ( .DIN1(_52394), .DIN2(_52395), .Q(_51990) );
  nnd2s1 _53089_inst ( .DIN1(_52270), .DIN2(_51888), .Q(_52395) );
  hi1s1 _53090_inst ( .DIN(_52043), .Q(_52270) );
  nor2s1 _53091_inst ( .DIN1(_52060), .DIN2(_52183), .Q(_52393) );
  nnd2s1 _53092_inst ( .DIN1(_52396), .DIN2(_52397), .Q(_52183) );
  nor2s1 _53093_inst ( .DIN1(_51807), .DIN2(_52398), .Q(_52397) );
  hi1s1 _53094_inst ( .DIN(_52399), .Q(_51807) );
  nor2s1 _53095_inst ( .DIN1(_52400), .DIN2(_52401), .Q(_52396) );
  nor2s1 _53096_inst ( .DIN1(_51794), .DIN2(_51861), .Q(_52400) );
  nnd2s1 _53097_inst ( .DIN1(_52108), .DIN2(_52402), .Q(_52060) );
  or2s1 _53098_inst ( .DIN1(_52172), .DIN2(_26289), .Q(_52402) );
  nnd2s1 _53099_inst ( .DIN1(_52403), .DIN2(_52404), .Q(____0___________0[11])
         );
  nor2s1 _53100_inst ( .DIN1(_52405), .DIN2(_52406), .Q(_52404) );
  nnd2s1 _53101_inst ( .DIN1(_52407), .DIN2(_52408), .Q(_52406) );
  nnd2s1 _53102_inst ( .DIN1(_52041), .DIN2(_51818), .Q(_52408) );
  hi1s1 _53103_inst ( .DIN(_52247), .Q(_52041) );
  nnd2s1 _53104_inst ( .DIN1(_52409), .DIN2(_44283), .Q(_52247) );
  hi1s1 _53105_inst ( .DIN(_46028), .Q(_44283) );
  nor2s1 _53106_inst ( .DIN1(_51931), .DIN2(_52410), .Q(_52407) );
  nor2s1 _53107_inst ( .DIN1(_52411), .DIN2(_26847), .Q(_52410) );
  nor2s1 _53108_inst ( .DIN1(_52412), .DIN2(_52413), .Q(_52411) );
  nnd2s1 _53109_inst ( .DIN1(_52055), .DIN2(_51873), .Q(_52413) );
  nnd2s1 _53110_inst ( .DIN1(_52414), .DIN2(_52415), .Q(_51873) );
  nor2s1 _53111_inst ( .DIN1(_52416), .DIN2(_52417), .Q(_52415) );
  nor2s1 _53112_inst ( .DIN1(_33865), .DIN2(_52418), .Q(_52414) );
  nnd2s1 _53113_inst ( .DIN1(_51963), .DIN2(_51923), .Q(_52412) );
  hi1s1 _53114_inst ( .DIN(_52419), .Q(_51931) );
  nnd2s1 _53115_inst ( .DIN1(_52420), .DIN2(_52421), .Q(_52405) );
  and2s1 _53116_inst ( .DIN1(_52422), .DIN2(_52223), .Q(_52421) );
  nor2s1 _53117_inst ( .DIN1(_52147), .DIN2(_52275), .Q(_52420) );
  nor2s1 _53118_inst ( .DIN1(_52423), .DIN2(_52424), .Q(_52403) );
  nnd2s1 _53119_inst ( .DIN1(_52425), .DIN2(_52426), .Q(_52424) );
  nor2s1 _53120_inst ( .DIN1(_52427), .DIN2(_52428), .Q(_52426) );
  nor2s1 _53121_inst ( .DIN1(_51802), .DIN2(_52429), .Q(_52428) );
  nor2s1 _53122_inst ( .DIN1(_51888), .DIN2(_52043), .Q(_52427) );
  nor2s1 _53123_inst ( .DIN1(_52263), .DIN2(_52430), .Q(_52425) );
  nnd2s1 _53124_inst ( .DIN1(_52431), .DIN2(_52432), .Q(_52263) );
  nor2s1 _53125_inst ( .DIN1(_52433), .DIN2(_52434), .Q(_52432) );
  nnd2s1 _53126_inst ( .DIN1(_51962), .DIN2(_52208), .Q(_52434) );
  nnd2s1 _53127_inst ( .DIN1(_52435), .DIN2(_51817), .Q(_52433) );
  nor2s1 _53128_inst ( .DIN1(_51913), .DIN2(_52359), .Q(_52435) );
  nor2s1 _53129_inst ( .DIN1(_52436), .DIN2(_52437), .Q(_52431) );
  nnd2s1 _53130_inst ( .DIN1(_52438), .DIN2(_51940), .Q(_52437) );
  nnd2s1 _53131_inst ( .DIN1(_52187), .DIN2(_26848), .Q(_51940) );
  hi1s1 _53132_inst ( .DIN(_52439), .Q(_52187) );
  hi1s1 _53133_inst ( .DIN(_52440), .Q(_52438) );
  nnd2s1 _53134_inst ( .DIN1(_52441), .DIN2(_52442), .Q(_52436) );
  nnd2s1 _53135_inst ( .DIN1(_52443), .DIN2(_26807), .Q(_52442) );
  nnd2s1 _53136_inst ( .DIN1(_51898), .DIN2(_51843), .Q(_52443) );
  nnd2s1 _53137_inst ( .DIN1(_52444), .DIN2(_45099), .Q(_51843) );
  or2s1 _53138_inst ( .DIN1(_52015), .DIN2(_51888), .Q(_52441) );
  nnd2s1 _53139_inst ( .DIN1(_52445), .DIN2(_52008), .Q(_52423) );
  nor2s1 _53140_inst ( .DIN1(_52123), .DIN2(_51887), .Q(_52008) );
  nor2s1 _53141_inst ( .DIN1(_52368), .DIN2(_51796), .Q(_51887) );
  nnd2s1 _53142_inst ( .DIN1(_52446), .DIN2(_52447), .Q(_52123) );
  nor2s1 _53143_inst ( .DIN1(_52448), .DIN2(_52449), .Q(_52447) );
  nnd2s1 _53144_inst ( .DIN1(_52450), .DIN2(_52097), .Q(_52449) );
  nor2s1 _53145_inst ( .DIN1(_52261), .DIN2(_52254), .Q(_52450) );
  hi1s1 _53146_inst ( .DIN(_52373), .Q(_52254) );
  nnd2s1 _53147_inst ( .DIN1(_52451), .DIN2(_52080), .Q(_52448) );
  and2s1 _53148_inst ( .DIN1(_51819), .DIN2(_52061), .Q(_52451) );
  nor2s1 _53149_inst ( .DIN1(_52452), .DIN2(_52453), .Q(_52446) );
  nnd2s1 _53150_inst ( .DIN1(_52454), .DIN2(_52455), .Q(_52453) );
  nor2s1 _53151_inst ( .DIN1(_52388), .DIN2(_52456), .Q(_52454) );
  nnd2s1 _53152_inst ( .DIN1(_52457), .DIN2(_52308), .Q(_52452) );
  hi1s1 _53153_inst ( .DIN(_51852), .Q(_52308) );
  nor2s1 _53154_inst ( .DIN1(_52271), .DIN2(_51798), .Q(_52457) );
  nnd2s1 _53155_inst ( .DIN1(_52360), .DIN2(_52458), .Q(_51798) );
  nor2s1 _53156_inst ( .DIN1(_51802), .DIN2(_51889), .Q(_52271) );
  nnd2s1 _53157_inst ( .DIN1(_52459), .DIN2(_45819), .Q(_51889) );
  nor2s1 _53158_inst ( .DIN1(_44600), .DIN2(_52418), .Q(_52459) );
  nor2s1 _53159_inst ( .DIN1(_52460), .DIN2(_51838), .Q(_52445) );
  nnd2s1 _53160_inst ( .DIN1(_52461), .DIN2(_52462), .Q(_51838) );
  nnd2s1 _53161_inst ( .DIN1(_52398), .DIN2(_51818), .Q(_52462) );
  hi1s1 _53162_inst ( .DIN(_52242), .Q(_52398) );
  nor2s1 _53163_inst ( .DIN1(_51970), .DIN2(_52463), .Q(_52461) );
  nnd2s1 _53164_inst ( .DIN1(_52464), .DIN2(_52465), .Q(____0___________0[10])
         );
  nor2s1 _53165_inst ( .DIN1(_52466), .DIN2(_52467), .Q(_52465) );
  nnd2s1 _53166_inst ( .DIN1(_52468), .DIN2(_52469), .Q(_52467) );
  nor2s1 _53167_inst ( .DIN1(_52058), .DIN2(_51864), .Q(_52469) );
  nnd2s1 _53168_inst ( .DIN1(_52470), .DIN2(_52471), .Q(_51864) );
  or2s1 _53169_inst ( .DIN1(_52391), .DIN2(_51794), .Q(_52471) );
  nor2s1 _53170_inst ( .DIN1(_52472), .DIN2(_52473), .Q(_52470) );
  nor2s1 _53171_inst ( .DIN1(_51888), .DIN2(_52392), .Q(_52473) );
  nor2s1 _53172_inst ( .DIN1(_51796), .DIN2(_52367), .Q(_52472) );
  nnd2s1 _53173_inst ( .DIN1(_52474), .DIN2(_52475), .Q(_52058) );
  nnd2s1 _53174_inst ( .DIN1(_52275), .DIN2(_51794), .Q(_52475) );
  hi1s1 _53175_inst ( .DIN(_52142), .Q(_52275) );
  nnd2s1 _53176_inst ( .DIN1(_44980), .DIN2(_52476), .Q(_52142) );
  and2s1 _53177_inst ( .DIN1(_52196), .DIN2(_52193), .Q(_52474) );
  nor2s1 _53178_inst ( .DIN1(_52175), .DIN2(_51936), .Q(_52468) );
  nnd2s1 _53179_inst ( .DIN1(_52477), .DIN2(_52061), .Q(_51936) );
  nnd2s1 _53180_inst ( .DIN1(_52478), .DIN2(_52479), .Q(_52061) );
  nor2s1 _53181_inst ( .DIN1(_52480), .DIN2(_52481), .Q(_52479) );
  nnd2s1 _53182_inst ( .DIN1(_52482), .DIN2(_45103), .Q(_52480) );
  nor2s1 _53183_inst ( .DIN1(_53525), .DIN2(_53526), .Q(_52482) );
  nor2s1 _53184_inst ( .DIN1(_52483), .DIN2(_52484), .Q(_52478) );
  nnd2s1 _53185_inst ( .DIN1(_52485), .DIN2(_1860), .Q(_52484) );
  nnd2s1 _53186_inst ( .DIN1(_52486), .DIN2(_1863), .Q(_52483) );
  nor2s1 _53187_inst ( .DIN1(_45104), .DIN2(_52487), .Q(_52486) );
  nor2s1 _53188_inst ( .DIN1(_52488), .DIN2(_52489), .Q(_52477) );
  nor2s1 _53189_inst ( .DIN1(_26807), .DIN2(_51846), .Q(_52489) );
  nor2s1 _53190_inst ( .DIN1(_51818), .DIN2(_52064), .Q(_52488) );
  nnd2s1 _53191_inst ( .DIN1(_52490), .DIN2(_52491), .Q(_52175) );
  nor2s1 _53192_inst ( .DIN1(_52262), .DIN2(_52492), .Q(_52491) );
  nnd2s1 _53193_inst ( .DIN1(_52422), .DIN2(_51923), .Q(_52492) );
  nnd2s1 _53194_inst ( .DIN1(_52444), .DIN2(_46026), .Q(_51923) );
  nnd2s1 _53195_inst ( .DIN1(_52286), .DIN2(_52493), .Q(_52422) );
  nnd2s1 _53196_inst ( .DIN1(_52330), .DIN2(_52494), .Q(_52493) );
  hi1s1 _53197_inst ( .DIN(_52331), .Q(_52286) );
  nnd2s1 _53198_inst ( .DIN1(_46030), .DIN2(_51818), .Q(_52331) );
  and2s1 _53199_inst ( .DIN1(_44317), .DIN2(_52495), .Q(_52262) );
  nor2s1 _53200_inst ( .DIN1(_52075), .DIN2(_52496), .Q(_52490) );
  nor2s1 _53201_inst ( .DIN1(_51888), .DIN2(_51281), .Q(_52496) );
  nnd2s1 _53202_inst ( .DIN1(_52497), .DIN2(_52498), .Q(_52466) );
  nor2s1 _53203_inst ( .DIN1(_51877), .DIN2(_52207), .Q(_52498) );
  nor2s1 _53204_inst ( .DIN1(_52499), .DIN2(_52500), .Q(_52497) );
  nor2s1 _53205_inst ( .DIN1(_51794), .DIN2(_52253), .Q(_52500) );
  nor2s1 _53206_inst ( .DIN1(_26807), .DIN2(_52202), .Q(_52499) );
  nnd2s1 _53207_inst ( .DIN1(_52501), .DIN2(_52502), .Q(_52202) );
  nor2s1 _53208_inst ( .DIN1(_44657), .DIN2(_42923), .Q(_52502) );
  nor2s1 _53209_inst ( .DIN1(_52503), .DIN2(_52504), .Q(_52464) );
  nnd2s1 _53210_inst ( .DIN1(_52505), .DIN2(_52506), .Q(_52504) );
  nor2s1 _53211_inst ( .DIN1(_52507), .DIN2(_52508), .Q(_52506) );
  nor2s1 _53212_inst ( .DIN1(_51802), .DIN2(_52043), .Q(_52508) );
  nnd2s1 _53213_inst ( .DIN1(_52509), .DIN2(_52510), .Q(_52043) );
  nor2s1 _53214_inst ( .DIN1(_43029), .DIN2(_52418), .Q(_52509) );
  hi1s1 _53215_inst ( .DIN(_52511), .Q(_52418) );
  nor2s1 _53216_inst ( .DIN1(_51888), .DIN2(_52097), .Q(_52507) );
  nor2s1 _53217_inst ( .DIN1(_52512), .DIN2(_52513), .Q(_52505) );
  nnd2s1 _53218_inst ( .DIN1(_52514), .DIN2(_52515), .Q(_52513) );
  nnd2s1 _53219_inst ( .DIN1(_52288), .DIN2(_26289), .Q(_52515) );
  nnd2s1 _53220_inst ( .DIN1(_52149), .DIN2(_26848), .Q(_52514) );
  hi1s1 _53221_inst ( .DIN(_52053), .Q(_52149) );
  nnd2s1 _53222_inst ( .DIN1(_52516), .DIN2(_52517), .Q(_52503) );
  nor2s1 _53223_inst ( .DIN1(_52081), .DIN2(_52124), .Q(_52517) );
  nnd2s1 _53224_inst ( .DIN1(_52518), .DIN2(_52519), .Q(_52124) );
  nnd2s1 _53225_inst ( .DIN1(_52224), .DIN2(_26848), .Q(_52519) );
  hi1s1 _53226_inst ( .DIN(_52368), .Q(_52224) );
  nnd2s1 _53227_inst ( .DIN1(_52520), .DIN2(_52521), .Q(_52368) );
  nor2s1 _53228_inst ( .DIN1(_45596), .DIN2(_46021), .Q(_52520) );
  nnd2s1 _53229_inst ( .DIN1(_52194), .DIN2(_51888), .Q(_52518) );
  nnd2s1 _53230_inst ( .DIN1(_52522), .DIN2(_52523), .Q(_52081) );
  nor2s1 _53231_inst ( .DIN1(_52524), .DIN2(_52525), .Q(_52523) );
  nnd2s1 _53232_inst ( .DIN1(_52526), .DIN2(_52215), .Q(_52525) );
  hi1s1 _53233_inst ( .DIN(_51955), .Q(_52215) );
  nor2s1 _53234_inst ( .DIN1(_52527), .DIN2(_52528), .Q(_51955) );
  nnd2s1 _53235_inst ( .DIN1(_31462), .DIN2(_42797), .Q(_52527) );
  hi1s1 _53236_inst ( .DIN(_33865), .Q(_31462) );
  nnd2s1 _53237_inst ( .DIN1(_51929), .DIN2(_51858), .Q(_52526) );
  hi1s1 _53238_inst ( .DIN(_51795), .Q(_51929) );
  nnd2s1 _53239_inst ( .DIN1(_52495), .DIN2(_42921), .Q(_51795) );
  nnd2s1 _53240_inst ( .DIN1(_52107), .DIN2(_52206), .Q(_52524) );
  nnd2s1 _53241_inst ( .DIN1(_52510), .DIN2(_52409), .Q(_52206) );
  hi1s1 _53242_inst ( .DIN(_42927), .Q(_52510) );
  nnd2s1 _53243_inst ( .DIN1(_52529), .DIN2(_52530), .Q(_42927) );
  nor2s1 _53244_inst ( .DIN1(_52531), .DIN2(_52532), .Q(_52522) );
  or2s1 _53245_inst ( .DIN1(_51938), .DIN2(_52388), .Q(_52532) );
  nnd2s1 _53246_inst ( .DIN1(_52533), .DIN2(_52534), .Q(_52388) );
  nnd2s1 _53247_inst ( .DIN1(_52535), .DIN2(_52536), .Q(_52534) );
  nor2s1 _53248_inst ( .DIN1(_1863), .DIN2(_52537), .Q(_52535) );
  nnd2s1 _53249_inst ( .DIN1(_52538), .DIN2(_52539), .Q(_51938) );
  nor2s1 _53250_inst ( .DIN1(_51972), .DIN2(_52540), .Q(_52539) );
  nor2s1 _53251_inst ( .DIN1(_52541), .DIN2(_52542), .Q(_52540) );
  nnd2s1 _53252_inst ( .DIN1(_51858), .DIN2(_52485), .Q(_52542) );
  hi1s1 _53253_inst ( .DIN(_52132), .Q(_51972) );
  nnd2s1 _53254_inst ( .DIN1(_51809), .DIN2(_26847), .Q(_52132) );
  nor2s1 _53255_inst ( .DIN1(_52543), .DIN2(_52544), .Q(_52538) );
  nor2s1 _53256_inst ( .DIN1(_51796), .DIN2(_52165), .Q(_52544) );
  hi1s1 _53257_inst ( .DIN(_52322), .Q(_52165) );
  nor2s1 _53258_inst ( .DIN1(_51802), .DIN2(_52293), .Q(_52543) );
  nnd2s1 _53259_inst ( .DIN1(_52545), .DIN2(_52546), .Q(_52531) );
  nnd2s1 _53260_inst ( .DIN1(_51930), .DIN2(_51888), .Q(_52546) );
  or2s1 _53261_inst ( .DIN1(_52292), .DIN2(_26848), .Q(_52545) );
  nor2s1 _53262_inst ( .DIN1(_52264), .DIN2(_52303), .Q(_52516) );
  nnd2s1 _53263_inst ( .DIN1(_52024), .DIN2(_52547), .Q(_52303) );
  nnd2s1 _53264_inst ( .DIN1(_52463), .DIN2(_26289), .Q(_52547) );
  nnd2s1 _53265_inst ( .DIN1(_52548), .DIN2(_52549), .Q(_52264) );
  nor2s1 _53266_inst ( .DIN1(_51996), .DIN2(_52550), .Q(_52549) );
  nnd2s1 _53267_inst ( .DIN1(_52040), .DIN2(_51819), .Q(_52550) );
  nnd2s1 _53268_inst ( .DIN1(_52551), .DIN2(_44287), .Q(_52040) );
  and2s1 _53269_inst ( .DIN1(_51970), .DIN2(_51794), .Q(_51996) );
  nor2s1 _53270_inst ( .DIN1(_51851), .DIN2(_52552), .Q(_52548) );
  nnd2s1 _53271_inst ( .DIN1(_52553), .DIN2(_52554), .Q(_52552) );
  nnd2s1 _53272_inst ( .DIN1(_52555), .DIN2(_51802), .Q(_52554) );
  nnd2s1 _53273_inst ( .DIN1(_52213), .DIN2(_52016), .Q(_52555) );
  nnd2s1 _53274_inst ( .DIN1(_52556), .DIN2(_52557), .Q(_52016) );
  nor2s1 _53275_inst ( .DIN1(_44600), .DIN2(_52558), .Q(_52557) );
  nnd2s1 _53276_inst ( .DIN1(_51971), .DIN2(_51818), .Q(_52553) );
  hi1s1 _53277_inst ( .DIN(_52108), .Q(_51971) );
  nnd2s1 _53278_inst ( .DIN1(_52559), .DIN2(_52560), .Q(_52108) );
  nor2s1 _53279_inst ( .DIN1(_52561), .DIN2(_46016), .Q(_52559) );
  nnd2s1 _53280_inst ( .DIN1(_52562), .DIN2(_52563), .Q(_51851) );
  nor2s1 _53281_inst ( .DIN1(_52156), .DIN2(_52564), .Q(_52563) );
  nnd2s1 _53282_inst ( .DIN1(_52399), .DIN2(_52166), .Q(_52564) );
  nnd2s1 _53283_inst ( .DIN1(_52565), .DIN2(_52566), .Q(_52166) );
  nnd2s1 _53284_inst ( .DIN1(_52567), .DIN2(_52568), .Q(_52566) );
  nnd2s1 _53285_inst ( .DIN1(_52569), .DIN2(_41915), .Q(_52568) );
  nor2s1 _53286_inst ( .DIN1(_44316), .DIN2(_26289), .Q(_52569) );
  nnd2s1 _53287_inst ( .DIN1(_52570), .DIN2(_41912), .Q(_52567) );
  nor2s1 _53288_inst ( .DIN1(_51802), .DIN2(_45813), .Q(_52570) );
  nnd2s1 _53289_inst ( .DIN1(_52571), .DIN2(_51888), .Q(_52399) );
  nor2s1 _53290_inst ( .DIN1(_44316), .DIN2(_52494), .Q(_52571) );
  nor2s1 _53291_inst ( .DIN1(_52460), .DIN2(_52572), .Q(_52562) );
  nnd2s1 _53292_inst ( .DIN1(_52182), .DIN2(_52074), .Q(_52572) );
  nnd2s1 _53293_inst ( .DIN1(_52573), .DIN2(_52574), .Q(_52074) );
  nnd2s1 _53294_inst ( .DIN1(_52575), .DIN2(_52576), .Q(_52460) );
  nor2s1 _53295_inst ( .DIN1(_52017), .DIN2(_52577), .Q(_52576) );
  nnd2s1 _53296_inst ( .DIN1(_52195), .DIN2(_52385), .Q(_52577) );
  nnd2s1 _53297_inst ( .DIN1(_51858), .DIN2(_52578), .Q(_52385) );
  or2s1 _53298_inst ( .DIN1(_52579), .DIN2(_26847), .Q(_52195) );
  nnd2s1 _53299_inst ( .DIN1(_52580), .DIN2(_52581), .Q(_52017) );
  nnd2s1 _53300_inst ( .DIN1(_52143), .DIN2(_26847), .Q(_52581) );
  hi1s1 _53301_inst ( .DIN(_52582), .Q(_52143) );
  nnd2s1 _53302_inst ( .DIN1(_52144), .DIN2(_26848), .Q(_52580) );
  nor2s1 _53303_inst ( .DIN1(_52188), .DIN2(_52583), .Q(_52575) );
  nnd2s1 _53304_inst ( .DIN1(_52353), .DIN2(_52584), .Q(_52188) );
  nnd2s1 _53305_inst ( .DIN1(_26848), .DIN2(_52585), .Q(_52584) );
  nnd2s1 _53306_inst ( .DIN1(_52586), .DIN2(_52587), .Q(____0___________0[0])
         );
  nor2s1 _53307_inst ( .DIN1(_52588), .DIN2(_52589), .Q(_52587) );
  nnd2s1 _53308_inst ( .DIN1(_52590), .DIN2(_52591), .Q(_52589) );
  nor2s1 _53309_inst ( .DIN1(_51919), .DIN2(_51853), .Q(_52591) );
  nnd2s1 _53310_inst ( .DIN1(_52592), .DIN2(_52593), .Q(_51853) );
  nor2s1 _53311_inst ( .DIN1(_52147), .DIN2(_52594), .Q(_52593) );
  or2s1 _53312_inst ( .DIN1(_52296), .DIN2(_51913), .Q(_52594) );
  and2s1 _53313_inst ( .DIN1(_52595), .DIN2(_26807), .Q(_51913) );
  nnd2s1 _53314_inst ( .DIN1(_52107), .DIN2(_52024), .Q(_52595) );
  nnd2s1 _53315_inst ( .DIN1(_52596), .DIN2(_42797), .Q(_52024) );
  nnd2s1 _53316_inst ( .DIN1(_52597), .DIN2(_52560), .Q(_52107) );
  nor2s1 _53317_inst ( .DIN1(_45823), .DIN2(_52561), .Q(_52597) );
  nor2s1 _53318_inst ( .DIN1(_52455), .DIN2(_51858), .Q(_52296) );
  and2s1 _53319_inst ( .DIN1(_52253), .DIN2(_52598), .Q(_52455) );
  nnd2s1 _53320_inst ( .DIN1(_52599), .DIN2(_52485), .Q(_52598) );
  nnd2s1 _53321_inst ( .DIN1(_52600), .DIN2(_52601), .Q(_52253) );
  hi1s1 _53322_inst ( .DIN(_52023), .Q(_52147) );
  nnd2s1 _53323_inst ( .DIN1(_52495), .DIN2(_44314), .Q(_52023) );
  hi1s1 _53324_inst ( .DIN(_42924), .Q(_44314) );
  nor2s1 _53325_inst ( .DIN1(_52602), .DIN2(_52603), .Q(_52592) );
  nnd2s1 _53326_inst ( .DIN1(_52604), .DIN2(_52439), .Q(_52603) );
  nnd2s1 _53327_inst ( .DIN1(_52605), .DIN2(_52556), .Q(_52439) );
  nor2s1 _53328_inst ( .DIN1(_43029), .DIN2(_45822), .Q(_52605) );
  nnd2s1 _53329_inst ( .DIN1(_52322), .DIN2(_26848), .Q(_52604) );
  nor2s1 _53330_inst ( .DIN1(_52606), .DIN2(_52607), .Q(_52322) );
  nnd2s1 _53331_inst ( .DIN1(_52608), .DIN2(_46027), .Q(_52606) );
  and2s1 _53332_inst ( .DIN1(_26807), .DIN2(_51964), .Q(_52602) );
  nor2s1 _53333_inst ( .DIN1(_46016), .DIN2(_52609), .Q(_51964) );
  nnd2s1 _53334_inst ( .DIN1(_52610), .DIN2(_52611), .Q(_46016) );
  and2s1 _53335_inst ( .DIN1(_1824), .DIN2(_52612), .Q(_52610) );
  nnd2s1 _53336_inst ( .DIN1(_52613), .DIN2(_52614), .Q(_51919) );
  nnd2s1 _53337_inst ( .DIN1(_51970), .DIN2(_51858), .Q(_52614) );
  and2s1 _53338_inst ( .DIN1(_52615), .DIN2(_52616), .Q(_51970) );
  nor2s1 _53339_inst ( .DIN1(_44600), .DIN2(_44377), .Q(_52616) );
  nor2s1 _53340_inst ( .DIN1(_44658), .DIN2(_46021), .Q(_52615) );
  and2s1 _53341_inst ( .DIN1(_52182), .DIN2(_52053), .Q(_52613) );
  nnd2s1 _53342_inst ( .DIN1(_42921), .DIN2(_52617), .Q(_52053) );
  nnd2s1 _53343_inst ( .DIN1(_52618), .DIN2(_52495), .Q(_52182) );
  nor2s1 _53344_inst ( .DIN1(_26289), .DIN2(_52619), .Q(_52618) );
  nor2s1 _53345_inst ( .DIN1(_52456), .DIN2(_52112), .Q(_52590) );
  nnd2s1 _53346_inst ( .DIN1(_52582), .DIN2(_52172), .Q(_52112) );
  nnd2s1 _53347_inst ( .DIN1(_52620), .DIN2(_52621), .Q(_52172) );
  nor2s1 _53348_inst ( .DIN1(_52622), .DIN2(_52623), .Q(_52621) );
  nnd2s1 _53349_inst ( .DIN1(_52624), .DIN2(_45102), .Q(_52623) );
  nnd2s1 _53350_inst ( .DIN1(_52625), .DIN2(_52626), .Q(_52582) );
  nor2s1 _53351_inst ( .DIN1(_44376), .DIN2(_45814), .Q(_52625) );
  nnd2s1 _53352_inst ( .DIN1(_52627), .DIN2(_52628), .Q(_52456) );
  nor2s1 _53353_inst ( .DIN1(_52629), .DIN2(_52630), .Q(_52628) );
  nnd2s1 _53354_inst ( .DIN1(_52391), .DIN2(_52099), .Q(_52630) );
  nnd2s1 _53355_inst ( .DIN1(_52631), .DIN2(_52600), .Q(_52099) );
  nnd2s1 _53356_inst ( .DIN1(_52632), .DIN2(_52633), .Q(_52391) );
  nor2s1 _53357_inst ( .DIN1(_52634), .DIN2(_52635), .Q(_52633) );
  nnd2s1 _53358_inst ( .DIN1(_52530), .DIN2(_1825), .Q(_52635) );
  nor2s1 _53359_inst ( .DIN1(_52636), .DIN2(_52637), .Q(_52632) );
  hi1s1 _53360_inst ( .DIN(_52600), .Q(_52637) );
  nnd2s1 _53361_inst ( .DIN1(_52638), .DIN2(_51846), .Q(_52629) );
  nnd2s1 _53362_inst ( .DIN1(_52639), .DIN2(_52640), .Q(_51846) );
  and2s1 _53363_inst ( .DIN1(_51281), .DIN2(_52293), .Q(_52638) );
  nnd2s1 _53364_inst ( .DIN1(_52641), .DIN2(_52601), .Q(_52293) );
  nnd2s1 _53365_inst ( .DIN1(_42797), .DIN2(_52642), .Q(_51281) );
  hi1s1 _53366_inst ( .DIN(_45823), .Q(_42797) );
  nor2s1 _53367_inst ( .DIN1(_52643), .DIN2(_52644), .Q(_52627) );
  nnd2s1 _53368_inst ( .DIN1(_52645), .DIN2(_51860), .Q(_52644) );
  nnd2s1 _53369_inst ( .DIN1(_52601), .DIN2(_52485), .Q(_51860) );
  and2s1 _53370_inst ( .DIN1(_52646), .DIN2(_52647), .Q(_52601) );
  hi1s1 _53371_inst ( .DIN(_51948), .Q(_52645) );
  nnd2s1 _53372_inst ( .DIN1(_52292), .DIN2(_52648), .Q(_51948) );
  nnd2s1 _53373_inst ( .DIN1(_52207), .DIN2(_26848), .Q(_52648) );
  hi1s1 _53374_inst ( .DIN(_51967), .Q(_52207) );
  nnd2s1 _53375_inst ( .DIN1(_52649), .DIN2(_52650), .Q(_51967) );
  nor2s1 _53376_inst ( .DIN1(_45407), .DIN2(_44657), .Q(_52650) );
  nor2s1 _53377_inst ( .DIN1(_44376), .DIN2(_52651), .Q(_52649) );
  nnd2s1 _53378_inst ( .DIN1(_52652), .DIN2(_52653), .Q(_52292) );
  nor2s1 _53379_inst ( .DIN1(_52634), .DIN2(_52654), .Q(_52653) );
  nnd2s1 _53380_inst ( .DIN1(_52624), .DIN2(_26438), .Q(_52654) );
  nor2s1 _53381_inst ( .DIN1(_52636), .DIN2(_52655), .Q(_52652) );
  nnd2s1 _53382_inst ( .DIN1(_52064), .DIN2(_52392), .Q(_52643) );
  nnd2s1 _53383_inst ( .DIN1(_52631), .DIN2(_52640), .Q(_52392) );
  nnd2s1 _53384_inst ( .DIN1(_52631), .DIN2(_52485), .Q(_52064) );
  and2s1 _53385_inst ( .DIN1(_52656), .DIN2(_52536), .Q(_52631) );
  nor2s1 _53386_inst ( .DIN1(_26438), .DIN2(_52634), .Q(_52656) );
  nnd2s1 _53387_inst ( .DIN1(_52657), .DIN2(_52658), .Q(_52588) );
  nor2s1 _53388_inst ( .DIN1(_52578), .DIN2(_52659), .Q(_52658) );
  nnd2s1 _53389_inst ( .DIN1(_52173), .DIN2(_52579), .Q(_52659) );
  nnd2s1 _53390_inst ( .DIN1(_52660), .DIN2(_52661), .Q(_52579) );
  nor2s1 _53391_inst ( .DIN1(_52622), .DIN2(_44077), .Q(_52661) );
  nor2s1 _53392_inst ( .DIN1(_52662), .DIN2(_44925), .Q(_52660) );
  nnd2s1 _53393_inst ( .DIN1(_52663), .DIN2(_41915), .Q(_52173) );
  nor2s1 _53394_inst ( .DIN1(_52664), .DIN2(_45813), .Q(_52663) );
  and2s1 _53395_inst ( .DIN1(_52665), .DIN2(_46019), .Q(_52578) );
  nor2s1 _53396_inst ( .DIN1(_52487), .DIN2(_52666), .Q(_46019) );
  nor2s1 _53397_inst ( .DIN1(_52664), .DIN2(_44657), .Q(_52665) );
  nor2s1 _53398_inst ( .DIN1(_52667), .DIN2(_52668), .Q(_52657) );
  nor2s1 _53399_inst ( .DIN1(_51858), .DIN2(_52669), .Q(_52668) );
  nor2s1 _53400_inst ( .DIN1(_52670), .DIN2(_52671), .Q(_52669) );
  hi1s1 _53401_inst ( .DIN(_51861), .Q(_52671) );
  nnd2s1 _53402_inst ( .DIN1(_52672), .DIN2(_44601), .Q(_51861) );
  nor2s1 _53403_inst ( .DIN1(_42924), .DIN2(_52381), .Q(_52670) );
  nnd2s1 _53404_inst ( .DIN1(_52626), .DIN2(_45664), .Q(_52381) );
  nor2s1 _53405_inst ( .DIN1(_44078), .DIN2(_52622), .Q(_52626) );
  nnd2s1 _53406_inst ( .DIN1(_52529), .DIN2(_52673), .Q(_42924) );
  nor2s1 _53407_inst ( .DIN1(_45103), .DIN2(_26414), .Q(_52529) );
  hi1s1 _53408_inst ( .DIN(_52353), .Q(_52667) );
  nnd2s1 _53409_inst ( .DIN1(_46026), .DIN2(_52617), .Q(_52353) );
  hi1s1 _53410_inst ( .DIN(_42923), .Q(_46026) );
  nor2s1 _53411_inst ( .DIN1(_52674), .DIN2(_52675), .Q(_52586) );
  nnd2s1 _53412_inst ( .DIN1(_52676), .DIN2(_52677), .Q(_52675) );
  nor2s1 _53413_inst ( .DIN1(_52512), .DIN2(_52678), .Q(_52677) );
  nnd2s1 _53414_inst ( .DIN1(_52679), .DIN2(_52680), .Q(_52678) );
  nnd2s1 _53415_inst ( .DIN1(_51888), .DIN2(_52681), .Q(_52680) );
  nnd2s1 _53416_inst ( .DIN1(_52213), .DIN2(_52533), .Q(_52681) );
  nnd2s1 _53417_inst ( .DIN1(_52599), .DIN2(_52600), .Q(_52533) );
  nnd2s1 _53418_inst ( .DIN1(_52551), .DIN2(_52682), .Q(_52213) );
  nnd2s1 _53419_inst ( .DIN1(_52683), .DIN2(_51802), .Q(_52679) );
  nor2s1 _53420_inst ( .DIN1(_52684), .DIN2(_52685), .Q(_52683) );
  nnd2s1 _53421_inst ( .DIN1(_41912), .DIN2(_44977), .Q(_52685) );
  nnd2s1 _53422_inst ( .DIN1(_52686), .DIN2(_52687), .Q(_52512) );
  nor2s1 _53423_inst ( .DIN1(_52688), .DIN2(_52689), .Q(_52687) );
  nnd2s1 _53424_inst ( .DIN1(_52690), .DIN2(_52373), .Q(_52689) );
  nnd2s1 _53425_inst ( .DIN1(_52691), .DIN2(_52692), .Q(_52373) );
  nor2s1 _53426_inst ( .DIN1(_52693), .DIN2(_52694), .Q(_52691) );
  nnd2s1 _53427_inst ( .DIN1(_51858), .DIN2(_51852), .Q(_52690) );
  nnd2s1 _53428_inst ( .DIN1(_52695), .DIN2(_52696), .Q(_51852) );
  nnd2s1 _53429_inst ( .DIN1(_52697), .DIN2(_52692), .Q(_52696) );
  nor2s1 _53430_inst ( .DIN1(_1824), .DIN2(_52634), .Q(_52692) );
  nor2s1 _53431_inst ( .DIN1(_52537), .DIN2(_52693), .Q(_52697) );
  nnd2s1 _53432_inst ( .DIN1(_52599), .DIN2(_52640), .Q(_52695) );
  hi1s1 _53433_inst ( .DIN(_52541), .Q(_52599) );
  nnd2s1 _53434_inst ( .DIN1(_52698), .DIN2(_52699), .Q(_52541) );
  nor2s1 _53435_inst ( .DIN1(_1863), .DIN2(_45103), .Q(_52699) );
  nor2s1 _53436_inst ( .DIN1(_52700), .DIN2(_52636), .Q(_52698) );
  hi1s1 _53437_inst ( .DIN(_51794), .Q(_51858) );
  nnd2s1 _53438_inst ( .DIN1(_52015), .DIN2(_52242), .Q(_52688) );
  nnd2s1 _53439_inst ( .DIN1(_46027), .DIN2(_52287), .Q(_52242) );
  nnd2s1 _53440_inst ( .DIN1(_45819), .DIN2(_52409), .Q(_52015) );
  nor2s1 _53441_inst ( .DIN1(_52528), .DIN2(_43029), .Q(_52409) );
  nor2s1 _53442_inst ( .DIN1(_52701), .DIN2(_52702), .Q(_52686) );
  nnd2s1 _53443_inst ( .DIN1(_52117), .DIN2(_52703), .Q(_52702) );
  nnd2s1 _53444_inst ( .DIN1(_51928), .DIN2(_51802), .Q(_52703) );
  hi1s1 _53445_inst ( .DIN(_51803), .Q(_51928) );
  nnd2s1 _53446_inst ( .DIN1(_52596), .DIN2(_44287), .Q(_51803) );
  hi1s1 _53447_inst ( .DIN(_52558), .Q(_44287) );
  and2s1 _53448_inst ( .DIN1(_52704), .DIN2(_52705), .Q(_52117) );
  nor2s1 _53449_inst ( .DIN1(_52706), .DIN2(_52707), .Q(_52705) );
  nnd2s1 _53450_inst ( .DIN1(_52223), .DIN2(_52203), .Q(_52707) );
  nnd2s1 _53451_inst ( .DIN1(_52708), .DIN2(_52709), .Q(_52203) );
  nor2s1 _53452_inst ( .DIN1(_26847), .DIN2(_42923), .Q(_52709) );
  nor2s1 _53453_inst ( .DIN1(_44077), .DIN2(_52684), .Q(_52708) );
  nnd2s1 _53454_inst ( .DIN1(_52240), .DIN2(_26807), .Q(_52223) );
  hi1s1 _53455_inst ( .DIN(_51876), .Q(_52240) );
  nnd2s1 _53456_inst ( .DIN1(_52710), .DIN2(_52511), .Q(_51876) );
  nor2s1 _53457_inst ( .DIN1(_33865), .DIN2(_45822), .Q(_52710) );
  nor2s1 _53458_inst ( .DIN1(_51796), .DIN2(_52201), .Q(_52706) );
  nnd2s1 _53459_inst ( .DIN1(_52573), .DIN2(_44602), .Q(_52201) );
  and2s1 _53460_inst ( .DIN1(_52711), .DIN2(_45818), .Q(_52573) );
  hi1s1 _53461_inst ( .DIN(_52651), .Q(_45818) );
  nnd2s1 _53462_inst ( .DIN1(_52712), .DIN2(_53524), .Q(_52651) );
  nor2s1 _53463_inst ( .DIN1(_44378), .DIN2(_44077), .Q(_52711) );
  nor2s1 _53464_inst ( .DIN1(_52401), .DIN2(_51946), .Q(_52704) );
  nnd2s1 _53465_inst ( .DIN1(_52713), .DIN2(_52714), .Q(_51946) );
  nnd2s1 _53466_inst ( .DIN1(_52092), .DIN2(_26289), .Q(_52714) );
  hi1s1 _53467_inst ( .DIN(_51962), .Q(_52092) );
  nnd2s1 _53468_inst ( .DIN1(_52715), .DIN2(_52511), .Q(_51962) );
  nor2s1 _53469_inst ( .DIN1(_44658), .DIN2(_44929), .Q(_52511) );
  nor2s1 _53470_inst ( .DIN1(_45823), .DIN2(_43029), .Q(_52715) );
  nnd2s1 _53471_inst ( .DIN1(_52716), .DIN2(_46025), .Q(_45823) );
  hi1s1 _53472_inst ( .DIN(_52416), .Q(_46025) );
  nnd2s1 _53473_inst ( .DIN1(_52148), .DIN2(_26848), .Q(_52713) );
  hi1s1 _53474_inst ( .DIN(_51963), .Q(_52148) );
  nnd2s1 _53475_inst ( .DIN1(_44286), .DIN2(_52717), .Q(_51963) );
  hi1s1 _53476_inst ( .DIN(_45814), .Q(_44286) );
  nnd2s1 _53477_inst ( .DIN1(_52718), .DIN2(_52719), .Q(_45814) );
  nor2s1 _53478_inst ( .DIN1(_52416), .DIN2(_52647), .Q(_52719) );
  nor2s1 _53479_inst ( .DIN1(_45103), .DIN2(_26421), .Q(_52718) );
  nnd2s1 _53480_inst ( .DIN1(_52243), .DIN2(_52720), .Q(_52401) );
  nnd2s1 _53481_inst ( .DIN1(_51808), .DIN2(_51802), .Q(_52720) );
  hi1s1 _53482_inst ( .DIN(_52235), .Q(_51808) );
  nnd2s1 _53483_inst ( .DIN1(_52721), .DIN2(_52722), .Q(_52235) );
  nor2s1 _53484_inst ( .DIN1(_44377), .DIN2(_52561), .Q(_52722) );
  nor2s1 _53485_inst ( .DIN1(_43029), .DIN2(_46028), .Q(_52721) );
  nnd2s1 _53486_inst ( .DIN1(_52723), .DIN2(_52724), .Q(_46028) );
  nor2s1 _53487_inst ( .DIN1(_52416), .DIN2(_45103), .Q(_52723) );
  nnd2s1 _53488_inst ( .DIN1(_52725), .DIN2(_52444), .Q(_52243) );
  hi1s1 _53489_inst ( .DIN(_52330), .Q(_52444) );
  nnd2s1 _53490_inst ( .DIN1(_52726), .DIN2(_52574), .Q(_52330) );
  hi1s1 _53491_inst ( .DIN(_52622), .Q(_52574) );
  nor2s1 _53492_inst ( .DIN1(_44378), .DIN2(_44078), .Q(_52726) );
  nor2s1 _53493_inst ( .DIN1(_26289), .DIN2(_52662), .Q(_52725) );
  nnd2s1 _53494_inst ( .DIN1(_52727), .DIN2(_52728), .Q(_52701) );
  nnd2s1 _53495_inst ( .DIN1(_52076), .DIN2(_51818), .Q(_52728) );
  hi1s1 _53496_inst ( .DIN(_51898), .Q(_52076) );
  nnd2s1 _53497_inst ( .DIN1(_52476), .DIN2(_42796), .Q(_51898) );
  and2s1 _53498_inst ( .DIN1(_52560), .DIN2(_41913), .Q(_52476) );
  hi1s1 _53499_inst ( .DIN(_44658), .Q(_41913) );
  nor2s1 _53500_inst ( .DIN1(_33865), .DIN2(_44377), .Q(_52560) );
  nnd2s1 _53501_inst ( .DIN1(_52729), .DIN2(_26807), .Q(_52727) );
  nnd2s1 _53502_inst ( .DIN1(_52080), .DIN2(_51817), .Q(_52729) );
  nnd2s1 _53503_inst ( .DIN1(_52730), .DIN2(_52731), .Q(_51817) );
  nor2s1 _53504_inst ( .DIN1(_52732), .DIN2(_44078), .Q(_52731) );
  nor2s1 _53505_inst ( .DIN1(_44376), .DIN2(_52733), .Q(_52730) );
  nnd2s1 _53506_inst ( .DIN1(_52639), .DIN2(_52600), .Q(_52080) );
  nor2s1 _53507_inst ( .DIN1(_52734), .DIN2(_52735), .Q(_52676) );
  nnd2s1 _53508_inst ( .DIN1(_52736), .DIN2(_52737), .Q(_52735) );
  nnd2s1 _53509_inst ( .DIN1(_52738), .DIN2(_26847), .Q(_52737) );
  nnd2s1 _53510_inst ( .DIN1(_52739), .DIN2(_52740), .Q(_52738) );
  nor2s1 _53511_inst ( .DIN1(_51942), .DIN2(_52741), .Q(_52740) );
  nnd2s1 _53512_inst ( .DIN1(_52360), .DIN2(_52208), .Q(_52741) );
  nnd2s1 _53513_inst ( .DIN1(_52551), .DIN2(_42796), .Q(_52208) );
  hi1s1 _53514_inst ( .DIN(_46021), .Q(_42796) );
  and2s1 _53515_inst ( .DIN1(_52742), .DIN2(_44928), .Q(_52551) );
  nor2s1 _53516_inst ( .DIN1(_44079), .DIN2(_43029), .Q(_52742) );
  nnd2s1 _53517_inst ( .DIN1(_52743), .DIN2(_52647), .Q(_52360) );
  hi1s1 _53518_inst ( .DIN(_52055), .Q(_51942) );
  nnd2s1 _53519_inst ( .DIN1(_52744), .DIN2(_52640), .Q(_52055) );
  hi1s1 _53520_inst ( .DIN(_52655), .Q(_52640) );
  nnd2s1 _53521_inst ( .DIN1(_52745), .DIN2(_1851), .Q(_52655) );
  nor2s1 _53522_inst ( .DIN1(_1853), .DIN2(_26409), .Q(_52745) );
  nor2s1 _53523_inst ( .DIN1(_52585), .DIN2(_52746), .Q(_52739) );
  nnd2s1 _53524_inst ( .DIN1(_52747), .DIN2(_52748), .Q(_52746) );
  nnd2s1 _53525_inst ( .DIN1(_52749), .DIN2(_52565), .Q(_52748) );
  hi1s1 _53526_inst ( .DIN(_52684), .Q(_52565) );
  nor2s1 _53527 ( .DIN1(_44316), .DIN2(_44077), .Q(_52749) );
  nnd2s1 _53528 ( .DIN1(_45098), .DIN2(_52384), .Q(_52747) );
  hi1s1 _53529 ( .DIN(_46022), .Q(_45098) );
  nnd2s1 _53530 ( .DIN1(_52750), .DIN2(_46024), .Q(_46022) );
  nnd2s1 _53531 ( .DIN1(_52751), .DIN2(_52752), .Q(_52585) );
  nnd2s1 _53532 ( .DIN1(_52753), .DIN2(_52754), .Q(_52752) );
  nor2s1 _53533 ( .DIN1(_44378), .DIN2(_44657), .Q(_52754) );
  nor2s1 _53534 ( .DIN1(_52622), .DIN2(_52755), .Q(_52753) );
  nnd2s1 _53535 ( .DIN1(_52756), .DIN2(_46030), .Q(_52751) );
  nor2s1 _53536 ( .DIN1(_52607), .DIN2(_44925), .Q(_52756) );
  nnd2s1 _53537 ( .DIN1(_51796), .DIN2(_52757), .Q(_52736) );
  nnd2s1 _53538 ( .DIN1(_52758), .DIN2(_52759), .Q(_52757) );
  nor2s1 _53539 ( .DIN1(_51809), .DIN2(_52288), .Q(_52759) );
  hi1s1 _53540 ( .DIN(_52458), .Q(_52288) );
  nnd2s1 _53541 ( .DIN1(_52760), .DIN2(_1863), .Q(_52458) );
  and2s1 _53542 ( .DIN1(_52682), .DIN2(_52642), .Q(_51809) );
  hi1s1 _53543 ( .DIN(_45822), .Q(_52682) );
  nor2s1 _53544 ( .DIN1(_51995), .DIN2(_52463), .Q(_52758) );
  hi1s1 _53545 ( .DIN(_52181), .Q(_52463) );
  nnd2s1 _53546 ( .DIN1(_52717), .DIN2(_46029), .Q(_52181) );
  hi1s1 _53547 ( .DIN(_52094), .Q(_51995) );
  nnd2s1 _53548 ( .DIN1(_45819), .DIN2(_52642), .Q(_52094) );
  and2s1 _53549 ( .DIN1(_52521), .DIN2(_44927), .Q(_52642) );
  hi1s1 _53550 ( .DIN(_44377), .Q(_44927) );
  nor2s1 _53551 ( .DIN1(_44600), .DIN2(_44079), .Q(_52521) );
  nnd2s1 _53552 ( .DIN1(_52761), .DIN2(_1852), .Q(_44079) );
  nor2s1 _53553 ( .DIN1(_26652), .DIN2(_26312), .Q(_52761) );
  hi1s1 _53554 ( .DIN(_42928), .Q(_45819) );
  nnd2s1 _53555 ( .DIN1(_52762), .DIN2(_52530), .Q(_42928) );
  nnd2s1 _53556 ( .DIN1(_52763), .DIN2(_52764), .Q(_52734) );
  nnd2s1 _53557 ( .DIN1(_51818), .DIN2(_52765), .Q(_52764) );
  nnd2s1 _53558 ( .DIN1(_52766), .DIN2(_52767), .Q(_52765) );
  hi1s1 _53559 ( .DIN(_51945), .Q(_52767) );
  nnd2s1 _53560 ( .DIN1(_51819), .DIN2(_52174), .Q(_51945) );
  nnd2s1 _53561 ( .DIN1(_52768), .DIN2(_42921), .Q(_52174) );
  nor2s1 _53562 ( .DIN1(_44376), .DIN2(_52607), .Q(_52768) );
  nnd2s1 _53563 ( .DIN1(_52639), .DIN2(_52485), .Q(_51819) );
  and2s1 _53564 ( .DIN1(_52646), .DIN2(_1824), .Q(_52639) );
  nor2s1 _53565 ( .DIN1(_52693), .DIN2(_1863), .Q(_52646) );
  nor2s1 _53566 ( .DIN1(_52131), .DIN2(_52261), .Q(_52766) );
  and2s1 _53567 ( .DIN1(_52744), .DIN2(_52485), .Q(_52261) );
  and2s1 _53568 ( .DIN1(_52769), .DIN2(_52770), .Q(_52744) );
  nor2s1 _53569 ( .DIN1(_1863), .DIN2(_1825), .Q(_52770) );
  nor2s1 _53570 ( .DIN1(_52771), .DIN2(_52636), .Q(_52769) );
  hi1s1 _53571 ( .DIN(_52005), .Q(_52131) );
  nnd2s1 _53572 ( .DIN1(_52772), .DIN2(_52773), .Q(_52005) );
  nor2s1 _53573 ( .DIN1(_44377), .DIN2(_43029), .Q(_52773) );
  nnd2s1 _53574 ( .DIN1(_52774), .DIN2(_1860), .Q(_43029) );
  nor2s1 _53575 ( .DIN1(_52634), .DIN2(_26541), .Q(_52774) );
  nnd2s1 _53576 ( .DIN1(_52775), .DIN2(_1877), .Q(_44377) );
  nor2s1 _53577 ( .DIN1(_53526), .DIN2(_1876), .Q(_52775) );
  nor2s1 _53578 ( .DIN1(_45822), .DIN2(_44658), .Q(_52772) );
  nnd2s1 _53579 ( .DIN1(_45102), .DIN2(_46024), .Q(_45822) );
  nnd2s1 _53580 ( .DIN1(_52776), .DIN2(_26807), .Q(_52763) );
  nnd2s1 _53581 ( .DIN1(_52777), .DIN2(_52778), .Q(_52776) );
  nnd2s1 _53582 ( .DIN1(_46030), .DIN2(_52287), .Q(_52778) );
  nor2s1 _53583 ( .DIN1(_52666), .DIN2(_52416), .Q(_46030) );
  nnd2s1 _53584 ( .DIN1(_1827), .DIN2(_26414), .Q(_52416) );
  nor2s1 _53585 ( .DIN1(_52237), .DIN2(_52779), .Q(_52777) );
  nor2s1 _53586 ( .DIN1(_52780), .DIN2(_52781), .Q(_52779) );
  nnd2s1 _53587 ( .DIN1(_52485), .DIN2(_1827), .Q(_52781) );
  hi1s1 _53588 ( .DIN(_52537), .Q(_52485) );
  nnd2s1 _53589 ( .DIN1(_52782), .DIN2(_1851), .Q(_52537) );
  nor2s1 _53590 ( .DIN1(_1877), .DIN2(_1853), .Q(_52782) );
  and2s1 _53591 ( .DIN1(_52358), .DIN2(_42921), .Q(_52237) );
  hi1s1 _53592 ( .DIN(_52755), .Q(_42921) );
  nnd2s1 _53593 ( .DIN1(_46024), .DIN2(_52612), .Q(_52755) );
  hi1s1 _53594 ( .DIN(_52417), .Q(_46024) );
  nnd2s1 _53595 ( .DIN1(_52783), .DIN2(_1825), .Q(_52417) );
  nor2s1 _53596 ( .DIN1(_53524), .DIN2(_52647), .Q(_52783) );
  nor2s1 _53597 ( .DIN1(_44378), .DIN2(_52607), .Q(_52358) );
  nnd2s1 _53598 ( .DIN1(_52784), .DIN2(_52785), .Q(_52674) );
  nor2s1 _53599 ( .DIN1(_52119), .DIN2(_52440), .Q(_52785) );
  nnd2s1 _53600 ( .DIN1(_52786), .DIN2(_52787), .Q(_52440) );
  nnd2s1 _53601 ( .DIN1(_52194), .DIN2(_51802), .Q(_52787) );
  nor2s1 _53602 ( .DIN1(_46021), .DIN2(_52609), .Q(_52194) );
  nnd2s1 _53603 ( .DIN1(_52788), .DIN2(_44928), .Q(_52609) );
  nor2s1 _53604 ( .DIN1(_44600), .DIN2(_44658), .Q(_52788) );
  nnd2s1 _53605 ( .DIN1(_52789), .DIN2(_1852), .Q(_44658) );
  nor2s1 _53606 ( .DIN1(_1853), .DIN2(_1851), .Q(_52789) );
  nnd2s1 _53607 ( .DIN1(_52762), .DIN2(_52673), .Q(_46021) );
  nor2s1 _53608 ( .DIN1(_1825), .DIN2(_26414), .Q(_52762) );
  nnd2s1 _53609 ( .DIN1(_52356), .DIN2(_26807), .Q(_52786) );
  hi1s1 _53610 ( .DIN(_52193), .Q(_52356) );
  nnd2s1 _53611 ( .DIN1(_52790), .DIN2(_45664), .Q(_52193) );
  nor2s1 _53612 ( .DIN1(_42923), .DIN2(_52607), .Q(_52790) );
  nnd2s1 _53613 ( .DIN1(_44601), .DIN2(_43949), .Q(_52607) );
  hi1s1 _53614 ( .DIN(_45407), .Q(_44601) );
  nnd2s1 _53615 ( .DIN1(_52624), .DIN2(_52612), .Q(_42923) );
  hi1s1 _53616 ( .DIN(_52666), .Q(_52624) );
  nnd2s1 _53617 ( .DIN1(_52791), .DIN2(_1825), .Q(_52666) );
  nor2s1 _53618 ( .DIN1(_53524), .DIN2(_1824), .Q(_52791) );
  nnd2s1 _53619 ( .DIN1(_52792), .DIN2(_52793), .Q(_52119) );
  nor2s1 _53620 ( .DIN1(_52158), .DIN2(_52794), .Q(_52793) );
  or2s1 _53621 ( .DIN1(_52359), .DIN2(_51806), .Q(_52794) );
  hi1s1 _53622 ( .DIN(_52133), .Q(_51806) );
  nnd2s1 _53623 ( .DIN1(_51877), .DIN2(_51794), .Q(_52133) );
  nnd2s1 _53624 ( .DIN1(______[9]), .DIN2(______[16]), .Q(_51794) );
  and2s1 _53625 ( .DIN1(_52556), .DIN2(_52795), .Q(_51877) );
  nor2s1 _53626 ( .DIN1(_33865), .DIN2(_52558), .Q(_52795) );
  nnd2s1 _53627 ( .DIN1(_52796), .DIN2(_52797), .Q(_52558) );
  nor2s1 _53628 ( .DIN1(_52647), .DIN2(_45103), .Q(_52797) );
  nor2s1 _53629 ( .DIN1(_26421), .DIN2(_52487), .Q(_52796) );
  nnd2s1 _53630 ( .DIN1(_52798), .DIN2(_53525), .Q(_33865) );
  nor2s1 _53631 ( .DIN1(_1860), .DIN2(_52634), .Q(_52798) );
  nor2s1 _53632 ( .DIN1(_52561), .DIN2(_44929), .Q(_52556) );
  nnd2s1 _53633 ( .DIN1(_52799), .DIN2(_1876), .Q(_44929) );
  nor2s1 _53634 ( .DIN1(_1877), .DIN2(_26245), .Q(_52799) );
  nor2s1 _53635 ( .DIN1(_52196), .DIN2(_51796), .Q(_52359) );
  hi1s1 _53636 ( .DIN(_26289), .Q(_51796) );
  nnd2s1 _53637 ( .DIN1(_52717), .DIN2(_46027), .Q(_52196) );
  hi1s1 _53638 ( .DIN(_52619), .Q(_46027) );
  nnd2s1 _53639 ( .DIN1(_52800), .DIN2(_52673), .Q(_52619) );
  hi1s1 _53640 ( .DIN(_52771), .Q(_52673) );
  nnd2s1 _53641 ( .DIN1(_52724), .DIN2(_26438), .Q(_52771) );
  hi1s1 _53642 ( .DIN(_45104), .Q(_52724) );
  nnd2s1 _53643 ( .DIN1(_53524), .DIN2(_52647), .Q(_45104) );
  nor2s1 _53644 ( .DIN1(_1826), .DIN2(_45103), .Q(_52800) );
  hi1s1 _53645 ( .DIN(_1825), .Q(_45103) );
  nor2s1 _53646 ( .DIN1(_52684), .DIN2(_44078), .Q(_52717) );
  nnd2s1 _53647 ( .DIN1(_45664), .DIN2(_44602), .Q(_52684) );
  hi1s1 _53648 ( .DIN(_44925), .Q(_45664) );
  hi1s1 _53649 ( .DIN(_52367), .Q(_52158) );
  nnd2s1 _53650 ( .DIN1(_46029), .DIN2(_52617), .Q(_52367) );
  and2s1 _53651 ( .DIN1(_52801), .DIN2(_41912), .Q(_52617) );
  hi1s1 _53652 ( .DIN(_44657), .Q(_41912) );
  nor2s1 _53653 ( .DIN1(_44378), .DIN2(_45407), .Q(_52801) );
  hi1s1 _53654 ( .DIN(_52662), .Q(_46029) );
  nor2s1 _53655 ( .DIN1(_52583), .DIN2(_52802), .Q(_52792) );
  nnd2s1 _53656 ( .DIN1(_52376), .DIN2(_52419), .Q(_52802) );
  nnd2s1 _53657 ( .DIN1(_52156), .DIN2(_26807), .Q(_52419) );
  hi1s1 _53658 ( .DIN(_51966), .Q(_52156) );
  nnd2s1 _53659 ( .DIN1(_52495), .DIN2(_45099), .Q(_51966) );
  hi1s1 _53660 ( .DIN(_44316), .Q(_45099) );
  nnd2s1 _53661 ( .DIN1(_52803), .DIN2(_52530), .Q(_44316) );
  hi1s1 _53662 ( .DIN(_52700), .Q(_52530) );
  nnd2s1 _53663 ( .DIN1(_52804), .DIN2(_53524), .Q(_52700) );
  nor2s1 _53664 ( .DIN1(_1827), .DIN2(_52647), .Q(_52804) );
  nor2s1 _53665 ( .DIN1(_1826), .DIN2(_1825), .Q(_52803) );
  and2s1 _53666 ( .DIN1(_52805), .DIN2(_41915), .Q(_52495) );
  hi1s1 _53667 ( .DIN(_44077), .Q(_41915) );
  nor2s1 _53668 ( .DIN1(_45407), .DIN2(_44376), .Q(_52805) );
  nnd2s1 _53669 ( .DIN1(_52806), .DIN2(_1860), .Q(_45407) );
  nor2s1 _53670 ( .DIN1(_1863), .DIN2(_26541), .Q(_52806) );
  nnd2s1 _53671 ( .DIN1(_52144), .DIN2(_26289), .Q(_52376) );
  and2s1 _53672 ( .DIN1(_52672), .DIN2(_44602), .Q(_52144) );
  hi1s1 _53673 ( .DIN(_52732), .Q(_44602) );
  and2s1 _53674 ( .DIN1(_52620), .DIN2(_44317), .Q(_52672) );
  hi1s1 _53675 ( .DIN(_52733), .Q(_44317) );
  nnd2s1 _53676 ( .DIN1(_52750), .DIN2(_52716), .Q(_52733) );
  nor2s1 _53677 ( .DIN1(_1827), .DIN2(_1826), .Q(_52750) );
  nor2s1 _53678 ( .DIN1(_44077), .DIN2(_44925), .Q(_52620) );
  nnd2s1 _53679 ( .DIN1(_52807), .DIN2(_53526), .Q(_44925) );
  nor2s1 _53680 ( .DIN1(_1877), .DIN2(_1876), .Q(_52807) );
  nnd2s1 _53681 ( .DIN1(_52350), .DIN2(_52808), .Q(_52583) );
  nnd2s1 _53682 ( .DIN1(_52155), .DIN2(_26847), .Q(_52808) );
  nor2s1 _53683 ( .DIN1(_45813), .DIN2(_52494), .Q(_52155) );
  hi1s1 _53684 ( .DIN(_52287), .Q(_52494) );
  nor2s1 _53685 ( .DIN1(_52664), .DIN2(_44078), .Q(_52287) );
  hi1s1 _53686 ( .DIN(_43949), .Q(_44078) );
  nor2s1 _53687 ( .DIN1(_52809), .DIN2(_1852), .Q(_43949) );
  or2s1 _53688 ( .DIN1(_44378), .DIN2(_52732), .Q(_52664) );
  nnd2s1 _53689 ( .DIN1(_52810), .DIN2(_1877), .Q(_44378) );
  nor2s1 _53690 ( .DIN1(_1876), .DIN2(_26245), .Q(_52810) );
  nnd2s1 _53691 ( .DIN1(_52811), .DIN2(_52501), .Q(_52350) );
  nor2s1 _53692 ( .DIN1(_52622), .DIN2(_44376), .Q(_52501) );
  hi1s1 _53693 ( .DIN(_52608), .Q(_44376) );
  nnd2s1 _53694 ( .DIN1(_52812), .DIN2(_53525), .Q(_52622) );
  nor2s1 _53695 ( .DIN1(_1863), .DIN2(_1860), .Q(_52812) );
  nor2s1 _53696 ( .DIN1(_44077), .DIN2(_52662), .Q(_52811) );
  nnd2s1 _53697 ( .DIN1(_52712), .DIN2(_26421), .Q(_52662) );
  and2s1 _53698 ( .DIN1(_52813), .DIN2(_45102), .Q(_52712) );
  nor2s1 _53699 ( .DIN1(_1825), .DIN2(_52647), .Q(_52813) );
  nnd2s1 _53700 ( .DIN1(_52814), .DIN2(_26312), .Q(_44077) );
  nor2s1 _53701 ( .DIN1(_52430), .DIN2(_52310), .Q(_52784) );
  nnd2s1 _53702 ( .DIN1(_52815), .DIN2(_52816), .Q(_52310) );
  nnd2s1 _53703 ( .DIN1(_51930), .DIN2(_51802), .Q(_52816) );
  hi1s1 _53704 ( .DIN(_52429), .Q(_51930) );
  nnd2s1 _53705 ( .DIN1(_52760), .DIN2(_52634), .Q(_52429) );
  and2s1 _53706 ( .DIN1(_52817), .DIN2(_52536), .Q(_52760) );
  hi1s1 _53707 ( .DIN(_52780), .Q(_52536) );
  nnd2s1 _53708 ( .DIN1(_52818), .DIN2(_52611), .Q(_52780) );
  nor2s1 _53709 ( .DIN1(_52647), .DIN2(_52636), .Q(_52818) );
  nor2s1 _53710 ( .DIN1(_1827), .DIN2(_52694), .Q(_52817) );
  hi1s1 _53711 ( .DIN(_52641), .Q(_52694) );
  nor2s1 _53712 ( .DIN1(_52809), .DIN2(_26409), .Q(_52641) );
  or2s1 _53713 ( .DIN1(_52097), .DIN2(_26835), .Q(_52815) );
  nnd2s1 _53714 ( .DIN1(______[16]), .DIN2(_39002), .Q(_51802) );
  nnd2s1 _53715 ( .DIN1(_52743), .DIN2(_1824), .Q(_52097) );
  and2s1 _53716 ( .DIN1(_52819), .DIN2(_52600), .Q(_52743) );
  nor2s1 _53717 ( .DIN1(_52809), .DIN2(_1877), .Q(_52600) );
  nnd2s1 _53718 ( .DIN1(_1853), .DIN2(_26312), .Q(_52809) );
  nor2s1 _53719 ( .DIN1(_52634), .DIN2(_52693), .Q(_52819) );
  nnd2s1 _53720 ( .DIN1(_52820), .DIN2(_52821), .Q(_52693) );
  nor2s1 _53721 ( .DIN1(_1825), .DIN2(_26438), .Q(_52821) );
  nor2s1 _53722 ( .DIN1(_26421), .DIN2(_52636), .Q(_52820) );
  nnd2s1 _53723 ( .DIN1(_52822), .DIN2(_52823), .Q(_52636) );
  nor2s1 _53724 ( .DIN1(_1826), .DIN2(_52824), .Q(_52823) );
  nnd2s1 _53725 ( .DIN1(_26245), .DIN2(_26541), .Q(_52824) );
  nor2s1 _53726 ( .DIN1(_26697), .DIN2(_52481), .Q(_52822) );
  nnd2s1 _53727 ( .DIN1(_1852), .DIN2(_1876), .Q(_52481) );
  hi1s1 _53728 ( .DIN(_1863), .Q(_52634) );
  nnd2s1 _53729 ( .DIN1(_52394), .DIN2(_52095), .Q(_52430) );
  nnd2s1 _53730 ( .DIN1(_52221), .DIN2(_26289), .Q(_52095) );
  hi1s1 _53731 ( .DIN(______[9]), .Q(_39002) );
  hi1s1 _53732 ( .DIN(_51922), .Q(_52221) );
  nnd2s1 _53733 ( .DIN1(_44980), .DIN2(_52596), .Q(_51922) );
  nor2s1 _53734 ( .DIN1(_52528), .DIN2(_44600), .Q(_52596) );
  nnd2s1 _53735 ( .DIN1(_52825), .DIN2(_26697), .Q(_44600) );
  nor2s1 _53736 ( .DIN1(_53525), .DIN2(_1863), .Q(_52825) );
  nnd2s1 _53737 ( .DIN1(_44928), .DIN2(_41914), .Q(_52528) );
  hi1s1 _53738 ( .DIN(_52561), .Q(_41914) );
  nnd2s1 _53739 ( .DIN1(_52826), .DIN2(_1851), .Q(_52561) );
  nor2s1 _53740 ( .DIN1(_1852), .DIN2(_26652), .Q(_52826) );
  hi1s1 _53741 ( .DIN(_45596), .Q(_44928) );
  nnd2s1 _53742 ( .DIN1(_52827), .DIN2(_1876), .Q(_45596) );
  nor2s1 _53743 ( .DIN1(_26245), .DIN2(_26409), .Q(_52827) );
  hi1s1 _53744 ( .DIN(_45812), .Q(_44980) );
  nnd2s1 _53745 ( .DIN1(_45102), .DIN2(_52716), .Q(_45812) );
  hi1s1 _53746 ( .DIN(_52487), .Q(_45102) );
  nnd2s1 _53747 ( .DIN1(_1826), .DIN2(_1827), .Q(_52487) );
  nnd2s1 _53748 ( .DIN1(_52075), .DIN2(_51818), .Q(_52394) );
  and2s1 _53749 ( .DIN1(_52384), .DIN2(_44977), .Q(_52075) );
  hi1s1 _53750 ( .DIN(_45813), .Q(_44977) );
  nnd2s1 _53751 ( .DIN1(_52716), .DIN2(_52612), .Q(_45813) );
  nor2s1 _53752 ( .DIN1(_26414), .DIN2(_1827), .Q(_52612) );
  and2s1 _53753 ( .DIN1(_52611), .DIN2(_52647), .Q(_52716) );
  hi1s1 _53754 ( .DIN(_1824), .Q(_52647) );
  nor2s1 _53755 ( .DIN1(_53524), .DIN2(_1825), .Q(_52611) );
  and2s1 _53756 ( .DIN1(_52828), .DIN2(_52608), .Q(_52384) );
  nor2s1 _53757 ( .DIN1(_52829), .DIN2(_1876), .Q(_52608) );
  nnd2s1 _53758 ( .DIN1(_26245), .DIN2(_26409), .Q(_52829) );
  nor2s1 _53759 ( .DIN1(_52732), .DIN2(_44657), .Q(_52828) );
  nnd2s1 _53760 ( .DIN1(_52814), .DIN2(_1851), .Q(_44657) );
  nor2s1 _53761 ( .DIN1(_1853), .DIN2(_1852), .Q(_52814) );
  nnd2s1 _53762 ( .DIN1(_52830), .DIN2(_1863), .Q(_52732) );
  nor2s1 _53763 ( .DIN1(_53525), .DIN2(_1860), .Q(_52830) );
endmodule

